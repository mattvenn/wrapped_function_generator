magic
tech sky130A
magscale 1 2
timestamp 1646413238
<< viali >>
rect 1869 49249 1903 49283
rect 8125 49249 8159 49283
rect 11989 49249 12023 49283
rect 15761 49249 15795 49283
rect 17877 49249 17911 49283
rect 22017 49249 22051 49283
rect 24409 49249 24443 49283
rect 27629 49249 27663 49283
rect 43177 49249 43211 49283
rect 47041 49249 47075 49283
rect 1409 49181 1443 49215
rect 4261 49181 4295 49215
rect 6561 49181 6595 49215
rect 7481 49181 7515 49215
rect 10977 49181 11011 49215
rect 11529 49181 11563 49215
rect 14933 49181 14967 49215
rect 17141 49181 17175 49215
rect 18153 49181 18187 49215
rect 19349 49181 19383 49215
rect 20177 49181 20211 49215
rect 22293 49181 22327 49215
rect 23857 49181 23891 49215
rect 24685 49181 24719 49215
rect 26433 49181 26467 49215
rect 26985 49181 27019 49215
rect 30021 49181 30055 49215
rect 31033 49181 31067 49215
rect 33793 49181 33827 49215
rect 35633 49181 35667 49215
rect 36277 49181 36311 49215
rect 38117 49181 38151 49215
rect 40785 49181 40819 49215
rect 41613 49181 41647 49215
rect 42441 49181 42475 49215
rect 45201 49181 45235 49215
rect 47777 49181 47811 49215
rect 1593 49113 1627 49147
rect 4629 49113 4663 49147
rect 5181 49113 5215 49147
rect 11713 49113 11747 49147
rect 27169 49113 27203 49147
rect 42625 49113 42659 49147
rect 45385 49113 45419 49147
rect 5273 49045 5307 49079
rect 6745 49045 6779 49079
rect 10149 49045 10183 49079
rect 15025 49045 15059 49079
rect 17233 49045 17267 49079
rect 19533 49045 19567 49079
rect 20269 49045 20303 49079
rect 30113 49045 30147 49079
rect 32137 49045 32171 49079
rect 38301 49045 38335 49079
rect 40877 49045 40911 49079
rect 41797 49045 41831 49079
rect 47869 49045 47903 49079
rect 5549 48773 5583 48807
rect 14749 48773 14783 48807
rect 31585 48773 31619 48807
rect 47961 48773 47995 48807
rect 1409 48705 1443 48739
rect 2329 48705 2363 48739
rect 6745 48705 6779 48739
rect 11621 48705 11655 48739
rect 12357 48705 12391 48739
rect 19257 48705 19291 48739
rect 25973 48705 26007 48739
rect 27445 48705 27479 48739
rect 29745 48705 29779 48739
rect 32137 48705 32171 48739
rect 34897 48705 34931 48739
rect 42441 48705 42475 48739
rect 43269 48705 43303 48739
rect 43729 48705 43763 48739
rect 46765 48705 46799 48739
rect 1593 48637 1627 48671
rect 3157 48637 3191 48671
rect 3341 48637 3375 48671
rect 4169 48637 4203 48671
rect 6929 48637 6963 48671
rect 7205 48637 7239 48671
rect 9137 48637 9171 48671
rect 9321 48637 9355 48671
rect 10517 48637 10551 48671
rect 12541 48637 12575 48671
rect 12817 48637 12851 48671
rect 16129 48637 16163 48671
rect 16681 48637 16715 48671
rect 16865 48637 16899 48671
rect 17141 48637 17175 48671
rect 19441 48637 19475 48671
rect 20729 48637 20763 48671
rect 22109 48637 22143 48671
rect 22569 48637 22603 48671
rect 22753 48637 22787 48671
rect 23489 48637 23523 48671
rect 25513 48637 25547 48671
rect 27629 48637 27663 48671
rect 27905 48637 27939 48671
rect 29929 48637 29963 48671
rect 32321 48637 32355 48671
rect 32873 48637 32907 48671
rect 35081 48637 35115 48671
rect 36093 48637 36127 48671
rect 38853 48637 38887 48671
rect 39313 48637 39347 48671
rect 39497 48637 39531 48671
rect 40049 48637 40083 48671
rect 44465 48637 44499 48671
rect 44649 48637 44683 48671
rect 45845 48637 45879 48671
rect 2513 48569 2547 48603
rect 5641 48501 5675 48535
rect 11805 48501 11839 48535
rect 14841 48501 14875 48535
rect 26157 48501 26191 48535
rect 41889 48501 41923 48535
rect 42533 48501 42567 48535
rect 43913 48501 43947 48535
rect 46949 48501 46983 48535
rect 48053 48501 48087 48535
rect 3985 48297 4019 48331
rect 7113 48297 7147 48331
rect 9321 48297 9355 48331
rect 16865 48297 16899 48331
rect 39957 48297 39991 48331
rect 45109 48297 45143 48331
rect 19441 48229 19475 48263
rect 41337 48229 41371 48263
rect 2789 48161 2823 48195
rect 4721 48161 4755 48195
rect 10149 48161 10183 48195
rect 10609 48161 10643 48195
rect 14933 48161 14967 48195
rect 22569 48161 22603 48195
rect 24409 48161 24443 48195
rect 24869 48161 24903 48195
rect 28365 48161 28399 48195
rect 29561 48161 29595 48195
rect 30021 48161 30055 48195
rect 32321 48161 32355 48195
rect 36001 48161 36035 48195
rect 36737 48161 36771 48195
rect 41797 48161 41831 48195
rect 42533 48161 42567 48195
rect 46305 48161 46339 48195
rect 46857 48161 46891 48195
rect 1409 48093 1443 48127
rect 7021 48093 7055 48127
rect 7849 48093 7883 48127
rect 13093 48093 13127 48127
rect 14473 48093 14507 48127
rect 16773 48093 16807 48127
rect 21373 48093 21407 48127
rect 21833 48093 21867 48127
rect 27157 48093 27191 48127
rect 31861 48093 31895 48127
rect 35449 48093 35483 48127
rect 39865 48093 39899 48127
rect 44097 48093 44131 48127
rect 45017 48093 45051 48127
rect 45661 48093 45695 48127
rect 1593 48025 1627 48059
rect 4905 48025 4939 48059
rect 6561 48025 6595 48059
rect 10333 48025 10367 48059
rect 14657 48025 14691 48059
rect 22017 48025 22051 48059
rect 24593 48025 24627 48059
rect 27353 48025 27387 48059
rect 29745 48025 29779 48059
rect 32045 48025 32079 48059
rect 36185 48025 36219 48059
rect 41981 48025 42015 48059
rect 46489 48025 46523 48059
rect 13185 47957 13219 47991
rect 35449 47957 35483 47991
rect 44281 47957 44315 47991
rect 45753 47957 45787 47991
rect 3249 47753 3283 47787
rect 4169 47753 4203 47787
rect 10241 47753 10275 47787
rect 10885 47753 10919 47787
rect 13369 47753 13403 47787
rect 14381 47753 14415 47787
rect 18613 47753 18647 47787
rect 22293 47753 22327 47787
rect 22937 47753 22971 47787
rect 24225 47753 24259 47787
rect 26341 47753 26375 47787
rect 27353 47753 27387 47787
rect 30573 47753 30607 47787
rect 31217 47753 31251 47787
rect 32229 47753 32263 47787
rect 35909 47753 35943 47787
rect 36553 47753 36587 47787
rect 41797 47753 41831 47787
rect 2605 47685 2639 47719
rect 6837 47685 6871 47719
rect 7573 47685 7607 47719
rect 17785 47685 17819 47719
rect 32965 47685 32999 47719
rect 33701 47685 33735 47719
rect 42625 47685 42659 47719
rect 1869 47617 1903 47651
rect 2513 47617 2547 47651
rect 3157 47617 3191 47651
rect 4077 47617 4111 47651
rect 4905 47617 4939 47651
rect 5549 47617 5583 47651
rect 6745 47617 6779 47651
rect 7389 47617 7423 47651
rect 10149 47617 10183 47651
rect 10793 47617 10827 47651
rect 11529 47617 11563 47651
rect 13277 47617 13311 47651
rect 14289 47617 14323 47651
rect 15485 47617 15519 47651
rect 17509 47617 17543 47651
rect 18521 47617 18555 47651
rect 22201 47617 22235 47651
rect 22845 47617 22879 47651
rect 24133 47617 24167 47651
rect 24961 47617 24995 47651
rect 25513 47617 25547 47651
rect 26249 47617 26283 47651
rect 27261 47617 27295 47651
rect 28181 47617 28215 47651
rect 30481 47617 30515 47651
rect 31125 47617 31159 47651
rect 32137 47617 32171 47651
rect 32873 47617 32907 47651
rect 33517 47617 33551 47651
rect 35817 47617 35851 47651
rect 36461 47617 36495 47651
rect 41705 47617 41739 47651
rect 42441 47617 42475 47651
rect 47869 47617 47903 47651
rect 7849 47549 7883 47583
rect 12357 47549 12391 47583
rect 25697 47549 25731 47583
rect 28365 47549 28399 47583
rect 28641 47549 28675 47583
rect 34713 47549 34747 47583
rect 44005 47549 44039 47583
rect 44741 47549 44775 47583
rect 44925 47549 44959 47583
rect 45201 47549 45235 47583
rect 2053 47481 2087 47515
rect 4997 47413 5031 47447
rect 5641 47413 5675 47447
rect 48053 47413 48087 47447
rect 1777 47209 1811 47243
rect 3985 47209 4019 47243
rect 25421 47209 25455 47243
rect 26065 47209 26099 47243
rect 26893 47209 26927 47243
rect 27905 47209 27939 47243
rect 29653 47209 29687 47243
rect 30481 47209 30515 47243
rect 45109 47209 45143 47243
rect 45753 47209 45787 47243
rect 4813 47073 4847 47107
rect 4997 47073 5031 47107
rect 5549 47073 5583 47107
rect 28549 47073 28583 47107
rect 42625 47073 42659 47107
rect 44465 47073 44499 47107
rect 46765 47073 46799 47107
rect 2237 47005 2271 47039
rect 3065 47005 3099 47039
rect 10241 47005 10275 47039
rect 10517 47005 10551 47039
rect 25605 47005 25639 47039
rect 26249 47005 26283 47039
rect 27813 47005 27847 47039
rect 28457 47005 28491 47039
rect 29561 47005 29595 47039
rect 45017 47005 45051 47039
rect 45661 47005 45695 47039
rect 46305 47005 46339 47039
rect 11161 46937 11195 46971
rect 12909 46937 12943 46971
rect 42809 46937 42843 46971
rect 46489 46937 46523 46971
rect 2329 46869 2363 46903
rect 10885 46665 10919 46699
rect 13185 46665 13219 46699
rect 47685 46665 47719 46699
rect 11897 46597 11931 46631
rect 1777 46529 1811 46563
rect 10701 46529 10735 46563
rect 43177 46529 43211 46563
rect 44005 46529 44039 46563
rect 44649 46529 44683 46563
rect 47593 46529 47627 46563
rect 1961 46461 1995 46495
rect 2789 46461 2823 46495
rect 38117 46461 38151 46495
rect 38301 46461 38335 46495
rect 38669 46461 38703 46495
rect 45201 46461 45235 46495
rect 45385 46461 45419 46495
rect 46857 46461 46891 46495
rect 4261 46325 4295 46359
rect 38485 46121 38519 46155
rect 44465 46121 44499 46155
rect 45293 46121 45327 46155
rect 1409 45985 1443 46019
rect 1593 45985 1627 46019
rect 2789 45985 2823 46019
rect 48145 45985 48179 46019
rect 11161 45917 11195 45951
rect 38393 45917 38427 45951
rect 45201 45917 45235 45951
rect 46305 45917 46339 45951
rect 11897 45849 11931 45883
rect 46489 45849 46523 45883
rect 46949 45509 46983 45543
rect 1409 45441 1443 45475
rect 2237 45441 2271 45475
rect 46857 45441 46891 45475
rect 47593 45441 47627 45475
rect 45109 45373 45143 45407
rect 45753 45373 45787 45407
rect 46397 45373 46431 45407
rect 47685 45373 47719 45407
rect 1593 45305 1627 45339
rect 2421 45237 2455 45271
rect 2237 45033 2271 45067
rect 45845 45033 45879 45067
rect 31953 44897 31987 44931
rect 33793 44897 33827 44931
rect 48145 44897 48179 44931
rect 1409 44829 1443 44863
rect 2145 44829 2179 44863
rect 2973 44829 3007 44863
rect 17049 44829 17083 44863
rect 46305 44829 46339 44863
rect 32137 44761 32171 44795
rect 46489 44761 46523 44795
rect 1593 44693 1627 44727
rect 17233 44693 17267 44727
rect 47685 44489 47719 44523
rect 2053 44353 2087 44387
rect 47041 44353 47075 44387
rect 47593 44353 47627 44387
rect 2237 44285 2271 44319
rect 3065 44285 3099 44319
rect 2973 43945 3007 43979
rect 1409 43741 1443 43775
rect 2881 43741 2915 43775
rect 36369 43741 36403 43775
rect 47317 43741 47351 43775
rect 48145 43741 48179 43775
rect 1685 43673 1719 43707
rect 36553 43673 36587 43707
rect 38209 43673 38243 43707
rect 47409 43605 47443 43639
rect 36553 43401 36587 43435
rect 36461 43265 36495 43299
rect 47869 43265 47903 43299
rect 48053 43061 48087 43095
rect 46489 42721 46523 42755
rect 48145 42721 48179 42755
rect 46305 42653 46339 42687
rect 47961 42177 47995 42211
rect 48145 42041 48179 42075
rect 2053 41973 2087 42007
rect 47041 41973 47075 42007
rect 1409 41633 1443 41667
rect 1869 41633 1903 41667
rect 46305 41633 46339 41667
rect 1593 41497 1627 41531
rect 46489 41497 46523 41531
rect 48145 41497 48179 41531
rect 2237 41225 2271 41259
rect 46857 41225 46891 41259
rect 1409 41089 1443 41123
rect 2145 41089 2179 41123
rect 46765 41089 46799 41123
rect 47869 41089 47903 41123
rect 1593 40885 1627 40919
rect 48053 40885 48087 40919
rect 46305 40545 46339 40579
rect 1869 40409 1903 40443
rect 2053 40409 2087 40443
rect 46489 40409 46523 40443
rect 48145 40409 48179 40443
rect 47041 40001 47075 40035
rect 47593 40001 47627 40035
rect 47685 40001 47719 40035
rect 2053 39797 2087 39831
rect 1409 39457 1443 39491
rect 2789 39457 2823 39491
rect 6837 39389 6871 39423
rect 7481 39389 7515 39423
rect 24685 39389 24719 39423
rect 24777 39389 24811 39423
rect 24869 39389 24903 39423
rect 25053 39389 25087 39423
rect 47317 39389 47351 39423
rect 47593 39389 47627 39423
rect 1593 39321 1627 39355
rect 7573 39253 7607 39287
rect 24409 39253 24443 39287
rect 2145 39049 2179 39083
rect 6837 38981 6871 39015
rect 21097 38981 21131 39015
rect 2053 38913 2087 38947
rect 6653 38913 6687 38947
rect 20913 38913 20947 38947
rect 24205 38913 24239 38947
rect 7113 38845 7147 38879
rect 23949 38845 23983 38879
rect 21281 38709 21315 38743
rect 25329 38709 25363 38743
rect 47777 38709 47811 38743
rect 46305 38369 46339 38403
rect 48145 38369 48179 38403
rect 20729 38301 20763 38335
rect 20818 38301 20852 38335
rect 20913 38301 20947 38335
rect 21097 38301 21131 38335
rect 21557 38301 21591 38335
rect 24409 38301 24443 38335
rect 24676 38301 24710 38335
rect 26985 38301 27019 38335
rect 20453 38233 20487 38267
rect 21802 38233 21836 38267
rect 27230 38233 27264 38267
rect 46489 38233 46523 38267
rect 22937 38165 22971 38199
rect 25789 38165 25823 38199
rect 28365 38165 28399 38199
rect 21833 37961 21867 37995
rect 24041 37961 24075 37995
rect 26341 37961 26375 37995
rect 46949 37961 46983 37995
rect 29929 37893 29963 37927
rect 30145 37893 30179 37927
rect 47961 37893 47995 37927
rect 19349 37825 19383 37859
rect 19533 37825 19567 37859
rect 20913 37825 20947 37859
rect 21005 37825 21039 37859
rect 21097 37825 21131 37859
rect 21281 37825 21315 37859
rect 22201 37825 22235 37859
rect 24317 37825 24351 37859
rect 24406 37831 24440 37865
rect 24501 37825 24535 37859
rect 24685 37825 24719 37859
rect 25145 37825 25179 37859
rect 25329 37825 25363 37859
rect 25973 37825 26007 37859
rect 26157 37825 26191 37859
rect 27537 37825 27571 37859
rect 27804 37825 27838 37859
rect 46857 37825 46891 37859
rect 1409 37757 1443 37791
rect 1685 37757 1719 37791
rect 22293 37757 22327 37791
rect 22477 37757 22511 37791
rect 25513 37757 25547 37791
rect 19717 37621 19751 37655
rect 20637 37621 20671 37655
rect 28917 37621 28951 37655
rect 30113 37621 30147 37655
rect 30297 37621 30331 37655
rect 48053 37621 48087 37655
rect 19625 37417 19659 37451
rect 24961 37417 24995 37451
rect 26709 37417 26743 37451
rect 32413 37417 32447 37451
rect 20177 37281 20211 37315
rect 25513 37281 25547 37315
rect 28365 37281 28399 37315
rect 18337 37213 18371 37247
rect 18426 37210 18460 37244
rect 18521 37213 18555 37247
rect 18705 37213 18739 37247
rect 20821 37213 20855 37247
rect 21088 37213 21122 37247
rect 26939 37213 26973 37247
rect 27058 37213 27092 37247
rect 27169 37213 27203 37247
rect 27353 37213 27387 37247
rect 29561 37213 29595 37247
rect 31953 37213 31987 37247
rect 47685 37213 47719 37247
rect 1869 37145 1903 37179
rect 2053 37145 2087 37179
rect 25329 37145 25363 37179
rect 29828 37145 29862 37179
rect 32229 37145 32263 37179
rect 18061 37077 18095 37111
rect 19993 37077 20027 37111
rect 20085 37077 20119 37111
rect 22201 37077 22235 37111
rect 25421 37077 25455 37111
rect 27813 37077 27847 37111
rect 28181 37077 28215 37111
rect 28273 37077 28307 37111
rect 30941 37077 30975 37111
rect 32429 37077 32463 37111
rect 32597 37077 32631 37111
rect 22201 36873 22235 36907
rect 24685 36873 24719 36907
rect 27629 36873 27663 36907
rect 29193 36873 29227 36907
rect 25053 36805 25087 36839
rect 26065 36805 26099 36839
rect 28825 36805 28859 36839
rect 18317 36737 18351 36771
rect 20453 36737 20487 36771
rect 20637 36737 20671 36771
rect 21833 36737 21867 36771
rect 22017 36737 22051 36771
rect 25145 36737 25179 36771
rect 26249 36737 26283 36771
rect 27997 36737 28031 36771
rect 28089 36737 28123 36771
rect 29009 36737 29043 36771
rect 29745 36737 29779 36771
rect 30012 36737 30046 36771
rect 32393 36737 32427 36771
rect 47593 36737 47627 36771
rect 18061 36669 18095 36703
rect 25329 36669 25363 36703
rect 28181 36669 28215 36703
rect 32137 36669 32171 36703
rect 2237 36533 2271 36567
rect 19441 36533 19475 36567
rect 20821 36533 20855 36567
rect 26433 36533 26467 36567
rect 31125 36533 31159 36567
rect 33517 36533 33551 36567
rect 47685 36533 47719 36567
rect 22477 36329 22511 36363
rect 27905 36329 27939 36363
rect 29837 36329 29871 36363
rect 31217 36329 31251 36363
rect 31953 36329 31987 36363
rect 30665 36261 30699 36295
rect 19625 36193 19659 36227
rect 20637 36193 20671 36227
rect 23029 36193 23063 36227
rect 24777 36193 24811 36227
rect 26893 36193 26927 36227
rect 30113 36193 30147 36227
rect 30297 36193 30331 36227
rect 32321 36193 32355 36227
rect 32413 36193 32447 36227
rect 46305 36193 46339 36227
rect 46489 36193 46523 36227
rect 48145 36193 48179 36227
rect 2789 36125 2823 36159
rect 18337 36125 18371 36159
rect 18429 36125 18463 36159
rect 18521 36125 18555 36159
rect 18705 36125 18739 36159
rect 26617 36125 26651 36159
rect 28181 36125 28215 36159
rect 28273 36125 28307 36159
rect 28365 36125 28399 36159
rect 28549 36125 28583 36159
rect 30021 36125 30055 36159
rect 30205 36125 30239 36159
rect 32137 36125 32171 36159
rect 32229 36125 32263 36159
rect 19257 36057 19291 36091
rect 19441 36057 19475 36091
rect 20882 36057 20916 36091
rect 25022 36057 25056 36091
rect 31033 36057 31067 36091
rect 31233 36057 31267 36091
rect 2881 35989 2915 36023
rect 18061 35989 18095 36023
rect 22017 35989 22051 36023
rect 22845 35989 22879 36023
rect 22937 35989 22971 36023
rect 26157 35989 26191 36023
rect 31401 35989 31435 36023
rect 20085 35785 20119 35819
rect 22109 35785 22143 35819
rect 24593 35785 24627 35819
rect 26985 35785 27019 35819
rect 30113 35785 30147 35819
rect 2145 35717 2179 35751
rect 22569 35717 22603 35751
rect 26065 35717 26099 35751
rect 28457 35717 28491 35751
rect 47961 35717 47995 35751
rect 1961 35649 1995 35683
rect 18153 35649 18187 35683
rect 18409 35649 18443 35683
rect 20315 35649 20349 35683
rect 20434 35649 20468 35683
rect 20545 35649 20579 35683
rect 20729 35649 20763 35683
rect 22477 35649 22511 35683
rect 23397 35649 23431 35683
rect 24869 35649 24903 35683
rect 24961 35649 24995 35683
rect 25053 35649 25087 35683
rect 25237 35649 25271 35683
rect 26249 35649 26283 35683
rect 27353 35649 27387 35683
rect 28273 35649 28307 35683
rect 29009 35649 29043 35683
rect 29285 35649 29319 35683
rect 30297 35649 30331 35683
rect 30389 35649 30423 35683
rect 30573 35649 30607 35683
rect 32393 35649 32427 35683
rect 46765 35649 46799 35683
rect 2789 35581 2823 35615
rect 22661 35581 22695 35615
rect 23581 35581 23615 35615
rect 26433 35581 26467 35615
rect 27445 35581 27479 35615
rect 27537 35581 27571 35615
rect 29193 35581 29227 35615
rect 30481 35581 30515 35615
rect 32137 35581 32171 35615
rect 48145 35513 48179 35547
rect 19533 35445 19567 35479
rect 29285 35445 29319 35479
rect 29469 35445 29503 35479
rect 33517 35445 33551 35479
rect 46305 35445 46339 35479
rect 46857 35445 46891 35479
rect 19441 35241 19475 35275
rect 21005 35241 21039 35275
rect 24685 35241 24719 35275
rect 25513 35241 25547 35275
rect 29561 35241 29595 35275
rect 30573 35241 30607 35275
rect 31953 35241 31987 35275
rect 21833 35173 21867 35207
rect 2053 35105 2087 35139
rect 20085 35105 20119 35139
rect 24501 35105 24535 35139
rect 32229 35105 32263 35139
rect 46305 35105 46339 35139
rect 46489 35105 46523 35139
rect 48145 35105 48179 35139
rect 2697 35037 2731 35071
rect 24685 35037 24719 35071
rect 25421 35037 25455 35071
rect 29561 35037 29595 35071
rect 29745 35037 29779 35071
rect 32137 35037 32171 35071
rect 32321 35037 32355 35071
rect 32413 35037 32447 35071
rect 1869 34969 1903 35003
rect 19809 34969 19843 35003
rect 20913 34969 20947 35003
rect 21649 34969 21683 35003
rect 24409 34969 24443 35003
rect 30389 34969 30423 35003
rect 30589 34969 30623 35003
rect 19901 34901 19935 34935
rect 24869 34901 24903 34935
rect 29929 34901 29963 34935
rect 30757 34901 30791 34935
rect 23581 34697 23615 34731
rect 24409 34697 24443 34731
rect 28733 34697 28767 34731
rect 32521 34697 32555 34731
rect 32689 34697 32723 34731
rect 1961 34629 1995 34663
rect 32321 34629 32355 34663
rect 1777 34561 1811 34595
rect 19717 34561 19751 34595
rect 20361 34561 20395 34595
rect 20545 34561 20579 34595
rect 22201 34561 22235 34595
rect 22468 34561 22502 34595
rect 24501 34561 24535 34595
rect 25513 34561 25547 34595
rect 25789 34561 25823 34595
rect 28273 34561 28307 34595
rect 28549 34561 28583 34595
rect 29193 34561 29227 34595
rect 29469 34561 29503 34595
rect 30849 34561 30883 34595
rect 30941 34561 30975 34595
rect 46765 34561 46799 34595
rect 2789 34493 2823 34527
rect 20729 34493 20763 34527
rect 24593 34493 24627 34527
rect 25605 34493 25639 34527
rect 28365 34493 28399 34527
rect 30665 34493 30699 34527
rect 30757 34493 30791 34527
rect 19809 34357 19843 34391
rect 24041 34357 24075 34391
rect 25513 34357 25547 34391
rect 25973 34357 26007 34391
rect 28273 34357 28307 34391
rect 30481 34357 30515 34391
rect 32505 34357 32539 34391
rect 46857 34357 46891 34391
rect 47777 34357 47811 34391
rect 20453 34153 20487 34187
rect 22017 34153 22051 34187
rect 24777 34153 24811 34187
rect 20913 34017 20947 34051
rect 21097 34017 21131 34051
rect 23857 34017 23891 34051
rect 28089 34017 28123 34051
rect 29561 34017 29595 34051
rect 32045 34017 32079 34051
rect 46305 34017 46339 34051
rect 46489 34017 46523 34051
rect 48145 34017 48179 34051
rect 19625 33949 19659 33983
rect 22293 33949 22327 33983
rect 22382 33943 22416 33977
rect 22498 33949 22532 33983
rect 22661 33949 22695 33983
rect 23489 33949 23523 33983
rect 25421 33949 25455 33983
rect 25605 33949 25639 33983
rect 25789 33949 25823 33983
rect 25973 33949 26007 33983
rect 26709 33949 26743 33983
rect 27905 33949 27939 33983
rect 29828 33949 29862 33983
rect 31769 33949 31803 33983
rect 19809 33881 19843 33915
rect 20821 33881 20855 33915
rect 23673 33881 23707 33915
rect 24685 33881 24719 33915
rect 26893 33881 26927 33915
rect 1869 33813 1903 33847
rect 19993 33813 20027 33847
rect 25881 33813 25915 33847
rect 27077 33813 27111 33847
rect 27537 33813 27571 33847
rect 27997 33813 28031 33847
rect 30941 33813 30975 33847
rect 20545 33609 20579 33643
rect 23305 33609 23339 33643
rect 25697 33609 25731 33643
rect 26249 33609 26283 33643
rect 28365 33609 28399 33643
rect 31125 33609 31159 33643
rect 21833 33541 21867 33575
rect 25605 33541 25639 33575
rect 32321 33541 32355 33575
rect 1777 33473 1811 33507
rect 18061 33473 18095 33507
rect 18328 33473 18362 33507
rect 20913 33473 20947 33507
rect 22109 33473 22143 33507
rect 22201 33473 22235 33507
rect 22293 33473 22327 33507
rect 22477 33473 22511 33507
rect 22937 33473 22971 33507
rect 24685 33473 24719 33507
rect 24777 33473 24811 33507
rect 26433 33473 26467 33507
rect 26985 33473 27019 33507
rect 27241 33473 27275 33507
rect 29653 33473 29687 33507
rect 31033 33473 31067 33507
rect 32137 33473 32171 33507
rect 46489 33473 46523 33507
rect 1961 33405 1995 33439
rect 2789 33405 2823 33439
rect 21005 33405 21039 33439
rect 21189 33405 21223 33439
rect 23029 33405 23063 33439
rect 24869 33405 24903 33439
rect 29377 33405 29411 33439
rect 46213 33405 46247 33439
rect 19441 33269 19475 33303
rect 23121 33269 23155 33303
rect 24317 33269 24351 33303
rect 32505 33269 32539 33303
rect 47777 33269 47811 33303
rect 2145 33065 2179 33099
rect 20545 33065 20579 33099
rect 20729 33065 20763 33099
rect 23029 33065 23063 33099
rect 26801 33065 26835 33099
rect 30297 33065 30331 33099
rect 30481 33065 30515 33099
rect 25789 32997 25823 33031
rect 16037 32929 16071 32963
rect 20361 32929 20395 32963
rect 21189 32929 21223 32963
rect 24409 32929 24443 32963
rect 28825 32929 28859 32963
rect 30205 32929 30239 32963
rect 31677 32929 31711 32963
rect 32597 32929 32631 32963
rect 46305 32929 46339 32963
rect 48053 32929 48087 32963
rect 1593 32861 1627 32895
rect 2053 32861 2087 32895
rect 2697 32861 2731 32895
rect 15577 32861 15611 32895
rect 20269 32861 20303 32895
rect 20545 32861 20579 32895
rect 21465 32861 21499 32895
rect 22661 32861 22695 32895
rect 23673 32861 23707 32895
rect 27077 32861 27111 32895
rect 27169 32861 27203 32895
rect 27261 32861 27295 32895
rect 27445 32861 27479 32895
rect 28733 32861 28767 32895
rect 30113 32861 30147 32895
rect 31493 32861 31527 32895
rect 36093 32861 36127 32895
rect 15761 32793 15795 32827
rect 19625 32793 19659 32827
rect 22845 32793 22879 32827
rect 23489 32793 23523 32827
rect 24654 32793 24688 32827
rect 31585 32793 31619 32827
rect 32842 32793 32876 32827
rect 46489 32793 46523 32827
rect 2789 32725 2823 32759
rect 19717 32725 19751 32759
rect 23857 32725 23891 32759
rect 28273 32725 28307 32759
rect 28641 32725 28675 32759
rect 31125 32725 31159 32759
rect 33977 32725 34011 32759
rect 36277 32725 36311 32759
rect 15669 32521 15703 32555
rect 19625 32521 19659 32555
rect 23213 32521 23247 32555
rect 24317 32521 24351 32555
rect 24685 32521 24719 32555
rect 24777 32521 24811 32555
rect 28733 32521 28767 32555
rect 30849 32521 30883 32555
rect 33977 32521 34011 32555
rect 36461 32521 36495 32555
rect 2145 32453 2179 32487
rect 19533 32453 19567 32487
rect 22569 32453 22603 32487
rect 22753 32453 22787 32487
rect 39129 32453 39163 32487
rect 1961 32385 1995 32419
rect 15577 32385 15611 32419
rect 18245 32385 18279 32419
rect 18429 32385 18463 32419
rect 20453 32385 20487 32419
rect 20545 32385 20579 32419
rect 20637 32385 20671 32419
rect 20821 32385 20855 32419
rect 21833 32385 21867 32419
rect 23469 32385 23503 32419
rect 23581 32385 23615 32419
rect 23673 32388 23707 32422
rect 23857 32385 23891 32419
rect 25605 32385 25639 32419
rect 26433 32385 26467 32419
rect 27353 32385 27387 32419
rect 27609 32385 27643 32419
rect 31217 32385 31251 32419
rect 32597 32385 32631 32419
rect 32853 32385 32887 32419
rect 36369 32385 36403 32419
rect 46397 32385 46431 32419
rect 2789 32317 2823 32351
rect 24869 32317 24903 32351
rect 31309 32317 31343 32351
rect 31401 32317 31435 32351
rect 37289 32317 37323 32351
rect 37473 32317 37507 32351
rect 46673 32317 46707 32351
rect 26249 32249 26283 32283
rect 18613 32181 18647 32215
rect 20177 32181 20211 32215
rect 21925 32181 21959 32215
rect 25697 32181 25731 32215
rect 16681 31977 16715 32011
rect 27077 31977 27111 32011
rect 35725 31977 35759 32011
rect 46765 31977 46799 32011
rect 21189 31909 21223 31943
rect 22385 31909 22419 31943
rect 26617 31909 26651 31943
rect 32413 31909 32447 31943
rect 1593 31841 1627 31875
rect 2881 31841 2915 31875
rect 28549 31841 28583 31875
rect 38577 31841 38611 31875
rect 47593 31841 47627 31875
rect 1409 31773 1443 31807
rect 15301 31773 15335 31807
rect 17141 31773 17175 31807
rect 19809 31773 19843 31807
rect 22201 31773 22235 31807
rect 23489 31773 23523 31807
rect 24685 31773 24719 31807
rect 24777 31773 24811 31807
rect 24869 31773 24903 31807
rect 25053 31773 25087 31807
rect 25697 31773 25731 31807
rect 27353 31773 27387 31807
rect 27445 31773 27479 31807
rect 27537 31773 27571 31807
rect 27721 31773 27755 31807
rect 28181 31773 28215 31807
rect 28365 31773 28399 31807
rect 31585 31773 31619 31807
rect 31769 31773 31803 31807
rect 32689 31773 32723 31807
rect 32778 31770 32812 31804
rect 32873 31773 32907 31807
rect 33057 31773 33091 31807
rect 33609 31773 33643 31807
rect 35633 31773 35667 31807
rect 36277 31773 36311 31807
rect 36553 31773 36587 31807
rect 37197 31773 37231 31807
rect 46673 31773 46707 31807
rect 47317 31773 47351 31807
rect 15568 31705 15602 31739
rect 17386 31705 17420 31739
rect 20076 31705 20110 31739
rect 23305 31705 23339 31739
rect 26433 31705 26467 31739
rect 33793 31705 33827 31739
rect 37381 31705 37415 31739
rect 18521 31637 18555 31671
rect 24409 31637 24443 31671
rect 25789 31637 25823 31671
rect 31953 31637 31987 31671
rect 2789 31433 2823 31467
rect 16865 31433 16899 31467
rect 18521 31433 18555 31467
rect 18981 31433 19015 31467
rect 28457 31433 28491 31467
rect 31493 31433 31527 31467
rect 32413 31433 32447 31467
rect 37381 31433 37415 31467
rect 20269 31365 20303 31399
rect 20729 31365 20763 31399
rect 23213 31365 23247 31399
rect 27813 31365 27847 31399
rect 28013 31365 28047 31399
rect 28825 31365 28859 31399
rect 29025 31365 29059 31399
rect 39773 31365 39807 31399
rect 1409 31297 1443 31331
rect 1685 31297 1719 31331
rect 2697 31297 2731 31331
rect 17141 31297 17175 31331
rect 17233 31297 17267 31331
rect 17325 31297 17359 31331
rect 17509 31297 17543 31331
rect 18889 31297 18923 31331
rect 20545 31297 20579 31331
rect 22293 31297 22327 31331
rect 25145 31297 25179 31331
rect 29929 31297 29963 31331
rect 31401 31297 31435 31331
rect 32689 31297 32723 31331
rect 32781 31297 32815 31331
rect 32873 31297 32907 31331
rect 33057 31297 33091 31331
rect 37289 31297 37323 31331
rect 19165 31229 19199 31263
rect 29837 31229 29871 31263
rect 30021 31229 30055 31263
rect 30113 31229 30147 31263
rect 35909 31229 35943 31263
rect 36185 31229 36219 31263
rect 37933 31229 37967 31263
rect 38117 31229 38151 31263
rect 28181 31161 28215 31195
rect 20913 31093 20947 31127
rect 22385 31093 22419 31127
rect 23305 31093 23339 31127
rect 24961 31093 24995 31127
rect 27997 31093 28031 31127
rect 29009 31093 29043 31127
rect 29193 31093 29227 31127
rect 29653 31093 29687 31127
rect 35541 31093 35575 31127
rect 2053 30889 2087 30923
rect 29009 30889 29043 30923
rect 31309 30889 31343 30923
rect 38025 30889 38059 30923
rect 17969 30821 18003 30855
rect 16589 30753 16623 30787
rect 24409 30753 24443 30787
rect 27629 30753 27663 30787
rect 20801 30685 20835 30719
rect 20910 30685 20944 30719
rect 21005 30685 21039 30719
rect 21189 30685 21223 30719
rect 22017 30685 22051 30719
rect 22937 30685 22971 30719
rect 24665 30685 24699 30719
rect 29929 30685 29963 30719
rect 30185 30685 30219 30719
rect 35633 30685 35667 30719
rect 36553 30685 36587 30719
rect 37933 30685 37967 30719
rect 16834 30617 16868 30651
rect 19257 30617 19291 30651
rect 19441 30617 19475 30651
rect 22201 30617 22235 30651
rect 22385 30617 22419 30651
rect 23121 30617 23155 30651
rect 27896 30617 27930 30651
rect 36001 30617 36035 30651
rect 36921 30617 36955 30651
rect 19625 30549 19659 30583
rect 20545 30549 20579 30583
rect 25789 30549 25823 30583
rect 16681 30277 16715 30311
rect 18613 30277 18647 30311
rect 21005 30277 21039 30311
rect 48145 30277 48179 30311
rect 2145 30209 2179 30243
rect 16957 30209 16991 30243
rect 17046 30209 17080 30243
rect 17146 30209 17180 30243
rect 17325 30209 17359 30243
rect 18521 30209 18555 30243
rect 19717 30209 19751 30243
rect 19809 30209 19843 30243
rect 20913 30209 20947 30243
rect 21833 30209 21867 30243
rect 22017 30209 22051 30243
rect 23213 30209 23247 30243
rect 24685 30209 24719 30243
rect 24869 30209 24903 30243
rect 25605 30209 25639 30243
rect 27445 30209 27479 30243
rect 28917 30209 28951 30243
rect 29101 30209 29135 30243
rect 29929 30209 29963 30243
rect 30185 30209 30219 30243
rect 37289 30209 37323 30243
rect 47961 30209 47995 30243
rect 18797 30141 18831 30175
rect 19993 30141 20027 30175
rect 21189 30141 21223 30175
rect 22201 30141 22235 30175
rect 23305 30141 23339 30175
rect 23397 30141 23431 30175
rect 28641 30141 28675 30175
rect 28825 30141 28859 30175
rect 29009 30141 29043 30175
rect 18153 30073 18187 30107
rect 20545 30073 20579 30107
rect 25789 30073 25823 30107
rect 31309 30073 31343 30107
rect 1685 30005 1719 30039
rect 2237 30005 2271 30039
rect 19349 30005 19383 30039
rect 22845 30005 22879 30039
rect 25053 30005 25087 30039
rect 27537 30005 27571 30039
rect 37473 30005 37507 30039
rect 18153 29801 18187 29835
rect 27537 29801 27571 29835
rect 29837 29801 29871 29835
rect 31033 29801 31067 29835
rect 34805 29801 34839 29835
rect 38669 29801 38703 29835
rect 23581 29733 23615 29767
rect 26341 29733 26375 29767
rect 35081 29733 35115 29767
rect 1409 29665 1443 29699
rect 1593 29665 1627 29699
rect 2789 29665 2823 29699
rect 22201 29665 22235 29699
rect 30021 29665 30055 29699
rect 30113 29665 30147 29699
rect 37289 29665 37323 29699
rect 16773 29597 16807 29631
rect 20177 29597 20211 29631
rect 20444 29597 20478 29631
rect 24961 29597 24995 29631
rect 30205 29597 30239 29631
rect 30297 29597 30331 29631
rect 32137 29597 32171 29631
rect 32321 29597 32355 29631
rect 32781 29597 32815 29631
rect 34713 29597 34747 29631
rect 34897 29597 34931 29631
rect 47685 29597 47719 29631
rect 17018 29529 17052 29563
rect 22446 29529 22480 29563
rect 25206 29529 25240 29563
rect 27445 29529 27479 29563
rect 28365 29529 28399 29563
rect 30941 29529 30975 29563
rect 32229 29529 32263 29563
rect 33026 29529 33060 29563
rect 37556 29529 37590 29563
rect 21557 29461 21591 29495
rect 28457 29461 28491 29495
rect 34161 29461 34195 29495
rect 16681 29257 16715 29291
rect 22017 29257 22051 29291
rect 24317 29257 24351 29291
rect 28733 29257 28767 29291
rect 29945 29257 29979 29291
rect 30113 29257 30147 29291
rect 32689 29257 32723 29291
rect 18153 29189 18187 29223
rect 27445 29189 27479 29223
rect 29745 29189 29779 29223
rect 35817 29189 35851 29223
rect 36645 29189 36679 29223
rect 37473 29189 37507 29223
rect 16911 29121 16945 29155
rect 17030 29124 17064 29158
rect 17141 29124 17175 29158
rect 17325 29121 17359 29155
rect 17785 29121 17819 29155
rect 17969 29121 18003 29155
rect 22293 29121 22327 29155
rect 22385 29121 22419 29155
rect 22477 29121 22511 29155
rect 22661 29121 22695 29155
rect 24593 29121 24627 29155
rect 24685 29121 24719 29155
rect 24777 29121 24811 29155
rect 24961 29121 24995 29155
rect 28457 29121 28491 29155
rect 28733 29121 28767 29155
rect 32597 29121 32631 29155
rect 33609 29121 33643 29155
rect 33876 29121 33910 29155
rect 35449 29121 35483 29155
rect 35633 29121 35667 29155
rect 35909 29121 35943 29155
rect 36553 29121 36587 29155
rect 37289 29121 37323 29155
rect 47593 29121 47627 29155
rect 27629 29053 27663 29087
rect 39129 29053 39163 29087
rect 47685 28985 47719 29019
rect 2053 28917 2087 28951
rect 29929 28917 29963 28951
rect 34989 28917 35023 28951
rect 26893 28713 26927 28747
rect 27997 28713 28031 28747
rect 28917 28645 28951 28679
rect 38761 28645 38795 28679
rect 1409 28577 1443 28611
rect 2789 28577 2823 28611
rect 27629 28577 27663 28611
rect 36461 28577 36495 28611
rect 38301 28577 38335 28611
rect 48145 28577 48179 28611
rect 19257 28509 19291 28543
rect 22201 28509 22235 28543
rect 24685 28509 24719 28543
rect 24777 28509 24811 28543
rect 24869 28509 24903 28543
rect 25053 28509 25087 28543
rect 25513 28509 25547 28543
rect 26801 28509 26835 28543
rect 27077 28509 27111 28543
rect 27813 28509 27847 28543
rect 28733 28509 28767 28543
rect 31710 28509 31744 28543
rect 32137 28509 32171 28543
rect 32229 28509 32263 28543
rect 32873 28509 32907 28543
rect 33057 28509 33091 28543
rect 33885 28509 33919 28543
rect 34069 28509 34103 28543
rect 34161 28509 34195 28543
rect 34713 28509 34747 28543
rect 34897 28509 34931 28543
rect 35265 28509 35299 28543
rect 38945 28509 38979 28543
rect 39037 28509 39071 28543
rect 46305 28509 46339 28543
rect 1593 28441 1627 28475
rect 17693 28441 17727 28475
rect 17877 28441 17911 28475
rect 23489 28441 23523 28475
rect 25697 28441 25731 28475
rect 35173 28441 35207 28475
rect 36645 28441 36679 28475
rect 38761 28441 38795 28475
rect 46489 28441 46523 28475
rect 18061 28373 18095 28407
rect 19349 28373 19383 28407
rect 22293 28373 22327 28407
rect 23581 28373 23615 28407
rect 24409 28373 24443 28407
rect 25881 28373 25915 28407
rect 31585 28373 31619 28407
rect 31769 28373 31803 28407
rect 32965 28373 32999 28407
rect 33701 28373 33735 28407
rect 2329 28169 2363 28203
rect 26433 28169 26467 28203
rect 36553 28169 36587 28203
rect 37565 28169 37599 28203
rect 17592 28101 17626 28135
rect 19165 28101 19199 28135
rect 20269 28101 20303 28135
rect 25298 28101 25332 28135
rect 34345 28101 34379 28135
rect 38669 28101 38703 28135
rect 39405 28101 39439 28135
rect 2237 28033 2271 28067
rect 12633 28033 12667 28067
rect 19395 28033 19429 28067
rect 19530 28033 19564 28067
rect 19625 28033 19659 28067
rect 19809 28033 19843 28067
rect 20453 28033 20487 28067
rect 22569 28033 22603 28067
rect 22661 28033 22695 28067
rect 22753 28033 22787 28067
rect 22937 28033 22971 28067
rect 23673 28033 23707 28067
rect 23765 28033 23799 28067
rect 23857 28033 23891 28067
rect 24041 28033 24075 28067
rect 25053 28033 25087 28067
rect 28457 28033 28491 28067
rect 30001 28033 30035 28067
rect 32137 28033 32171 28067
rect 32321 28033 32355 28067
rect 34253 28033 34287 28067
rect 36461 28033 36495 28067
rect 37473 28033 37507 28067
rect 37657 28033 37691 28067
rect 38577 28033 38611 28067
rect 47869 28033 47903 28067
rect 17325 27965 17359 27999
rect 29745 27965 29779 27999
rect 39221 27965 39255 27999
rect 41061 27965 41095 27999
rect 45201 27965 45235 27999
rect 45385 27965 45419 27999
rect 46029 27965 46063 27999
rect 31125 27897 31159 27931
rect 12725 27829 12759 27863
rect 18705 27829 18739 27863
rect 20637 27829 20671 27863
rect 22293 27829 22327 27863
rect 23397 27829 23431 27863
rect 28549 27829 28583 27863
rect 28917 27829 28951 27863
rect 32137 27829 32171 27863
rect 48053 27829 48087 27863
rect 24777 27625 24811 27659
rect 29561 27625 29595 27659
rect 33241 27625 33275 27659
rect 17325 27557 17359 27591
rect 20821 27557 20855 27591
rect 32505 27557 32539 27591
rect 45569 27557 45603 27591
rect 23305 27489 23339 27523
rect 39865 27489 39899 27523
rect 46305 27489 46339 27523
rect 46489 27489 46523 27523
rect 48145 27489 48179 27523
rect 1777 27421 1811 27455
rect 2237 27421 2271 27455
rect 3065 27421 3099 27455
rect 15945 27421 15979 27455
rect 18291 27421 18325 27455
rect 18429 27421 18463 27455
rect 18521 27421 18555 27455
rect 18705 27421 18739 27455
rect 19441 27421 19475 27455
rect 21603 27421 21637 27455
rect 21741 27421 21775 27455
rect 21854 27421 21888 27455
rect 22017 27421 22051 27455
rect 23029 27421 23063 27455
rect 25973 27421 26007 27455
rect 26065 27421 26099 27455
rect 26157 27421 26191 27455
rect 26341 27421 26375 27455
rect 26801 27421 26835 27455
rect 28641 27421 28675 27455
rect 29837 27421 29871 27455
rect 31125 27421 31159 27455
rect 31392 27421 31426 27455
rect 33057 27421 33091 27455
rect 36001 27421 36035 27455
rect 39129 27421 39163 27455
rect 45477 27421 45511 27455
rect 16212 27353 16246 27387
rect 19686 27353 19720 27387
rect 24409 27353 24443 27387
rect 24593 27353 24627 27387
rect 25697 27353 25731 27387
rect 27046 27353 27080 27387
rect 29561 27353 29595 27387
rect 29745 27353 29779 27387
rect 33885 27353 33919 27387
rect 34069 27353 34103 27387
rect 35173 27353 35207 27387
rect 35357 27353 35391 27387
rect 36268 27353 36302 27387
rect 39221 27353 39255 27387
rect 40049 27353 40083 27387
rect 41705 27353 41739 27387
rect 2329 27285 2363 27319
rect 18061 27285 18095 27319
rect 21373 27285 21407 27319
rect 28181 27285 28215 27319
rect 28825 27285 28859 27319
rect 35541 27285 35575 27319
rect 37381 27285 37415 27319
rect 26157 27081 26191 27115
rect 37289 27081 37323 27115
rect 46581 27081 46615 27115
rect 1961 27013 1995 27047
rect 11989 27013 12023 27047
rect 18429 27013 18463 27047
rect 21097 27013 21131 27047
rect 21281 27013 21315 27047
rect 1777 26945 1811 26979
rect 15761 26945 15795 26979
rect 16681 26945 16715 26979
rect 18245 26945 18279 26979
rect 20913 26945 20947 26979
rect 21833 26945 21867 26979
rect 22089 26945 22123 26979
rect 23857 26945 23891 26979
rect 24113 26945 24147 26979
rect 25881 26945 25915 26979
rect 25973 26945 26007 26979
rect 27169 26945 27203 26979
rect 28089 26945 28123 26979
rect 28457 26945 28491 26979
rect 30021 26945 30055 26979
rect 30113 26945 30147 26979
rect 30205 26945 30239 26979
rect 30389 26945 30423 26979
rect 33241 26945 33275 26979
rect 33508 26945 33542 26979
rect 35265 26945 35299 26979
rect 35449 26945 35483 26979
rect 36323 26945 36357 26979
rect 36461 26945 36495 26979
rect 36574 26945 36608 26979
rect 36737 26945 36771 26979
rect 37565 26945 37599 26979
rect 37654 26951 37688 26985
rect 37749 26945 37783 26979
rect 37933 26945 37967 26979
rect 38577 26945 38611 26979
rect 46489 26945 46523 26979
rect 2789 26877 2823 26911
rect 11805 26877 11839 26911
rect 12265 26877 12299 26911
rect 17049 26877 17083 26911
rect 18705 26877 18739 26911
rect 26157 26877 26191 26911
rect 35633 26877 35667 26911
rect 39221 26877 39255 26911
rect 39405 26877 39439 26911
rect 41061 26877 41095 26911
rect 25237 26809 25271 26843
rect 15853 26741 15887 26775
rect 23213 26741 23247 26775
rect 26985 26741 27019 26775
rect 29745 26741 29779 26775
rect 34621 26741 34655 26775
rect 36093 26741 36127 26775
rect 38669 26741 38703 26775
rect 19257 26537 19291 26571
rect 20729 26537 20763 26571
rect 24961 26537 24995 26571
rect 26065 26537 26099 26571
rect 32321 26537 32355 26571
rect 37749 26537 37783 26571
rect 39221 26537 39255 26571
rect 18613 26469 18647 26503
rect 23857 26469 23891 26503
rect 47961 26469 47995 26503
rect 1409 26401 1443 26435
rect 2789 26401 2823 26435
rect 15669 26401 15703 26435
rect 15853 26401 15887 26435
rect 30205 26401 30239 26435
rect 34713 26401 34747 26435
rect 39865 26401 39899 26435
rect 40049 26401 40083 26435
rect 18245 26333 18279 26367
rect 18429 26333 18463 26367
rect 19533 26333 19567 26367
rect 19625 26333 19659 26367
rect 19717 26333 19751 26367
rect 19901 26333 19935 26367
rect 20637 26333 20671 26367
rect 22477 26333 22511 26367
rect 24869 26333 24903 26367
rect 30461 26333 30495 26367
rect 33701 26333 33735 26367
rect 33885 26333 33919 26367
rect 34969 26333 35003 26367
rect 35078 26333 35112 26367
rect 35173 26330 35207 26364
rect 35351 26333 35385 26367
rect 36369 26333 36403 26367
rect 36625 26333 36659 26367
rect 39129 26333 39163 26367
rect 48145 26333 48179 26367
rect 1593 26265 1627 26299
rect 17509 26265 17543 26299
rect 22744 26265 22778 26299
rect 25973 26265 26007 26299
rect 32229 26265 32263 26299
rect 41705 26265 41739 26299
rect 31585 26197 31619 26231
rect 34069 26197 34103 26231
rect 2789 25993 2823 26027
rect 23765 25925 23799 25959
rect 29653 25925 29687 25959
rect 30021 25925 30055 25959
rect 30757 25925 30791 25959
rect 34989 25925 35023 25959
rect 35173 25925 35207 25959
rect 1409 25857 1443 25891
rect 2697 25857 2731 25891
rect 15577 25857 15611 25891
rect 15945 25857 15979 25891
rect 16681 25857 16715 25891
rect 20361 25857 20395 25891
rect 20545 25857 20579 25891
rect 23397 25857 23431 25891
rect 23581 25857 23615 25891
rect 29837 25857 29871 25891
rect 30573 25857 30607 25891
rect 33195 25857 33229 25891
rect 33330 25857 33364 25891
rect 33425 25857 33459 25891
rect 33609 25857 33643 25891
rect 36323 25857 36357 25891
rect 36461 25857 36495 25891
rect 36553 25860 36587 25894
rect 36737 25857 36771 25891
rect 1685 25789 1719 25823
rect 17141 25789 17175 25823
rect 45201 25789 45235 25823
rect 45385 25789 45419 25823
rect 46857 25789 46891 25823
rect 16037 25653 16071 25687
rect 20729 25653 20763 25687
rect 32965 25653 32999 25687
rect 36093 25653 36127 25687
rect 47777 25653 47811 25687
rect 19993 25449 20027 25483
rect 20729 25449 20763 25483
rect 35817 25449 35851 25483
rect 45753 25449 45787 25483
rect 47133 25449 47167 25483
rect 47869 25449 47903 25483
rect 19901 25313 19935 25347
rect 20821 25313 20855 25347
rect 29009 25313 29043 25347
rect 47501 25313 47535 25347
rect 15117 25245 15151 25279
rect 16589 25245 16623 25279
rect 17601 25245 17635 25279
rect 19717 25245 19751 25279
rect 19993 25245 20027 25279
rect 21005 25245 21039 25279
rect 25329 25245 25363 25279
rect 25421 25245 25455 25279
rect 25513 25245 25547 25279
rect 25697 25245 25731 25279
rect 30343 25245 30377 25279
rect 30481 25245 30515 25279
rect 30594 25245 30628 25279
rect 30751 25245 30785 25279
rect 33425 25245 33459 25279
rect 33517 25245 33551 25279
rect 33609 25245 33643 25279
rect 33793 25245 33827 25279
rect 36277 25245 36311 25279
rect 36533 25245 36567 25279
rect 40325 25245 40359 25279
rect 45661 25245 45695 25279
rect 47869 25245 47903 25279
rect 15853 25177 15887 25211
rect 20729 25177 20763 25211
rect 28089 25177 28123 25211
rect 28825 25177 28859 25211
rect 31217 25177 31251 25211
rect 31401 25177 31435 25211
rect 35449 25177 35483 25211
rect 35633 25177 35667 25211
rect 20177 25109 20211 25143
rect 21189 25109 21223 25143
rect 25053 25109 25087 25143
rect 28181 25109 28215 25143
rect 30113 25109 30147 25143
rect 31585 25109 31619 25143
rect 33149 25109 33183 25143
rect 37657 25109 37691 25143
rect 40141 25109 40175 25143
rect 47685 25109 47719 25143
rect 20177 24905 20211 24939
rect 21097 24905 21131 24939
rect 32781 24905 32815 24939
rect 33508 24837 33542 24871
rect 2145 24769 2179 24803
rect 15761 24769 15795 24803
rect 16129 24769 16163 24803
rect 16681 24769 16715 24803
rect 18797 24769 18831 24803
rect 19073 24769 19107 24803
rect 19717 24769 19751 24803
rect 19993 24769 20027 24803
rect 20637 24769 20671 24803
rect 20913 24769 20947 24803
rect 22753 24769 22787 24803
rect 22937 24769 22971 24803
rect 23029 24769 23063 24803
rect 23489 24769 23523 24803
rect 24961 24769 24995 24803
rect 25228 24769 25262 24803
rect 27997 24769 28031 24803
rect 28273 24769 28307 24803
rect 29193 24769 29227 24803
rect 30472 24769 30506 24803
rect 32413 24769 32447 24803
rect 32597 24769 32631 24803
rect 39764 24769 39798 24803
rect 41889 24769 41923 24803
rect 42441 24769 42475 24803
rect 42697 24769 42731 24803
rect 46857 24769 46891 24803
rect 47869 24769 47903 24803
rect 17141 24701 17175 24735
rect 18889 24701 18923 24735
rect 19901 24701 19935 24735
rect 20821 24701 20855 24735
rect 28181 24701 28215 24735
rect 28917 24701 28951 24735
rect 30205 24701 30239 24735
rect 33241 24701 33275 24735
rect 39497 24701 39531 24735
rect 19257 24633 19291 24667
rect 34621 24633 34655 24667
rect 41705 24633 41739 24667
rect 48053 24633 48087 24667
rect 2237 24565 2271 24599
rect 19073 24565 19107 24599
rect 19993 24565 20027 24599
rect 20913 24565 20947 24599
rect 22569 24565 22603 24599
rect 23581 24565 23615 24599
rect 26341 24565 26375 24599
rect 28273 24565 28307 24599
rect 28457 24565 28491 24599
rect 31585 24565 31619 24599
rect 40877 24565 40911 24599
rect 43821 24565 43855 24599
rect 46949 24565 46983 24599
rect 19717 24361 19751 24395
rect 20177 24361 20211 24395
rect 20913 24361 20947 24395
rect 28549 24361 28583 24395
rect 29653 24361 29687 24395
rect 38853 24361 38887 24395
rect 40325 24361 40359 24395
rect 41797 24361 41831 24395
rect 41981 24361 42015 24395
rect 42533 24361 42567 24395
rect 27445 24293 27479 24327
rect 29009 24293 29043 24327
rect 40509 24293 40543 24327
rect 40969 24293 41003 24327
rect 43269 24293 43303 24327
rect 16865 24225 16899 24259
rect 17877 24225 17911 24259
rect 19809 24225 19843 24259
rect 20821 24225 20855 24259
rect 21925 24225 21959 24259
rect 27537 24225 27571 24259
rect 29837 24225 29871 24259
rect 32781 24225 32815 24259
rect 34713 24225 34747 24259
rect 46305 24225 46339 24259
rect 46489 24225 46523 24259
rect 48145 24225 48179 24259
rect 1409 24157 1443 24191
rect 1685 24157 1719 24191
rect 2881 24157 2915 24191
rect 15761 24157 15795 24191
rect 16221 24157 16255 24191
rect 16405 24157 16439 24191
rect 19993 24157 20027 24191
rect 20913 24157 20947 24191
rect 22192 24157 22226 24191
rect 24501 24157 24535 24191
rect 24685 24157 24719 24191
rect 25329 24157 25363 24191
rect 27169 24157 27203 24191
rect 27316 24157 27350 24191
rect 28641 24157 28675 24191
rect 28825 24157 28859 24191
rect 30021 24157 30055 24191
rect 31953 24157 31987 24191
rect 32042 24157 32076 24191
rect 32137 24157 32171 24191
rect 32321 24157 32355 24191
rect 34969 24157 35003 24191
rect 37105 24157 37139 24191
rect 38117 24157 38151 24191
rect 38761 24157 38795 24191
rect 39957 24157 39991 24191
rect 41153 24157 41187 24191
rect 42605 24157 42639 24191
rect 42729 24135 42763 24169
rect 43177 24157 43211 24191
rect 43361 24157 43395 24191
rect 44005 24157 44039 24191
rect 17049 24089 17083 24123
rect 19717 24089 19751 24123
rect 20637 24089 20671 24123
rect 25596 24089 25630 24123
rect 28365 24089 28399 24123
rect 29561 24089 29595 24123
rect 30849 24089 30883 24123
rect 31033 24089 31067 24123
rect 31677 24089 31711 24123
rect 33026 24089 33060 24123
rect 38301 24089 38335 24123
rect 41613 24089 41647 24123
rect 42441 24089 42475 24123
rect 16313 24021 16347 24055
rect 21097 24021 21131 24055
rect 23305 24021 23339 24055
rect 24685 24021 24719 24055
rect 26709 24021 26743 24055
rect 27813 24021 27847 24055
rect 30205 24021 30239 24055
rect 31217 24021 31251 24055
rect 34161 24021 34195 24055
rect 36093 24021 36127 24055
rect 37289 24021 37323 24055
rect 39221 24021 39255 24055
rect 40325 24021 40359 24055
rect 41813 24021 41847 24055
rect 43821 24021 43855 24055
rect 21097 23817 21131 23851
rect 24961 23817 24995 23851
rect 26433 23817 26467 23851
rect 29101 23817 29135 23851
rect 33149 23817 33183 23851
rect 36645 23817 36679 23851
rect 38853 23817 38887 23851
rect 38945 23817 38979 23851
rect 40141 23817 40175 23851
rect 40969 23817 41003 23851
rect 48053 23817 48087 23851
rect 1961 23749 1995 23783
rect 15945 23749 15979 23783
rect 19717 23749 19751 23783
rect 35725 23749 35759 23783
rect 37289 23749 37323 23783
rect 37505 23749 37539 23783
rect 41613 23749 41647 23783
rect 43168 23749 43202 23783
rect 47961 23749 47995 23783
rect 1777 23681 1811 23715
rect 15669 23681 15703 23715
rect 16957 23681 16991 23715
rect 19993 23681 20027 23715
rect 20637 23681 20671 23715
rect 20821 23681 20855 23715
rect 20913 23681 20947 23715
rect 22385 23681 22419 23715
rect 22652 23681 22686 23715
rect 24317 23681 24351 23715
rect 24501 23681 24535 23715
rect 25237 23681 25271 23715
rect 25326 23681 25360 23715
rect 25442 23681 25476 23715
rect 25605 23681 25639 23715
rect 26065 23681 26099 23715
rect 26249 23681 26283 23715
rect 28181 23681 28215 23715
rect 28549 23681 28583 23715
rect 29377 23681 29411 23715
rect 29561 23681 29595 23715
rect 30297 23681 30331 23715
rect 32781 23681 32815 23715
rect 32965 23681 32999 23715
rect 35909 23681 35943 23715
rect 36369 23681 36403 23715
rect 39681 23681 39715 23715
rect 40601 23681 40635 23715
rect 40785 23681 40819 23715
rect 41429 23681 41463 23715
rect 2789 23613 2823 23647
rect 17141 23613 17175 23647
rect 17509 23613 17543 23647
rect 19809 23613 19843 23647
rect 28089 23613 28123 23647
rect 36645 23613 36679 23647
rect 39037 23613 39071 23647
rect 41797 23613 41831 23647
rect 42901 23613 42935 23647
rect 20177 23545 20211 23579
rect 28733 23545 28767 23579
rect 29745 23545 29779 23579
rect 44281 23545 44315 23579
rect 19901 23477 19935 23511
rect 20913 23477 20947 23511
rect 23765 23477 23799 23511
rect 24409 23477 24443 23511
rect 28457 23477 28491 23511
rect 29377 23477 29411 23511
rect 30389 23477 30423 23511
rect 36461 23477 36495 23511
rect 37473 23477 37507 23511
rect 37657 23477 37691 23511
rect 38485 23477 38519 23511
rect 39957 23477 39991 23511
rect 17601 23273 17635 23307
rect 18153 23273 18187 23307
rect 20177 23273 20211 23307
rect 20361 23273 20395 23307
rect 28365 23273 28399 23307
rect 35725 23273 35759 23307
rect 37197 23273 37231 23307
rect 40233 23273 40267 23307
rect 28549 23205 28583 23239
rect 30205 23205 30239 23239
rect 35265 23205 35299 23239
rect 38761 23205 38795 23239
rect 19993 23137 20027 23171
rect 37289 23137 37323 23171
rect 38485 23137 38519 23171
rect 41521 23137 41555 23171
rect 41705 23137 41739 23171
rect 42349 23137 42383 23171
rect 43637 23137 43671 23171
rect 16221 23069 16255 23103
rect 18061 23069 18095 23103
rect 20177 23069 20211 23103
rect 23489 23069 23523 23103
rect 28181 23069 28215 23103
rect 28365 23069 28399 23103
rect 30849 23069 30883 23103
rect 32137 23069 32171 23103
rect 35081 23069 35115 23103
rect 35725 23069 35759 23103
rect 35909 23069 35943 23103
rect 36001 23069 36035 23103
rect 37381 23069 37415 23103
rect 38393 23069 38427 23103
rect 39865 23069 39899 23103
rect 40049 23069 40083 23103
rect 41613 23069 41647 23103
rect 41797 23069 41831 23103
rect 42625 23069 42659 23103
rect 43913 23069 43947 23103
rect 16466 23001 16500 23035
rect 19901 23001 19935 23035
rect 23305 23001 23339 23035
rect 23673 23001 23707 23035
rect 27537 23001 27571 23035
rect 30021 23001 30055 23035
rect 31033 23001 31067 23035
rect 32321 23001 32355 23035
rect 37105 23001 37139 23035
rect 27629 22933 27663 22967
rect 31217 22933 31251 22967
rect 32505 22933 32539 22967
rect 36185 22933 36219 22967
rect 37565 22933 37599 22967
rect 41337 22933 41371 22967
rect 16865 22729 16899 22763
rect 20085 22729 20119 22763
rect 23397 22729 23431 22763
rect 27813 22729 27847 22763
rect 40325 22729 40359 22763
rect 40509 22729 40543 22763
rect 48053 22729 48087 22763
rect 2053 22661 2087 22695
rect 17785 22661 17819 22695
rect 27629 22661 27663 22695
rect 38117 22661 38151 22695
rect 42441 22661 42475 22695
rect 1869 22593 1903 22627
rect 3433 22593 3467 22627
rect 15485 22593 15519 22627
rect 16773 22593 16807 22627
rect 17417 22593 17451 22627
rect 17601 22593 17635 22627
rect 18501 22593 18535 22627
rect 18610 22599 18644 22633
rect 18705 22596 18739 22630
rect 18889 22593 18923 22627
rect 19625 22593 19659 22627
rect 19901 22593 19935 22627
rect 23213 22593 23247 22627
rect 23489 22593 23523 22627
rect 24869 22593 24903 22627
rect 24961 22593 24995 22627
rect 25053 22593 25087 22627
rect 25237 22593 25271 22627
rect 27445 22593 27479 22627
rect 28457 22593 28491 22627
rect 28733 22593 28767 22627
rect 29469 22593 29503 22627
rect 31217 22593 31251 22627
rect 31309 22593 31343 22627
rect 31401 22593 31435 22627
rect 31585 22593 31619 22627
rect 32505 22593 32539 22627
rect 32597 22593 32631 22627
rect 32689 22593 32723 22627
rect 32873 22593 32907 22627
rect 33609 22593 33643 22627
rect 33701 22593 33735 22627
rect 33793 22593 33827 22627
rect 33977 22593 34011 22627
rect 35817 22593 35851 22627
rect 36001 22593 36035 22627
rect 37289 22593 37323 22627
rect 38301 22593 38335 22627
rect 38393 22593 38427 22627
rect 40417 22593 40451 22627
rect 41797 22593 41831 22627
rect 42717 22593 42751 22627
rect 45293 22593 45327 22627
rect 45477 22593 45511 22627
rect 47961 22593 47995 22627
rect 15761 22525 15795 22559
rect 19717 22525 19751 22559
rect 28917 22525 28951 22559
rect 37381 22525 37415 22559
rect 41521 22525 41555 22559
rect 41613 22525 41647 22559
rect 41705 22525 41739 22559
rect 42625 22525 42659 22559
rect 23213 22457 23247 22491
rect 38117 22457 38151 22491
rect 40141 22457 40175 22491
rect 3525 22389 3559 22423
rect 18245 22389 18279 22423
rect 19625 22389 19659 22423
rect 24593 22389 24627 22423
rect 29561 22389 29595 22423
rect 30941 22389 30975 22423
rect 32229 22389 32263 22423
rect 33333 22389 33367 22423
rect 35909 22389 35943 22423
rect 36185 22389 36219 22423
rect 37381 22389 37415 22423
rect 37657 22389 37691 22423
rect 40693 22389 40727 22423
rect 41337 22389 41371 22423
rect 42441 22389 42475 22423
rect 42901 22389 42935 22423
rect 45661 22389 45695 22423
rect 34069 22185 34103 22219
rect 40509 22185 40543 22219
rect 42073 22185 42107 22219
rect 18245 22117 18279 22151
rect 31769 22117 31803 22151
rect 41153 22117 41187 22151
rect 42257 22117 42291 22151
rect 4261 22049 4295 22083
rect 14105 22049 14139 22083
rect 15485 22049 15519 22083
rect 24685 22049 24719 22083
rect 28457 22049 28491 22083
rect 36829 22049 36863 22083
rect 45109 22049 45143 22083
rect 3065 21981 3099 22015
rect 3801 21981 3835 22015
rect 16865 21981 16899 22015
rect 19257 21981 19291 22015
rect 27215 21981 27249 22015
rect 27353 21981 27387 22015
rect 27445 21981 27479 22015
rect 27629 21981 27663 22015
rect 28181 21981 28215 22015
rect 32689 21981 32723 22015
rect 36185 21981 36219 22015
rect 36369 21981 36403 22015
rect 37105 21981 37139 22015
rect 40417 21981 40451 22015
rect 41153 21981 41187 22015
rect 41337 21981 41371 22015
rect 43223 21981 43257 22015
rect 43361 21981 43395 22015
rect 43458 21981 43492 22015
rect 43637 21981 43671 22015
rect 48145 21981 48179 22015
rect 3157 21913 3191 21947
rect 3985 21913 4019 21947
rect 14289 21913 14323 21947
rect 17132 21913 17166 21947
rect 19441 21913 19475 21947
rect 24952 21913 24986 21947
rect 30481 21913 30515 21947
rect 32934 21913 32968 21947
rect 41889 21913 41923 21947
rect 42089 21913 42123 21947
rect 45354 21913 45388 21947
rect 47961 21913 47995 21947
rect 19625 21845 19659 21879
rect 26065 21845 26099 21879
rect 26985 21845 27019 21879
rect 36369 21845 36403 21879
rect 42993 21845 43027 21879
rect 46489 21845 46523 21879
rect 13921 21641 13955 21675
rect 31493 21641 31527 21675
rect 37867 21641 37901 21675
rect 46857 21641 46891 21675
rect 3525 21573 3559 21607
rect 17049 21573 17083 21607
rect 19502 21573 19536 21607
rect 30380 21573 30414 21607
rect 32781 21573 32815 21607
rect 34130 21573 34164 21607
rect 37657 21573 37691 21607
rect 38669 21573 38703 21607
rect 40969 21573 41003 21607
rect 13829 21505 13863 21539
rect 14933 21505 14967 21539
rect 19257 21505 19291 21539
rect 21833 21505 21867 21539
rect 22089 21505 22123 21539
rect 23857 21505 23891 21539
rect 24041 21505 24075 21539
rect 24133 21505 24167 21539
rect 25053 21505 25087 21539
rect 25320 21505 25354 21539
rect 27353 21505 27387 21539
rect 27609 21505 27643 21539
rect 29193 21505 29227 21539
rect 29377 21505 29411 21539
rect 30113 21505 30147 21539
rect 32321 21505 32355 21539
rect 33011 21505 33045 21539
rect 33149 21505 33183 21539
rect 33241 21505 33275 21539
rect 33425 21505 33459 21539
rect 38485 21505 38519 21539
rect 38770 21527 38804 21561
rect 43801 21505 43835 21539
rect 45477 21505 45511 21539
rect 45744 21505 45778 21539
rect 3341 21437 3375 21471
rect 5181 21437 5215 21471
rect 15945 21437 15979 21471
rect 33885 21437 33919 21471
rect 43545 21437 43579 21471
rect 20637 21369 20671 21403
rect 35265 21369 35299 21403
rect 38485 21369 38519 21403
rect 40601 21369 40635 21403
rect 18337 21301 18371 21335
rect 23213 21301 23247 21335
rect 23673 21301 23707 21335
rect 26433 21301 26467 21335
rect 28733 21301 28767 21335
rect 29561 21301 29595 21335
rect 32137 21301 32171 21335
rect 37841 21301 37875 21335
rect 38025 21301 38059 21335
rect 40969 21301 41003 21335
rect 41153 21301 41187 21335
rect 44925 21301 44959 21335
rect 47777 21301 47811 21335
rect 19257 21097 19291 21131
rect 21189 21097 21223 21131
rect 21925 21097 21959 21131
rect 35081 21097 35115 21131
rect 37657 21097 37691 21131
rect 37749 21097 37783 21131
rect 41245 21097 41279 21131
rect 44465 21097 44499 21131
rect 45017 21097 45051 21131
rect 22845 21029 22879 21063
rect 25053 21029 25087 21063
rect 27353 21029 27387 21063
rect 16589 20961 16623 20995
rect 23397 20961 23431 20995
rect 26525 20961 26559 20995
rect 32781 20961 32815 20995
rect 37841 20961 37875 20995
rect 42625 20961 42659 20995
rect 42901 20961 42935 20995
rect 46305 20961 46339 20995
rect 46949 20961 46983 20995
rect 14933 20893 14967 20927
rect 16037 20893 16071 20927
rect 18521 20893 18555 20927
rect 19533 20893 19567 20927
rect 19625 20893 19659 20927
rect 19717 20893 19751 20927
rect 19901 20893 19935 20927
rect 22109 20893 22143 20927
rect 22293 20893 22327 20927
rect 22385 20893 22419 20927
rect 24409 20893 24443 20927
rect 25283 20893 25317 20927
rect 25421 20893 25455 20927
rect 25513 20893 25547 20927
rect 25697 20893 25731 20927
rect 26157 20893 26191 20927
rect 26985 20893 27019 20927
rect 27169 20893 27203 20927
rect 28365 20893 28399 20927
rect 28549 20893 28583 20927
rect 29561 20893 29595 20927
rect 31401 20893 31435 20927
rect 31677 20893 31711 20927
rect 33048 20893 33082 20927
rect 34713 20893 34747 20927
rect 34897 20893 34931 20927
rect 38117 20893 38151 20927
rect 39865 20893 39899 20927
rect 41889 20893 41923 20927
rect 44097 20893 44131 20927
rect 45247 20893 45281 20927
rect 45366 20890 45400 20924
rect 45498 20893 45532 20927
rect 45661 20893 45695 20927
rect 15485 20825 15519 20859
rect 16221 20825 16255 20859
rect 18337 20825 18371 20859
rect 21097 20825 21131 20859
rect 23305 20825 23339 20859
rect 26341 20825 26375 20859
rect 29817 20825 29851 20859
rect 40132 20825 40166 20859
rect 44281 20825 44315 20859
rect 46489 20825 46523 20859
rect 18705 20757 18739 20791
rect 23213 20757 23247 20791
rect 24501 20757 24535 20791
rect 28549 20757 28583 20791
rect 30941 20757 30975 20791
rect 34161 20757 34195 20791
rect 37381 20757 37415 20791
rect 38025 20757 38059 20791
rect 41705 20757 41739 20791
rect 14841 20553 14875 20587
rect 16865 20553 16899 20587
rect 19395 20553 19429 20587
rect 22753 20553 22787 20587
rect 24225 20553 24259 20587
rect 25237 20553 25271 20587
rect 28825 20553 28859 20587
rect 29929 20553 29963 20587
rect 36737 20553 36771 20587
rect 43269 20553 43303 20587
rect 44465 20553 44499 20587
rect 47685 20553 47719 20587
rect 24869 20485 24903 20519
rect 31493 20485 31527 20519
rect 32321 20485 32355 20519
rect 36277 20485 36311 20519
rect 40141 20485 40175 20519
rect 40325 20485 40359 20519
rect 45937 20485 45971 20519
rect 11713 20417 11747 20451
rect 14749 20417 14783 20451
rect 15485 20417 15519 20451
rect 16681 20417 16715 20451
rect 18225 20417 18259 20451
rect 18318 20417 18352 20451
rect 18429 20417 18463 20451
rect 18613 20417 18647 20451
rect 23029 20417 23063 20451
rect 23213 20417 23247 20451
rect 23765 20417 23799 20451
rect 24041 20417 24075 20451
rect 25053 20417 25087 20451
rect 28641 20417 28675 20451
rect 30205 20417 30239 20451
rect 30294 20423 30328 20457
rect 30389 20417 30423 20451
rect 30573 20417 30607 20451
rect 31401 20417 31435 20451
rect 36553 20417 36587 20451
rect 37473 20417 37507 20451
rect 38301 20417 38335 20451
rect 38485 20417 38519 20451
rect 40785 20417 40819 20451
rect 43453 20417 43487 20451
rect 44741 20417 44775 20451
rect 44830 20417 44864 20451
rect 44925 20417 44959 20451
rect 45109 20417 45143 20451
rect 45569 20417 45603 20451
rect 45753 20417 45787 20451
rect 46857 20417 46891 20451
rect 47593 20417 47627 20451
rect 11897 20349 11931 20383
rect 12173 20349 12207 20383
rect 15945 20349 15979 20383
rect 19165 20349 19199 20383
rect 22937 20349 22971 20383
rect 23121 20349 23155 20383
rect 23857 20349 23891 20383
rect 32137 20349 32171 20383
rect 33977 20349 34011 20383
rect 36369 20349 36403 20383
rect 37565 20349 37599 20383
rect 37841 20349 37875 20383
rect 41061 20349 41095 20383
rect 17969 20213 18003 20247
rect 23765 20213 23799 20247
rect 36277 20213 36311 20247
rect 38301 20213 38335 20247
rect 46949 20213 46983 20247
rect 11897 20009 11931 20043
rect 17141 20009 17175 20043
rect 22845 20009 22879 20043
rect 25789 20009 25823 20043
rect 28641 20009 28675 20043
rect 30481 20009 30515 20043
rect 32321 20009 32355 20043
rect 38209 20009 38243 20043
rect 40785 20009 40819 20043
rect 41245 20009 41279 20043
rect 19257 19941 19291 19975
rect 20637 19873 20671 19907
rect 22707 19873 22741 19907
rect 26617 19873 26651 19907
rect 37105 19873 37139 19907
rect 37381 19873 37415 19907
rect 40877 19873 40911 19907
rect 46305 19873 46339 19907
rect 11805 19805 11839 19839
rect 15761 19805 15795 19839
rect 16028 19805 16062 19839
rect 18225 19805 18259 19839
rect 18318 19805 18352 19839
rect 18434 19805 18468 19839
rect 18613 19805 18647 19839
rect 19441 19805 19475 19839
rect 22569 19805 22603 19839
rect 23029 19805 23063 19839
rect 25605 19805 25639 19839
rect 26341 19805 26375 19839
rect 26433 19805 26467 19839
rect 30113 19805 30147 19839
rect 31953 19805 31987 19839
rect 32137 19805 32171 19839
rect 37013 19805 37047 19839
rect 41061 19805 41095 19839
rect 48145 19805 48179 19839
rect 20904 19737 20938 19771
rect 28549 19737 28583 19771
rect 30297 19737 30331 19771
rect 31033 19737 31067 19771
rect 31217 19737 31251 19771
rect 38025 19737 38059 19771
rect 38225 19737 38259 19771
rect 40785 19737 40819 19771
rect 41705 19737 41739 19771
rect 41889 19737 41923 19771
rect 45109 19737 45143 19771
rect 45293 19737 45327 19771
rect 46489 19737 46523 19771
rect 17969 19669 18003 19703
rect 22017 19669 22051 19703
rect 23029 19669 23063 19703
rect 26617 19669 26651 19703
rect 38393 19669 38427 19703
rect 42073 19669 42107 19703
rect 45477 19669 45511 19703
rect 22293 19465 22327 19499
rect 27083 19465 27117 19499
rect 29285 19465 29319 19499
rect 39227 19465 39261 19499
rect 39313 19465 39347 19499
rect 46949 19465 46983 19499
rect 17141 19397 17175 19431
rect 34437 19397 34471 19431
rect 37565 19397 37599 19431
rect 41429 19397 41463 19431
rect 2237 19329 2271 19363
rect 17325 19329 17359 19363
rect 18199 19329 18233 19363
rect 18318 19329 18352 19363
rect 18434 19329 18468 19363
rect 18625 19329 18659 19363
rect 19993 19329 20027 19363
rect 21833 19329 21867 19363
rect 22293 19329 22327 19363
rect 23121 19329 23155 19363
rect 25513 19329 25547 19363
rect 26985 19329 27019 19363
rect 27169 19329 27203 19363
rect 27261 19329 27295 19363
rect 29193 19329 29227 19363
rect 30849 19329 30883 19363
rect 33425 19329 33459 19363
rect 33517 19329 33551 19363
rect 33609 19329 33643 19363
rect 33793 19329 33827 19363
rect 34253 19329 34287 19363
rect 37289 19329 37323 19363
rect 38209 19329 38243 19363
rect 38393 19329 38427 19363
rect 38485 19329 38519 19363
rect 39129 19329 39163 19363
rect 39405 19329 39439 19363
rect 40325 19329 40359 19363
rect 40417 19329 40451 19363
rect 42625 19329 42659 19363
rect 43361 19329 43395 19363
rect 44824 19329 44858 19363
rect 46857 19329 46891 19363
rect 47961 19329 47995 19363
rect 17509 19261 17543 19295
rect 23213 19261 23247 19295
rect 23397 19261 23431 19295
rect 25605 19261 25639 19295
rect 25789 19261 25823 19295
rect 37565 19261 37599 19295
rect 43085 19261 43119 19295
rect 44557 19261 44591 19295
rect 22109 19193 22143 19227
rect 22753 19193 22787 19227
rect 37381 19193 37415 19227
rect 40601 19193 40635 19227
rect 41061 19193 41095 19227
rect 41613 19193 41647 19227
rect 1777 19125 1811 19159
rect 2329 19125 2363 19159
rect 17969 19125 18003 19159
rect 19809 19125 19843 19159
rect 21971 19125 22005 19159
rect 25145 19125 25179 19159
rect 30941 19125 30975 19159
rect 33149 19125 33183 19159
rect 34621 19125 34655 19159
rect 38485 19125 38519 19159
rect 38669 19125 38703 19159
rect 41429 19125 41463 19159
rect 42441 19125 42475 19159
rect 45937 19125 45971 19159
rect 48053 19125 48087 19159
rect 18521 18921 18555 18955
rect 25559 18921 25593 18955
rect 32413 18921 32447 18955
rect 36093 18921 36127 18955
rect 37841 18921 37875 18955
rect 39129 18921 39163 18955
rect 40417 18921 40451 18955
rect 41429 18921 41463 18955
rect 22293 18853 22327 18887
rect 26985 18853 27019 18887
rect 37473 18853 37507 18887
rect 40601 18853 40635 18887
rect 41061 18853 41095 18887
rect 1409 18785 1443 18819
rect 1593 18785 1627 18819
rect 2789 18785 2823 18819
rect 22385 18785 22419 18819
rect 23121 18785 23155 18819
rect 31033 18785 31067 18819
rect 38761 18785 38795 18819
rect 46489 18785 46523 18819
rect 47133 18785 47167 18819
rect 16313 18717 16347 18751
rect 19349 18717 19383 18751
rect 19616 18717 19650 18751
rect 22109 18717 22143 18751
rect 22845 18717 22879 18751
rect 23029 18717 23063 18751
rect 23213 18717 23247 18751
rect 23397 18717 23431 18751
rect 24593 18717 24627 18751
rect 24777 18717 24811 18751
rect 24869 18717 24903 18751
rect 25329 18717 25363 18751
rect 26617 18717 26651 18751
rect 27445 18717 27479 18751
rect 29745 18717 29779 18751
rect 30021 18717 30055 18751
rect 33609 18717 33643 18751
rect 33701 18717 33735 18751
rect 33793 18717 33827 18751
rect 33977 18717 34011 18751
rect 34713 18717 34747 18751
rect 37749 18717 37783 18751
rect 37933 18717 37967 18751
rect 38025 18717 38059 18751
rect 38209 18717 38243 18751
rect 38853 18717 38887 18751
rect 42073 18717 42107 18751
rect 45247 18717 45281 18751
rect 45382 18717 45416 18751
rect 45477 18717 45511 18751
rect 45661 18717 45695 18751
rect 46305 18717 46339 18751
rect 16580 18649 16614 18683
rect 18153 18649 18187 18683
rect 18337 18649 18371 18683
rect 21925 18649 21959 18683
rect 26801 18649 26835 18683
rect 27712 18649 27746 18683
rect 31278 18649 31312 18683
rect 33333 18649 33367 18683
rect 34958 18649 34992 18683
rect 40233 18649 40267 18683
rect 42340 18649 42374 18683
rect 44097 18649 44131 18683
rect 44281 18649 44315 18683
rect 17693 18581 17727 18615
rect 20729 18581 20763 18615
rect 23581 18581 23615 18615
rect 24409 18581 24443 18615
rect 28825 18581 28859 18615
rect 40443 18581 40477 18615
rect 41429 18581 41463 18615
rect 41613 18581 41647 18615
rect 43453 18581 43487 18615
rect 44465 18581 44499 18615
rect 45017 18581 45051 18615
rect 20269 18377 20303 18411
rect 22017 18377 22051 18411
rect 22385 18377 22419 18411
rect 25697 18377 25731 18411
rect 27905 18377 27939 18411
rect 28549 18377 28583 18411
rect 30941 18377 30975 18411
rect 38669 18377 38703 18411
rect 41521 18377 41555 18411
rect 43821 18377 43855 18411
rect 46489 18377 46523 18411
rect 15301 18309 15335 18343
rect 15393 18309 15427 18343
rect 17040 18309 17074 18343
rect 20729 18309 20763 18343
rect 22937 18309 22971 18343
rect 32505 18309 32539 18343
rect 34222 18309 34256 18343
rect 41153 18309 41187 18343
rect 45354 18309 45388 18343
rect 2053 18241 2087 18275
rect 20637 18241 20671 18275
rect 22201 18241 22235 18275
rect 22477 18241 22511 18275
rect 23121 18241 23155 18275
rect 23213 18241 23247 18275
rect 23857 18241 23891 18275
rect 24961 18241 24995 18275
rect 26065 18241 26099 18275
rect 27169 18241 27203 18275
rect 27353 18241 27387 18275
rect 27537 18241 27571 18275
rect 27721 18241 27755 18275
rect 28365 18241 28399 18275
rect 30021 18241 30055 18275
rect 31217 18241 31251 18275
rect 31309 18241 31343 18275
rect 31401 18241 31435 18275
rect 31585 18241 31619 18275
rect 32137 18241 32171 18275
rect 32321 18241 32355 18275
rect 37473 18241 37507 18275
rect 38485 18241 38519 18275
rect 41337 18241 41371 18275
rect 42697 18241 42731 18275
rect 45109 18241 45143 18275
rect 47593 18241 47627 18275
rect 15577 18173 15611 18207
rect 16773 18173 16807 18207
rect 20913 18173 20947 18207
rect 25237 18173 25271 18207
rect 26157 18173 26191 18207
rect 26249 18173 26283 18207
rect 27445 18173 27479 18207
rect 29837 18173 29871 18207
rect 33977 18173 34011 18207
rect 37565 18173 37599 18207
rect 37841 18173 37875 18207
rect 38301 18173 38335 18207
rect 42441 18173 42475 18207
rect 18153 18105 18187 18139
rect 2145 18037 2179 18071
rect 2881 18037 2915 18071
rect 23121 18037 23155 18071
rect 23397 18037 23431 18071
rect 24041 18037 24075 18071
rect 25053 18037 25087 18071
rect 25145 18037 25179 18071
rect 30205 18037 30239 18071
rect 35357 18037 35391 18071
rect 47685 18037 47719 18071
rect 15853 17833 15887 17867
rect 23397 17833 23431 17867
rect 23673 17833 23707 17867
rect 25237 17833 25271 17867
rect 25697 17833 25731 17867
rect 28917 17833 28951 17867
rect 32873 17833 32907 17867
rect 34161 17833 34195 17867
rect 37933 17833 37967 17867
rect 41981 17833 42015 17867
rect 45017 17833 45051 17867
rect 19993 17765 20027 17799
rect 27629 17765 27663 17799
rect 1409 17697 1443 17731
rect 1593 17697 1627 17731
rect 2789 17697 2823 17731
rect 20637 17697 20671 17731
rect 31401 17697 31435 17731
rect 39957 17697 39991 17731
rect 46305 17697 46339 17731
rect 46489 17697 46523 17731
rect 48145 17697 48179 17731
rect 15761 17629 15795 17663
rect 23213 17629 23247 17663
rect 23397 17629 23431 17663
rect 23489 17629 23523 17663
rect 25421 17629 25455 17663
rect 25513 17629 25547 17663
rect 25789 17629 25823 17663
rect 26341 17629 26375 17663
rect 27445 17629 27479 17663
rect 28733 17629 28767 17663
rect 29561 17629 29595 17663
rect 31677 17629 31711 17663
rect 32781 17629 32815 17663
rect 37933 17629 37967 17663
rect 38117 17629 38151 17663
rect 40233 17629 40267 17663
rect 41245 17629 41279 17663
rect 41429 17629 41463 17663
rect 42165 17629 42199 17663
rect 43269 17629 43303 17663
rect 45247 17629 45281 17663
rect 45385 17629 45419 17663
rect 45482 17629 45516 17663
rect 45661 17629 45695 17663
rect 17509 17561 17543 17595
rect 17877 17561 17911 17595
rect 22569 17561 22603 17595
rect 22753 17561 22787 17595
rect 26525 17561 26559 17595
rect 29828 17561 29862 17595
rect 33793 17561 33827 17595
rect 33977 17561 34011 17595
rect 20361 17493 20395 17527
rect 20453 17493 20487 17527
rect 30941 17493 30975 17527
rect 41429 17493 41463 17527
rect 43085 17493 43119 17527
rect 23029 17289 23063 17323
rect 29837 17289 29871 17323
rect 36001 17289 36035 17323
rect 40969 17289 41003 17323
rect 41629 17289 41663 17323
rect 2053 17221 2087 17255
rect 16037 17221 16071 17255
rect 16865 17221 16899 17255
rect 23949 17221 23983 17255
rect 26249 17221 26283 17255
rect 31125 17221 31159 17255
rect 33885 17221 33919 17255
rect 34069 17221 34103 17255
rect 39865 17221 39899 17255
rect 40601 17221 40635 17255
rect 41429 17221 41463 17255
rect 45385 17221 45419 17255
rect 47685 17221 47719 17255
rect 1869 17153 1903 17187
rect 15945 17153 15979 17187
rect 16681 17153 16715 17187
rect 19248 17153 19282 17187
rect 22937 17153 22971 17187
rect 23765 17153 23799 17187
rect 25513 17153 25547 17187
rect 25697 17153 25731 17187
rect 27721 17153 27755 17187
rect 30021 17153 30055 17187
rect 30113 17153 30147 17187
rect 30297 17153 30331 17187
rect 30389 17153 30423 17187
rect 30941 17153 30975 17187
rect 35909 17153 35943 17187
rect 37749 17153 37783 17187
rect 40049 17153 40083 17187
rect 40141 17153 40175 17187
rect 40785 17153 40819 17187
rect 47593 17153 47627 17187
rect 18337 17085 18371 17119
rect 18981 17085 19015 17119
rect 45201 17085 45235 17119
rect 46857 17085 46891 17119
rect 37933 17017 37967 17051
rect 40141 17017 40175 17051
rect 2697 16949 2731 16983
rect 20361 16949 20395 16983
rect 25605 16949 25639 16983
rect 26341 16949 26375 16983
rect 27997 16949 28031 16983
rect 34253 16949 34287 16983
rect 41613 16949 41647 16983
rect 41797 16949 41831 16983
rect 17877 16745 17911 16779
rect 23121 16745 23155 16779
rect 25145 16745 25179 16779
rect 26157 16745 26191 16779
rect 42165 16745 42199 16779
rect 45845 16745 45879 16779
rect 23305 16677 23339 16711
rect 26985 16677 27019 16711
rect 27905 16677 27939 16711
rect 37657 16677 37691 16711
rect 1409 16609 1443 16643
rect 2237 16609 2271 16643
rect 20269 16609 20303 16643
rect 23213 16609 23247 16643
rect 40141 16609 40175 16643
rect 46305 16609 46339 16643
rect 15945 16541 15979 16575
rect 19257 16541 19291 16575
rect 22109 16541 22143 16575
rect 22293 16541 22327 16575
rect 23029 16541 23063 16575
rect 23489 16541 23523 16575
rect 25053 16541 25087 16575
rect 25697 16541 25731 16575
rect 25881 16541 25915 16575
rect 25973 16541 26007 16575
rect 26249 16541 26283 16575
rect 27721 16541 27755 16575
rect 30757 16541 30791 16575
rect 31585 16541 31619 16575
rect 33701 16541 33735 16575
rect 33793 16541 33827 16575
rect 33885 16541 33919 16575
rect 34069 16541 34103 16575
rect 38669 16541 38703 16575
rect 39221 16541 39255 16575
rect 1593 16473 1627 16507
rect 16589 16473 16623 16507
rect 19533 16473 19567 16507
rect 20536 16473 20570 16507
rect 26801 16473 26835 16507
rect 30941 16473 30975 16507
rect 31852 16473 31886 16507
rect 36369 16473 36403 16507
rect 40408 16473 40442 16507
rect 41981 16473 42015 16507
rect 46489 16473 46523 16507
rect 48145 16473 48179 16507
rect 16037 16405 16071 16439
rect 21649 16405 21683 16439
rect 22201 16405 22235 16439
rect 22753 16405 22787 16439
rect 31125 16405 31159 16439
rect 32965 16405 32999 16439
rect 33425 16405 33459 16439
rect 41521 16405 41555 16439
rect 42181 16405 42215 16439
rect 42349 16405 42383 16439
rect 2237 16201 2271 16235
rect 20637 16201 20671 16235
rect 23673 16201 23707 16235
rect 32137 16201 32171 16235
rect 35541 16201 35575 16235
rect 40693 16201 40727 16235
rect 41245 16201 41279 16235
rect 46489 16201 46523 16235
rect 17049 16133 17083 16167
rect 33701 16133 33735 16167
rect 2145 16065 2179 16099
rect 14013 16065 14047 16099
rect 19257 16065 19291 16099
rect 20821 16065 20855 16099
rect 21833 16065 21867 16099
rect 22005 16065 22039 16099
rect 22118 16065 22152 16099
rect 22339 16065 22373 16099
rect 23489 16065 23523 16099
rect 24133 16065 24167 16099
rect 24317 16065 24351 16099
rect 24961 16065 24995 16099
rect 29469 16065 29503 16099
rect 30573 16065 30607 16099
rect 30665 16065 30699 16099
rect 30757 16065 30791 16099
rect 30941 16065 30975 16099
rect 32413 16065 32447 16099
rect 32505 16065 32539 16099
rect 32597 16065 32631 16099
rect 32781 16065 32815 16099
rect 33517 16065 33551 16099
rect 34417 16065 34451 16099
rect 37473 16065 37507 16099
rect 39037 16065 39071 16099
rect 39126 16068 39160 16102
rect 39221 16065 39255 16099
rect 39405 16065 39439 16099
rect 40509 16065 40543 16099
rect 40785 16065 40819 16099
rect 41429 16065 41463 16099
rect 42625 16065 42659 16099
rect 46397 16065 46431 16099
rect 47593 16065 47627 16099
rect 14197 15997 14231 16031
rect 14473 15997 14507 16031
rect 16865 15997 16899 16031
rect 18245 15997 18279 16031
rect 19901 15997 19935 16031
rect 22201 15997 22235 16031
rect 22569 15997 22603 16031
rect 23305 15997 23339 16031
rect 25053 15997 25087 16031
rect 29653 15997 29687 16031
rect 34161 15997 34195 16031
rect 40325 15997 40359 16031
rect 24501 15929 24535 15963
rect 37657 15929 37691 15963
rect 30297 15861 30331 15895
rect 38761 15861 38795 15895
rect 42441 15861 42475 15895
rect 45937 15861 45971 15895
rect 47685 15861 47719 15895
rect 14197 15657 14231 15691
rect 21925 15657 21959 15691
rect 31953 15657 31987 15691
rect 39037 15657 39071 15691
rect 24685 15589 24719 15623
rect 25329 15589 25363 15623
rect 16773 15521 16807 15555
rect 18153 15521 18187 15555
rect 20637 15521 20671 15555
rect 26525 15521 26559 15555
rect 38117 15521 38151 15555
rect 40325 15521 40359 15555
rect 46305 15521 46339 15555
rect 46489 15521 46523 15555
rect 48145 15521 48179 15555
rect 14105 15453 14139 15487
rect 15393 15453 15427 15487
rect 16037 15453 16071 15487
rect 22477 15453 22511 15487
rect 22744 15453 22778 15487
rect 24409 15453 24443 15487
rect 24593 15453 24627 15487
rect 25237 15453 25271 15487
rect 25421 15453 25455 15487
rect 26341 15453 26375 15487
rect 27629 15453 27663 15487
rect 30573 15453 30607 15487
rect 30829 15453 30863 15487
rect 36921 15453 36955 15487
rect 37013 15453 37047 15487
rect 37105 15453 37139 15487
rect 37289 15453 37323 15487
rect 37749 15453 37783 15487
rect 38669 15453 38703 15487
rect 40592 15453 40626 15487
rect 15485 15385 15519 15419
rect 16957 15385 16991 15419
rect 20453 15385 20487 15419
rect 21833 15385 21867 15419
rect 27896 15385 27930 15419
rect 34713 15385 34747 15419
rect 34897 15385 34931 15419
rect 37933 15385 37967 15419
rect 38853 15385 38887 15419
rect 16221 15317 16255 15351
rect 19993 15317 20027 15351
rect 20361 15317 20395 15351
rect 23857 15317 23891 15351
rect 25973 15317 26007 15351
rect 26433 15317 26467 15351
rect 29009 15317 29043 15351
rect 35081 15317 35115 15351
rect 36645 15317 36679 15351
rect 41705 15317 41739 15351
rect 27445 15113 27479 15147
rect 30297 15113 30331 15147
rect 46857 15113 46891 15147
rect 16037 15045 16071 15079
rect 16865 15045 16899 15079
rect 18981 15045 19015 15079
rect 21833 15045 21867 15079
rect 22845 15045 22879 15079
rect 24869 15045 24903 15079
rect 25053 15045 25087 15079
rect 27905 15045 27939 15079
rect 28641 15045 28675 15079
rect 30113 15045 30147 15079
rect 36645 15045 36679 15079
rect 37473 15045 37507 15079
rect 15945 14977 15979 15011
rect 22017 14977 22051 15011
rect 22109 14977 22143 15011
rect 22385 14977 22419 15011
rect 23029 14977 23063 15011
rect 23213 14977 23247 15011
rect 23305 14977 23339 15011
rect 24041 14977 24075 15011
rect 26065 14977 26099 15011
rect 27813 14977 27847 15011
rect 28917 14977 28951 15011
rect 29929 14977 29963 15011
rect 31197 14977 31231 15011
rect 31306 14980 31340 15014
rect 31406 14977 31440 15011
rect 31585 14977 31619 15011
rect 32137 14977 32171 15011
rect 32393 14977 32427 15011
rect 34345 14977 34379 15011
rect 34612 14977 34646 15011
rect 36553 14977 36587 15011
rect 39589 14977 39623 15011
rect 39845 14977 39879 15011
rect 47041 14977 47075 15011
rect 16681 14909 16715 14943
rect 18245 14909 18279 14943
rect 26157 14909 26191 14943
rect 27997 14909 28031 14943
rect 28733 14909 28767 14943
rect 37289 14909 37323 14943
rect 39037 14909 39071 14943
rect 30573 14841 30607 14875
rect 30941 14841 30975 14875
rect 35725 14841 35759 14875
rect 20269 14773 20303 14807
rect 22293 14773 22327 14807
rect 24225 14773 24259 14807
rect 26157 14773 26191 14807
rect 26433 14773 26467 14807
rect 28733 14773 28767 14807
rect 29101 14773 29135 14807
rect 33517 14773 33551 14807
rect 40969 14773 41003 14807
rect 47777 14773 47811 14807
rect 16957 14569 16991 14603
rect 25421 14569 25455 14603
rect 26709 14569 26743 14603
rect 31493 14569 31527 14603
rect 34713 14569 34747 14603
rect 37841 14569 37875 14603
rect 20637 14501 20671 14535
rect 22017 14501 22051 14535
rect 26985 14501 27019 14535
rect 32689 14501 32723 14535
rect 34161 14501 34195 14535
rect 19257 14433 19291 14467
rect 22477 14433 22511 14467
rect 22661 14433 22695 14467
rect 25697 14433 25731 14467
rect 27813 14433 27847 14467
rect 36461 14433 36495 14467
rect 46305 14433 46339 14467
rect 2053 14365 2087 14399
rect 16865 14365 16899 14399
rect 17693 14365 17727 14399
rect 21281 14365 21315 14399
rect 22385 14365 22419 14399
rect 24777 14365 24811 14399
rect 25605 14365 25639 14399
rect 25789 14365 25823 14399
rect 25881 14365 25915 14399
rect 26433 14365 26467 14399
rect 26709 14365 26743 14399
rect 27537 14365 27571 14399
rect 27721 14365 27755 14399
rect 27905 14365 27939 14399
rect 28089 14365 28123 14399
rect 28273 14365 28307 14399
rect 32505 14365 32539 14399
rect 34943 14365 34977 14399
rect 35081 14365 35115 14399
rect 35178 14362 35212 14396
rect 35357 14365 35391 14399
rect 36728 14365 36762 14399
rect 38393 14365 38427 14399
rect 18521 14297 18555 14331
rect 19524 14297 19558 14331
rect 21465 14297 21499 14331
rect 31125 14297 31159 14331
rect 31309 14297 31343 14331
rect 33977 14297 34011 14331
rect 46489 14297 46523 14331
rect 48145 14297 48179 14331
rect 24869 14229 24903 14263
rect 38485 14229 38519 14263
rect 20085 14025 20119 14059
rect 21189 14025 21223 14059
rect 23213 14025 23247 14059
rect 46765 14025 46799 14059
rect 48053 14025 48087 14059
rect 19625 13957 19659 13991
rect 25053 13957 25087 13991
rect 28917 13957 28951 13991
rect 32873 13957 32907 13991
rect 33517 13957 33551 13991
rect 33885 13957 33919 13991
rect 35633 13957 35667 13991
rect 38485 13957 38519 13991
rect 1777 13889 1811 13923
rect 16681 13889 16715 13923
rect 17693 13889 17727 13923
rect 19257 13889 19291 13923
rect 20269 13889 20303 13923
rect 21097 13889 21131 13923
rect 21281 13889 21315 13923
rect 22201 13889 22235 13923
rect 23121 13889 23155 13923
rect 24409 13889 24443 13923
rect 25329 13889 25363 13923
rect 26157 13889 26191 13923
rect 27721 13889 27755 13923
rect 32137 13889 32171 13923
rect 33701 13889 33735 13923
rect 34575 13889 34609 13923
rect 34694 13889 34728 13923
rect 34805 13892 34839 13926
rect 34989 13889 35023 13923
rect 35449 13889 35483 13923
rect 46673 13889 46707 13923
rect 47869 13889 47903 13923
rect 1961 13821 1995 13855
rect 2789 13821 2823 13855
rect 18061 13821 18095 13855
rect 22293 13821 22327 13855
rect 22477 13821 22511 13855
rect 25237 13821 25271 13855
rect 26433 13821 26467 13855
rect 27813 13821 27847 13855
rect 27905 13821 27939 13855
rect 29101 13821 29135 13855
rect 30113 13821 30147 13855
rect 30389 13821 30423 13855
rect 33057 13821 33091 13855
rect 35817 13821 35851 13855
rect 38301 13821 38335 13855
rect 39957 13821 39991 13855
rect 21833 13753 21867 13787
rect 24593 13753 24627 13787
rect 25973 13753 26007 13787
rect 16773 13685 16807 13719
rect 25329 13685 25363 13719
rect 25513 13685 25547 13719
rect 26341 13685 26375 13719
rect 27353 13685 27387 13719
rect 32229 13685 32263 13719
rect 34345 13685 34379 13719
rect 2145 13481 2179 13515
rect 21465 13481 21499 13515
rect 22569 13481 22603 13515
rect 23581 13481 23615 13515
rect 29009 13481 29043 13515
rect 31769 13481 31803 13515
rect 26985 13413 27019 13447
rect 19257 13345 19291 13379
rect 21373 13345 21407 13379
rect 24869 13345 24903 13379
rect 24961 13345 24995 13379
rect 26525 13345 26559 13379
rect 27721 13345 27755 13379
rect 27813 13345 27847 13379
rect 30665 13345 30699 13379
rect 32321 13345 32355 13379
rect 32505 13345 32539 13379
rect 33701 13345 33735 13379
rect 34713 13345 34747 13379
rect 2053 13277 2087 13311
rect 18337 13277 18371 13311
rect 18429 13277 18463 13311
rect 18521 13277 18555 13311
rect 18705 13277 18739 13311
rect 19533 13277 19567 13311
rect 21281 13277 21315 13311
rect 22109 13277 22143 13311
rect 22385 13277 22419 13311
rect 22569 13277 22603 13311
rect 23397 13277 23431 13311
rect 26617 13277 26651 13311
rect 27445 13277 27479 13311
rect 27629 13277 27663 13311
rect 27997 13277 28031 13311
rect 30481 13277 30515 13311
rect 31677 13277 31711 13311
rect 23213 13209 23247 13243
rect 28641 13209 28675 13243
rect 28825 13209 28859 13243
rect 34958 13209 34992 13243
rect 18061 13141 18095 13175
rect 21649 13141 21683 13175
rect 22753 13141 22787 13175
rect 24409 13141 24443 13175
rect 24777 13141 24811 13175
rect 28181 13141 28215 13175
rect 36093 13141 36127 13175
rect 1593 12937 1627 12971
rect 26249 12937 26283 12971
rect 29653 12937 29687 12971
rect 16865 12869 16899 12903
rect 25053 12869 25087 12903
rect 26157 12869 26191 12903
rect 34682 12869 34716 12903
rect 1409 12801 1443 12835
rect 20637 12801 20671 12835
rect 22017 12801 22051 12835
rect 22293 12801 22327 12835
rect 23121 12801 23155 12835
rect 25329 12801 25363 12835
rect 26985 12801 27019 12835
rect 28529 12801 28563 12835
rect 30389 12801 30423 12835
rect 32137 12801 32171 12835
rect 32393 12801 32427 12835
rect 34437 12801 34471 12835
rect 16681 12733 16715 12767
rect 17141 12733 17175 12767
rect 19349 12733 19383 12767
rect 19625 12733 19659 12767
rect 22201 12733 22235 12767
rect 23397 12733 23431 12767
rect 25237 12733 25271 12767
rect 27261 12733 27295 12767
rect 28273 12733 28307 12767
rect 30665 12733 30699 12767
rect 20729 12597 20763 12631
rect 21833 12597 21867 12631
rect 25053 12597 25087 12631
rect 25513 12597 25547 12631
rect 27077 12597 27111 12631
rect 27537 12597 27571 12631
rect 33517 12597 33551 12631
rect 35817 12597 35851 12631
rect 17877 12393 17911 12427
rect 18705 12393 18739 12427
rect 21649 12393 21683 12427
rect 22937 12393 22971 12427
rect 25329 12393 25363 12427
rect 25789 12393 25823 12427
rect 31309 12393 31343 12427
rect 34713 12393 34747 12427
rect 19441 12257 19475 12291
rect 22293 12257 22327 12291
rect 27813 12257 27847 12291
rect 32781 12257 32815 12291
rect 16497 12189 16531 12223
rect 18521 12189 18555 12223
rect 19257 12189 19291 12223
rect 22109 12189 22143 12223
rect 22845 12189 22879 12223
rect 23213 12189 23247 12223
rect 24685 12189 24719 12223
rect 24869 12189 24903 12223
rect 25513 12189 25547 12223
rect 25645 12189 25679 12223
rect 27721 12189 27755 12223
rect 30481 12189 30515 12223
rect 31585 12189 31619 12223
rect 31677 12189 31711 12223
rect 31769 12189 31803 12223
rect 31953 12189 31987 12223
rect 32597 12189 32631 12223
rect 33241 12189 33275 12223
rect 34989 12189 35023 12223
rect 35081 12189 35115 12223
rect 35173 12189 35207 12223
rect 35357 12189 35391 12223
rect 35909 12189 35943 12223
rect 16764 12121 16798 12155
rect 18337 12121 18371 12155
rect 21097 12121 21131 12155
rect 25329 12121 25363 12155
rect 30665 12121 30699 12155
rect 32413 12121 32447 12155
rect 22017 12053 22051 12087
rect 23397 12053 23431 12087
rect 27261 12053 27295 12087
rect 27629 12053 27663 12087
rect 33333 12053 33367 12087
rect 36093 12053 36127 12087
rect 19165 11849 19199 11883
rect 25513 11849 25547 11883
rect 29193 11849 29227 11883
rect 18052 11781 18086 11815
rect 19625 11781 19659 11815
rect 32505 11781 32539 11815
rect 33333 11781 33367 11815
rect 2053 11713 2087 11747
rect 19901 11713 19935 11747
rect 19993 11713 20027 11747
rect 20085 11713 20119 11747
rect 20269 11713 20303 11747
rect 21833 11713 21867 11747
rect 22017 11713 22051 11747
rect 22109 11713 22143 11747
rect 22385 11713 22419 11747
rect 23213 11713 23247 11747
rect 23489 11713 23523 11747
rect 25697 11713 25731 11747
rect 28080 11713 28114 11747
rect 30297 11713 30331 11747
rect 31171 11713 31205 11747
rect 31309 11713 31343 11747
rect 31422 11713 31456 11747
rect 31585 11713 31619 11747
rect 32137 11713 32171 11747
rect 32321 11713 32355 11747
rect 33149 11713 33183 11747
rect 17785 11645 17819 11679
rect 22201 11645 22235 11679
rect 25973 11645 26007 11679
rect 27813 11645 27847 11679
rect 34345 11645 34379 11679
rect 30481 11577 30515 11611
rect 2145 11509 2179 11543
rect 22569 11509 22603 11543
rect 23029 11509 23063 11543
rect 23397 11509 23431 11543
rect 25881 11509 25915 11543
rect 30941 11509 30975 11543
rect 47777 11509 47811 11543
rect 19625 11305 19659 11339
rect 21833 11305 21867 11339
rect 23765 11305 23799 11339
rect 25789 11305 25823 11339
rect 27997 11305 28031 11339
rect 32873 11237 32907 11271
rect 1593 11169 1627 11203
rect 2789 11169 2823 11203
rect 26617 11169 26651 11203
rect 27537 11169 27571 11203
rect 46305 11169 46339 11203
rect 1409 11101 1443 11135
rect 19441 11101 19475 11135
rect 20453 11101 20487 11135
rect 22385 11101 22419 11135
rect 25605 11101 25639 11135
rect 25881 11101 25915 11135
rect 27261 11101 27295 11135
rect 27445 11101 27479 11135
rect 27629 11101 27663 11135
rect 27813 11101 27847 11135
rect 28549 11101 28583 11135
rect 30021 11101 30055 11135
rect 31493 11101 31527 11135
rect 31760 11101 31794 11135
rect 19257 11033 19291 11067
rect 20720 11033 20754 11067
rect 22652 11033 22686 11067
rect 24593 11033 24627 11067
rect 24777 11033 24811 11067
rect 24961 11033 24995 11067
rect 26433 11033 26467 11067
rect 28733 11033 28767 11067
rect 46489 11033 46523 11067
rect 48145 11033 48179 11067
rect 25421 10965 25455 10999
rect 30113 10965 30147 10999
rect 23397 10761 23431 10795
rect 24041 10761 24075 10795
rect 46949 10761 46983 10795
rect 23121 10693 23155 10727
rect 25237 10693 25271 10727
rect 26065 10693 26099 10727
rect 26249 10693 26283 10727
rect 1409 10625 1443 10659
rect 2329 10625 2363 10659
rect 18797 10625 18831 10659
rect 18889 10625 18923 10659
rect 18981 10625 19015 10659
rect 19165 10625 19199 10659
rect 22845 10625 22879 10659
rect 23029 10625 23063 10659
rect 23213 10625 23247 10659
rect 23857 10625 23891 10659
rect 24133 10625 24167 10659
rect 24961 10625 24995 10659
rect 25145 10625 25179 10659
rect 25329 10625 25363 10659
rect 26341 10625 26375 10659
rect 26985 10625 27019 10659
rect 27169 10625 27203 10659
rect 28549 10625 28583 10659
rect 30067 10625 30101 10659
rect 30202 10625 30236 10659
rect 30297 10625 30331 10659
rect 30481 10625 30515 10659
rect 32597 10625 32631 10659
rect 46857 10625 46891 10659
rect 47869 10625 47903 10659
rect 28825 10557 28859 10591
rect 33241 10557 33275 10591
rect 33425 10557 33459 10591
rect 34621 10557 34655 10591
rect 1593 10489 1627 10523
rect 26065 10489 26099 10523
rect 32689 10489 32723 10523
rect 48053 10489 48087 10523
rect 18521 10421 18555 10455
rect 23857 10421 23891 10455
rect 25513 10421 25547 10455
rect 27077 10421 27111 10455
rect 29837 10421 29871 10455
rect 23029 10217 23063 10251
rect 25421 10217 25455 10251
rect 26249 10217 26283 10251
rect 27353 10217 27387 10251
rect 29009 10217 29043 10251
rect 32965 10217 32999 10251
rect 25421 10081 25455 10115
rect 26341 10081 26375 10115
rect 31585 10081 31619 10115
rect 2053 10013 2087 10047
rect 16865 10013 16899 10047
rect 19349 10013 19383 10047
rect 19717 10013 19751 10047
rect 22937 10013 22971 10047
rect 23121 10013 23155 10047
rect 24593 10013 24627 10047
rect 25513 10013 25547 10047
rect 26525 10013 26559 10047
rect 28825 10013 28859 10047
rect 29561 10013 29595 10047
rect 17132 9945 17166 9979
rect 19533 9945 19567 9979
rect 22017 9945 22051 9979
rect 23673 9945 23707 9979
rect 24777 9945 24811 9979
rect 25237 9945 25271 9979
rect 26249 9945 26283 9979
rect 27261 9945 27295 9979
rect 28641 9945 28675 9979
rect 29828 9945 29862 9979
rect 31830 9945 31864 9979
rect 18245 9877 18279 9911
rect 22109 9877 22143 9911
rect 23765 9877 23799 9911
rect 25697 9877 25731 9911
rect 26709 9877 26743 9911
rect 30941 9877 30975 9911
rect 18429 9673 18463 9707
rect 22569 9673 22603 9707
rect 25697 9673 25731 9707
rect 26157 9673 26191 9707
rect 27169 9673 27203 9707
rect 30941 9673 30975 9707
rect 27537 9605 27571 9639
rect 32321 9605 32355 9639
rect 1777 9537 1811 9571
rect 17417 9537 17451 9571
rect 18061 9537 18095 9571
rect 18245 9537 18279 9571
rect 19717 9537 19751 9571
rect 19809 9537 19843 9571
rect 19901 9537 19935 9571
rect 20085 9537 20119 9571
rect 22385 9537 22419 9571
rect 22661 9537 22695 9571
rect 23765 9537 23799 9571
rect 23949 9537 23983 9571
rect 24409 9537 24443 9571
rect 26065 9537 26099 9571
rect 31217 9537 31251 9571
rect 31306 9543 31340 9577
rect 31406 9537 31440 9571
rect 31597 9537 31631 9571
rect 32137 9537 32171 9571
rect 1961 9469 1995 9503
rect 2789 9469 2823 9503
rect 24685 9469 24719 9503
rect 26341 9469 26375 9503
rect 27629 9469 27663 9503
rect 27721 9469 27755 9503
rect 32505 9469 32539 9503
rect 17509 9333 17543 9367
rect 19441 9333 19475 9367
rect 22385 9333 22419 9367
rect 23765 9333 23799 9367
rect 24501 9333 24535 9367
rect 24961 9333 24995 9367
rect 2237 9129 2271 9163
rect 23397 9129 23431 9163
rect 25605 9129 25639 9163
rect 47869 9129 47903 9163
rect 21373 9061 21407 9095
rect 22753 9061 22787 9095
rect 26985 9061 27019 9095
rect 16865 8993 16899 9027
rect 17049 8993 17083 9027
rect 17325 8993 17359 9027
rect 21557 8993 21591 9027
rect 22293 8993 22327 9027
rect 27445 8993 27479 9027
rect 2145 8925 2179 8959
rect 19257 8925 19291 8959
rect 19524 8925 19558 8959
rect 21281 8925 21315 8959
rect 22017 8925 22051 8959
rect 22201 8925 22235 8959
rect 22385 8925 22419 8959
rect 22569 8925 22603 8959
rect 23581 8925 23615 8959
rect 23765 8925 23799 8959
rect 23857 8925 23891 8959
rect 24409 8925 24443 8959
rect 24593 8925 24627 8959
rect 24685 8925 24719 8959
rect 24777 8925 24811 8959
rect 24972 8925 25006 8959
rect 25789 8925 25823 8959
rect 25881 8925 25915 8959
rect 26065 8925 26099 8959
rect 26167 8925 26201 8959
rect 30895 8925 30929 8959
rect 31033 8925 31067 8959
rect 31130 8925 31164 8959
rect 31309 8925 31343 8959
rect 26617 8857 26651 8891
rect 26801 8857 26835 8891
rect 27712 8857 27746 8891
rect 47777 8857 47811 8891
rect 20637 8789 20671 8823
rect 21557 8789 21591 8823
rect 25145 8789 25179 8823
rect 28825 8789 28859 8823
rect 30665 8789 30699 8823
rect 24041 8585 24075 8619
rect 24409 8585 24443 8619
rect 25697 8585 25731 8619
rect 27905 8585 27939 8619
rect 31585 8585 31619 8619
rect 32505 8585 32539 8619
rect 2237 8517 2271 8551
rect 22100 8517 22134 8551
rect 24501 8517 24535 8551
rect 30472 8517 30506 8551
rect 1869 8449 1903 8483
rect 17601 8449 17635 8483
rect 17868 8449 17902 8483
rect 25237 8449 25271 8483
rect 25513 8449 25547 8483
rect 27169 8449 27203 8483
rect 27353 8449 27387 8483
rect 27721 8449 27755 8483
rect 29377 8449 29411 8483
rect 29466 8455 29500 8489
rect 29561 8452 29595 8486
rect 29745 8449 29779 8483
rect 30205 8449 30239 8483
rect 32137 8449 32171 8483
rect 32321 8449 32355 8483
rect 47869 8449 47903 8483
rect 19441 8381 19475 8415
rect 19625 8381 19659 8415
rect 21281 8381 21315 8415
rect 21833 8381 21867 8415
rect 24593 8381 24627 8415
rect 25329 8381 25363 8415
rect 27445 8381 27479 8415
rect 27537 8381 27571 8415
rect 48053 8313 48087 8347
rect 18981 8245 19015 8279
rect 23213 8245 23247 8279
rect 25329 8245 25363 8279
rect 29101 8245 29135 8279
rect 30021 8041 30055 8075
rect 22109 7973 22143 8007
rect 26617 7973 26651 8007
rect 2145 7905 2179 7939
rect 19257 7905 19291 7939
rect 19717 7905 19751 7939
rect 22753 7905 22787 7939
rect 30481 7905 30515 7939
rect 31861 7905 31895 7939
rect 18337 7837 18371 7871
rect 18521 7837 18555 7871
rect 22569 7837 22603 7871
rect 25237 7837 25271 7871
rect 29653 7837 29687 7871
rect 46305 7837 46339 7871
rect 1869 7769 1903 7803
rect 19441 7769 19475 7803
rect 25504 7769 25538 7803
rect 29837 7769 29871 7803
rect 30665 7769 30699 7803
rect 46489 7769 46523 7803
rect 48145 7769 48179 7803
rect 18705 7701 18739 7735
rect 22477 7701 22511 7735
rect 18521 7497 18555 7531
rect 19349 7497 19383 7531
rect 24869 7497 24903 7531
rect 30941 7497 30975 7531
rect 46765 7497 46799 7531
rect 29254 7429 29288 7463
rect 18429 7361 18463 7395
rect 19625 7361 19659 7395
rect 19730 7361 19764 7395
rect 19830 7361 19864 7395
rect 19993 7361 20027 7395
rect 23489 7361 23523 7395
rect 23756 7361 23790 7395
rect 28365 7361 28399 7395
rect 30849 7361 30883 7395
rect 46673 7361 46707 7395
rect 47777 7361 47811 7395
rect 29009 7293 29043 7327
rect 2329 7157 2363 7191
rect 28457 7157 28491 7191
rect 30389 7157 30423 7191
rect 19441 6953 19475 6987
rect 29561 6817 29595 6851
rect 29745 6817 29779 6851
rect 30941 6817 30975 6851
rect 45661 6817 45695 6851
rect 46857 6817 46891 6851
rect 2973 6749 3007 6783
rect 19349 6749 19383 6783
rect 21097 6749 21131 6783
rect 20913 6681 20947 6715
rect 45845 6681 45879 6715
rect 3065 6613 3099 6647
rect 21281 6613 21315 6647
rect 45937 6409 45971 6443
rect 2237 6341 2271 6375
rect 20821 6341 20855 6375
rect 21005 6341 21039 6375
rect 27629 6341 27663 6375
rect 2053 6273 2087 6307
rect 23673 6273 23707 6307
rect 23765 6273 23799 6307
rect 23857 6273 23891 6307
rect 24041 6273 24075 6307
rect 27813 6273 27847 6307
rect 45845 6273 45879 6307
rect 2789 6205 2823 6239
rect 1593 6069 1627 6103
rect 21189 6069 21223 6103
rect 23397 6069 23431 6103
rect 27997 6069 28031 6103
rect 47777 6069 47811 6103
rect 28549 5865 28583 5899
rect 22017 5797 22051 5831
rect 25789 5797 25823 5831
rect 24409 5729 24443 5763
rect 27169 5729 27203 5763
rect 46305 5729 46339 5763
rect 1777 5661 1811 5695
rect 2237 5661 2271 5695
rect 2881 5661 2915 5695
rect 20637 5661 20671 5695
rect 22707 5661 22741 5695
rect 22845 5661 22879 5695
rect 22937 5661 22971 5695
rect 23121 5661 23155 5695
rect 24665 5661 24699 5695
rect 20904 5593 20938 5627
rect 22477 5593 22511 5627
rect 27436 5593 27470 5627
rect 46489 5593 46523 5627
rect 48145 5593 48179 5627
rect 2329 5525 2363 5559
rect 2973 5525 3007 5559
rect 23213 5321 23247 5355
rect 24041 5321 24075 5355
rect 27721 5321 27755 5355
rect 46949 5321 46983 5355
rect 1961 5253 1995 5287
rect 20637 5253 20671 5287
rect 22078 5253 22112 5287
rect 23673 5253 23707 5287
rect 1777 5185 1811 5219
rect 20867 5185 20901 5219
rect 21005 5185 21039 5219
rect 21118 5188 21152 5222
rect 21281 5185 21315 5219
rect 21833 5185 21867 5219
rect 23857 5185 23891 5219
rect 27997 5185 28031 5219
rect 28089 5185 28123 5219
rect 28181 5185 28215 5219
rect 28365 5185 28399 5219
rect 46857 5185 46891 5219
rect 47869 5185 47903 5219
rect 2789 5117 2823 5151
rect 48053 5049 48087 5083
rect 1409 4641 1443 4675
rect 2789 4641 2823 4675
rect 30941 4641 30975 4675
rect 6469 4573 6503 4607
rect 13369 4573 13403 4607
rect 30297 4573 30331 4607
rect 41981 4573 42015 4607
rect 45845 4573 45879 4607
rect 46305 4573 46339 4607
rect 1593 4505 1627 4539
rect 30481 4505 30515 4539
rect 46489 4505 46523 4539
rect 48145 4505 48179 4539
rect 22017 4165 22051 4199
rect 47961 4165 47995 4199
rect 1593 4097 1627 4131
rect 2237 4097 2271 4131
rect 3065 4097 3099 4131
rect 6377 4097 6411 4131
rect 7021 4097 7055 4131
rect 13185 4097 13219 4131
rect 20913 4097 20947 4131
rect 21005 4097 21039 4131
rect 29653 4097 29687 4131
rect 30573 4097 30607 4131
rect 36369 4097 36403 4131
rect 38025 4097 38059 4131
rect 39497 4097 39531 4131
rect 42441 4097 42475 4131
rect 44189 4097 44223 4131
rect 45845 4097 45879 4131
rect 46857 4097 46891 4131
rect 46949 4097 46983 4131
rect 13369 4029 13403 4063
rect 13645 4029 13679 4063
rect 21833 4029 21867 4063
rect 22293 4029 22327 4063
rect 48145 4029 48179 4063
rect 12725 3961 12759 3995
rect 43729 3961 43763 3995
rect 1685 3893 1719 3927
rect 2329 3893 2363 3927
rect 3157 3893 3191 3927
rect 3893 3893 3927 3927
rect 6469 3893 6503 3927
rect 7113 3893 7147 3927
rect 12081 3893 12115 3927
rect 20453 3893 20487 3927
rect 29745 3893 29779 3927
rect 30665 3893 30699 3927
rect 31401 3893 31435 3927
rect 32965 3893 32999 3927
rect 36461 3893 36495 3927
rect 38117 3893 38151 3927
rect 39589 3893 39623 3927
rect 41705 3893 41739 3927
rect 42533 3893 42567 3927
rect 44281 3893 44315 3927
rect 45385 3893 45419 3927
rect 45937 3893 45971 3927
rect 13093 3621 13127 3655
rect 1409 3553 1443 3587
rect 1593 3553 1627 3587
rect 1869 3553 1903 3587
rect 3985 3553 4019 3587
rect 4261 3553 4295 3587
rect 6193 3553 6227 3587
rect 6377 3553 6411 3587
rect 7205 3553 7239 3587
rect 20177 3553 20211 3587
rect 20361 3553 20395 3587
rect 20637 3553 20671 3587
rect 26065 3553 26099 3587
rect 26433 3553 26467 3587
rect 31585 3553 31619 3587
rect 36185 3553 36219 3587
rect 36737 3553 36771 3587
rect 41429 3553 41463 3587
rect 41889 3553 41923 3587
rect 46029 3553 46063 3587
rect 46213 3553 46247 3587
rect 46489 3553 46523 3587
rect 3801 3485 3835 3519
rect 11621 3485 11655 3519
rect 12265 3485 12299 3519
rect 13001 3485 13035 3519
rect 14657 3485 14691 3519
rect 15117 3485 15151 3519
rect 17601 3485 17635 3519
rect 18429 3485 18463 3519
rect 22753 3485 22787 3519
rect 23213 3485 23247 3519
rect 25881 3485 25915 3519
rect 29009 3485 29043 3519
rect 29561 3485 29595 3519
rect 30389 3485 30423 3519
rect 33149 3485 33183 3519
rect 36001 3485 36035 3519
rect 38945 3485 38979 3519
rect 40785 3485 40819 3519
rect 44005 3485 44039 3519
rect 45017 3485 45051 3519
rect 30573 3417 30607 3451
rect 40877 3417 40911 3451
rect 41613 3417 41647 3451
rect 11713 3349 11747 3383
rect 12357 3349 12391 3383
rect 15209 3349 15243 3383
rect 17693 3349 17727 3383
rect 23305 3349 23339 3383
rect 29653 3349 29687 3383
rect 33241 3349 33275 3383
rect 40141 3349 40175 3383
rect 45109 3349 45143 3383
rect 20177 3145 20211 3179
rect 46305 3145 46339 3179
rect 1961 3077 1995 3111
rect 6561 3077 6595 3111
rect 12173 3077 12207 3111
rect 14473 3077 14507 3111
rect 17969 3077 18003 3111
rect 23673 3077 23707 3111
rect 29929 3077 29963 3111
rect 32965 3077 32999 3111
rect 35081 3077 35115 3111
rect 35817 3077 35851 3111
rect 37933 3077 37967 3111
rect 40233 3077 40267 3111
rect 44005 3077 44039 3111
rect 4261 3009 4295 3043
rect 8677 3009 8711 3043
rect 11989 3009 12023 3043
rect 14289 3009 14323 3043
rect 17785 3009 17819 3043
rect 20085 3009 20119 3043
rect 21189 3009 21223 3043
rect 23489 3009 23523 3043
rect 26065 3009 26099 3043
rect 29745 3009 29779 3043
rect 32781 3009 32815 3043
rect 36461 3009 36495 3043
rect 37749 3009 37783 3043
rect 40049 3009 40083 3043
rect 42993 3009 43027 3043
rect 43821 3009 43855 3043
rect 46213 3009 46247 3043
rect 47869 3009 47903 3043
rect 1777 2941 1811 2975
rect 3157 2941 3191 2975
rect 5457 2941 5491 2975
rect 6377 2941 6411 2975
rect 6837 2941 6871 2975
rect 12909 2941 12943 2975
rect 15485 2941 15519 2975
rect 18245 2941 18279 2975
rect 23949 2941 23983 2975
rect 30297 2941 30331 2975
rect 33517 2941 33551 2975
rect 35449 2941 35483 2975
rect 39589 2941 39623 2975
rect 41245 2941 41279 2975
rect 44465 2941 44499 2975
rect 8861 2873 8895 2907
rect 48053 2873 48087 2907
rect 35219 2805 35253 2839
rect 35357 2805 35391 2839
rect 43085 2805 43119 2839
rect 3065 2601 3099 2635
rect 9183 2601 9217 2635
rect 20269 2601 20303 2635
rect 22845 2601 22879 2635
rect 23397 2601 23431 2635
rect 27353 2601 27387 2635
rect 1593 2533 1627 2567
rect 14749 2533 14783 2567
rect 24685 2533 24719 2567
rect 33149 2533 33183 2567
rect 33977 2533 34011 2567
rect 34897 2533 34931 2567
rect 38761 2533 38795 2567
rect 11713 2465 11747 2499
rect 11897 2465 11931 2499
rect 25513 2465 25547 2499
rect 30481 2465 30515 2499
rect 42441 2465 42475 2499
rect 42625 2465 42659 2499
rect 42901 2465 42935 2499
rect 45017 2465 45051 2499
rect 45201 2465 45235 2499
rect 45569 2465 45603 2499
rect 1409 2397 1443 2431
rect 2145 2397 2179 2431
rect 7205 2397 7239 2431
rect 7481 2397 7515 2431
rect 8953 2397 8987 2431
rect 10241 2397 10275 2431
rect 17509 2397 17543 2431
rect 17785 2397 17819 2431
rect 20085 2397 20119 2431
rect 23581 2397 23615 2431
rect 27169 2397 27203 2431
rect 32965 2397 32999 2431
rect 34161 2397 34195 2431
rect 35081 2397 35115 2431
rect 38945 2397 38979 2431
rect 4721 2329 4755 2363
rect 13553 2329 13587 2363
rect 14565 2329 14599 2363
rect 22753 2329 22787 2363
rect 24501 2329 24535 2363
rect 25329 2329 25363 2363
rect 27997 2329 28031 2363
rect 36277 2329 36311 2363
rect 47777 2329 47811 2363
rect 2329 2261 2363 2295
rect 4997 2261 5031 2295
rect 10425 2261 10459 2295
rect 28089 2261 28123 2295
rect 36369 2261 36403 2295
rect 47869 2261 47903 2295
<< metal1 >>
rect 3418 49852 3424 49904
rect 3476 49892 3482 49904
rect 8202 49892 8208 49904
rect 3476 49864 8208 49892
rect 3476 49852 3482 49864
rect 8202 49852 8208 49864
rect 8260 49852 8266 49904
rect 43990 49716 43996 49768
rect 44048 49756 44054 49768
rect 46750 49756 46756 49768
rect 44048 49728 46756 49756
rect 44048 49716 44054 49728
rect 46750 49716 46756 49728
rect 46808 49716 46814 49768
rect 1104 49530 48852 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 48852 49530
rect 1104 49456 48852 49478
rect 1302 49240 1308 49292
rect 1360 49280 1366 49292
rect 1857 49283 1915 49289
rect 1857 49280 1869 49283
rect 1360 49252 1869 49280
rect 1360 49240 1366 49252
rect 1857 49249 1869 49252
rect 1903 49249 1915 49283
rect 1857 49243 1915 49249
rect 5810 49240 5816 49292
rect 5868 49280 5874 49292
rect 8113 49283 8171 49289
rect 8113 49280 8125 49283
rect 5868 49252 8125 49280
rect 5868 49240 5874 49252
rect 8113 49249 8125 49252
rect 8159 49249 8171 49283
rect 8113 49243 8171 49249
rect 10318 49240 10324 49292
rect 10376 49280 10382 49292
rect 11977 49283 12035 49289
rect 11977 49280 11989 49283
rect 10376 49252 11989 49280
rect 10376 49240 10382 49252
rect 11977 49249 11989 49252
rect 12023 49249 12035 49283
rect 11977 49243 12035 49249
rect 12342 49240 12348 49292
rect 12400 49280 12406 49292
rect 15749 49283 15807 49289
rect 15749 49280 15761 49283
rect 12400 49252 15761 49280
rect 12400 49240 12406 49252
rect 15749 49249 15761 49252
rect 15795 49249 15807 49283
rect 15749 49243 15807 49249
rect 17865 49283 17923 49289
rect 17865 49249 17877 49283
rect 17911 49280 17923 49283
rect 18046 49280 18052 49292
rect 17911 49252 18052 49280
rect 17911 49249 17923 49252
rect 17865 49243 17923 49249
rect 18046 49240 18052 49252
rect 18104 49240 18110 49292
rect 22002 49280 22008 49292
rect 21963 49252 22008 49280
rect 22002 49240 22008 49252
rect 22060 49240 22066 49292
rect 24210 49240 24216 49292
rect 24268 49280 24274 49292
rect 24397 49283 24455 49289
rect 24397 49280 24409 49283
rect 24268 49252 24409 49280
rect 24268 49240 24274 49252
rect 24397 49249 24409 49252
rect 24443 49249 24455 49283
rect 27614 49280 27620 49292
rect 27575 49252 27620 49280
rect 24397 49243 24455 49249
rect 27614 49240 27620 49252
rect 27672 49240 27678 49292
rect 43162 49280 43168 49292
rect 43123 49252 43168 49280
rect 43162 49240 43168 49252
rect 43220 49240 43226 49292
rect 47029 49283 47087 49289
rect 47029 49249 47041 49283
rect 47075 49280 47087 49283
rect 48314 49280 48320 49292
rect 47075 49252 48320 49280
rect 47075 49249 47087 49252
rect 47029 49243 47087 49249
rect 48314 49240 48320 49252
rect 48372 49240 48378 49292
rect 1397 49215 1455 49221
rect 1397 49181 1409 49215
rect 1443 49181 1455 49215
rect 1397 49175 1455 49181
rect 1412 49076 1440 49175
rect 3602 49172 3608 49224
rect 3660 49212 3666 49224
rect 4249 49215 4307 49221
rect 4249 49212 4261 49215
rect 3660 49184 4261 49212
rect 3660 49172 3666 49184
rect 4249 49181 4261 49184
rect 4295 49181 4307 49215
rect 6546 49212 6552 49224
rect 6507 49184 6552 49212
rect 4249 49175 4307 49181
rect 6546 49172 6552 49184
rect 6604 49172 6610 49224
rect 7466 49212 7472 49224
rect 7427 49184 7472 49212
rect 7466 49172 7472 49184
rect 7524 49172 7530 49224
rect 10965 49215 11023 49221
rect 10965 49181 10977 49215
rect 11011 49212 11023 49215
rect 11517 49215 11575 49221
rect 11517 49212 11529 49215
rect 11011 49184 11529 49212
rect 11011 49181 11023 49184
rect 10965 49175 11023 49181
rect 11517 49181 11529 49184
rect 11563 49181 11575 49215
rect 11517 49175 11575 49181
rect 14182 49172 14188 49224
rect 14240 49212 14246 49224
rect 14921 49215 14979 49221
rect 14921 49212 14933 49215
rect 14240 49184 14933 49212
rect 14240 49172 14246 49184
rect 14921 49181 14933 49184
rect 14967 49181 14979 49215
rect 14921 49175 14979 49181
rect 16574 49172 16580 49224
rect 16632 49212 16638 49224
rect 17129 49215 17187 49221
rect 17129 49212 17141 49215
rect 16632 49184 17141 49212
rect 16632 49172 16638 49184
rect 17129 49181 17141 49184
rect 17175 49181 17187 49215
rect 17129 49175 17187 49181
rect 18141 49215 18199 49221
rect 18141 49181 18153 49215
rect 18187 49181 18199 49215
rect 19334 49212 19340 49224
rect 19295 49184 19340 49212
rect 18141 49175 18199 49181
rect 1581 49147 1639 49153
rect 1581 49113 1593 49147
rect 1627 49144 1639 49147
rect 2590 49144 2596 49156
rect 1627 49116 2596 49144
rect 1627 49113 1639 49116
rect 1581 49107 1639 49113
rect 2590 49104 2596 49116
rect 2648 49104 2654 49156
rect 4614 49144 4620 49156
rect 4575 49116 4620 49144
rect 4614 49104 4620 49116
rect 4672 49104 4678 49156
rect 5166 49144 5172 49156
rect 5127 49116 5172 49144
rect 5166 49104 5172 49116
rect 5224 49104 5230 49156
rect 11698 49144 11704 49156
rect 11659 49116 11704 49144
rect 11698 49104 11704 49116
rect 11756 49104 11762 49156
rect 18156 49144 18184 49175
rect 19334 49172 19340 49184
rect 19392 49172 19398 49224
rect 20162 49212 20168 49224
rect 20123 49184 20168 49212
rect 20162 49172 20168 49184
rect 20220 49172 20226 49224
rect 22278 49212 22284 49224
rect 22239 49184 22284 49212
rect 22278 49172 22284 49184
rect 22336 49172 22342 49224
rect 23842 49212 23848 49224
rect 23803 49184 23848 49212
rect 23842 49172 23848 49184
rect 23900 49172 23906 49224
rect 24670 49212 24676 49224
rect 24631 49184 24676 49212
rect 24670 49172 24676 49184
rect 24728 49172 24734 49224
rect 26418 49212 26424 49224
rect 26379 49184 26424 49212
rect 26418 49172 26424 49184
rect 26476 49172 26482 49224
rect 26970 49212 26976 49224
rect 26931 49184 26976 49212
rect 26970 49172 26976 49184
rect 27028 49172 27034 49224
rect 28994 49172 29000 49224
rect 29052 49212 29058 49224
rect 30009 49215 30067 49221
rect 30009 49212 30021 49215
rect 29052 49184 30021 49212
rect 29052 49172 29058 49184
rect 30009 49181 30021 49184
rect 30055 49181 30067 49215
rect 30009 49175 30067 49181
rect 31021 49215 31079 49221
rect 31021 49181 31033 49215
rect 31067 49181 31079 49215
rect 31021 49175 31079 49181
rect 24486 49144 24492 49156
rect 18156 49116 24492 49144
rect 24486 49104 24492 49116
rect 24544 49104 24550 49156
rect 27154 49144 27160 49156
rect 27115 49116 27160 49144
rect 27154 49104 27160 49116
rect 27212 49104 27218 49156
rect 29730 49104 29736 49156
rect 29788 49144 29794 49156
rect 31036 49144 31064 49175
rect 33502 49172 33508 49224
rect 33560 49212 33566 49224
rect 33781 49215 33839 49221
rect 33781 49212 33793 49215
rect 33560 49184 33793 49212
rect 33560 49172 33566 49184
rect 33781 49181 33793 49184
rect 33827 49181 33839 49215
rect 33781 49175 33839 49181
rect 34882 49172 34888 49224
rect 34940 49212 34946 49224
rect 35621 49215 35679 49221
rect 35621 49212 35633 49215
rect 34940 49184 35633 49212
rect 34940 49172 34946 49184
rect 35621 49181 35633 49184
rect 35667 49181 35679 49215
rect 36262 49212 36268 49224
rect 36223 49184 36268 49212
rect 35621 49175 35679 49181
rect 36262 49172 36268 49184
rect 36320 49172 36326 49224
rect 38102 49212 38108 49224
rect 38063 49184 38108 49212
rect 38102 49172 38108 49184
rect 38160 49172 38166 49224
rect 40770 49212 40776 49224
rect 40731 49184 40776 49212
rect 40770 49172 40776 49184
rect 40828 49172 40834 49224
rect 41598 49212 41604 49224
rect 41559 49184 41604 49212
rect 41598 49172 41604 49184
rect 41656 49172 41662 49224
rect 42426 49212 42432 49224
rect 42387 49184 42432 49212
rect 42426 49172 42432 49184
rect 42484 49172 42490 49224
rect 45189 49215 45247 49221
rect 45189 49181 45201 49215
rect 45235 49181 45247 49215
rect 47762 49212 47768 49224
rect 47723 49184 47768 49212
rect 45189 49175 45247 49181
rect 29788 49116 31064 49144
rect 29788 49104 29794 49116
rect 41414 49104 41420 49156
rect 41472 49144 41478 49156
rect 42613 49147 42671 49153
rect 42613 49144 42625 49147
rect 41472 49116 42625 49144
rect 41472 49104 41478 49116
rect 42613 49113 42625 49116
rect 42659 49113 42671 49147
rect 42613 49107 42671 49113
rect 3970 49076 3976 49088
rect 1412 49048 3976 49076
rect 3970 49036 3976 49048
rect 4028 49036 4034 49088
rect 5258 49076 5264 49088
rect 5219 49048 5264 49076
rect 5258 49036 5264 49048
rect 5316 49036 5322 49088
rect 6730 49076 6736 49088
rect 6691 49048 6736 49076
rect 6730 49036 6736 49048
rect 6788 49036 6794 49088
rect 10134 49076 10140 49088
rect 10095 49048 10140 49076
rect 10134 49036 10140 49048
rect 10192 49036 10198 49088
rect 15010 49076 15016 49088
rect 14971 49048 15016 49076
rect 15010 49036 15016 49048
rect 15068 49036 15074 49088
rect 17218 49076 17224 49088
rect 17179 49048 17224 49076
rect 17218 49036 17224 49048
rect 17276 49036 17282 49088
rect 19521 49079 19579 49085
rect 19521 49045 19533 49079
rect 19567 49076 19579 49079
rect 20070 49076 20076 49088
rect 19567 49048 20076 49076
rect 19567 49045 19579 49048
rect 19521 49039 19579 49045
rect 20070 49036 20076 49048
rect 20128 49036 20134 49088
rect 20254 49076 20260 49088
rect 20215 49048 20260 49076
rect 20254 49036 20260 49048
rect 20312 49036 20318 49088
rect 29270 49036 29276 49088
rect 29328 49076 29334 49088
rect 30101 49079 30159 49085
rect 30101 49076 30113 49079
rect 29328 49048 30113 49076
rect 29328 49036 29334 49048
rect 30101 49045 30113 49048
rect 30147 49045 30159 49079
rect 32122 49076 32128 49088
rect 32083 49048 32128 49076
rect 30101 49039 30159 49045
rect 32122 49036 32128 49048
rect 32180 49036 32186 49088
rect 38286 49076 38292 49088
rect 38247 49048 38292 49076
rect 38286 49036 38292 49048
rect 38344 49036 38350 49088
rect 40862 49076 40868 49088
rect 40823 49048 40868 49076
rect 40862 49036 40868 49048
rect 40920 49036 40926 49088
rect 41598 49036 41604 49088
rect 41656 49076 41662 49088
rect 41785 49079 41843 49085
rect 41785 49076 41797 49079
rect 41656 49048 41797 49076
rect 41656 49036 41662 49048
rect 41785 49045 41797 49048
rect 41831 49045 41843 49079
rect 45204 49076 45232 49175
rect 47762 49172 47768 49184
rect 47820 49172 47826 49224
rect 45373 49147 45431 49153
rect 45373 49113 45385 49147
rect 45419 49144 45431 49147
rect 45738 49144 45744 49156
rect 45419 49116 45744 49144
rect 45419 49113 45431 49116
rect 45373 49107 45431 49113
rect 45738 49104 45744 49116
rect 45796 49104 45802 49156
rect 45278 49076 45284 49088
rect 45204 49048 45284 49076
rect 41785 49039 41843 49045
rect 45278 49036 45284 49048
rect 45336 49036 45342 49088
rect 47118 49036 47124 49088
rect 47176 49076 47182 49088
rect 47857 49079 47915 49085
rect 47857 49076 47869 49079
rect 47176 49048 47869 49076
rect 47176 49036 47182 49048
rect 47857 49045 47869 49048
rect 47903 49045 47915 49079
rect 47857 49039 47915 49045
rect 1104 48986 48852 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 48852 48986
rect 1104 48912 48852 48934
rect 24670 48832 24676 48884
rect 24728 48872 24734 48884
rect 30006 48872 30012 48884
rect 24728 48844 30012 48872
rect 24728 48832 24734 48844
rect 30006 48832 30012 48844
rect 30064 48832 30070 48884
rect 46290 48872 46296 48884
rect 43272 48844 46296 48872
rect 14 48764 20 48816
rect 72 48804 78 48816
rect 72 48776 2360 48804
rect 72 48764 78 48776
rect 658 48696 664 48748
rect 716 48736 722 48748
rect 2332 48745 2360 48776
rect 3878 48764 3884 48816
rect 3936 48804 3942 48816
rect 3936 48776 4844 48804
rect 3936 48764 3942 48776
rect 1397 48739 1455 48745
rect 1397 48736 1409 48739
rect 716 48708 1409 48736
rect 716 48696 722 48708
rect 1397 48705 1409 48708
rect 1443 48705 1455 48739
rect 1397 48699 1455 48705
rect 2317 48739 2375 48745
rect 2317 48705 2329 48739
rect 2363 48705 2375 48739
rect 2317 48699 2375 48705
rect 1486 48628 1492 48680
rect 1544 48668 1550 48680
rect 1581 48671 1639 48677
rect 1581 48668 1593 48671
rect 1544 48640 1593 48668
rect 1544 48628 1550 48640
rect 1581 48637 1593 48640
rect 1627 48637 1639 48671
rect 3142 48668 3148 48680
rect 3103 48640 3148 48668
rect 1581 48631 1639 48637
rect 3142 48628 3148 48640
rect 3200 48628 3206 48680
rect 3329 48671 3387 48677
rect 3329 48637 3341 48671
rect 3375 48668 3387 48671
rect 4062 48668 4068 48680
rect 3375 48640 4068 48668
rect 3375 48637 3387 48640
rect 3329 48631 3387 48637
rect 4062 48628 4068 48640
rect 4120 48628 4126 48680
rect 4154 48628 4160 48680
rect 4212 48668 4218 48680
rect 4816 48668 4844 48776
rect 4890 48764 4896 48816
rect 4948 48804 4954 48816
rect 5537 48807 5595 48813
rect 5537 48804 5549 48807
rect 4948 48776 5549 48804
rect 4948 48764 4954 48776
rect 5537 48773 5549 48776
rect 5583 48773 5595 48807
rect 7466 48804 7472 48816
rect 5537 48767 5595 48773
rect 6748 48776 7472 48804
rect 6748 48745 6776 48776
rect 7466 48764 7472 48776
rect 7524 48764 7530 48816
rect 8202 48764 8208 48816
rect 8260 48804 8266 48816
rect 8260 48776 10548 48804
rect 8260 48764 8266 48776
rect 6733 48739 6791 48745
rect 6733 48705 6745 48739
rect 6779 48705 6791 48739
rect 6733 48699 6791 48705
rect 5534 48668 5540 48680
rect 4212 48640 4257 48668
rect 4816 48640 5540 48668
rect 4212 48628 4218 48640
rect 5534 48628 5540 48640
rect 5592 48628 5598 48680
rect 6914 48628 6920 48680
rect 6972 48668 6978 48680
rect 7190 48668 7196 48680
rect 6972 48640 7017 48668
rect 7151 48640 7196 48668
rect 6972 48628 6978 48640
rect 7190 48628 7196 48640
rect 7248 48628 7254 48680
rect 9122 48668 9128 48680
rect 9083 48640 9128 48668
rect 9122 48628 9128 48640
rect 9180 48628 9186 48680
rect 9309 48671 9367 48677
rect 9309 48637 9321 48671
rect 9355 48668 9367 48671
rect 10226 48668 10232 48680
rect 9355 48640 10232 48668
rect 9355 48637 9367 48640
rect 9309 48631 9367 48637
rect 10226 48628 10232 48640
rect 10284 48628 10290 48680
rect 10520 48677 10548 48776
rect 13814 48764 13820 48816
rect 13872 48804 13878 48816
rect 14737 48807 14795 48813
rect 14737 48804 14749 48807
rect 13872 48776 14749 48804
rect 13872 48764 13878 48776
rect 14737 48773 14749 48776
rect 14783 48773 14795 48807
rect 19426 48804 19432 48816
rect 14737 48767 14795 48773
rect 19260 48776 19432 48804
rect 11606 48736 11612 48748
rect 11567 48708 11612 48736
rect 11606 48696 11612 48708
rect 11664 48696 11670 48748
rect 12342 48736 12348 48748
rect 12303 48708 12348 48736
rect 12342 48696 12348 48708
rect 12400 48696 12406 48748
rect 19260 48745 19288 48776
rect 19426 48764 19432 48776
rect 19484 48764 19490 48816
rect 31573 48807 31631 48813
rect 31573 48773 31585 48807
rect 31619 48804 31631 48807
rect 31938 48804 31944 48816
rect 31619 48776 31944 48804
rect 31619 48773 31631 48776
rect 31573 48767 31631 48773
rect 31938 48764 31944 48776
rect 31996 48764 32002 48816
rect 19245 48739 19303 48745
rect 19245 48705 19257 48739
rect 19291 48705 19303 48739
rect 19245 48699 19303 48705
rect 25406 48696 25412 48748
rect 25464 48736 25470 48748
rect 25961 48739 26019 48745
rect 25961 48736 25973 48739
rect 25464 48708 25973 48736
rect 25464 48696 25470 48708
rect 25961 48705 25973 48708
rect 26007 48705 26019 48739
rect 25961 48699 26019 48705
rect 26418 48696 26424 48748
rect 26476 48736 26482 48748
rect 27433 48739 27491 48745
rect 27433 48736 27445 48739
rect 26476 48708 27445 48736
rect 26476 48696 26482 48708
rect 27433 48705 27445 48708
rect 27479 48705 27491 48739
rect 29730 48736 29736 48748
rect 29691 48708 29736 48736
rect 27433 48699 27491 48705
rect 29730 48696 29736 48708
rect 29788 48696 29794 48748
rect 32122 48736 32128 48748
rect 32083 48708 32128 48736
rect 32122 48696 32128 48708
rect 32180 48696 32186 48748
rect 34882 48736 34888 48748
rect 34843 48708 34888 48736
rect 34882 48696 34888 48708
rect 34940 48696 34946 48748
rect 42334 48696 42340 48748
rect 42392 48736 42398 48748
rect 43272 48745 43300 48844
rect 46290 48832 46296 48844
rect 46348 48832 46354 48884
rect 44450 48804 44456 48816
rect 43732 48776 44456 48804
rect 43732 48745 43760 48776
rect 44450 48764 44456 48776
rect 44508 48764 44514 48816
rect 47949 48807 48007 48813
rect 47949 48773 47961 48807
rect 47995 48804 48007 48807
rect 48958 48804 48964 48816
rect 47995 48776 48964 48804
rect 47995 48773 48007 48776
rect 47949 48767 48007 48773
rect 48958 48764 48964 48776
rect 49016 48764 49022 48816
rect 42429 48739 42487 48745
rect 42429 48736 42441 48739
rect 42392 48708 42441 48736
rect 42392 48696 42398 48708
rect 42429 48705 42441 48708
rect 42475 48705 42487 48739
rect 42429 48699 42487 48705
rect 43257 48739 43315 48745
rect 43257 48705 43269 48739
rect 43303 48705 43315 48739
rect 43257 48699 43315 48705
rect 43717 48739 43775 48745
rect 43717 48705 43729 48739
rect 43763 48705 43775 48739
rect 46750 48736 46756 48748
rect 46711 48708 46756 48736
rect 43717 48699 43775 48705
rect 46750 48696 46756 48708
rect 46808 48696 46814 48748
rect 10505 48671 10563 48677
rect 10505 48637 10517 48671
rect 10551 48637 10563 48671
rect 12526 48668 12532 48680
rect 12487 48640 12532 48668
rect 10505 48631 10563 48637
rect 12526 48628 12532 48640
rect 12584 48628 12590 48680
rect 12618 48628 12624 48680
rect 12676 48668 12682 48680
rect 12805 48671 12863 48677
rect 12805 48668 12817 48671
rect 12676 48640 12817 48668
rect 12676 48628 12682 48640
rect 12805 48637 12817 48640
rect 12851 48637 12863 48671
rect 12805 48631 12863 48637
rect 16117 48671 16175 48677
rect 16117 48637 16129 48671
rect 16163 48668 16175 48671
rect 16669 48671 16727 48677
rect 16669 48668 16681 48671
rect 16163 48640 16681 48668
rect 16163 48637 16175 48640
rect 16117 48631 16175 48637
rect 16669 48637 16681 48640
rect 16715 48637 16727 48671
rect 16850 48668 16856 48680
rect 16811 48640 16856 48668
rect 16669 48631 16727 48637
rect 16850 48628 16856 48640
rect 16908 48628 16914 48680
rect 16942 48628 16948 48680
rect 17000 48668 17006 48680
rect 17129 48671 17187 48677
rect 17129 48668 17141 48671
rect 17000 48640 17141 48668
rect 17000 48628 17006 48640
rect 17129 48637 17141 48640
rect 17175 48637 17187 48671
rect 17129 48631 17187 48637
rect 19429 48671 19487 48677
rect 19429 48637 19441 48671
rect 19475 48668 19487 48671
rect 19518 48668 19524 48680
rect 19475 48640 19524 48668
rect 19475 48637 19487 48640
rect 19429 48631 19487 48637
rect 19518 48628 19524 48640
rect 19576 48628 19582 48680
rect 20622 48628 20628 48680
rect 20680 48668 20686 48680
rect 20717 48671 20775 48677
rect 20717 48668 20729 48671
rect 20680 48640 20729 48668
rect 20680 48628 20686 48640
rect 20717 48637 20729 48640
rect 20763 48637 20775 48671
rect 20717 48631 20775 48637
rect 22097 48671 22155 48677
rect 22097 48637 22109 48671
rect 22143 48668 22155 48671
rect 22557 48671 22615 48677
rect 22557 48668 22569 48671
rect 22143 48640 22569 48668
rect 22143 48637 22155 48640
rect 22097 48631 22155 48637
rect 22557 48637 22569 48640
rect 22603 48637 22615 48671
rect 22738 48668 22744 48680
rect 22699 48640 22744 48668
rect 22557 48631 22615 48637
rect 22738 48628 22744 48640
rect 22796 48628 22802 48680
rect 23474 48668 23480 48680
rect 23435 48640 23480 48668
rect 23474 48628 23480 48640
rect 23532 48628 23538 48680
rect 25501 48671 25559 48677
rect 25501 48637 25513 48671
rect 25547 48668 25559 48671
rect 26510 48668 26516 48680
rect 25547 48640 26516 48668
rect 25547 48637 25559 48640
rect 25501 48631 25559 48637
rect 26510 48628 26516 48640
rect 26568 48628 26574 48680
rect 27614 48668 27620 48680
rect 27575 48640 27620 48668
rect 27614 48628 27620 48640
rect 27672 48628 27678 48680
rect 27890 48668 27896 48680
rect 27851 48640 27896 48668
rect 27890 48628 27896 48640
rect 27948 48628 27954 48680
rect 29917 48671 29975 48677
rect 29917 48637 29929 48671
rect 29963 48668 29975 48671
rect 30558 48668 30564 48680
rect 29963 48640 30564 48668
rect 29963 48637 29975 48640
rect 29917 48631 29975 48637
rect 30558 48628 30564 48640
rect 30616 48628 30622 48680
rect 32306 48668 32312 48680
rect 32267 48640 32312 48668
rect 32306 48628 32312 48640
rect 32364 48628 32370 48680
rect 32858 48668 32864 48680
rect 32819 48640 32864 48668
rect 32858 48628 32864 48640
rect 32916 48628 32922 48680
rect 35069 48671 35127 48677
rect 35069 48637 35081 48671
rect 35115 48668 35127 48671
rect 36078 48668 36084 48680
rect 35115 48640 35894 48668
rect 36039 48640 36084 48668
rect 35115 48637 35127 48640
rect 35069 48631 35127 48637
rect 2501 48603 2559 48609
rect 2501 48569 2513 48603
rect 2547 48600 2559 48603
rect 30742 48600 30748 48612
rect 2547 48572 30748 48600
rect 2547 48569 2559 48572
rect 2501 48563 2559 48569
rect 30742 48560 30748 48572
rect 30800 48560 30806 48612
rect 5626 48532 5632 48544
rect 5587 48504 5632 48532
rect 5626 48492 5632 48504
rect 5684 48492 5690 48544
rect 11790 48532 11796 48544
rect 11751 48504 11796 48532
rect 11790 48492 11796 48504
rect 11848 48492 11854 48544
rect 14826 48532 14832 48544
rect 14787 48504 14832 48532
rect 14826 48492 14832 48504
rect 14884 48492 14890 48544
rect 26145 48535 26203 48541
rect 26145 48501 26157 48535
rect 26191 48532 26203 48535
rect 27522 48532 27528 48544
rect 26191 48504 27528 48532
rect 26191 48501 26203 48504
rect 26145 48495 26203 48501
rect 27522 48492 27528 48504
rect 27580 48492 27586 48544
rect 35866 48532 35894 48640
rect 36078 48628 36084 48640
rect 36136 48628 36142 48680
rect 38841 48671 38899 48677
rect 38841 48637 38853 48671
rect 38887 48668 38899 48671
rect 39301 48671 39359 48677
rect 39301 48668 39313 48671
rect 38887 48640 39313 48668
rect 38887 48637 38899 48640
rect 38841 48631 38899 48637
rect 39301 48637 39313 48640
rect 39347 48637 39359 48671
rect 39482 48668 39488 48680
rect 39443 48640 39488 48668
rect 39301 48631 39359 48637
rect 39482 48628 39488 48640
rect 39540 48628 39546 48680
rect 40034 48668 40040 48680
rect 39995 48640 40040 48668
rect 40034 48628 40040 48640
rect 40092 48628 40098 48680
rect 44450 48668 44456 48680
rect 44411 48640 44456 48668
rect 44450 48628 44456 48640
rect 44508 48628 44514 48680
rect 44634 48668 44640 48680
rect 44595 48640 44640 48668
rect 44634 48628 44640 48640
rect 44692 48628 44698 48680
rect 45830 48668 45836 48680
rect 45791 48640 45836 48668
rect 45830 48628 45836 48640
rect 45888 48628 45894 48680
rect 35986 48532 35992 48544
rect 35866 48504 35992 48532
rect 35986 48492 35992 48504
rect 36044 48492 36050 48544
rect 37642 48492 37648 48544
rect 37700 48532 37706 48544
rect 38562 48532 38568 48544
rect 37700 48504 38568 48532
rect 37700 48492 37706 48504
rect 38562 48492 38568 48504
rect 38620 48492 38626 48544
rect 41782 48492 41788 48544
rect 41840 48532 41846 48544
rect 41877 48535 41935 48541
rect 41877 48532 41889 48535
rect 41840 48504 41889 48532
rect 41840 48492 41846 48504
rect 41877 48501 41889 48504
rect 41923 48501 41935 48535
rect 41877 48495 41935 48501
rect 42521 48535 42579 48541
rect 42521 48501 42533 48535
rect 42567 48532 42579 48535
rect 42794 48532 42800 48544
rect 42567 48504 42800 48532
rect 42567 48501 42579 48504
rect 42521 48495 42579 48501
rect 42794 48492 42800 48504
rect 42852 48492 42858 48544
rect 43898 48532 43904 48544
rect 43859 48504 43904 48532
rect 43898 48492 43904 48504
rect 43956 48492 43962 48544
rect 46934 48532 46940 48544
rect 46895 48504 46940 48532
rect 46934 48492 46940 48504
rect 46992 48492 46998 48544
rect 47210 48492 47216 48544
rect 47268 48532 47274 48544
rect 48041 48535 48099 48541
rect 48041 48532 48053 48535
rect 47268 48504 48053 48532
rect 47268 48492 47274 48504
rect 48041 48501 48053 48504
rect 48087 48501 48099 48535
rect 48041 48495 48099 48501
rect 1104 48442 48852 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 48852 48442
rect 1104 48368 48852 48390
rect 3142 48288 3148 48340
rect 3200 48328 3206 48340
rect 3973 48331 4031 48337
rect 3973 48328 3985 48331
rect 3200 48300 3985 48328
rect 3200 48288 3206 48300
rect 3973 48297 3985 48300
rect 4019 48297 4031 48331
rect 3973 48291 4031 48297
rect 6914 48288 6920 48340
rect 6972 48328 6978 48340
rect 7101 48331 7159 48337
rect 7101 48328 7113 48331
rect 6972 48300 7113 48328
rect 6972 48288 6978 48300
rect 7101 48297 7113 48300
rect 7147 48297 7159 48331
rect 7101 48291 7159 48297
rect 9122 48288 9128 48340
rect 9180 48328 9186 48340
rect 9309 48331 9367 48337
rect 9309 48328 9321 48331
rect 9180 48300 9321 48328
rect 9180 48288 9186 48300
rect 9309 48297 9321 48300
rect 9355 48297 9367 48331
rect 16850 48328 16856 48340
rect 16811 48300 16856 48328
rect 9309 48291 9367 48297
rect 16850 48288 16856 48300
rect 16908 48288 16914 48340
rect 39482 48288 39488 48340
rect 39540 48328 39546 48340
rect 39945 48331 40003 48337
rect 39945 48328 39957 48331
rect 39540 48300 39957 48328
rect 39540 48288 39546 48300
rect 39945 48297 39957 48300
rect 39991 48297 40003 48331
rect 39945 48291 40003 48297
rect 44634 48288 44640 48340
rect 44692 48328 44698 48340
rect 45097 48331 45155 48337
rect 45097 48328 45109 48331
rect 44692 48300 45109 48328
rect 44692 48288 44698 48300
rect 45097 48297 45109 48300
rect 45143 48297 45155 48331
rect 45097 48291 45155 48297
rect 1946 48220 1952 48272
rect 2004 48260 2010 48272
rect 5166 48260 5172 48272
rect 2004 48232 5172 48260
rect 2004 48220 2010 48232
rect 5166 48220 5172 48232
rect 5224 48220 5230 48272
rect 9674 48220 9680 48272
rect 9732 48260 9738 48272
rect 9732 48232 10640 48260
rect 9732 48220 9738 48232
rect 2774 48192 2780 48204
rect 2735 48164 2780 48192
rect 2774 48152 2780 48164
rect 2832 48152 2838 48204
rect 4709 48195 4767 48201
rect 4709 48161 4721 48195
rect 4755 48192 4767 48195
rect 5810 48192 5816 48204
rect 4755 48164 5816 48192
rect 4755 48161 4767 48164
rect 4709 48155 4767 48161
rect 5810 48152 5816 48164
rect 5868 48152 5874 48204
rect 10134 48192 10140 48204
rect 10095 48164 10140 48192
rect 10134 48152 10140 48164
rect 10192 48152 10198 48204
rect 10612 48201 10640 48232
rect 11698 48220 11704 48272
rect 11756 48260 11762 48272
rect 19426 48260 19432 48272
rect 11756 48232 16574 48260
rect 19387 48232 19432 48260
rect 11756 48220 11762 48232
rect 10597 48195 10655 48201
rect 10597 48161 10609 48195
rect 10643 48161 10655 48195
rect 14918 48192 14924 48204
rect 14879 48164 14924 48192
rect 10597 48155 10655 48161
rect 14918 48152 14924 48164
rect 14976 48152 14982 48204
rect 1394 48124 1400 48136
rect 1355 48096 1400 48124
rect 1394 48084 1400 48096
rect 1452 48084 1458 48136
rect 7006 48124 7012 48136
rect 6967 48096 7012 48124
rect 7006 48084 7012 48096
rect 7064 48084 7070 48136
rect 7374 48084 7380 48136
rect 7432 48124 7438 48136
rect 7837 48127 7895 48133
rect 7837 48124 7849 48127
rect 7432 48096 7849 48124
rect 7432 48084 7438 48096
rect 7837 48093 7849 48096
rect 7883 48093 7895 48127
rect 13078 48124 13084 48136
rect 13039 48096 13084 48124
rect 7837 48087 7895 48093
rect 13078 48084 13084 48096
rect 13136 48084 13142 48136
rect 14458 48124 14464 48136
rect 14419 48096 14464 48124
rect 14458 48084 14464 48096
rect 14516 48084 14522 48136
rect 1578 48056 1584 48068
rect 1539 48028 1584 48056
rect 1578 48016 1584 48028
rect 1636 48016 1642 48068
rect 4893 48059 4951 48065
rect 4893 48025 4905 48059
rect 4939 48056 4951 48059
rect 6178 48056 6184 48068
rect 4939 48028 6184 48056
rect 4939 48025 4951 48028
rect 4893 48019 4951 48025
rect 6178 48016 6184 48028
rect 6236 48016 6242 48068
rect 6549 48059 6607 48065
rect 6549 48025 6561 48059
rect 6595 48025 6607 48059
rect 6549 48019 6607 48025
rect 10321 48059 10379 48065
rect 10321 48025 10333 48059
rect 10367 48056 10379 48059
rect 10870 48056 10876 48068
rect 10367 48028 10876 48056
rect 10367 48025 10379 48028
rect 10321 48019 10379 48025
rect 3786 47948 3792 48000
rect 3844 47988 3850 48000
rect 6564 47988 6592 48019
rect 10870 48016 10876 48028
rect 10928 48016 10934 48068
rect 14366 48016 14372 48068
rect 14424 48056 14430 48068
rect 14645 48059 14703 48065
rect 14645 48056 14657 48059
rect 14424 48028 14657 48056
rect 14424 48016 14430 48028
rect 14645 48025 14657 48028
rect 14691 48025 14703 48059
rect 14645 48019 14703 48025
rect 3844 47960 6592 47988
rect 3844 47948 3850 47960
rect 6638 47948 6644 48000
rect 6696 47988 6702 48000
rect 10502 47988 10508 48000
rect 6696 47960 10508 47988
rect 6696 47948 6702 47960
rect 10502 47948 10508 47960
rect 10560 47948 10566 48000
rect 13173 47991 13231 47997
rect 13173 47957 13185 47991
rect 13219 47988 13231 47991
rect 14918 47988 14924 48000
rect 13219 47960 14924 47988
rect 13219 47957 13231 47960
rect 13173 47951 13231 47957
rect 14918 47948 14924 47960
rect 14976 47948 14982 48000
rect 16546 47988 16574 48232
rect 19426 48220 19432 48232
rect 19484 48220 19490 48272
rect 19978 48220 19984 48272
rect 20036 48260 20042 48272
rect 20036 48232 36860 48260
rect 20036 48220 20042 48232
rect 17586 48192 17592 48204
rect 16776 48164 17592 48192
rect 16776 48133 16804 48164
rect 17586 48152 17592 48164
rect 17644 48192 17650 48204
rect 22094 48192 22100 48204
rect 17644 48164 22100 48192
rect 17644 48152 17650 48164
rect 22094 48152 22100 48164
rect 22152 48152 22158 48204
rect 22554 48192 22560 48204
rect 22515 48164 22560 48192
rect 22554 48152 22560 48164
rect 22612 48152 22618 48204
rect 23842 48152 23848 48204
rect 23900 48192 23906 48204
rect 24397 48195 24455 48201
rect 24397 48192 24409 48195
rect 23900 48164 24409 48192
rect 23900 48152 23906 48164
rect 24397 48161 24409 48164
rect 24443 48161 24455 48195
rect 24397 48155 24455 48161
rect 24578 48152 24584 48204
rect 24636 48192 24642 48204
rect 24857 48195 24915 48201
rect 24857 48192 24869 48195
rect 24636 48164 24869 48192
rect 24636 48152 24642 48164
rect 24857 48161 24869 48164
rect 24903 48161 24915 48195
rect 28074 48192 28080 48204
rect 24857 48155 24915 48161
rect 26206 48164 28080 48192
rect 16761 48127 16819 48133
rect 16761 48093 16773 48127
rect 16807 48093 16819 48127
rect 16761 48087 16819 48093
rect 21361 48127 21419 48133
rect 21361 48093 21373 48127
rect 21407 48124 21419 48127
rect 21821 48127 21879 48133
rect 21821 48124 21833 48127
rect 21407 48096 21833 48124
rect 21407 48093 21419 48096
rect 21361 48087 21419 48093
rect 21821 48093 21833 48096
rect 21867 48093 21879 48127
rect 24302 48124 24308 48136
rect 21821 48087 21879 48093
rect 23216 48096 24308 48124
rect 22002 48056 22008 48068
rect 21963 48028 22008 48056
rect 22002 48016 22008 48028
rect 22060 48016 22066 48068
rect 22094 48016 22100 48068
rect 22152 48056 22158 48068
rect 23216 48056 23244 48096
rect 24302 48084 24308 48096
rect 24360 48084 24366 48136
rect 22152 48028 23244 48056
rect 22152 48016 22158 48028
rect 24210 48016 24216 48068
rect 24268 48056 24274 48068
rect 24581 48059 24639 48065
rect 24581 48056 24593 48059
rect 24268 48028 24593 48056
rect 24268 48016 24274 48028
rect 24581 48025 24593 48028
rect 24627 48025 24639 48059
rect 24581 48019 24639 48025
rect 24670 48016 24676 48068
rect 24728 48056 24734 48068
rect 26206 48056 26234 48164
rect 28074 48152 28080 48164
rect 28132 48152 28138 48204
rect 28350 48192 28356 48204
rect 28311 48164 28356 48192
rect 28350 48152 28356 48164
rect 28408 48152 28414 48204
rect 29549 48195 29607 48201
rect 29549 48161 29561 48195
rect 29595 48192 29607 48195
rect 29822 48192 29828 48204
rect 29595 48164 29828 48192
rect 29595 48161 29607 48164
rect 29549 48155 29607 48161
rect 26510 48084 26516 48136
rect 26568 48124 26574 48136
rect 27145 48127 27203 48133
rect 27145 48124 27157 48127
rect 26568 48096 27157 48124
rect 26568 48084 26574 48096
rect 27145 48093 27157 48096
rect 27191 48093 27203 48127
rect 27145 48087 27203 48093
rect 24728 48028 26234 48056
rect 27341 48059 27399 48065
rect 24728 48016 24734 48028
rect 27341 48025 27353 48059
rect 27387 48056 27399 48059
rect 27890 48056 27896 48068
rect 27387 48028 27896 48056
rect 27387 48025 27399 48028
rect 27341 48019 27399 48025
rect 27890 48016 27896 48028
rect 27948 48016 27954 48068
rect 28166 48016 28172 48068
rect 28224 48056 28230 48068
rect 29564 48056 29592 48155
rect 29822 48152 29828 48164
rect 29880 48152 29886 48204
rect 29914 48152 29920 48204
rect 29972 48192 29978 48204
rect 30009 48195 30067 48201
rect 30009 48192 30021 48195
rect 29972 48164 30021 48192
rect 29972 48152 29978 48164
rect 30009 48161 30021 48164
rect 30055 48161 30067 48195
rect 30009 48155 30067 48161
rect 30926 48152 30932 48204
rect 30984 48192 30990 48204
rect 32309 48195 32367 48201
rect 32309 48192 32321 48195
rect 30984 48164 32321 48192
rect 30984 48152 30990 48164
rect 32309 48161 32321 48164
rect 32355 48161 32367 48195
rect 32309 48155 32367 48161
rect 35989 48195 36047 48201
rect 35989 48161 36001 48195
rect 36035 48192 36047 48195
rect 36262 48192 36268 48204
rect 36035 48164 36268 48192
rect 36035 48161 36047 48164
rect 35989 48155 36047 48161
rect 36262 48152 36268 48164
rect 36320 48152 36326 48204
rect 36722 48192 36728 48204
rect 36683 48164 36728 48192
rect 36722 48152 36728 48164
rect 36780 48152 36786 48204
rect 36832 48192 36860 48232
rect 37274 48220 37280 48272
rect 37332 48260 37338 48272
rect 41230 48260 41236 48272
rect 37332 48232 41236 48260
rect 37332 48220 37338 48232
rect 41230 48220 41236 48232
rect 41288 48220 41294 48272
rect 41325 48263 41383 48269
rect 41325 48229 41337 48263
rect 41371 48260 41383 48263
rect 42426 48260 42432 48272
rect 41371 48232 42432 48260
rect 41371 48229 41383 48232
rect 41325 48223 41383 48229
rect 42426 48220 42432 48232
rect 42484 48220 42490 48272
rect 41414 48192 41420 48204
rect 36832 48164 41420 48192
rect 41414 48152 41420 48164
rect 41472 48152 41478 48204
rect 41782 48192 41788 48204
rect 41743 48164 41788 48192
rect 41782 48152 41788 48164
rect 41840 48152 41846 48204
rect 42518 48192 42524 48204
rect 42479 48164 42524 48192
rect 42518 48152 42524 48164
rect 42576 48152 42582 48204
rect 46290 48192 46296 48204
rect 46251 48164 46296 48192
rect 46290 48152 46296 48164
rect 46348 48152 46354 48204
rect 46842 48192 46848 48204
rect 46803 48164 46848 48192
rect 46842 48152 46848 48164
rect 46900 48152 46906 48204
rect 31846 48124 31852 48136
rect 31807 48096 31852 48124
rect 31846 48084 31852 48096
rect 31904 48084 31910 48136
rect 35437 48127 35495 48133
rect 35437 48093 35449 48127
rect 35483 48124 35495 48127
rect 35802 48124 35808 48136
rect 35483 48096 35808 48124
rect 35483 48093 35495 48096
rect 35437 48087 35495 48093
rect 35802 48084 35808 48096
rect 35860 48084 35866 48136
rect 39853 48127 39911 48133
rect 39853 48093 39865 48127
rect 39899 48093 39911 48127
rect 44082 48124 44088 48136
rect 44043 48096 44088 48124
rect 39853 48087 39911 48093
rect 29730 48056 29736 48068
rect 28224 48028 29592 48056
rect 29691 48028 29736 48056
rect 28224 48016 28230 48028
rect 29730 48016 29736 48028
rect 29788 48016 29794 48068
rect 29822 48016 29828 48068
rect 29880 48056 29886 48068
rect 31754 48056 31760 48068
rect 29880 48028 31760 48056
rect 29880 48016 29886 48028
rect 31754 48016 31760 48028
rect 31812 48016 31818 48068
rect 32030 48056 32036 48068
rect 31991 48028 32036 48056
rect 32030 48016 32036 48028
rect 32088 48016 32094 48068
rect 36173 48059 36231 48065
rect 36173 48025 36185 48059
rect 36219 48056 36231 48059
rect 36538 48056 36544 48068
rect 36219 48028 36544 48056
rect 36219 48025 36231 48028
rect 36173 48019 36231 48025
rect 36538 48016 36544 48028
rect 36596 48016 36602 48068
rect 35437 47991 35495 47997
rect 35437 47988 35449 47991
rect 16546 47960 35449 47988
rect 35437 47957 35449 47960
rect 35483 47957 35495 47991
rect 35437 47951 35495 47957
rect 35894 47948 35900 48000
rect 35952 47988 35958 48000
rect 36446 47988 36452 48000
rect 35952 47960 36452 47988
rect 35952 47948 35958 47960
rect 36446 47948 36452 47960
rect 36504 47988 36510 48000
rect 39868 47988 39896 48087
rect 44082 48084 44088 48096
rect 44140 48084 44146 48136
rect 45005 48127 45063 48133
rect 45005 48093 45017 48127
rect 45051 48093 45063 48127
rect 45646 48124 45652 48136
rect 45607 48096 45652 48124
rect 45005 48087 45063 48093
rect 41782 48016 41788 48068
rect 41840 48056 41846 48068
rect 41969 48059 42027 48065
rect 41969 48056 41981 48059
rect 41840 48028 41981 48056
rect 41840 48016 41846 48028
rect 41969 48025 41981 48028
rect 42015 48025 42027 48059
rect 45020 48056 45048 48087
rect 45646 48084 45652 48096
rect 45704 48084 45710 48136
rect 41969 48019 42027 48025
rect 42076 48028 45048 48056
rect 46477 48059 46535 48065
rect 42076 47988 42104 48028
rect 46477 48025 46489 48059
rect 46523 48056 46535 48059
rect 47670 48056 47676 48068
rect 46523 48028 47676 48056
rect 46523 48025 46535 48028
rect 46477 48019 46535 48025
rect 47670 48016 47676 48028
rect 47728 48016 47734 48068
rect 36504 47960 42104 47988
rect 36504 47948 36510 47960
rect 44174 47948 44180 48000
rect 44232 47988 44238 48000
rect 44269 47991 44327 47997
rect 44269 47988 44281 47991
rect 44232 47960 44281 47988
rect 44232 47948 44238 47960
rect 44269 47957 44281 47960
rect 44315 47957 44327 47991
rect 44269 47951 44327 47957
rect 44358 47948 44364 48000
rect 44416 47988 44422 48000
rect 45741 47991 45799 47997
rect 45741 47988 45753 47991
rect 44416 47960 45753 47988
rect 44416 47948 44422 47960
rect 45741 47957 45753 47960
rect 45787 47957 45799 47991
rect 45741 47951 45799 47957
rect 1104 47898 48852 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 48852 47898
rect 1104 47824 48852 47846
rect 1578 47744 1584 47796
rect 1636 47784 1642 47796
rect 3237 47787 3295 47793
rect 3237 47784 3249 47787
rect 1636 47756 3249 47784
rect 1636 47744 1642 47756
rect 3237 47753 3249 47756
rect 3283 47753 3295 47787
rect 4154 47784 4160 47796
rect 4115 47756 4160 47784
rect 3237 47747 3295 47753
rect 4154 47744 4160 47756
rect 4212 47744 4218 47796
rect 5442 47744 5448 47796
rect 5500 47784 5506 47796
rect 10226 47784 10232 47796
rect 5500 47756 10088 47784
rect 10187 47756 10232 47784
rect 5500 47744 5506 47756
rect 2590 47716 2596 47728
rect 2551 47688 2596 47716
rect 2590 47676 2596 47688
rect 2648 47676 2654 47728
rect 2682 47676 2688 47728
rect 2740 47716 2746 47728
rect 6638 47716 6644 47728
rect 2740 47688 6644 47716
rect 2740 47676 2746 47688
rect 1854 47648 1860 47660
rect 1815 47620 1860 47648
rect 1854 47608 1860 47620
rect 1912 47608 1918 47660
rect 2498 47648 2504 47660
rect 2459 47620 2504 47648
rect 2498 47608 2504 47620
rect 2556 47608 2562 47660
rect 3142 47648 3148 47660
rect 3103 47620 3148 47648
rect 3142 47608 3148 47620
rect 3200 47608 3206 47660
rect 4062 47648 4068 47660
rect 4023 47620 4068 47648
rect 4062 47608 4068 47620
rect 4120 47608 4126 47660
rect 4908 47657 4936 47688
rect 6638 47676 6644 47688
rect 6696 47676 6702 47728
rect 6825 47719 6883 47725
rect 6825 47685 6837 47719
rect 6871 47716 6883 47719
rect 7561 47719 7619 47725
rect 7561 47716 7573 47719
rect 6871 47688 7573 47716
rect 6871 47685 6883 47688
rect 6825 47679 6883 47685
rect 7561 47685 7573 47688
rect 7607 47685 7619 47719
rect 7561 47679 7619 47685
rect 4893 47651 4951 47657
rect 4893 47617 4905 47651
rect 4939 47617 4951 47651
rect 4893 47611 4951 47617
rect 5537 47651 5595 47657
rect 5537 47617 5549 47651
rect 5583 47617 5595 47651
rect 5537 47611 5595 47617
rect 6733 47651 6791 47657
rect 6733 47617 6745 47651
rect 6779 47648 6791 47651
rect 7374 47648 7380 47660
rect 6779 47620 6868 47648
rect 7335 47620 7380 47648
rect 6779 47617 6791 47620
rect 6733 47611 6791 47617
rect 2041 47515 2099 47521
rect 2041 47481 2053 47515
rect 2087 47512 2099 47515
rect 2406 47512 2412 47524
rect 2087 47484 2412 47512
rect 2087 47481 2099 47484
rect 2041 47475 2099 47481
rect 2406 47472 2412 47484
rect 2464 47472 2470 47524
rect 4798 47472 4804 47524
rect 4856 47512 4862 47524
rect 5552 47512 5580 47611
rect 6840 47592 6868 47620
rect 7374 47608 7380 47620
rect 7432 47608 7438 47660
rect 6822 47540 6828 47592
rect 6880 47540 6886 47592
rect 7834 47580 7840 47592
rect 7795 47552 7840 47580
rect 7834 47540 7840 47552
rect 7892 47540 7898 47592
rect 9950 47512 9956 47524
rect 4856 47484 9956 47512
rect 4856 47472 4862 47484
rect 9950 47472 9956 47484
rect 10008 47472 10014 47524
rect 10060 47512 10088 47756
rect 10226 47744 10232 47756
rect 10284 47744 10290 47796
rect 10870 47784 10876 47796
rect 10831 47756 10876 47784
rect 10870 47744 10876 47756
rect 10928 47744 10934 47796
rect 12526 47744 12532 47796
rect 12584 47784 12590 47796
rect 13357 47787 13415 47793
rect 13357 47784 13369 47787
rect 12584 47756 13369 47784
rect 12584 47744 12590 47756
rect 13357 47753 13369 47756
rect 13403 47753 13415 47787
rect 14366 47784 14372 47796
rect 14327 47756 14372 47784
rect 13357 47747 13415 47753
rect 14366 47744 14372 47756
rect 14424 47744 14430 47796
rect 14918 47744 14924 47796
rect 14976 47784 14982 47796
rect 18506 47784 18512 47796
rect 14976 47756 18512 47784
rect 14976 47744 14982 47756
rect 18506 47744 18512 47756
rect 18564 47744 18570 47796
rect 18601 47787 18659 47793
rect 18601 47753 18613 47787
rect 18647 47784 18659 47787
rect 19426 47784 19432 47796
rect 18647 47756 19432 47784
rect 18647 47753 18659 47756
rect 18601 47747 18659 47753
rect 19426 47744 19432 47756
rect 19484 47744 19490 47796
rect 22002 47744 22008 47796
rect 22060 47784 22066 47796
rect 22281 47787 22339 47793
rect 22281 47784 22293 47787
rect 22060 47756 22293 47784
rect 22060 47744 22066 47756
rect 22281 47753 22293 47756
rect 22327 47753 22339 47787
rect 22281 47747 22339 47753
rect 22738 47744 22744 47796
rect 22796 47784 22802 47796
rect 22925 47787 22983 47793
rect 22925 47784 22937 47787
rect 22796 47756 22937 47784
rect 22796 47744 22802 47756
rect 22925 47753 22937 47756
rect 22971 47753 22983 47787
rect 24210 47784 24216 47796
rect 24171 47756 24216 47784
rect 22925 47747 22983 47753
rect 24210 47744 24216 47756
rect 24268 47744 24274 47796
rect 24302 47744 24308 47796
rect 24360 47784 24366 47796
rect 26142 47784 26148 47796
rect 24360 47756 26148 47784
rect 24360 47744 24366 47756
rect 26142 47744 26148 47756
rect 26200 47744 26206 47796
rect 26329 47787 26387 47793
rect 26329 47753 26341 47787
rect 26375 47784 26387 47787
rect 27154 47784 27160 47796
rect 26375 47756 27160 47784
rect 26375 47753 26387 47756
rect 26329 47747 26387 47753
rect 27154 47744 27160 47756
rect 27212 47744 27218 47796
rect 27341 47787 27399 47793
rect 27341 47753 27353 47787
rect 27387 47784 27399 47787
rect 27614 47784 27620 47796
rect 27387 47756 27620 47784
rect 27387 47753 27399 47756
rect 27341 47747 27399 47753
rect 27614 47744 27620 47756
rect 27672 47744 27678 47796
rect 28074 47744 28080 47796
rect 28132 47784 28138 47796
rect 30374 47784 30380 47796
rect 28132 47756 30380 47784
rect 28132 47744 28138 47756
rect 30374 47744 30380 47756
rect 30432 47744 30438 47796
rect 30558 47784 30564 47796
rect 30519 47756 30564 47784
rect 30558 47744 30564 47756
rect 30616 47744 30622 47796
rect 31205 47787 31263 47793
rect 31205 47753 31217 47787
rect 31251 47784 31263 47787
rect 32030 47784 32036 47796
rect 31251 47756 32036 47784
rect 31251 47753 31263 47756
rect 31205 47747 31263 47753
rect 32030 47744 32036 47756
rect 32088 47744 32094 47796
rect 32217 47787 32275 47793
rect 32217 47753 32229 47787
rect 32263 47784 32275 47787
rect 32306 47784 32312 47796
rect 32263 47756 32312 47784
rect 32263 47753 32275 47756
rect 32217 47747 32275 47753
rect 32306 47744 32312 47756
rect 32364 47744 32370 47796
rect 35897 47787 35955 47793
rect 35897 47753 35909 47787
rect 35943 47784 35955 47787
rect 35986 47784 35992 47796
rect 35943 47756 35992 47784
rect 35943 47753 35955 47756
rect 35897 47747 35955 47753
rect 35986 47744 35992 47756
rect 36044 47744 36050 47796
rect 36538 47784 36544 47796
rect 36499 47756 36544 47784
rect 36538 47744 36544 47756
rect 36596 47744 36602 47796
rect 41782 47784 41788 47796
rect 41743 47756 41788 47784
rect 41782 47744 41788 47756
rect 41840 47744 41846 47796
rect 45462 47784 45468 47796
rect 42444 47756 45468 47784
rect 13170 47716 13176 47728
rect 10152 47688 13176 47716
rect 10152 47657 10180 47688
rect 13170 47676 13176 47688
rect 13228 47676 13234 47728
rect 17773 47719 17831 47725
rect 17773 47685 17785 47719
rect 17819 47716 17831 47719
rect 19978 47716 19984 47728
rect 17819 47688 19984 47716
rect 17819 47685 17831 47688
rect 17773 47679 17831 47685
rect 19978 47676 19984 47688
rect 20036 47676 20042 47728
rect 32953 47719 33011 47725
rect 21376 47688 32904 47716
rect 10137 47651 10195 47657
rect 10137 47617 10149 47651
rect 10183 47617 10195 47651
rect 10778 47648 10784 47660
rect 10739 47620 10784 47648
rect 10137 47611 10195 47617
rect 10778 47608 10784 47620
rect 10836 47608 10842 47660
rect 10962 47608 10968 47660
rect 11020 47648 11026 47660
rect 11517 47651 11575 47657
rect 11517 47648 11529 47651
rect 11020 47620 11529 47648
rect 11020 47608 11026 47620
rect 11517 47617 11529 47620
rect 11563 47617 11575 47651
rect 13262 47648 13268 47660
rect 11517 47611 11575 47617
rect 12084 47620 13124 47648
rect 13223 47620 13268 47648
rect 10502 47540 10508 47592
rect 10560 47580 10566 47592
rect 12084 47580 12112 47620
rect 12342 47580 12348 47592
rect 10560 47552 12112 47580
rect 12303 47552 12348 47580
rect 10560 47540 10566 47552
rect 12342 47540 12348 47552
rect 12400 47540 12406 47592
rect 13096 47580 13124 47620
rect 13262 47608 13268 47620
rect 13320 47608 13326 47660
rect 14277 47651 14335 47657
rect 14277 47617 14289 47651
rect 14323 47617 14335 47651
rect 14277 47611 14335 47617
rect 14292 47580 14320 47611
rect 14458 47608 14464 47660
rect 14516 47648 14522 47660
rect 15473 47651 15531 47657
rect 15473 47648 15485 47651
rect 14516 47620 15485 47648
rect 14516 47608 14522 47620
rect 15473 47617 15485 47620
rect 15519 47617 15531 47651
rect 15473 47611 15531 47617
rect 15838 47608 15844 47660
rect 15896 47648 15902 47660
rect 17497 47651 17555 47657
rect 17497 47648 17509 47651
rect 15896 47620 17509 47648
rect 15896 47608 15902 47620
rect 17497 47617 17509 47620
rect 17543 47617 17555 47651
rect 17497 47611 17555 47617
rect 18046 47608 18052 47660
rect 18104 47648 18110 47660
rect 18509 47651 18567 47657
rect 18509 47648 18521 47651
rect 18104 47620 18521 47648
rect 18104 47608 18110 47620
rect 18509 47617 18521 47620
rect 18555 47617 18567 47651
rect 18509 47611 18567 47617
rect 21376 47580 21404 47688
rect 22189 47651 22247 47657
rect 22189 47617 22201 47651
rect 22235 47617 22247 47651
rect 22830 47648 22836 47660
rect 22791 47620 22836 47648
rect 22189 47611 22247 47617
rect 13096 47552 21404 47580
rect 22204 47580 22232 47611
rect 22830 47608 22836 47620
rect 22888 47608 22894 47660
rect 23658 47608 23664 47660
rect 23716 47648 23722 47660
rect 24121 47651 24179 47657
rect 24121 47648 24133 47651
rect 23716 47620 24133 47648
rect 23716 47608 23722 47620
rect 24121 47617 24133 47620
rect 24167 47648 24179 47651
rect 24670 47648 24676 47660
rect 24167 47620 24676 47648
rect 24167 47617 24179 47620
rect 24121 47611 24179 47617
rect 24670 47608 24676 47620
rect 24728 47608 24734 47660
rect 24946 47648 24952 47660
rect 24907 47620 24952 47648
rect 24946 47608 24952 47620
rect 25004 47608 25010 47660
rect 25501 47651 25559 47657
rect 25501 47617 25513 47651
rect 25547 47648 25559 47651
rect 26050 47648 26056 47660
rect 25547 47620 26056 47648
rect 25547 47617 25559 47620
rect 25501 47611 25559 47617
rect 26050 47608 26056 47620
rect 26108 47608 26114 47660
rect 26237 47651 26295 47657
rect 26237 47617 26249 47651
rect 26283 47648 26295 47651
rect 27246 47648 27252 47660
rect 26283 47620 26317 47648
rect 27207 47620 27252 47648
rect 26283 47617 26295 47620
rect 26237 47611 26295 47617
rect 23106 47580 23112 47592
rect 22204 47552 23112 47580
rect 23106 47540 23112 47552
rect 23164 47540 23170 47592
rect 25685 47583 25743 47589
rect 25685 47549 25697 47583
rect 25731 47580 25743 47583
rect 25866 47580 25872 47592
rect 25731 47552 25872 47580
rect 25731 47549 25743 47552
rect 25685 47543 25743 47549
rect 25866 47540 25872 47552
rect 25924 47540 25930 47592
rect 25958 47540 25964 47592
rect 26016 47580 26022 47592
rect 26252 47580 26280 47611
rect 27246 47608 27252 47620
rect 27304 47608 27310 47660
rect 28166 47648 28172 47660
rect 28127 47620 28172 47648
rect 28166 47608 28172 47620
rect 28224 47608 28230 47660
rect 30469 47651 30527 47657
rect 30469 47617 30481 47651
rect 30515 47617 30527 47651
rect 31110 47648 31116 47660
rect 31071 47620 31116 47648
rect 30469 47611 30527 47617
rect 27982 47580 27988 47592
rect 26016 47552 27988 47580
rect 26016 47540 26022 47552
rect 27982 47540 27988 47552
rect 28040 47540 28046 47592
rect 28353 47583 28411 47589
rect 28353 47549 28365 47583
rect 28399 47580 28411 47583
rect 28534 47580 28540 47592
rect 28399 47552 28540 47580
rect 28399 47549 28411 47552
rect 28353 47543 28411 47549
rect 28534 47540 28540 47552
rect 28592 47540 28598 47592
rect 28629 47583 28687 47589
rect 28629 47549 28641 47583
rect 28675 47549 28687 47583
rect 28629 47543 28687 47549
rect 28644 47512 28672 47543
rect 10060 47484 28672 47512
rect 4982 47444 4988 47456
rect 4943 47416 4988 47444
rect 4982 47404 4988 47416
rect 5040 47404 5046 47456
rect 5629 47447 5687 47453
rect 5629 47413 5641 47447
rect 5675 47444 5687 47447
rect 6178 47444 6184 47456
rect 5675 47416 6184 47444
rect 5675 47413 5687 47416
rect 5629 47407 5687 47413
rect 6178 47404 6184 47416
rect 6236 47404 6242 47456
rect 22094 47404 22100 47456
rect 22152 47444 22158 47456
rect 25958 47444 25964 47456
rect 22152 47416 25964 47444
rect 22152 47404 22158 47416
rect 25958 47404 25964 47416
rect 26016 47404 26022 47456
rect 26142 47404 26148 47456
rect 26200 47444 26206 47456
rect 27246 47444 27252 47456
rect 26200 47416 27252 47444
rect 26200 47404 26206 47416
rect 27246 47404 27252 47416
rect 27304 47444 27310 47456
rect 30484 47444 30512 47611
rect 31110 47608 31116 47620
rect 31168 47608 31174 47660
rect 32122 47648 32128 47660
rect 32083 47620 32128 47648
rect 32122 47608 32128 47620
rect 32180 47608 32186 47660
rect 32876 47657 32904 47688
rect 32953 47685 32965 47719
rect 32999 47716 33011 47719
rect 33689 47719 33747 47725
rect 33689 47716 33701 47719
rect 32999 47688 33701 47716
rect 32999 47685 33011 47688
rect 32953 47679 33011 47685
rect 33689 47685 33701 47688
rect 33735 47685 33747 47719
rect 33689 47679 33747 47685
rect 32861 47651 32919 47657
rect 32861 47617 32873 47651
rect 32907 47617 32919 47651
rect 33502 47648 33508 47660
rect 33463 47620 33508 47648
rect 32861 47611 32919 47617
rect 33502 47608 33508 47620
rect 33560 47608 33566 47660
rect 35802 47648 35808 47660
rect 35763 47620 35808 47648
rect 35802 47608 35808 47620
rect 35860 47608 35866 47660
rect 36446 47648 36452 47660
rect 36407 47620 36452 47648
rect 36446 47608 36452 47620
rect 36504 47608 36510 47660
rect 41690 47648 41696 47660
rect 41651 47620 41696 47648
rect 41690 47608 41696 47620
rect 41748 47608 41754 47660
rect 42444 47657 42472 47756
rect 45462 47744 45468 47756
rect 45520 47744 45526 47796
rect 42613 47719 42671 47725
rect 42613 47685 42625 47719
rect 42659 47716 42671 47719
rect 44358 47716 44364 47728
rect 42659 47688 44364 47716
rect 42659 47685 42671 47688
rect 42613 47679 42671 47685
rect 44358 47676 44364 47688
rect 44416 47676 44422 47728
rect 45646 47716 45652 47728
rect 44468 47688 45652 47716
rect 42429 47651 42487 47657
rect 42429 47617 42441 47651
rect 42475 47617 42487 47651
rect 42429 47611 42487 47617
rect 31754 47540 31760 47592
rect 31812 47580 31818 47592
rect 32490 47580 32496 47592
rect 31812 47552 32496 47580
rect 31812 47540 31818 47552
rect 32490 47540 32496 47552
rect 32548 47540 32554 47592
rect 34698 47580 34704 47592
rect 34659 47552 34704 47580
rect 34698 47540 34704 47552
rect 34756 47540 34762 47592
rect 43990 47580 43996 47592
rect 43951 47552 43996 47580
rect 43990 47540 43996 47552
rect 44048 47540 44054 47592
rect 30558 47472 30564 47524
rect 30616 47512 30622 47524
rect 44468 47512 44496 47688
rect 45646 47676 45652 47688
rect 45704 47676 45710 47728
rect 47854 47648 47860 47660
rect 47815 47620 47860 47648
rect 47854 47608 47860 47620
rect 47912 47608 47918 47660
rect 44726 47580 44732 47592
rect 44687 47552 44732 47580
rect 44726 47540 44732 47552
rect 44784 47540 44790 47592
rect 44913 47583 44971 47589
rect 44913 47549 44925 47583
rect 44959 47580 44971 47583
rect 45094 47580 45100 47592
rect 44959 47552 45100 47580
rect 44959 47549 44971 47552
rect 44913 47543 44971 47549
rect 45094 47540 45100 47552
rect 45152 47540 45158 47592
rect 45186 47540 45192 47592
rect 45244 47580 45250 47592
rect 45244 47552 45289 47580
rect 45244 47540 45250 47552
rect 30616 47484 44496 47512
rect 30616 47472 30622 47484
rect 48038 47444 48044 47456
rect 27304 47416 30512 47444
rect 47999 47416 48044 47444
rect 27304 47404 27310 47416
rect 48038 47404 48044 47416
rect 48096 47404 48102 47456
rect 1104 47354 48852 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 48852 47354
rect 1104 47280 48852 47302
rect 1394 47200 1400 47252
rect 1452 47240 1458 47252
rect 1765 47243 1823 47249
rect 1765 47240 1777 47243
rect 1452 47212 1777 47240
rect 1452 47200 1458 47212
rect 1765 47209 1777 47212
rect 1811 47209 1823 47243
rect 3970 47240 3976 47252
rect 3931 47212 3976 47240
rect 1765 47203 1823 47209
rect 3970 47200 3976 47212
rect 4028 47200 4034 47252
rect 18506 47200 18512 47252
rect 18564 47240 18570 47252
rect 24302 47240 24308 47252
rect 18564 47212 24308 47240
rect 18564 47200 18570 47212
rect 24302 47200 24308 47212
rect 24360 47200 24366 47252
rect 25406 47240 25412 47252
rect 25367 47212 25412 47240
rect 25406 47200 25412 47212
rect 25464 47200 25470 47252
rect 26050 47240 26056 47252
rect 26011 47212 26056 47240
rect 26050 47200 26056 47212
rect 26108 47200 26114 47252
rect 26881 47243 26939 47249
rect 26881 47209 26893 47243
rect 26927 47240 26939 47243
rect 26970 47240 26976 47252
rect 26927 47212 26976 47240
rect 26927 47209 26939 47212
rect 26881 47203 26939 47209
rect 26970 47200 26976 47212
rect 27028 47200 27034 47252
rect 27890 47240 27896 47252
rect 27851 47212 27896 47240
rect 27890 47200 27896 47212
rect 27948 47200 27954 47252
rect 27982 47200 27988 47252
rect 28040 47240 28046 47252
rect 29641 47243 29699 47249
rect 28040 47212 28488 47240
rect 28040 47200 28046 47212
rect 12342 47132 12348 47184
rect 12400 47172 12406 47184
rect 28460 47172 28488 47212
rect 29641 47209 29653 47243
rect 29687 47240 29699 47243
rect 29730 47240 29736 47252
rect 29687 47212 29736 47240
rect 29687 47209 29699 47212
rect 29641 47203 29699 47209
rect 29730 47200 29736 47212
rect 29788 47200 29794 47252
rect 30469 47243 30527 47249
rect 30469 47209 30481 47243
rect 30515 47240 30527 47243
rect 31846 47240 31852 47252
rect 30515 47212 31852 47240
rect 30515 47209 30527 47212
rect 30469 47203 30527 47209
rect 31846 47200 31852 47212
rect 31904 47200 31910 47252
rect 45094 47240 45100 47252
rect 45055 47212 45100 47240
rect 45094 47200 45100 47212
rect 45152 47200 45158 47252
rect 45738 47240 45744 47252
rect 45699 47212 45744 47240
rect 45738 47200 45744 47212
rect 45796 47200 45802 47252
rect 35802 47172 35808 47184
rect 12400 47144 28396 47172
rect 28460 47144 35808 47172
rect 12400 47132 12406 47144
rect 4798 47104 4804 47116
rect 4759 47076 4804 47104
rect 4798 47064 4804 47076
rect 4856 47064 4862 47116
rect 4982 47104 4988 47116
rect 4943 47076 4988 47104
rect 4982 47064 4988 47076
rect 5040 47064 5046 47116
rect 5534 47104 5540 47116
rect 5495 47076 5540 47104
rect 5534 47064 5540 47076
rect 5592 47064 5598 47116
rect 6886 47076 10640 47104
rect 2222 47036 2228 47048
rect 2135 47008 2228 47036
rect 2222 46996 2228 47008
rect 2280 47036 2286 47048
rect 2682 47036 2688 47048
rect 2280 47008 2688 47036
rect 2280 46996 2286 47008
rect 2682 46996 2688 47008
rect 2740 46996 2746 47048
rect 2866 46996 2872 47048
rect 2924 47036 2930 47048
rect 3053 47039 3111 47045
rect 3053 47036 3065 47039
rect 2924 47008 3065 47036
rect 2924 46996 2930 47008
rect 3053 47005 3065 47008
rect 3099 47005 3111 47039
rect 3053 46999 3111 47005
rect 6178 46996 6184 47048
rect 6236 47036 6242 47048
rect 6886 47036 6914 47076
rect 6236 47008 6914 47036
rect 10229 47039 10287 47045
rect 6236 46996 6242 47008
rect 10229 47005 10241 47039
rect 10275 47005 10287 47039
rect 10502 47036 10508 47048
rect 10463 47008 10508 47036
rect 10229 46999 10287 47005
rect 1578 46860 1584 46912
rect 1636 46900 1642 46912
rect 2317 46903 2375 46909
rect 2317 46900 2329 46903
rect 1636 46872 2329 46900
rect 1636 46860 1642 46872
rect 2317 46869 2329 46872
rect 2363 46869 2375 46903
rect 10244 46900 10272 46999
rect 10502 46996 10508 47008
rect 10560 46996 10566 47048
rect 10612 47036 10640 47076
rect 10778 47064 10784 47116
rect 10836 47104 10842 47116
rect 28368 47104 28396 47144
rect 35802 47132 35808 47144
rect 35860 47172 35866 47184
rect 45646 47172 45652 47184
rect 35860 47144 45652 47172
rect 35860 47132 35866 47144
rect 45646 47132 45652 47144
rect 45704 47132 45710 47184
rect 49602 47172 49608 47184
rect 45756 47144 49608 47172
rect 10836 47076 28304 47104
rect 28368 47076 28488 47104
rect 10836 47064 10842 47076
rect 24946 47036 24952 47048
rect 10612 47008 24952 47036
rect 24946 46996 24952 47008
rect 25004 46996 25010 47048
rect 25590 47036 25596 47048
rect 25551 47008 25596 47036
rect 25590 46996 25596 47008
rect 25648 46996 25654 47048
rect 26234 46996 26240 47048
rect 26292 47036 26298 47048
rect 27801 47039 27859 47045
rect 26292 47008 26337 47036
rect 26292 46996 26298 47008
rect 27801 47005 27813 47039
rect 27847 47005 27859 47039
rect 27801 46999 27859 47005
rect 10962 46928 10968 46980
rect 11020 46968 11026 46980
rect 11149 46971 11207 46977
rect 11149 46968 11161 46971
rect 11020 46940 11161 46968
rect 11020 46928 11026 46940
rect 11149 46937 11161 46940
rect 11195 46937 11207 46971
rect 11149 46931 11207 46937
rect 12250 46928 12256 46980
rect 12308 46968 12314 46980
rect 12897 46971 12955 46977
rect 12897 46968 12909 46971
rect 12308 46940 12909 46968
rect 12308 46928 12314 46940
rect 12897 46937 12909 46940
rect 12943 46968 12955 46971
rect 27816 46968 27844 46999
rect 12943 46940 27844 46968
rect 28276 46968 28304 47076
rect 28460 47045 28488 47076
rect 28534 47064 28540 47116
rect 28592 47104 28598 47116
rect 42613 47107 42671 47113
rect 28592 47076 28637 47104
rect 28592 47064 28598 47076
rect 42613 47073 42625 47107
rect 42659 47104 42671 47107
rect 43162 47104 43168 47116
rect 42659 47076 43168 47104
rect 42659 47073 42671 47076
rect 42613 47067 42671 47073
rect 43162 47064 43168 47076
rect 43220 47064 43226 47116
rect 44453 47107 44511 47113
rect 44453 47073 44465 47107
rect 44499 47104 44511 47107
rect 45756 47104 45784 47144
rect 49602 47132 49608 47144
rect 49660 47132 49666 47184
rect 44499 47076 45784 47104
rect 44499 47073 44511 47076
rect 44453 47067 44511 47073
rect 46658 47064 46664 47116
rect 46716 47104 46722 47116
rect 46753 47107 46811 47113
rect 46753 47104 46765 47107
rect 46716 47076 46765 47104
rect 46716 47064 46722 47076
rect 46753 47073 46765 47076
rect 46799 47073 46811 47107
rect 46753 47067 46811 47073
rect 28445 47039 28503 47045
rect 28445 47005 28457 47039
rect 28491 47036 28503 47039
rect 29549 47039 29607 47045
rect 29549 47036 29561 47039
rect 28491 47008 29561 47036
rect 28491 47005 28503 47008
rect 28445 46999 28503 47005
rect 29549 47005 29561 47008
rect 29595 47005 29607 47039
rect 29549 46999 29607 47005
rect 45005 47039 45063 47045
rect 45005 47005 45017 47039
rect 45051 47036 45063 47039
rect 45186 47036 45192 47048
rect 45051 47008 45192 47036
rect 45051 47005 45063 47008
rect 45005 46999 45063 47005
rect 45186 46996 45192 47008
rect 45244 46996 45250 47048
rect 45646 47036 45652 47048
rect 45607 47008 45652 47036
rect 45646 46996 45652 47008
rect 45704 46996 45710 47048
rect 46293 47039 46351 47045
rect 46293 47005 46305 47039
rect 46339 47005 46351 47039
rect 46293 46999 46351 47005
rect 32122 46968 32128 46980
rect 28276 46940 32128 46968
rect 12943 46937 12955 46940
rect 12897 46931 12955 46937
rect 32122 46928 32128 46940
rect 32180 46928 32186 46980
rect 42794 46968 42800 46980
rect 42755 46940 42800 46968
rect 42794 46928 42800 46940
rect 42852 46928 42858 46980
rect 44266 46928 44272 46980
rect 44324 46968 44330 46980
rect 46308 46968 46336 46999
rect 46474 46968 46480 46980
rect 44324 46940 46336 46968
rect 46435 46940 46480 46968
rect 44324 46928 44330 46940
rect 46474 46928 46480 46940
rect 46532 46928 46538 46980
rect 10980 46900 11008 46928
rect 10244 46872 11008 46900
rect 2317 46863 2375 46869
rect 1104 46810 48852 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 48852 46810
rect 1104 46736 48852 46758
rect 10873 46699 10931 46705
rect 10873 46665 10885 46699
rect 10919 46696 10931 46699
rect 10962 46696 10968 46708
rect 10919 46668 10968 46696
rect 10919 46665 10931 46668
rect 10873 46659 10931 46665
rect 10962 46656 10968 46668
rect 11020 46696 11026 46708
rect 13170 46696 13176 46708
rect 11020 46668 11928 46696
rect 13131 46668 13176 46696
rect 11020 46656 11026 46668
rect 2866 46628 2872 46640
rect 1780 46600 2872 46628
rect 1780 46569 1808 46600
rect 2866 46588 2872 46600
rect 2924 46588 2930 46640
rect 11900 46637 11928 46668
rect 13170 46656 13176 46668
rect 13228 46656 13234 46708
rect 38654 46696 38660 46708
rect 16546 46668 38660 46696
rect 11885 46631 11943 46637
rect 11885 46597 11897 46631
rect 11931 46597 11943 46631
rect 11885 46591 11943 46597
rect 1765 46563 1823 46569
rect 1765 46529 1777 46563
rect 1811 46529 1823 46563
rect 1765 46523 1823 46529
rect 9950 46520 9956 46572
rect 10008 46560 10014 46572
rect 10689 46563 10747 46569
rect 10689 46560 10701 46563
rect 10008 46532 10701 46560
rect 10008 46520 10014 46532
rect 10689 46529 10701 46532
rect 10735 46560 10747 46563
rect 15930 46560 15936 46572
rect 10735 46532 15936 46560
rect 10735 46529 10747 46532
rect 10689 46523 10747 46529
rect 15930 46520 15936 46532
rect 15988 46520 15994 46572
rect 1946 46492 1952 46504
rect 1907 46464 1952 46492
rect 1946 46452 1952 46464
rect 2004 46452 2010 46504
rect 2774 46492 2780 46504
rect 2735 46464 2780 46492
rect 2774 46452 2780 46464
rect 2832 46452 2838 46504
rect 10686 46384 10692 46436
rect 10744 46424 10750 46436
rect 16546 46424 16574 46668
rect 38654 46656 38660 46668
rect 38712 46656 38718 46708
rect 47670 46696 47676 46708
rect 47631 46668 47676 46696
rect 47670 46656 47676 46668
rect 47728 46656 47734 46708
rect 22830 46588 22836 46640
rect 22888 46628 22894 46640
rect 22888 46600 47624 46628
rect 22888 46588 22894 46600
rect 43162 46560 43168 46572
rect 43123 46532 43168 46560
rect 43162 46520 43168 46532
rect 43220 46520 43226 46572
rect 43993 46563 44051 46569
rect 43993 46529 44005 46563
rect 44039 46560 44051 46563
rect 44266 46560 44272 46572
rect 44039 46532 44272 46560
rect 44039 46529 44051 46532
rect 43993 46523 44051 46529
rect 44266 46520 44272 46532
rect 44324 46520 44330 46572
rect 44450 46520 44456 46572
rect 44508 46560 44514 46572
rect 47596 46569 47624 46600
rect 44637 46563 44695 46569
rect 44637 46560 44649 46563
rect 44508 46532 44649 46560
rect 44508 46520 44514 46532
rect 44637 46529 44649 46532
rect 44683 46529 44695 46563
rect 44637 46523 44695 46529
rect 47581 46563 47639 46569
rect 47581 46529 47593 46563
rect 47627 46529 47639 46563
rect 47581 46523 47639 46529
rect 38105 46495 38163 46501
rect 38105 46461 38117 46495
rect 38151 46461 38163 46495
rect 38105 46455 38163 46461
rect 38289 46495 38347 46501
rect 38289 46461 38301 46495
rect 38335 46492 38347 46495
rect 38470 46492 38476 46504
rect 38335 46464 38476 46492
rect 38335 46461 38347 46464
rect 38289 46455 38347 46461
rect 10744 46396 16574 46424
rect 10744 46384 10750 46396
rect 1394 46316 1400 46368
rect 1452 46356 1458 46368
rect 4249 46359 4307 46365
rect 4249 46356 4261 46359
rect 1452 46328 4261 46356
rect 1452 46316 1458 46328
rect 4249 46325 4261 46328
rect 4295 46325 4307 46359
rect 38120 46356 38148 46455
rect 38470 46452 38476 46464
rect 38528 46452 38534 46504
rect 38654 46492 38660 46504
rect 38615 46464 38660 46492
rect 38654 46452 38660 46464
rect 38712 46452 38718 46504
rect 45094 46452 45100 46504
rect 45152 46492 45158 46504
rect 45189 46495 45247 46501
rect 45189 46492 45201 46495
rect 45152 46464 45201 46492
rect 45152 46452 45158 46464
rect 45189 46461 45201 46464
rect 45235 46461 45247 46495
rect 45370 46492 45376 46504
rect 45331 46464 45376 46492
rect 45189 46455 45247 46461
rect 45370 46452 45376 46464
rect 45428 46452 45434 46504
rect 46842 46492 46848 46504
rect 46803 46464 46848 46492
rect 46842 46452 46848 46464
rect 46900 46452 46906 46504
rect 38654 46356 38660 46368
rect 38120 46328 38660 46356
rect 4249 46319 4307 46325
rect 38654 46316 38660 46328
rect 38712 46316 38718 46368
rect 1104 46266 48852 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 48852 46266
rect 1104 46192 48852 46214
rect 38470 46152 38476 46164
rect 38431 46124 38476 46152
rect 38470 46112 38476 46124
rect 38528 46112 38534 46164
rect 44453 46155 44511 46161
rect 44453 46121 44465 46155
rect 44499 46152 44511 46155
rect 44726 46152 44732 46164
rect 44499 46124 44732 46152
rect 44499 46121 44511 46124
rect 44453 46115 44511 46121
rect 44726 46112 44732 46124
rect 44784 46112 44790 46164
rect 45281 46155 45339 46161
rect 45281 46121 45293 46155
rect 45327 46152 45339 46155
rect 45370 46152 45376 46164
rect 45327 46124 45376 46152
rect 45327 46121 45339 46124
rect 45281 46115 45339 46121
rect 45370 46112 45376 46124
rect 45428 46112 45434 46164
rect 1394 46016 1400 46028
rect 1355 45988 1400 46016
rect 1394 45976 1400 45988
rect 1452 45976 1458 46028
rect 1578 46016 1584 46028
rect 1539 45988 1584 46016
rect 1578 45976 1584 45988
rect 1636 45976 1642 46028
rect 2774 46016 2780 46028
rect 2735 45988 2780 46016
rect 2774 45976 2780 45988
rect 2832 45976 2838 46028
rect 48130 46016 48136 46028
rect 48091 45988 48136 46016
rect 48130 45976 48136 45988
rect 48188 45976 48194 46028
rect 10962 45908 10968 45960
rect 11020 45948 11026 45960
rect 11149 45951 11207 45957
rect 11149 45948 11161 45951
rect 11020 45920 11161 45948
rect 11020 45908 11026 45920
rect 11149 45917 11161 45920
rect 11195 45917 11207 45951
rect 11149 45911 11207 45917
rect 38381 45951 38439 45957
rect 38381 45917 38393 45951
rect 38427 45948 38439 45951
rect 41690 45948 41696 45960
rect 38427 45920 41696 45948
rect 38427 45917 38439 45920
rect 38381 45911 38439 45917
rect 41690 45908 41696 45920
rect 41748 45908 41754 45960
rect 45186 45948 45192 45960
rect 45147 45920 45192 45948
rect 45186 45908 45192 45920
rect 45244 45908 45250 45960
rect 46290 45948 46296 45960
rect 46251 45920 46296 45948
rect 46290 45908 46296 45920
rect 46348 45908 46354 45960
rect 7466 45840 7472 45892
rect 7524 45880 7530 45892
rect 11885 45883 11943 45889
rect 11885 45880 11897 45883
rect 7524 45852 11897 45880
rect 7524 45840 7530 45852
rect 11885 45849 11897 45852
rect 11931 45880 11943 45883
rect 22094 45880 22100 45892
rect 11931 45852 22100 45880
rect 11931 45849 11943 45852
rect 11885 45843 11943 45849
rect 22094 45840 22100 45852
rect 22152 45840 22158 45892
rect 46477 45883 46535 45889
rect 46477 45849 46489 45883
rect 46523 45880 46535 45883
rect 47026 45880 47032 45892
rect 46523 45852 47032 45880
rect 46523 45849 46535 45852
rect 46477 45843 46535 45849
rect 47026 45840 47032 45852
rect 47084 45840 47090 45892
rect 1104 45722 48852 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 48852 45722
rect 1104 45648 48852 45670
rect 22094 45568 22100 45620
rect 22152 45608 22158 45620
rect 22830 45608 22836 45620
rect 22152 45580 22836 45608
rect 22152 45568 22158 45580
rect 22830 45568 22836 45580
rect 22888 45568 22894 45620
rect 46937 45543 46995 45549
rect 46937 45509 46949 45543
rect 46983 45540 46995 45543
rect 47026 45540 47032 45552
rect 46983 45512 47032 45540
rect 46983 45509 46995 45512
rect 46937 45503 46995 45509
rect 47026 45500 47032 45512
rect 47084 45500 47090 45552
rect 1394 45472 1400 45484
rect 1355 45444 1400 45472
rect 1394 45432 1400 45444
rect 1452 45432 1458 45484
rect 2222 45472 2228 45484
rect 2183 45444 2228 45472
rect 2222 45432 2228 45444
rect 2280 45432 2286 45484
rect 12986 45432 12992 45484
rect 13044 45472 13050 45484
rect 46845 45475 46903 45481
rect 46845 45472 46857 45475
rect 13044 45444 46857 45472
rect 13044 45432 13050 45444
rect 46845 45441 46857 45444
rect 46891 45441 46903 45475
rect 46845 45435 46903 45441
rect 47581 45475 47639 45481
rect 47581 45441 47593 45475
rect 47627 45472 47639 45475
rect 47762 45472 47768 45484
rect 47627 45444 47768 45472
rect 47627 45441 47639 45444
rect 47581 45435 47639 45441
rect 47762 45432 47768 45444
rect 47820 45432 47826 45484
rect 2406 45364 2412 45416
rect 2464 45404 2470 45416
rect 2590 45404 2596 45416
rect 2464 45376 2596 45404
rect 2464 45364 2470 45376
rect 2590 45364 2596 45376
rect 2648 45364 2654 45416
rect 45094 45404 45100 45416
rect 45055 45376 45100 45404
rect 45094 45364 45100 45376
rect 45152 45364 45158 45416
rect 45278 45364 45284 45416
rect 45336 45404 45342 45416
rect 45741 45407 45799 45413
rect 45741 45404 45753 45407
rect 45336 45376 45753 45404
rect 45336 45364 45342 45376
rect 45741 45373 45753 45376
rect 45787 45373 45799 45407
rect 45741 45367 45799 45373
rect 46290 45364 46296 45416
rect 46348 45404 46354 45416
rect 46385 45407 46443 45413
rect 46385 45404 46397 45407
rect 46348 45376 46397 45404
rect 46348 45364 46354 45376
rect 46385 45373 46397 45376
rect 46431 45373 46443 45407
rect 46385 45367 46443 45373
rect 46474 45364 46480 45416
rect 46532 45404 46538 45416
rect 47673 45407 47731 45413
rect 47673 45404 47685 45407
rect 46532 45376 47685 45404
rect 46532 45364 46538 45376
rect 47673 45373 47685 45376
rect 47719 45373 47731 45407
rect 47673 45367 47731 45373
rect 1581 45339 1639 45345
rect 1581 45305 1593 45339
rect 1627 45336 1639 45339
rect 1627 45308 6914 45336
rect 1627 45305 1639 45308
rect 1581 45299 1639 45305
rect 2406 45268 2412 45280
rect 2367 45240 2412 45268
rect 2406 45228 2412 45240
rect 2464 45228 2470 45280
rect 6886 45268 6914 45308
rect 19426 45268 19432 45280
rect 6886 45240 19432 45268
rect 19426 45228 19432 45240
rect 19484 45228 19490 45280
rect 1104 45178 48852 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 48852 45178
rect 1104 45104 48852 45126
rect 1946 45024 1952 45076
rect 2004 45064 2010 45076
rect 2225 45067 2283 45073
rect 2225 45064 2237 45067
rect 2004 45036 2237 45064
rect 2004 45024 2010 45036
rect 2225 45033 2237 45036
rect 2271 45033 2283 45067
rect 2225 45027 2283 45033
rect 45462 45024 45468 45076
rect 45520 45064 45526 45076
rect 45833 45067 45891 45073
rect 45833 45064 45845 45067
rect 45520 45036 45845 45064
rect 45520 45024 45526 45036
rect 45833 45033 45845 45036
rect 45879 45033 45891 45067
rect 45833 45027 45891 45033
rect 31941 44931 31999 44937
rect 31941 44897 31953 44931
rect 31987 44928 31999 44931
rect 32122 44928 32128 44940
rect 31987 44900 32128 44928
rect 31987 44897 31999 44900
rect 31941 44891 31999 44897
rect 32122 44888 32128 44900
rect 32180 44888 32186 44940
rect 33781 44931 33839 44937
rect 33781 44897 33793 44931
rect 33827 44928 33839 44931
rect 37274 44928 37280 44940
rect 33827 44900 37280 44928
rect 33827 44897 33839 44900
rect 33781 44891 33839 44897
rect 37274 44888 37280 44900
rect 37332 44888 37338 44940
rect 48130 44928 48136 44940
rect 48091 44900 48136 44928
rect 48130 44888 48136 44900
rect 48188 44888 48194 44940
rect 1394 44860 1400 44872
rect 1355 44832 1400 44860
rect 1394 44820 1400 44832
rect 1452 44820 1458 44872
rect 2133 44863 2191 44869
rect 2133 44829 2145 44863
rect 2179 44860 2191 44863
rect 2222 44860 2228 44872
rect 2179 44832 2228 44860
rect 2179 44829 2191 44832
rect 2133 44823 2191 44829
rect 2222 44820 2228 44832
rect 2280 44820 2286 44872
rect 2961 44863 3019 44869
rect 2961 44829 2973 44863
rect 3007 44829 3019 44863
rect 2961 44823 3019 44829
rect 2038 44752 2044 44804
rect 2096 44792 2102 44804
rect 2976 44792 3004 44823
rect 16758 44820 16764 44872
rect 16816 44860 16822 44872
rect 17037 44863 17095 44869
rect 17037 44860 17049 44863
rect 16816 44832 17049 44860
rect 16816 44820 16822 44832
rect 17037 44829 17049 44832
rect 17083 44829 17095 44863
rect 46290 44860 46296 44872
rect 46251 44832 46296 44860
rect 17037 44823 17095 44829
rect 46290 44820 46296 44832
rect 46348 44820 46354 44872
rect 32125 44795 32183 44801
rect 32125 44792 32137 44795
rect 2096 44764 3004 44792
rect 26206 44764 32137 44792
rect 2096 44752 2102 44764
rect 1581 44727 1639 44733
rect 1581 44693 1593 44727
rect 1627 44724 1639 44727
rect 1670 44724 1676 44736
rect 1627 44696 1676 44724
rect 1627 44693 1639 44696
rect 1581 44687 1639 44693
rect 1670 44684 1676 44696
rect 1728 44684 1734 44736
rect 17221 44727 17279 44733
rect 17221 44693 17233 44727
rect 17267 44724 17279 44727
rect 26206 44724 26234 44764
rect 32125 44761 32137 44764
rect 32171 44761 32183 44795
rect 32125 44755 32183 44761
rect 46477 44795 46535 44801
rect 46477 44761 46489 44795
rect 46523 44792 46535 44795
rect 47670 44792 47676 44804
rect 46523 44764 47676 44792
rect 46523 44761 46535 44764
rect 46477 44755 46535 44761
rect 47670 44752 47676 44764
rect 47728 44752 47734 44804
rect 17267 44696 26234 44724
rect 17267 44693 17279 44696
rect 17221 44687 17279 44693
rect 1104 44634 48852 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 48852 44634
rect 1104 44560 48852 44582
rect 47670 44520 47676 44532
rect 47631 44492 47676 44520
rect 47670 44480 47676 44492
rect 47728 44480 47734 44532
rect 2038 44384 2044 44396
rect 1999 44356 2044 44384
rect 2038 44344 2044 44356
rect 2096 44344 2102 44396
rect 46290 44344 46296 44396
rect 46348 44384 46354 44396
rect 47029 44387 47087 44393
rect 47029 44384 47041 44387
rect 46348 44356 47041 44384
rect 46348 44344 46354 44356
rect 47029 44353 47041 44356
rect 47075 44353 47087 44387
rect 47578 44384 47584 44396
rect 47539 44356 47584 44384
rect 47029 44347 47087 44353
rect 47578 44344 47584 44356
rect 47636 44344 47642 44396
rect 2225 44319 2283 44325
rect 2225 44285 2237 44319
rect 2271 44316 2283 44319
rect 2958 44316 2964 44328
rect 2271 44288 2964 44316
rect 2271 44285 2283 44288
rect 2225 44279 2283 44285
rect 2958 44276 2964 44288
rect 3016 44276 3022 44328
rect 3050 44276 3056 44328
rect 3108 44316 3114 44328
rect 3108 44288 3153 44316
rect 3108 44276 3114 44288
rect 17218 44140 17224 44192
rect 17276 44180 17282 44192
rect 26142 44180 26148 44192
rect 17276 44152 26148 44180
rect 17276 44140 17282 44152
rect 26142 44140 26148 44152
rect 26200 44140 26206 44192
rect 1104 44090 48852 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 48852 44090
rect 1104 44016 48852 44038
rect 2958 43976 2964 43988
rect 2919 43948 2964 43976
rect 2958 43936 2964 43948
rect 3016 43936 3022 43988
rect 1394 43772 1400 43784
rect 1355 43744 1400 43772
rect 1394 43732 1400 43744
rect 1452 43732 1458 43784
rect 2869 43775 2927 43781
rect 2869 43741 2881 43775
rect 2915 43772 2927 43775
rect 3326 43772 3332 43784
rect 2915 43744 3332 43772
rect 2915 43741 2927 43744
rect 2869 43735 2927 43741
rect 3326 43732 3332 43744
rect 3384 43732 3390 43784
rect 36078 43732 36084 43784
rect 36136 43772 36142 43784
rect 36357 43775 36415 43781
rect 36357 43772 36369 43775
rect 36136 43744 36369 43772
rect 36136 43732 36142 43744
rect 36357 43741 36369 43744
rect 36403 43741 36415 43775
rect 47302 43772 47308 43784
rect 47263 43744 47308 43772
rect 36357 43735 36415 43741
rect 47302 43732 47308 43744
rect 47360 43732 47366 43784
rect 47486 43732 47492 43784
rect 47544 43772 47550 43784
rect 48133 43775 48191 43781
rect 48133 43772 48145 43775
rect 47544 43744 48145 43772
rect 47544 43732 47550 43744
rect 48133 43741 48145 43744
rect 48179 43741 48191 43775
rect 48133 43735 48191 43741
rect 1673 43707 1731 43713
rect 1673 43673 1685 43707
rect 1719 43704 1731 43707
rect 1762 43704 1768 43716
rect 1719 43676 1768 43704
rect 1719 43673 1731 43676
rect 1673 43667 1731 43673
rect 1762 43664 1768 43676
rect 1820 43664 1826 43716
rect 36538 43704 36544 43716
rect 36499 43676 36544 43704
rect 36538 43664 36544 43676
rect 36596 43664 36602 43716
rect 38197 43707 38255 43713
rect 38197 43673 38209 43707
rect 38243 43704 38255 43707
rect 46842 43704 46848 43716
rect 38243 43676 46848 43704
rect 38243 43673 38255 43676
rect 38197 43667 38255 43673
rect 46842 43664 46848 43676
rect 46900 43664 46906 43716
rect 47394 43636 47400 43648
rect 47355 43608 47400 43636
rect 47394 43596 47400 43608
rect 47452 43596 47458 43648
rect 1104 43546 48852 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 48852 43546
rect 1104 43472 48852 43494
rect 36538 43432 36544 43444
rect 36499 43404 36544 43432
rect 36538 43392 36544 43404
rect 36596 43392 36602 43444
rect 36446 43296 36452 43308
rect 36407 43268 36452 43296
rect 36446 43256 36452 43268
rect 36504 43256 36510 43308
rect 47854 43296 47860 43308
rect 47815 43268 47860 43296
rect 47854 43256 47860 43268
rect 47912 43256 47918 43308
rect 47670 43052 47676 43104
rect 47728 43092 47734 43104
rect 48041 43095 48099 43101
rect 48041 43092 48053 43095
rect 47728 43064 48053 43092
rect 47728 43052 47734 43064
rect 48041 43061 48053 43064
rect 48087 43061 48099 43095
rect 48041 43055 48099 43061
rect 1104 43002 48852 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 48852 43002
rect 1104 42928 48852 42950
rect 46477 42755 46535 42761
rect 46477 42721 46489 42755
rect 46523 42752 46535 42755
rect 47394 42752 47400 42764
rect 46523 42724 47400 42752
rect 46523 42721 46535 42724
rect 46477 42715 46535 42721
rect 47394 42712 47400 42724
rect 47452 42712 47458 42764
rect 48130 42752 48136 42764
rect 48091 42724 48136 42752
rect 48130 42712 48136 42724
rect 48188 42712 48194 42764
rect 46293 42687 46351 42693
rect 46293 42653 46305 42687
rect 46339 42653 46351 42687
rect 46293 42647 46351 42653
rect 46308 42616 46336 42647
rect 47486 42616 47492 42628
rect 46308 42588 47492 42616
rect 47486 42576 47492 42588
rect 47544 42576 47550 42628
rect 1104 42458 48852 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 48852 42458
rect 1104 42384 48852 42406
rect 47946 42208 47952 42220
rect 47907 42180 47952 42208
rect 47946 42168 47952 42180
rect 48004 42168 48010 42220
rect 28442 42032 28448 42084
rect 28500 42072 28506 42084
rect 48133 42075 48191 42081
rect 48133 42072 48145 42075
rect 28500 42044 48145 42072
rect 28500 42032 28506 42044
rect 48133 42041 48145 42044
rect 48179 42041 48191 42075
rect 48133 42035 48191 42041
rect 1394 41964 1400 42016
rect 1452 42004 1458 42016
rect 2041 42007 2099 42013
rect 2041 42004 2053 42007
rect 1452 41976 2053 42004
rect 1452 41964 1458 41976
rect 2041 41973 2053 41976
rect 2087 41973 2099 42007
rect 2041 41967 2099 41973
rect 46290 41964 46296 42016
rect 46348 42004 46354 42016
rect 47029 42007 47087 42013
rect 47029 42004 47041 42007
rect 46348 41976 47041 42004
rect 46348 41964 46354 41976
rect 47029 41973 47041 41976
rect 47075 41973 47087 42007
rect 47029 41967 47087 41973
rect 1104 41914 48852 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 48852 41914
rect 1104 41840 48852 41862
rect 1394 41664 1400 41676
rect 1355 41636 1400 41664
rect 1394 41624 1400 41636
rect 1452 41624 1458 41676
rect 1854 41664 1860 41676
rect 1815 41636 1860 41664
rect 1854 41624 1860 41636
rect 1912 41624 1918 41676
rect 46290 41664 46296 41676
rect 46251 41636 46296 41664
rect 46290 41624 46296 41636
rect 46348 41624 46354 41676
rect 1578 41528 1584 41540
rect 1539 41500 1584 41528
rect 1578 41488 1584 41500
rect 1636 41488 1642 41540
rect 46474 41528 46480 41540
rect 46435 41500 46480 41528
rect 46474 41488 46480 41500
rect 46532 41488 46538 41540
rect 48130 41528 48136 41540
rect 48091 41500 48136 41528
rect 48130 41488 48136 41500
rect 48188 41488 48194 41540
rect 1104 41370 48852 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 48852 41370
rect 1104 41296 48852 41318
rect 1578 41216 1584 41268
rect 1636 41256 1642 41268
rect 2225 41259 2283 41265
rect 2225 41256 2237 41259
rect 1636 41228 2237 41256
rect 1636 41216 1642 41228
rect 2225 41225 2237 41228
rect 2271 41225 2283 41259
rect 2225 41219 2283 41225
rect 46474 41216 46480 41268
rect 46532 41256 46538 41268
rect 46845 41259 46903 41265
rect 46845 41256 46857 41259
rect 46532 41228 46857 41256
rect 46532 41216 46538 41228
rect 46845 41225 46857 41228
rect 46891 41225 46903 41259
rect 46845 41219 46903 41225
rect 1394 41120 1400 41132
rect 1355 41092 1400 41120
rect 1394 41080 1400 41092
rect 1452 41080 1458 41132
rect 2133 41123 2191 41129
rect 2133 41089 2145 41123
rect 2179 41120 2191 41123
rect 2314 41120 2320 41132
rect 2179 41092 2320 41120
rect 2179 41089 2191 41092
rect 2133 41083 2191 41089
rect 2314 41080 2320 41092
rect 2372 41080 2378 41132
rect 41690 41080 41696 41132
rect 41748 41120 41754 41132
rect 46658 41120 46664 41132
rect 41748 41092 46664 41120
rect 41748 41080 41754 41092
rect 46658 41080 46664 41092
rect 46716 41120 46722 41132
rect 46753 41123 46811 41129
rect 46753 41120 46765 41123
rect 46716 41092 46765 41120
rect 46716 41080 46722 41092
rect 46753 41089 46765 41092
rect 46799 41089 46811 41123
rect 47854 41120 47860 41132
rect 47815 41092 47860 41120
rect 46753 41083 46811 41089
rect 47854 41080 47860 41092
rect 47912 41080 47918 41132
rect 1581 40919 1639 40925
rect 1581 40885 1593 40919
rect 1627 40916 1639 40919
rect 1946 40916 1952 40928
rect 1627 40888 1952 40916
rect 1627 40885 1639 40888
rect 1581 40879 1639 40885
rect 1946 40876 1952 40888
rect 2004 40876 2010 40928
rect 48041 40919 48099 40925
rect 48041 40885 48053 40919
rect 48087 40916 48099 40919
rect 48222 40916 48228 40928
rect 48087 40888 48228 40916
rect 48087 40885 48099 40888
rect 48041 40879 48099 40885
rect 48222 40876 48228 40888
rect 48280 40876 48286 40928
rect 1104 40826 48852 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 48852 40826
rect 1104 40752 48852 40774
rect 46293 40579 46351 40585
rect 46293 40545 46305 40579
rect 46339 40576 46351 40579
rect 47026 40576 47032 40588
rect 46339 40548 47032 40576
rect 46339 40545 46351 40548
rect 46293 40539 46351 40545
rect 47026 40536 47032 40548
rect 47084 40536 47090 40588
rect 1854 40440 1860 40452
rect 1815 40412 1860 40440
rect 1854 40400 1860 40412
rect 1912 40400 1918 40452
rect 2041 40443 2099 40449
rect 2041 40409 2053 40443
rect 2087 40440 2099 40443
rect 3694 40440 3700 40452
rect 2087 40412 3700 40440
rect 2087 40409 2099 40412
rect 2041 40403 2099 40409
rect 3694 40400 3700 40412
rect 3752 40400 3758 40452
rect 46477 40443 46535 40449
rect 46477 40409 46489 40443
rect 46523 40440 46535 40443
rect 47670 40440 47676 40452
rect 46523 40412 47676 40440
rect 46523 40409 46535 40412
rect 46477 40403 46535 40409
rect 47670 40400 47676 40412
rect 47728 40400 47734 40452
rect 48130 40440 48136 40452
rect 48091 40412 48136 40440
rect 48130 40400 48136 40412
rect 48188 40400 48194 40452
rect 1104 40282 48852 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 48852 40282
rect 1104 40208 48852 40230
rect 47026 40032 47032 40044
rect 46987 40004 47032 40032
rect 47026 39992 47032 40004
rect 47084 39992 47090 40044
rect 47581 40035 47639 40041
rect 47581 40001 47593 40035
rect 47627 40001 47639 40035
rect 47581 39995 47639 40001
rect 45646 39924 45652 39976
rect 45704 39964 45710 39976
rect 47596 39964 47624 39995
rect 47670 39992 47676 40044
rect 47728 40032 47734 40044
rect 47728 40004 47773 40032
rect 47728 39992 47734 40004
rect 45704 39936 47624 39964
rect 45704 39924 45710 39936
rect 1394 39788 1400 39840
rect 1452 39828 1458 39840
rect 2041 39831 2099 39837
rect 2041 39828 2053 39831
rect 1452 39800 2053 39828
rect 1452 39788 1458 39800
rect 2041 39797 2053 39800
rect 2087 39797 2099 39831
rect 2041 39791 2099 39797
rect 1104 39738 48852 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 48852 39738
rect 1104 39664 48852 39686
rect 1394 39488 1400 39500
rect 1355 39460 1400 39488
rect 1394 39448 1400 39460
rect 1452 39448 1458 39500
rect 2774 39488 2780 39500
rect 2735 39460 2780 39488
rect 2774 39448 2780 39460
rect 2832 39448 2838 39500
rect 24394 39448 24400 39500
rect 24452 39488 24458 39500
rect 24452 39460 24808 39488
rect 24452 39448 24458 39460
rect 6638 39380 6644 39432
rect 6696 39420 6702 39432
rect 6825 39423 6883 39429
rect 6825 39420 6837 39423
rect 6696 39392 6837 39420
rect 6696 39380 6702 39392
rect 6825 39389 6837 39392
rect 6871 39389 6883 39423
rect 7466 39420 7472 39432
rect 7427 39392 7472 39420
rect 6825 39383 6883 39389
rect 7466 39380 7472 39392
rect 7524 39380 7530 39432
rect 24486 39380 24492 39432
rect 24544 39420 24550 39432
rect 24780 39429 24808 39460
rect 24673 39423 24731 39429
rect 24673 39420 24685 39423
rect 24544 39392 24685 39420
rect 24544 39380 24550 39392
rect 24673 39389 24685 39392
rect 24719 39389 24731 39423
rect 24673 39383 24731 39389
rect 24765 39423 24823 39429
rect 24765 39389 24777 39423
rect 24811 39389 24823 39423
rect 24765 39383 24823 39389
rect 24857 39423 24915 39429
rect 24857 39389 24869 39423
rect 24903 39389 24915 39423
rect 24857 39383 24915 39389
rect 1581 39355 1639 39361
rect 1581 39321 1593 39355
rect 1627 39352 1639 39355
rect 2130 39352 2136 39364
rect 1627 39324 2136 39352
rect 1627 39321 1639 39324
rect 1581 39315 1639 39321
rect 2130 39312 2136 39324
rect 2188 39312 2194 39364
rect 24872 39352 24900 39383
rect 24946 39380 24952 39432
rect 25004 39420 25010 39432
rect 25041 39423 25099 39429
rect 25041 39420 25053 39423
rect 25004 39392 25053 39420
rect 25004 39380 25010 39392
rect 25041 39389 25053 39392
rect 25087 39389 25099 39423
rect 25041 39383 25099 39389
rect 46842 39380 46848 39432
rect 46900 39420 46906 39432
rect 47305 39423 47363 39429
rect 47305 39420 47317 39423
rect 46900 39392 47317 39420
rect 46900 39380 46906 39392
rect 47305 39389 47317 39392
rect 47351 39389 47363 39423
rect 47305 39383 47363 39389
rect 47581 39423 47639 39429
rect 47581 39389 47593 39423
rect 47627 39389 47639 39423
rect 47581 39383 47639 39389
rect 26326 39352 26332 39364
rect 24872 39324 26332 39352
rect 26326 39312 26332 39324
rect 26384 39312 26390 39364
rect 32214 39312 32220 39364
rect 32272 39352 32278 39364
rect 47596 39352 47624 39383
rect 32272 39324 47624 39352
rect 32272 39312 32278 39324
rect 6822 39244 6828 39296
rect 6880 39284 6886 39296
rect 7561 39287 7619 39293
rect 7561 39284 7573 39287
rect 6880 39256 7573 39284
rect 6880 39244 6886 39256
rect 7561 39253 7573 39256
rect 7607 39253 7619 39287
rect 7561 39247 7619 39253
rect 24397 39287 24455 39293
rect 24397 39253 24409 39287
rect 24443 39284 24455 39287
rect 24486 39284 24492 39296
rect 24443 39256 24492 39284
rect 24443 39253 24455 39256
rect 24397 39247 24455 39253
rect 24486 39244 24492 39256
rect 24544 39244 24550 39296
rect 1104 39194 48852 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 48852 39194
rect 1104 39120 48852 39142
rect 2130 39080 2136 39092
rect 2091 39052 2136 39080
rect 2130 39040 2136 39052
rect 2188 39040 2194 39092
rect 6822 39012 6828 39024
rect 6783 38984 6828 39012
rect 6822 38972 6828 38984
rect 6880 38972 6886 39024
rect 20530 38972 20536 39024
rect 20588 39012 20594 39024
rect 21085 39015 21143 39021
rect 21085 39012 21097 39015
rect 20588 38984 21097 39012
rect 20588 38972 20594 38984
rect 21085 38981 21097 38984
rect 21131 38981 21143 39015
rect 21085 38975 21143 38981
rect 1394 38904 1400 38956
rect 1452 38944 1458 38956
rect 2041 38947 2099 38953
rect 2041 38944 2053 38947
rect 1452 38916 2053 38944
rect 1452 38904 1458 38916
rect 2041 38913 2053 38916
rect 2087 38913 2099 38947
rect 6638 38944 6644 38956
rect 6599 38916 6644 38944
rect 2041 38907 2099 38913
rect 6638 38904 6644 38916
rect 6696 38904 6702 38956
rect 20898 38944 20904 38956
rect 20859 38916 20904 38944
rect 20898 38904 20904 38916
rect 20956 38904 20962 38956
rect 24026 38904 24032 38956
rect 24084 38944 24090 38956
rect 24193 38947 24251 38953
rect 24193 38944 24205 38947
rect 24084 38916 24205 38944
rect 24084 38904 24090 38916
rect 24193 38913 24205 38916
rect 24239 38913 24251 38947
rect 24193 38907 24251 38913
rect 5534 38836 5540 38888
rect 5592 38876 5598 38888
rect 7101 38879 7159 38885
rect 7101 38876 7113 38879
rect 5592 38848 7113 38876
rect 5592 38836 5598 38848
rect 7101 38845 7113 38848
rect 7147 38845 7159 38879
rect 23934 38876 23940 38888
rect 23895 38848 23940 38876
rect 7101 38839 7159 38845
rect 23934 38836 23940 38848
rect 23992 38836 23998 38888
rect 21082 38700 21088 38752
rect 21140 38740 21146 38752
rect 21269 38743 21327 38749
rect 21269 38740 21281 38743
rect 21140 38712 21281 38740
rect 21140 38700 21146 38712
rect 21269 38709 21281 38712
rect 21315 38709 21327 38743
rect 21269 38703 21327 38709
rect 25038 38700 25044 38752
rect 25096 38740 25102 38752
rect 25317 38743 25375 38749
rect 25317 38740 25329 38743
rect 25096 38712 25329 38740
rect 25096 38700 25102 38712
rect 25317 38709 25329 38712
rect 25363 38709 25375 38743
rect 47762 38740 47768 38752
rect 47723 38712 47768 38740
rect 25317 38703 25375 38709
rect 47762 38700 47768 38712
rect 47820 38700 47826 38752
rect 1104 38650 48852 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 48852 38650
rect 1104 38576 48852 38598
rect 20806 38428 20812 38480
rect 20864 38428 20870 38480
rect 5626 38360 5632 38412
rect 5684 38400 5690 38412
rect 5684 38372 20760 38400
rect 5684 38360 5690 38372
rect 20732 38341 20760 38372
rect 20824 38341 20852 38428
rect 21450 38400 21456 38412
rect 20916 38372 21456 38400
rect 20916 38341 20944 38372
rect 21450 38360 21456 38372
rect 21508 38360 21514 38412
rect 46293 38403 46351 38409
rect 46293 38369 46305 38403
rect 46339 38400 46351 38403
rect 47762 38400 47768 38412
rect 46339 38372 47768 38400
rect 46339 38369 46351 38372
rect 46293 38363 46351 38369
rect 47762 38360 47768 38372
rect 47820 38360 47826 38412
rect 48130 38400 48136 38412
rect 48091 38372 48136 38400
rect 48130 38360 48136 38372
rect 48188 38360 48194 38412
rect 20717 38335 20775 38341
rect 20717 38301 20729 38335
rect 20763 38301 20775 38335
rect 20717 38295 20775 38301
rect 20806 38335 20864 38341
rect 20806 38301 20818 38335
rect 20852 38301 20864 38335
rect 20806 38295 20864 38301
rect 20901 38335 20959 38341
rect 20901 38301 20913 38335
rect 20947 38301 20959 38335
rect 20901 38295 20959 38301
rect 21085 38335 21143 38341
rect 21085 38301 21097 38335
rect 21131 38332 21143 38335
rect 21266 38332 21272 38344
rect 21131 38304 21272 38332
rect 21131 38301 21143 38304
rect 21085 38295 21143 38301
rect 21266 38292 21272 38304
rect 21324 38292 21330 38344
rect 21542 38332 21548 38344
rect 21503 38304 21548 38332
rect 21542 38292 21548 38304
rect 21600 38292 21606 38344
rect 23934 38292 23940 38344
rect 23992 38332 23998 38344
rect 24397 38335 24455 38341
rect 24397 38332 24409 38335
rect 23992 38304 24409 38332
rect 23992 38292 23998 38304
rect 24397 38301 24409 38304
rect 24443 38301 24455 38335
rect 24397 38295 24455 38301
rect 20441 38267 20499 38273
rect 20441 38233 20453 38267
rect 20487 38264 20499 38267
rect 21790 38267 21848 38273
rect 21790 38264 21802 38267
rect 20487 38236 21802 38264
rect 20487 38233 20499 38236
rect 20441 38227 20499 38233
rect 21790 38233 21802 38236
rect 21836 38233 21848 38267
rect 21790 38227 21848 38233
rect 22738 38156 22744 38208
rect 22796 38196 22802 38208
rect 22925 38199 22983 38205
rect 22925 38196 22937 38199
rect 22796 38168 22937 38196
rect 22796 38156 22802 38168
rect 22925 38165 22937 38168
rect 22971 38165 22983 38199
rect 24412 38196 24440 38295
rect 24486 38292 24492 38344
rect 24544 38332 24550 38344
rect 24664 38335 24722 38341
rect 24664 38332 24676 38335
rect 24544 38304 24676 38332
rect 24544 38292 24550 38304
rect 24664 38301 24676 38304
rect 24710 38301 24722 38335
rect 26973 38335 27031 38341
rect 26973 38332 26985 38335
rect 24664 38295 24722 38301
rect 24780 38304 26985 38332
rect 24780 38208 24808 38304
rect 26973 38301 26985 38304
rect 27019 38301 27031 38335
rect 26973 38295 27031 38301
rect 26694 38224 26700 38276
rect 26752 38264 26758 38276
rect 27218 38267 27276 38273
rect 27218 38264 27230 38267
rect 26752 38236 27230 38264
rect 26752 38224 26758 38236
rect 27218 38233 27230 38236
rect 27264 38233 27276 38267
rect 27218 38227 27276 38233
rect 46477 38267 46535 38273
rect 46477 38233 46489 38267
rect 46523 38264 46535 38267
rect 46934 38264 46940 38276
rect 46523 38236 46940 38264
rect 46523 38233 46535 38236
rect 46477 38227 46535 38233
rect 46934 38224 46940 38236
rect 46992 38224 46998 38276
rect 24762 38196 24768 38208
rect 24412 38168 24768 38196
rect 22925 38159 22983 38165
rect 24762 38156 24768 38168
rect 24820 38156 24826 38208
rect 25774 38196 25780 38208
rect 25735 38168 25780 38196
rect 25774 38156 25780 38168
rect 25832 38156 25838 38208
rect 27982 38156 27988 38208
rect 28040 38196 28046 38208
rect 28353 38199 28411 38205
rect 28353 38196 28365 38199
rect 28040 38168 28365 38196
rect 28040 38156 28046 38168
rect 28353 38165 28365 38168
rect 28399 38165 28411 38199
rect 28353 38159 28411 38165
rect 1104 38106 48852 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 48852 38106
rect 1104 38032 48852 38054
rect 20898 37952 20904 38004
rect 20956 37992 20962 38004
rect 21821 37995 21879 38001
rect 21821 37992 21833 37995
rect 20956 37964 21833 37992
rect 20956 37952 20962 37964
rect 21821 37961 21833 37964
rect 21867 37961 21879 37995
rect 24026 37992 24032 38004
rect 23987 37964 24032 37992
rect 21821 37955 21879 37961
rect 24026 37952 24032 37964
rect 24084 37952 24090 38004
rect 24394 37952 24400 38004
rect 24452 37952 24458 38004
rect 26326 37992 26332 38004
rect 26287 37964 26332 37992
rect 26326 37952 26332 37964
rect 26384 37952 26390 38004
rect 40862 37992 40868 38004
rect 26436 37964 40868 37992
rect 20916 37896 24164 37924
rect 19334 37856 19340 37868
rect 19295 37828 19340 37856
rect 19334 37816 19340 37828
rect 19392 37816 19398 37868
rect 19521 37859 19579 37865
rect 19521 37825 19533 37859
rect 19567 37856 19579 37859
rect 20530 37856 20536 37868
rect 19567 37828 20536 37856
rect 19567 37825 19579 37828
rect 19521 37819 19579 37825
rect 20530 37816 20536 37828
rect 20588 37816 20594 37868
rect 20916 37865 20944 37896
rect 20901 37859 20959 37865
rect 20901 37825 20913 37859
rect 20947 37825 20959 37859
rect 20901 37819 20959 37825
rect 20993 37859 21051 37865
rect 20993 37825 21005 37859
rect 21039 37825 21051 37859
rect 20993 37819 21051 37825
rect 1394 37788 1400 37800
rect 1355 37760 1400 37788
rect 1394 37748 1400 37760
rect 1452 37748 1458 37800
rect 1673 37791 1731 37797
rect 1673 37757 1685 37791
rect 1719 37788 1731 37791
rect 1719 37760 6914 37788
rect 1719 37757 1731 37760
rect 1673 37751 1731 37757
rect 6886 37720 6914 37760
rect 19794 37748 19800 37800
rect 19852 37788 19858 37800
rect 20806 37788 20812 37800
rect 19852 37760 20812 37788
rect 19852 37748 19858 37760
rect 20806 37748 20812 37760
rect 20864 37788 20870 37800
rect 21008 37788 21036 37819
rect 21082 37816 21088 37868
rect 21140 37856 21146 37868
rect 21140 37828 21185 37856
rect 21140 37816 21146 37828
rect 21266 37816 21272 37868
rect 21324 37856 21330 37868
rect 22189 37859 22247 37865
rect 21324 37828 21417 37856
rect 21324 37816 21330 37828
rect 22189 37825 22201 37859
rect 22235 37856 22247 37859
rect 22370 37856 22376 37868
rect 22235 37828 22376 37856
rect 22235 37825 22247 37828
rect 22189 37819 22247 37825
rect 22370 37816 22376 37828
rect 22428 37816 22434 37868
rect 20864 37760 21036 37788
rect 20864 37748 20870 37760
rect 17770 37720 17776 37732
rect 6886 37692 17776 37720
rect 17770 37680 17776 37692
rect 17828 37680 17834 37732
rect 20990 37680 20996 37732
rect 21048 37720 21054 37732
rect 21284 37720 21312 37816
rect 22281 37791 22339 37797
rect 22281 37757 22293 37791
rect 22327 37757 22339 37791
rect 22462 37788 22468 37800
rect 22423 37760 22468 37788
rect 22281 37751 22339 37757
rect 21048 37692 21312 37720
rect 22296 37720 22324 37751
rect 22462 37748 22468 37760
rect 22520 37748 22526 37800
rect 24136 37788 24164 37896
rect 24409 37871 24437 37952
rect 24302 37856 24308 37868
rect 24263 37828 24308 37856
rect 24302 37816 24308 37828
rect 24360 37816 24366 37868
rect 24394 37865 24452 37871
rect 24394 37831 24406 37865
rect 24440 37831 24452 37865
rect 24394 37825 24452 37831
rect 24489 37859 24547 37865
rect 24489 37825 24501 37859
rect 24535 37825 24547 37859
rect 24489 37819 24547 37825
rect 24673 37859 24731 37865
rect 24673 37825 24685 37859
rect 24719 37856 24731 37859
rect 24946 37856 24952 37868
rect 24719 37828 24952 37856
rect 24719 37825 24731 37828
rect 24673 37819 24731 37825
rect 24504 37788 24532 37819
rect 24946 37816 24952 37828
rect 25004 37816 25010 37868
rect 25130 37856 25136 37868
rect 25091 37828 25136 37856
rect 25130 37816 25136 37828
rect 25188 37816 25194 37868
rect 25317 37859 25375 37865
rect 25317 37825 25329 37859
rect 25363 37856 25375 37859
rect 25958 37856 25964 37868
rect 25363 37828 25636 37856
rect 25919 37828 25964 37856
rect 25363 37825 25375 37828
rect 25317 37819 25375 37825
rect 25501 37791 25559 37797
rect 25501 37788 25513 37791
rect 24136 37760 24440 37788
rect 24504 37760 25513 37788
rect 24118 37720 24124 37732
rect 22296 37692 24124 37720
rect 21048 37680 21054 37692
rect 24118 37680 24124 37692
rect 24176 37680 24182 37732
rect 24412 37720 24440 37760
rect 25501 37757 25513 37760
rect 25547 37757 25559 37791
rect 25608 37788 25636 37828
rect 25958 37816 25964 37828
rect 26016 37816 26022 37868
rect 26145 37859 26203 37865
rect 26145 37825 26157 37859
rect 26191 37825 26203 37859
rect 26145 37819 26203 37825
rect 26050 37788 26056 37800
rect 25608 37760 26056 37788
rect 25501 37751 25559 37757
rect 26050 37748 26056 37760
rect 26108 37788 26114 37800
rect 26160 37788 26188 37819
rect 26108 37760 26188 37788
rect 26108 37748 26114 37760
rect 26436 37720 26464 37964
rect 40862 37952 40868 37964
rect 40920 37952 40926 38004
rect 46934 37992 46940 38004
rect 46895 37964 46940 37992
rect 46934 37952 46940 37964
rect 46992 37952 46998 38004
rect 29546 37924 29552 37936
rect 27540 37896 29552 37924
rect 27540 37865 27568 37896
rect 29546 37884 29552 37896
rect 29604 37884 29610 37936
rect 29914 37924 29920 37936
rect 29875 37896 29920 37924
rect 29914 37884 29920 37896
rect 29972 37884 29978 37936
rect 30133 37927 30191 37933
rect 30133 37893 30145 37927
rect 30179 37924 30191 37927
rect 31110 37924 31116 37936
rect 30179 37896 31116 37924
rect 30179 37893 30191 37896
rect 30133 37887 30191 37893
rect 31110 37884 31116 37896
rect 31168 37884 31174 37936
rect 47946 37924 47952 37936
rect 47907 37896 47952 37924
rect 47946 37884 47952 37896
rect 48004 37884 48010 37936
rect 27798 37865 27804 37868
rect 27525 37859 27583 37865
rect 27525 37825 27537 37859
rect 27571 37825 27583 37859
rect 27525 37819 27583 37825
rect 27792 37819 27804 37865
rect 27856 37856 27862 37868
rect 27856 37828 27892 37856
rect 27798 37816 27804 37819
rect 27856 37816 27862 37828
rect 46566 37816 46572 37868
rect 46624 37856 46630 37868
rect 46845 37859 46903 37865
rect 46845 37856 46857 37859
rect 46624 37828 46857 37856
rect 46624 37816 46630 37828
rect 46845 37825 46857 37828
rect 46891 37825 46903 37859
rect 46845 37819 46903 37825
rect 47026 37748 47032 37800
rect 47084 37788 47090 37800
rect 47210 37788 47216 37800
rect 47084 37760 47216 37788
rect 47084 37748 47090 37760
rect 47210 37748 47216 37760
rect 47268 37748 47274 37800
rect 24412 37692 26464 37720
rect 19702 37652 19708 37664
rect 19663 37624 19708 37652
rect 19702 37612 19708 37624
rect 19760 37612 19766 37664
rect 20625 37655 20683 37661
rect 20625 37621 20637 37655
rect 20671 37652 20683 37655
rect 20898 37652 20904 37664
rect 20671 37624 20904 37652
rect 20671 37621 20683 37624
rect 20625 37615 20683 37621
rect 20898 37612 20904 37624
rect 20956 37612 20962 37664
rect 28166 37612 28172 37664
rect 28224 37652 28230 37664
rect 28905 37655 28963 37661
rect 28905 37652 28917 37655
rect 28224 37624 28917 37652
rect 28224 37612 28230 37624
rect 28905 37621 28917 37624
rect 28951 37621 28963 37655
rect 30098 37652 30104 37664
rect 30059 37624 30104 37652
rect 28905 37615 28963 37621
rect 30098 37612 30104 37624
rect 30156 37612 30162 37664
rect 30282 37652 30288 37664
rect 30243 37624 30288 37652
rect 30282 37612 30288 37624
rect 30340 37612 30346 37664
rect 47394 37612 47400 37664
rect 47452 37652 47458 37664
rect 48041 37655 48099 37661
rect 48041 37652 48053 37655
rect 47452 37624 48053 37652
rect 47452 37612 47458 37624
rect 48041 37621 48053 37624
rect 48087 37621 48099 37655
rect 48041 37615 48099 37621
rect 1104 37562 48852 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 48852 37562
rect 1104 37488 48852 37510
rect 19334 37408 19340 37460
rect 19392 37448 19398 37460
rect 19613 37451 19671 37457
rect 19613 37448 19625 37451
rect 19392 37420 19625 37448
rect 19392 37408 19398 37420
rect 19613 37417 19625 37420
rect 19659 37417 19671 37451
rect 19613 37411 19671 37417
rect 20070 37408 20076 37460
rect 20128 37448 20134 37460
rect 20346 37448 20352 37460
rect 20128 37420 20352 37448
rect 20128 37408 20134 37420
rect 20346 37408 20352 37420
rect 20404 37408 20410 37460
rect 21542 37448 21548 37460
rect 20824 37420 21548 37448
rect 20070 37272 20076 37324
rect 20128 37312 20134 37324
rect 20165 37315 20223 37321
rect 20165 37312 20177 37315
rect 20128 37284 20177 37312
rect 20128 37272 20134 37284
rect 20165 37281 20177 37284
rect 20211 37281 20223 37315
rect 20165 37275 20223 37281
rect 17770 37204 17776 37256
rect 17828 37244 17834 37256
rect 18325 37247 18383 37253
rect 18325 37244 18337 37247
rect 17828 37216 18337 37244
rect 17828 37204 17834 37216
rect 18325 37213 18337 37216
rect 18371 37213 18383 37247
rect 18325 37207 18383 37213
rect 18414 37244 18472 37250
rect 18414 37210 18426 37244
rect 18460 37210 18472 37244
rect 18414 37204 18472 37210
rect 18509 37247 18567 37253
rect 18509 37213 18521 37247
rect 18555 37213 18567 37247
rect 18509 37207 18567 37213
rect 18693 37247 18751 37253
rect 18693 37213 18705 37247
rect 18739 37244 18751 37247
rect 18739 37216 20300 37244
rect 18739 37213 18751 37216
rect 18693 37207 18751 37213
rect 1854 37176 1860 37188
rect 1815 37148 1860 37176
rect 1854 37136 1860 37148
rect 1912 37136 1918 37188
rect 2038 37176 2044 37188
rect 1999 37148 2044 37176
rect 2038 37136 2044 37148
rect 2096 37136 2102 37188
rect 18432 37176 18460 37204
rect 18340 37148 18460 37176
rect 18524 37176 18552 37207
rect 19702 37176 19708 37188
rect 18524 37148 19708 37176
rect 18049 37111 18107 37117
rect 18049 37077 18061 37111
rect 18095 37108 18107 37111
rect 18138 37108 18144 37120
rect 18095 37080 18144 37108
rect 18095 37077 18107 37080
rect 18049 37071 18107 37077
rect 18138 37068 18144 37080
rect 18196 37068 18202 37120
rect 18340 37108 18368 37148
rect 19702 37136 19708 37148
rect 19760 37136 19766 37188
rect 19794 37136 19800 37188
rect 19852 37136 19858 37188
rect 20272 37176 20300 37216
rect 20622 37204 20628 37256
rect 20680 37244 20686 37256
rect 20824 37253 20852 37420
rect 21542 37408 21548 37420
rect 21600 37408 21606 37460
rect 24949 37451 25007 37457
rect 24949 37417 24961 37451
rect 24995 37448 25007 37451
rect 25958 37448 25964 37460
rect 24995 37420 25964 37448
rect 24995 37417 25007 37420
rect 24949 37411 25007 37417
rect 25958 37408 25964 37420
rect 26016 37408 26022 37460
rect 26694 37448 26700 37460
rect 26655 37420 26700 37448
rect 26694 37408 26700 37420
rect 26752 37408 26758 37460
rect 30190 37408 30196 37460
rect 30248 37448 30254 37460
rect 32401 37451 32459 37457
rect 32401 37448 32413 37451
rect 30248 37420 32413 37448
rect 30248 37408 30254 37420
rect 32401 37417 32413 37420
rect 32447 37417 32459 37451
rect 32401 37411 32459 37417
rect 47210 37408 47216 37460
rect 47268 37448 47274 37460
rect 47670 37448 47676 37460
rect 47268 37420 47676 37448
rect 47268 37408 47274 37420
rect 47670 37408 47676 37420
rect 47728 37408 47734 37460
rect 24118 37340 24124 37392
rect 24176 37380 24182 37392
rect 27982 37380 27988 37392
rect 24176 37352 27988 37380
rect 24176 37340 24182 37352
rect 27982 37340 27988 37352
rect 28040 37340 28046 37392
rect 25498 37312 25504 37324
rect 25459 37284 25504 37312
rect 25498 37272 25504 37284
rect 25556 37272 25562 37324
rect 27246 37312 27252 37324
rect 27077 37284 27252 37312
rect 20809 37247 20867 37253
rect 20809 37244 20821 37247
rect 20680 37216 20821 37244
rect 20680 37204 20686 37216
rect 20809 37213 20821 37216
rect 20855 37213 20867 37247
rect 20809 37207 20867 37213
rect 20898 37204 20904 37256
rect 20956 37244 20962 37256
rect 21076 37247 21134 37253
rect 21076 37244 21088 37247
rect 20956 37216 21088 37244
rect 20956 37204 20962 37216
rect 21076 37213 21088 37216
rect 21122 37213 21134 37247
rect 21076 37207 21134 37213
rect 26510 37204 26516 37256
rect 26568 37244 26574 37256
rect 27077 37253 27105 37284
rect 27246 37272 27252 37284
rect 27304 37272 27310 37324
rect 28350 37312 28356 37324
rect 28311 37284 28356 37312
rect 28350 37272 28356 37284
rect 28408 37272 28414 37324
rect 34606 37272 34612 37324
rect 34664 37312 34670 37324
rect 46842 37312 46848 37324
rect 34664 37284 46848 37312
rect 34664 37272 34670 37284
rect 46842 37272 46848 37284
rect 46900 37272 46906 37324
rect 26927 37247 26985 37253
rect 26927 37244 26939 37247
rect 26568 37216 26939 37244
rect 26568 37204 26574 37216
rect 26927 37213 26939 37216
rect 26973 37213 26985 37247
rect 26927 37207 26985 37213
rect 27046 37247 27105 37253
rect 27046 37213 27058 37247
rect 27092 37216 27105 37247
rect 27157 37247 27215 37253
rect 27092 37213 27104 37216
rect 27046 37207 27104 37213
rect 27157 37213 27169 37247
rect 27203 37213 27215 37247
rect 27157 37207 27215 37213
rect 20990 37176 20996 37188
rect 20272 37148 20996 37176
rect 20990 37136 20996 37148
rect 21048 37136 21054 37188
rect 25317 37179 25375 37185
rect 25317 37176 25329 37179
rect 21192 37148 25329 37176
rect 19334 37108 19340 37120
rect 18340 37080 19340 37108
rect 19334 37068 19340 37080
rect 19392 37108 19398 37120
rect 19812 37108 19840 37136
rect 19978 37108 19984 37120
rect 19392 37080 19840 37108
rect 19939 37080 19984 37108
rect 19392 37068 19398 37080
rect 19978 37068 19984 37080
rect 20036 37068 20042 37120
rect 20073 37111 20131 37117
rect 20073 37077 20085 37111
rect 20119 37108 20131 37111
rect 21192 37108 21220 37148
rect 25317 37145 25329 37148
rect 25363 37176 25375 37179
rect 25774 37176 25780 37188
rect 25363 37148 25780 37176
rect 25363 37145 25375 37148
rect 25317 37139 25375 37145
rect 25774 37136 25780 37148
rect 25832 37136 25838 37188
rect 27172 37176 27200 37207
rect 27338 37204 27344 37256
rect 27396 37244 27402 37256
rect 27706 37244 27712 37256
rect 27396 37216 27712 37244
rect 27396 37204 27402 37216
rect 27706 37204 27712 37216
rect 27764 37204 27770 37256
rect 29546 37244 29552 37256
rect 29507 37216 29552 37244
rect 29546 37204 29552 37216
rect 29604 37204 29610 37256
rect 31941 37247 31999 37253
rect 31941 37213 31953 37247
rect 31987 37244 31999 37247
rect 47670 37244 47676 37256
rect 31987 37216 32260 37244
rect 47631 37216 47676 37244
rect 31987 37213 31999 37216
rect 31941 37207 31999 37213
rect 32232 37188 32260 37216
rect 47670 37204 47676 37216
rect 47728 37204 47734 37256
rect 29178 37176 29184 37188
rect 27172 37148 29184 37176
rect 29178 37136 29184 37148
rect 29236 37136 29242 37188
rect 29822 37185 29828 37188
rect 29816 37139 29828 37185
rect 29880 37176 29886 37188
rect 29880 37148 29916 37176
rect 29822 37136 29828 37139
rect 29880 37136 29886 37148
rect 31110 37136 31116 37188
rect 31168 37176 31174 37188
rect 32214 37176 32220 37188
rect 31168 37148 31984 37176
rect 32175 37148 32220 37176
rect 31168 37136 31174 37148
rect 20119 37080 21220 37108
rect 22189 37111 22247 37117
rect 20119 37077 20131 37080
rect 20073 37071 20131 37077
rect 22189 37077 22201 37111
rect 22235 37108 22247 37111
rect 22370 37108 22376 37120
rect 22235 37080 22376 37108
rect 22235 37077 22247 37080
rect 22189 37071 22247 37077
rect 22370 37068 22376 37080
rect 22428 37108 22434 37120
rect 23290 37108 23296 37120
rect 22428 37080 23296 37108
rect 22428 37068 22434 37080
rect 23290 37068 23296 37080
rect 23348 37068 23354 37120
rect 25409 37111 25467 37117
rect 25409 37077 25421 37111
rect 25455 37108 25467 37111
rect 26694 37108 26700 37120
rect 25455 37080 26700 37108
rect 25455 37077 25467 37080
rect 25409 37071 25467 37077
rect 26694 37068 26700 37080
rect 26752 37068 26758 37120
rect 26786 37068 26792 37120
rect 26844 37108 26850 37120
rect 27801 37111 27859 37117
rect 27801 37108 27813 37111
rect 26844 37080 27813 37108
rect 26844 37068 26850 37080
rect 27801 37077 27813 37080
rect 27847 37077 27859 37111
rect 27801 37071 27859 37077
rect 28074 37068 28080 37120
rect 28132 37108 28138 37120
rect 28169 37111 28227 37117
rect 28169 37108 28181 37111
rect 28132 37080 28181 37108
rect 28132 37068 28138 37080
rect 28169 37077 28181 37080
rect 28215 37077 28227 37111
rect 28169 37071 28227 37077
rect 28261 37111 28319 37117
rect 28261 37077 28273 37111
rect 28307 37108 28319 37111
rect 30098 37108 30104 37120
rect 28307 37080 30104 37108
rect 28307 37077 28319 37080
rect 28261 37071 28319 37077
rect 30098 37068 30104 37080
rect 30156 37108 30162 37120
rect 30929 37111 30987 37117
rect 30929 37108 30941 37111
rect 30156 37080 30941 37108
rect 30156 37068 30162 37080
rect 30929 37077 30941 37080
rect 30975 37077 30987 37111
rect 31956 37108 31984 37148
rect 32214 37136 32220 37148
rect 32272 37136 32278 37188
rect 32417 37111 32475 37117
rect 32417 37108 32429 37111
rect 31956 37080 32429 37108
rect 30929 37071 30987 37077
rect 32417 37077 32429 37080
rect 32463 37077 32475 37111
rect 32582 37108 32588 37120
rect 32543 37080 32588 37108
rect 32417 37071 32475 37077
rect 32582 37068 32588 37080
rect 32640 37068 32646 37120
rect 1104 37018 48852 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 48852 37018
rect 1104 36944 48852 36966
rect 21450 36864 21456 36916
rect 21508 36904 21514 36916
rect 22189 36907 22247 36913
rect 22189 36904 22201 36907
rect 21508 36876 22201 36904
rect 21508 36864 21514 36876
rect 22189 36873 22201 36876
rect 22235 36873 22247 36907
rect 22189 36867 22247 36873
rect 24673 36907 24731 36913
rect 24673 36873 24685 36907
rect 24719 36904 24731 36907
rect 25130 36904 25136 36916
rect 24719 36876 25136 36904
rect 24719 36873 24731 36876
rect 24673 36867 24731 36873
rect 25130 36864 25136 36876
rect 25188 36864 25194 36916
rect 25222 36864 25228 36916
rect 25280 36904 25286 36916
rect 27338 36904 27344 36916
rect 25280 36876 27344 36904
rect 25280 36864 25286 36876
rect 27338 36864 27344 36876
rect 27396 36864 27402 36916
rect 27617 36907 27675 36913
rect 27617 36873 27629 36907
rect 27663 36904 27675 36907
rect 29178 36904 29184 36916
rect 27663 36876 28856 36904
rect 29139 36876 29184 36904
rect 27663 36873 27675 36876
rect 27617 36867 27675 36873
rect 2038 36796 2044 36848
rect 2096 36836 2102 36848
rect 24578 36836 24584 36848
rect 2096 36808 24584 36836
rect 2096 36796 2102 36808
rect 24578 36796 24584 36808
rect 24636 36796 24642 36848
rect 25038 36836 25044 36848
rect 24999 36808 25044 36836
rect 25038 36796 25044 36808
rect 25096 36796 25102 36848
rect 26053 36839 26111 36845
rect 26053 36805 26065 36839
rect 26099 36836 26111 36839
rect 26786 36836 26792 36848
rect 26099 36808 26792 36836
rect 26099 36805 26111 36808
rect 26053 36799 26111 36805
rect 26786 36796 26792 36808
rect 26844 36796 26850 36848
rect 28828 36845 28856 36876
rect 29178 36864 29184 36876
rect 29236 36864 29242 36916
rect 28813 36839 28871 36845
rect 27172 36808 28488 36836
rect 18138 36728 18144 36780
rect 18196 36768 18202 36780
rect 18305 36771 18363 36777
rect 18305 36768 18317 36771
rect 18196 36740 18317 36768
rect 18196 36728 18202 36740
rect 18305 36737 18317 36740
rect 18351 36737 18363 36771
rect 18305 36731 18363 36737
rect 20441 36771 20499 36777
rect 20441 36737 20453 36771
rect 20487 36737 20499 36771
rect 20441 36731 20499 36737
rect 18046 36700 18052 36712
rect 18007 36672 18052 36700
rect 18046 36660 18052 36672
rect 18104 36660 18110 36712
rect 20456 36700 20484 36731
rect 20530 36728 20536 36780
rect 20588 36768 20594 36780
rect 20625 36771 20683 36777
rect 20625 36768 20637 36771
rect 20588 36740 20637 36768
rect 20588 36728 20594 36740
rect 20625 36737 20637 36740
rect 20671 36737 20683 36771
rect 21818 36768 21824 36780
rect 21779 36740 21824 36768
rect 20625 36731 20683 36737
rect 21818 36728 21824 36740
rect 21876 36728 21882 36780
rect 21910 36728 21916 36780
rect 21968 36768 21974 36780
rect 22005 36771 22063 36777
rect 22005 36768 22017 36771
rect 21968 36740 22017 36768
rect 21968 36728 21974 36740
rect 22005 36737 22017 36740
rect 22051 36737 22063 36771
rect 22005 36731 22063 36737
rect 25133 36771 25191 36777
rect 25133 36737 25145 36771
rect 25179 36768 25191 36771
rect 26234 36768 26240 36780
rect 25179 36740 26096 36768
rect 26147 36740 26240 36768
rect 25179 36737 25191 36740
rect 25133 36731 25191 36737
rect 21266 36700 21272 36712
rect 20456 36672 21272 36700
rect 21266 36660 21272 36672
rect 21324 36660 21330 36712
rect 25317 36703 25375 36709
rect 25317 36669 25329 36703
rect 25363 36700 25375 36703
rect 25498 36700 25504 36712
rect 25363 36672 25504 36700
rect 25363 36669 25375 36672
rect 25317 36663 25375 36669
rect 25498 36660 25504 36672
rect 25556 36660 25562 36712
rect 26068 36700 26096 36740
rect 26234 36728 26240 36740
rect 26292 36768 26298 36780
rect 27172 36768 27200 36808
rect 27982 36768 27988 36780
rect 26292 36740 27200 36768
rect 27943 36740 27988 36768
rect 26292 36728 26298 36740
rect 27982 36728 27988 36740
rect 28040 36728 28046 36780
rect 28077 36771 28135 36777
rect 28077 36737 28089 36771
rect 28123 36768 28135 36771
rect 28258 36768 28264 36780
rect 28123 36740 28264 36768
rect 28123 36737 28135 36740
rect 28077 36731 28135 36737
rect 28258 36728 28264 36740
rect 28316 36728 28322 36780
rect 27890 36700 27896 36712
rect 26068 36672 27896 36700
rect 27890 36660 27896 36672
rect 27948 36660 27954 36712
rect 28169 36703 28227 36709
rect 28169 36669 28181 36703
rect 28215 36700 28227 36703
rect 28350 36700 28356 36712
rect 28215 36672 28356 36700
rect 28215 36669 28227 36672
rect 28169 36663 28227 36669
rect 27614 36592 27620 36644
rect 27672 36632 27678 36644
rect 28184 36632 28212 36663
rect 28350 36660 28356 36672
rect 28408 36660 28414 36712
rect 28460 36700 28488 36808
rect 28813 36805 28825 36839
rect 28859 36805 28871 36839
rect 28813 36799 28871 36805
rect 28997 36771 29055 36777
rect 28997 36737 29009 36771
rect 29043 36737 29055 36771
rect 28997 36731 29055 36737
rect 29012 36700 29040 36731
rect 29546 36728 29552 36780
rect 29604 36768 29610 36780
rect 30006 36777 30012 36780
rect 29733 36771 29791 36777
rect 29733 36768 29745 36771
rect 29604 36740 29745 36768
rect 29604 36728 29610 36740
rect 29733 36737 29745 36740
rect 29779 36737 29791 36771
rect 29733 36731 29791 36737
rect 30000 36731 30012 36777
rect 30064 36768 30070 36780
rect 30064 36740 30100 36768
rect 30006 36728 30012 36731
rect 30064 36728 30070 36740
rect 31938 36728 31944 36780
rect 31996 36768 32002 36780
rect 32381 36771 32439 36777
rect 32381 36768 32393 36771
rect 31996 36740 32393 36768
rect 31996 36728 32002 36740
rect 32381 36737 32393 36740
rect 32427 36737 32439 36771
rect 47578 36768 47584 36780
rect 47539 36740 47584 36768
rect 32381 36731 32439 36737
rect 47578 36728 47584 36740
rect 47636 36728 47642 36780
rect 32122 36700 32128 36712
rect 28460 36672 29040 36700
rect 32083 36672 32128 36700
rect 32122 36660 32128 36672
rect 32180 36660 32186 36712
rect 27672 36604 28212 36632
rect 27672 36592 27678 36604
rect 1946 36524 1952 36576
rect 2004 36564 2010 36576
rect 2225 36567 2283 36573
rect 2225 36564 2237 36567
rect 2004 36536 2237 36564
rect 2004 36524 2010 36536
rect 2225 36533 2237 36536
rect 2271 36533 2283 36567
rect 2225 36527 2283 36533
rect 19429 36567 19487 36573
rect 19429 36533 19441 36567
rect 19475 36564 19487 36567
rect 19978 36564 19984 36576
rect 19475 36536 19984 36564
rect 19475 36533 19487 36536
rect 19429 36527 19487 36533
rect 19978 36524 19984 36536
rect 20036 36524 20042 36576
rect 20806 36564 20812 36576
rect 20767 36536 20812 36564
rect 20806 36524 20812 36536
rect 20864 36524 20870 36576
rect 24946 36524 24952 36576
rect 25004 36564 25010 36576
rect 25222 36564 25228 36576
rect 25004 36536 25228 36564
rect 25004 36524 25010 36536
rect 25222 36524 25228 36536
rect 25280 36524 25286 36576
rect 26421 36567 26479 36573
rect 26421 36533 26433 36567
rect 26467 36564 26479 36567
rect 28350 36564 28356 36576
rect 26467 36536 28356 36564
rect 26467 36533 26479 36536
rect 26421 36527 26479 36533
rect 28350 36524 28356 36536
rect 28408 36524 28414 36576
rect 30374 36524 30380 36576
rect 30432 36564 30438 36576
rect 31113 36567 31171 36573
rect 31113 36564 31125 36567
rect 30432 36536 31125 36564
rect 30432 36524 30438 36536
rect 31113 36533 31125 36536
rect 31159 36533 31171 36567
rect 33502 36564 33508 36576
rect 33463 36536 33508 36564
rect 31113 36527 31171 36533
rect 33502 36524 33508 36536
rect 33560 36524 33566 36576
rect 46474 36524 46480 36576
rect 46532 36564 46538 36576
rect 47673 36567 47731 36573
rect 47673 36564 47685 36567
rect 46532 36536 47685 36564
rect 46532 36524 46538 36536
rect 47673 36533 47685 36536
rect 47719 36533 47731 36567
rect 47673 36527 47731 36533
rect 1104 36474 48852 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 48852 36474
rect 1104 36400 48852 36422
rect 21818 36320 21824 36372
rect 21876 36360 21882 36372
rect 22465 36363 22523 36369
rect 22465 36360 22477 36363
rect 21876 36332 22477 36360
rect 21876 36320 21882 36332
rect 22465 36329 22477 36332
rect 22511 36329 22523 36363
rect 22465 36323 22523 36329
rect 24578 36320 24584 36372
rect 24636 36360 24642 36372
rect 24636 36332 27752 36360
rect 24636 36320 24642 36332
rect 27724 36292 27752 36332
rect 27798 36320 27804 36372
rect 27856 36360 27862 36372
rect 27893 36363 27951 36369
rect 27893 36360 27905 36363
rect 27856 36332 27905 36360
rect 27856 36320 27862 36332
rect 27893 36329 27905 36332
rect 27939 36329 27951 36363
rect 29822 36360 29828 36372
rect 29783 36332 29828 36360
rect 27893 36323 27951 36329
rect 29822 36320 29828 36332
rect 29880 36320 29886 36372
rect 30190 36320 30196 36372
rect 30248 36360 30254 36372
rect 31205 36363 31263 36369
rect 31205 36360 31217 36363
rect 30248 36332 31217 36360
rect 30248 36320 30254 36332
rect 31205 36329 31217 36332
rect 31251 36329 31263 36363
rect 31938 36360 31944 36372
rect 31899 36332 31944 36360
rect 31205 36323 31263 36329
rect 31938 36320 31944 36332
rect 31996 36320 32002 36372
rect 30653 36295 30711 36301
rect 30653 36292 30665 36295
rect 18524 36264 19656 36292
rect 27724 36264 30665 36292
rect 2590 36184 2596 36236
rect 2648 36224 2654 36236
rect 2648 36196 6914 36224
rect 2648 36184 2654 36196
rect 2777 36159 2835 36165
rect 2777 36125 2789 36159
rect 2823 36156 2835 36159
rect 3418 36156 3424 36168
rect 2823 36128 3424 36156
rect 2823 36125 2835 36128
rect 2777 36119 2835 36125
rect 3418 36116 3424 36128
rect 3476 36116 3482 36168
rect 6886 36156 6914 36196
rect 18524 36165 18552 36264
rect 19628 36233 19656 36264
rect 30653 36261 30665 36264
rect 30699 36261 30711 36295
rect 30653 36255 30711 36261
rect 19613 36227 19671 36233
rect 19613 36193 19625 36227
rect 19659 36193 19671 36227
rect 20622 36224 20628 36236
rect 20583 36196 20628 36224
rect 19613 36187 19671 36193
rect 20622 36184 20628 36196
rect 20680 36184 20686 36236
rect 22462 36184 22468 36236
rect 22520 36224 22526 36236
rect 22646 36224 22652 36236
rect 22520 36196 22652 36224
rect 22520 36184 22526 36196
rect 22646 36184 22652 36196
rect 22704 36224 22710 36236
rect 23017 36227 23075 36233
rect 23017 36224 23029 36227
rect 22704 36196 23029 36224
rect 22704 36184 22710 36196
rect 23017 36193 23029 36196
rect 23063 36193 23075 36227
rect 24762 36224 24768 36236
rect 24723 36196 24768 36224
rect 23017 36187 23075 36193
rect 24762 36184 24768 36196
rect 24820 36184 24826 36236
rect 26881 36227 26939 36233
rect 26881 36224 26893 36227
rect 25976 36196 26893 36224
rect 18325 36159 18383 36165
rect 18325 36156 18337 36159
rect 6886 36128 18337 36156
rect 18325 36125 18337 36128
rect 18371 36125 18383 36159
rect 18325 36119 18383 36125
rect 18417 36159 18475 36165
rect 18417 36125 18429 36159
rect 18463 36125 18475 36159
rect 18417 36119 18475 36125
rect 18509 36159 18567 36165
rect 18509 36125 18521 36159
rect 18555 36125 18567 36159
rect 18509 36119 18567 36125
rect 18693 36159 18751 36165
rect 18693 36125 18705 36159
rect 18739 36156 18751 36159
rect 18739 36128 21036 36156
rect 18739 36125 18751 36128
rect 18693 36119 18751 36125
rect 18432 36088 18460 36119
rect 21008 36100 21036 36128
rect 24394 36116 24400 36168
rect 24452 36156 24458 36168
rect 25976 36156 26004 36196
rect 26881 36193 26893 36196
rect 26927 36224 26939 36227
rect 27246 36224 27252 36236
rect 26927 36196 27252 36224
rect 26927 36193 26939 36196
rect 26881 36187 26939 36193
rect 27246 36184 27252 36196
rect 27304 36224 27310 36236
rect 30098 36224 30104 36236
rect 27304 36196 28304 36224
rect 30059 36196 30104 36224
rect 27304 36184 27310 36196
rect 26602 36156 26608 36168
rect 24452 36128 26004 36156
rect 26563 36128 26608 36156
rect 24452 36116 24458 36128
rect 26602 36116 26608 36128
rect 26660 36116 26666 36168
rect 27890 36116 27896 36168
rect 27948 36156 27954 36168
rect 28276 36165 28304 36196
rect 30098 36184 30104 36196
rect 30156 36184 30162 36236
rect 30282 36224 30288 36236
rect 30243 36196 30288 36224
rect 30282 36184 30288 36196
rect 30340 36184 30346 36236
rect 28169 36159 28227 36165
rect 28169 36156 28181 36159
rect 27948 36128 28181 36156
rect 27948 36116 27954 36128
rect 28169 36125 28181 36128
rect 28215 36125 28227 36159
rect 28169 36119 28227 36125
rect 28261 36159 28319 36165
rect 28261 36125 28273 36159
rect 28307 36125 28319 36159
rect 28261 36119 28319 36125
rect 28350 36116 28356 36168
rect 28408 36156 28414 36168
rect 28408 36128 28453 36156
rect 28408 36116 28414 36128
rect 28534 36116 28540 36168
rect 28592 36156 28598 36168
rect 28592 36128 28637 36156
rect 28592 36116 28598 36128
rect 29914 36116 29920 36168
rect 29972 36156 29978 36168
rect 30009 36159 30067 36165
rect 30009 36156 30021 36159
rect 29972 36128 30021 36156
rect 29972 36116 29978 36128
rect 30009 36125 30021 36128
rect 30055 36125 30067 36159
rect 30009 36119 30067 36125
rect 30193 36159 30251 36165
rect 30193 36125 30205 36159
rect 30239 36156 30251 36159
rect 30558 36156 30564 36168
rect 30239 36128 30564 36156
rect 30239 36125 30251 36128
rect 30193 36119 30251 36125
rect 30558 36116 30564 36128
rect 30616 36116 30622 36168
rect 19150 36088 19156 36100
rect 18432 36060 19156 36088
rect 19150 36048 19156 36060
rect 19208 36048 19214 36100
rect 19245 36091 19303 36097
rect 19245 36057 19257 36091
rect 19291 36088 19303 36091
rect 19334 36088 19340 36100
rect 19291 36060 19340 36088
rect 19291 36057 19303 36060
rect 19245 36051 19303 36057
rect 19334 36048 19340 36060
rect 19392 36048 19398 36100
rect 19429 36091 19487 36097
rect 19429 36057 19441 36091
rect 19475 36057 19487 36091
rect 19429 36051 19487 36057
rect 2866 36020 2872 36032
rect 2827 35992 2872 36020
rect 2866 35980 2872 35992
rect 2924 35980 2930 36032
rect 18049 36023 18107 36029
rect 18049 35989 18061 36023
rect 18095 36020 18107 36023
rect 18230 36020 18236 36032
rect 18095 35992 18236 36020
rect 18095 35989 18107 35992
rect 18049 35983 18107 35989
rect 18230 35980 18236 35992
rect 18288 35980 18294 36032
rect 19444 36020 19472 36051
rect 20714 36048 20720 36100
rect 20772 36088 20778 36100
rect 20870 36091 20928 36097
rect 20870 36088 20882 36091
rect 20772 36060 20882 36088
rect 20772 36048 20778 36060
rect 20870 36057 20882 36060
rect 20916 36057 20928 36091
rect 20870 36051 20928 36057
rect 20990 36048 20996 36100
rect 21048 36048 21054 36100
rect 24854 36048 24860 36100
rect 24912 36088 24918 36100
rect 25010 36091 25068 36097
rect 25010 36088 25022 36091
rect 24912 36060 25022 36088
rect 24912 36048 24918 36060
rect 25010 36057 25022 36060
rect 25056 36057 25068 36091
rect 30668 36088 30696 36255
rect 30834 36252 30840 36304
rect 30892 36292 30898 36304
rect 47670 36292 47676 36304
rect 30892 36264 32720 36292
rect 30892 36252 30898 36264
rect 31662 36184 31668 36236
rect 31720 36224 31726 36236
rect 32309 36227 32367 36233
rect 32309 36224 32321 36227
rect 31720 36196 32321 36224
rect 31720 36184 31726 36196
rect 32309 36193 32321 36196
rect 32355 36193 32367 36227
rect 32309 36187 32367 36193
rect 32401 36227 32459 36233
rect 32401 36193 32413 36227
rect 32447 36224 32459 36227
rect 32582 36224 32588 36236
rect 32447 36196 32588 36224
rect 32447 36193 32459 36196
rect 32401 36187 32459 36193
rect 32582 36184 32588 36196
rect 32640 36184 32646 36236
rect 32030 36116 32036 36168
rect 32088 36156 32094 36168
rect 32125 36159 32183 36165
rect 32125 36156 32137 36159
rect 32088 36128 32137 36156
rect 32088 36116 32094 36128
rect 32125 36125 32137 36128
rect 32171 36125 32183 36159
rect 32125 36119 32183 36125
rect 32217 36159 32275 36165
rect 32217 36125 32229 36159
rect 32263 36156 32275 36159
rect 32692 36156 32720 36264
rect 46308 36264 47676 36292
rect 46308 36233 46336 36264
rect 47670 36252 47676 36264
rect 47728 36252 47734 36304
rect 46293 36227 46351 36233
rect 46293 36193 46305 36227
rect 46339 36193 46351 36227
rect 46474 36224 46480 36236
rect 46435 36196 46480 36224
rect 46293 36187 46351 36193
rect 46474 36184 46480 36196
rect 46532 36184 46538 36236
rect 48130 36224 48136 36236
rect 48091 36196 48136 36224
rect 48130 36184 48136 36196
rect 48188 36184 48194 36236
rect 33502 36156 33508 36168
rect 32263 36128 33508 36156
rect 32263 36125 32275 36128
rect 32217 36119 32275 36125
rect 33502 36116 33508 36128
rect 33560 36116 33566 36168
rect 31021 36091 31079 36097
rect 31021 36088 31033 36091
rect 30668 36060 31033 36088
rect 25010 36051 25068 36057
rect 31021 36057 31033 36060
rect 31067 36057 31079 36091
rect 31021 36051 31079 36057
rect 31110 36048 31116 36100
rect 31168 36088 31174 36100
rect 31221 36091 31279 36097
rect 31221 36088 31233 36091
rect 31168 36060 31233 36088
rect 31168 36048 31174 36060
rect 31221 36057 31233 36060
rect 31267 36057 31279 36091
rect 31221 36051 31279 36057
rect 21450 36020 21456 36032
rect 19444 35992 21456 36020
rect 21450 35980 21456 35992
rect 21508 36020 21514 36032
rect 21910 36020 21916 36032
rect 21508 35992 21916 36020
rect 21508 35980 21514 35992
rect 21910 35980 21916 35992
rect 21968 35980 21974 36032
rect 22005 36023 22063 36029
rect 22005 35989 22017 36023
rect 22051 36020 22063 36023
rect 22462 36020 22468 36032
rect 22051 35992 22468 36020
rect 22051 35989 22063 35992
rect 22005 35983 22063 35989
rect 22462 35980 22468 35992
rect 22520 35980 22526 36032
rect 22738 35980 22744 36032
rect 22796 36020 22802 36032
rect 22833 36023 22891 36029
rect 22833 36020 22845 36023
rect 22796 35992 22845 36020
rect 22796 35980 22802 35992
rect 22833 35989 22845 35992
rect 22879 35989 22891 36023
rect 22833 35983 22891 35989
rect 22925 36023 22983 36029
rect 22925 35989 22937 36023
rect 22971 36020 22983 36023
rect 23566 36020 23572 36032
rect 22971 35992 23572 36020
rect 22971 35989 22983 35992
rect 22925 35983 22983 35989
rect 23566 35980 23572 35992
rect 23624 35980 23630 36032
rect 25314 35980 25320 36032
rect 25372 36020 25378 36032
rect 26145 36023 26203 36029
rect 26145 36020 26157 36023
rect 25372 35992 26157 36020
rect 25372 35980 25378 35992
rect 26145 35989 26157 35992
rect 26191 36020 26203 36023
rect 27338 36020 27344 36032
rect 26191 35992 27344 36020
rect 26191 35989 26203 35992
rect 26145 35983 26203 35989
rect 27338 35980 27344 35992
rect 27396 35980 27402 36032
rect 28258 35980 28264 36032
rect 28316 36020 28322 36032
rect 30834 36020 30840 36032
rect 28316 35992 30840 36020
rect 28316 35980 28322 35992
rect 30834 35980 30840 35992
rect 30892 35980 30898 36032
rect 31386 36020 31392 36032
rect 31347 35992 31392 36020
rect 31386 35980 31392 35992
rect 31444 35980 31450 36032
rect 1104 35930 48852 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 48852 35930
rect 1104 35856 48852 35878
rect 20073 35819 20131 35825
rect 20073 35785 20085 35819
rect 20119 35816 20131 35819
rect 20714 35816 20720 35828
rect 20119 35788 20720 35816
rect 20119 35785 20131 35788
rect 20073 35779 20131 35785
rect 20714 35776 20720 35788
rect 20772 35776 20778 35828
rect 21266 35776 21272 35828
rect 21324 35816 21330 35828
rect 22097 35819 22155 35825
rect 22097 35816 22109 35819
rect 21324 35788 22109 35816
rect 21324 35776 21330 35788
rect 22097 35785 22109 35788
rect 22143 35785 22155 35819
rect 22097 35779 22155 35785
rect 24581 35819 24639 35825
rect 24581 35785 24593 35819
rect 24627 35816 24639 35819
rect 24854 35816 24860 35828
rect 24627 35788 24860 35816
rect 24627 35785 24639 35788
rect 24581 35779 24639 35785
rect 24854 35776 24860 35788
rect 24912 35776 24918 35828
rect 25038 35776 25044 35828
rect 25096 35776 25102 35828
rect 26973 35819 27031 35825
rect 26973 35785 26985 35819
rect 27019 35785 27031 35819
rect 26973 35779 27031 35785
rect 2133 35751 2191 35757
rect 2133 35717 2145 35751
rect 2179 35748 2191 35751
rect 2866 35748 2872 35760
rect 2179 35720 2872 35748
rect 2179 35717 2191 35720
rect 2133 35711 2191 35717
rect 2866 35708 2872 35720
rect 2924 35708 2930 35760
rect 18046 35708 18052 35760
rect 18104 35748 18110 35760
rect 19702 35748 19708 35760
rect 18104 35720 19708 35748
rect 18104 35708 18110 35720
rect 1946 35680 1952 35692
rect 1907 35652 1952 35680
rect 1946 35640 1952 35652
rect 2004 35640 2010 35692
rect 18156 35689 18184 35720
rect 19702 35708 19708 35720
rect 19760 35708 19766 35760
rect 20806 35748 20812 35760
rect 20548 35720 20812 35748
rect 18141 35683 18199 35689
rect 18141 35649 18153 35683
rect 18187 35649 18199 35683
rect 18141 35643 18199 35649
rect 18230 35640 18236 35692
rect 18288 35680 18294 35692
rect 18397 35683 18455 35689
rect 18397 35680 18409 35683
rect 18288 35652 18409 35680
rect 18288 35640 18294 35652
rect 18397 35649 18409 35652
rect 18443 35649 18455 35683
rect 18397 35643 18455 35649
rect 20254 35640 20260 35692
rect 20312 35689 20318 35692
rect 20548 35689 20576 35720
rect 20806 35708 20812 35720
rect 20864 35708 20870 35760
rect 22557 35751 22615 35757
rect 22557 35717 22569 35751
rect 22603 35748 22615 35751
rect 25056 35748 25084 35776
rect 22603 35720 25084 35748
rect 26053 35751 26111 35757
rect 22603 35717 22615 35720
rect 22557 35711 22615 35717
rect 26053 35717 26065 35751
rect 26099 35748 26111 35751
rect 26988 35748 27016 35779
rect 27062 35776 27068 35828
rect 27120 35816 27126 35828
rect 27120 35788 29316 35816
rect 27120 35776 27126 35788
rect 27614 35748 27620 35760
rect 26099 35720 27016 35748
rect 27264 35720 27620 35748
rect 26099 35717 26111 35720
rect 26053 35711 26111 35717
rect 20312 35683 20361 35689
rect 20312 35649 20315 35683
rect 20349 35649 20361 35683
rect 20312 35643 20361 35649
rect 20422 35683 20480 35689
rect 20422 35649 20434 35683
rect 20468 35649 20480 35683
rect 20422 35643 20480 35649
rect 20533 35683 20591 35689
rect 20533 35649 20545 35683
rect 20579 35649 20591 35683
rect 20533 35643 20591 35649
rect 20717 35683 20775 35689
rect 20717 35649 20729 35683
rect 20763 35680 20775 35683
rect 20990 35680 20996 35692
rect 20763 35652 20996 35680
rect 20763 35649 20775 35652
rect 20717 35643 20775 35649
rect 20312 35640 20318 35643
rect 2774 35612 2780 35624
rect 2735 35584 2780 35612
rect 2774 35572 2780 35584
rect 2832 35572 2838 35624
rect 19150 35572 19156 35624
rect 19208 35612 19214 35624
rect 19610 35612 19616 35624
rect 19208 35584 19616 35612
rect 19208 35572 19214 35584
rect 19610 35572 19616 35584
rect 19668 35612 19674 35624
rect 20437 35612 20465 35643
rect 20990 35640 20996 35652
rect 21048 35640 21054 35692
rect 22462 35680 22468 35692
rect 22375 35652 22468 35680
rect 22462 35640 22468 35652
rect 22520 35680 22526 35692
rect 22830 35680 22836 35692
rect 22520 35652 22836 35680
rect 22520 35640 22526 35652
rect 22830 35640 22836 35652
rect 22888 35640 22894 35692
rect 23385 35683 23443 35689
rect 23385 35649 23397 35683
rect 23431 35680 23443 35683
rect 24210 35680 24216 35692
rect 23431 35652 24216 35680
rect 23431 35649 23443 35652
rect 23385 35643 23443 35649
rect 24210 35640 24216 35652
rect 24268 35640 24274 35692
rect 24302 35640 24308 35692
rect 24360 35680 24366 35692
rect 24857 35683 24915 35689
rect 24857 35680 24869 35683
rect 24360 35652 24869 35680
rect 24360 35640 24366 35652
rect 24857 35649 24869 35652
rect 24903 35649 24915 35683
rect 24857 35643 24915 35649
rect 24949 35683 25007 35689
rect 24949 35649 24961 35683
rect 24995 35649 25007 35683
rect 24949 35643 25007 35649
rect 25041 35683 25099 35689
rect 25041 35649 25053 35683
rect 25087 35649 25099 35683
rect 25222 35680 25228 35692
rect 25183 35652 25228 35680
rect 25041 35643 25099 35649
rect 19668 35584 20465 35612
rect 19668 35572 19674 35584
rect 22646 35572 22652 35624
rect 22704 35612 22710 35624
rect 23569 35615 23627 35621
rect 23569 35612 23581 35615
rect 22704 35584 23581 35612
rect 22704 35572 22710 35584
rect 23569 35581 23581 35584
rect 23615 35581 23627 35615
rect 23569 35575 23627 35581
rect 24394 35572 24400 35624
rect 24452 35612 24458 35624
rect 24964 35612 24992 35643
rect 24452 35584 24992 35612
rect 25056 35612 25084 35643
rect 25222 35640 25228 35652
rect 25280 35640 25286 35692
rect 26234 35680 26240 35692
rect 26195 35652 26240 35680
rect 26234 35640 26240 35652
rect 26292 35640 26298 35692
rect 27264 35680 27292 35720
rect 26712 35652 27292 35680
rect 26421 35615 26479 35621
rect 26421 35612 26433 35615
rect 25056 35584 26433 35612
rect 24452 35572 24458 35584
rect 26421 35581 26433 35584
rect 26467 35581 26479 35615
rect 26421 35575 26479 35581
rect 20070 35504 20076 35556
rect 20128 35544 20134 35556
rect 22664 35544 22692 35572
rect 20128 35516 22692 35544
rect 20128 35504 20134 35516
rect 25498 35504 25504 35556
rect 25556 35544 25562 35556
rect 26712 35544 26740 35652
rect 27338 35640 27344 35692
rect 27396 35680 27402 35692
rect 27396 35652 27441 35680
rect 27396 35640 27402 35652
rect 27540 35621 27568 35720
rect 27614 35708 27620 35720
rect 27672 35708 27678 35760
rect 27706 35708 27712 35760
rect 27764 35748 27770 35760
rect 28445 35751 28503 35757
rect 28445 35748 28457 35751
rect 27764 35720 28457 35748
rect 27764 35708 27770 35720
rect 28445 35717 28457 35720
rect 28491 35748 28503 35751
rect 28534 35748 28540 35760
rect 28491 35720 28540 35748
rect 28491 35717 28503 35720
rect 28445 35711 28503 35717
rect 28534 35708 28540 35720
rect 28592 35708 28598 35760
rect 28166 35640 28172 35692
rect 28224 35680 28230 35692
rect 28261 35683 28319 35689
rect 28261 35680 28273 35683
rect 28224 35652 28273 35680
rect 28224 35640 28230 35652
rect 28261 35649 28273 35652
rect 28307 35649 28319 35683
rect 28994 35680 29000 35692
rect 28955 35652 29000 35680
rect 28261 35643 28319 35649
rect 28994 35640 29000 35652
rect 29052 35640 29058 35692
rect 29288 35689 29316 35788
rect 30006 35776 30012 35828
rect 30064 35816 30070 35828
rect 30101 35819 30159 35825
rect 30101 35816 30113 35819
rect 30064 35788 30113 35816
rect 30064 35776 30070 35788
rect 30101 35785 30113 35788
rect 30147 35785 30159 35819
rect 30101 35779 30159 35785
rect 29914 35708 29920 35760
rect 29972 35748 29978 35760
rect 32030 35748 32036 35760
rect 29972 35720 32036 35748
rect 29972 35708 29978 35720
rect 29273 35683 29331 35689
rect 29273 35649 29285 35683
rect 29319 35680 29331 35683
rect 29362 35680 29368 35692
rect 29319 35652 29368 35680
rect 29319 35649 29331 35652
rect 29273 35643 29331 35649
rect 29362 35640 29368 35652
rect 29420 35640 29426 35692
rect 30208 35680 30236 35720
rect 32030 35708 32036 35720
rect 32088 35708 32094 35760
rect 47946 35748 47952 35760
rect 47907 35720 47952 35748
rect 47946 35708 47952 35720
rect 48004 35708 48010 35760
rect 30285 35683 30343 35689
rect 30285 35680 30297 35683
rect 30208 35652 30297 35680
rect 30285 35649 30297 35652
rect 30331 35649 30343 35683
rect 30285 35643 30343 35649
rect 30374 35640 30380 35692
rect 30432 35680 30438 35692
rect 30561 35683 30619 35689
rect 30432 35652 30477 35680
rect 30432 35640 30438 35652
rect 30561 35649 30573 35683
rect 30607 35680 30619 35683
rect 31386 35680 31392 35692
rect 30607 35652 31392 35680
rect 30607 35649 30619 35652
rect 30561 35643 30619 35649
rect 31386 35640 31392 35652
rect 31444 35640 31450 35692
rect 32214 35640 32220 35692
rect 32272 35680 32278 35692
rect 32381 35683 32439 35689
rect 32381 35680 32393 35683
rect 32272 35652 32393 35680
rect 32272 35640 32278 35652
rect 32381 35649 32393 35652
rect 32427 35649 32439 35683
rect 32381 35643 32439 35649
rect 45646 35640 45652 35692
rect 45704 35680 45710 35692
rect 46753 35683 46811 35689
rect 46753 35680 46765 35683
rect 45704 35652 46765 35680
rect 45704 35640 45710 35652
rect 46753 35649 46765 35652
rect 46799 35649 46811 35683
rect 46753 35643 46811 35649
rect 27433 35615 27491 35621
rect 27433 35581 27445 35615
rect 27479 35581 27491 35615
rect 27433 35575 27491 35581
rect 27525 35615 27583 35621
rect 27525 35581 27537 35615
rect 27571 35581 27583 35615
rect 27525 35575 27583 35581
rect 29181 35615 29239 35621
rect 29181 35581 29193 35615
rect 29227 35612 29239 35615
rect 30098 35612 30104 35624
rect 29227 35584 30104 35612
rect 29227 35581 29239 35584
rect 29181 35575 29239 35581
rect 25556 35516 26740 35544
rect 27448 35544 27476 35575
rect 30098 35572 30104 35584
rect 30156 35572 30162 35624
rect 30392 35544 30420 35640
rect 30469 35615 30527 35621
rect 30469 35581 30481 35615
rect 30515 35581 30527 35615
rect 32122 35612 32128 35624
rect 32083 35584 32128 35612
rect 30469 35575 30527 35581
rect 27448 35516 30420 35544
rect 30484 35544 30512 35575
rect 32122 35572 32128 35584
rect 32180 35572 32186 35624
rect 30558 35544 30564 35556
rect 30484 35516 30564 35544
rect 25556 35504 25562 35516
rect 19518 35476 19524 35488
rect 19479 35448 19524 35476
rect 19518 35436 19524 35448
rect 19576 35436 19582 35488
rect 19702 35436 19708 35488
rect 19760 35476 19766 35488
rect 20622 35476 20628 35488
rect 19760 35448 20628 35476
rect 19760 35436 19766 35448
rect 20622 35436 20628 35448
rect 20680 35436 20686 35488
rect 29288 35485 29316 35516
rect 30558 35504 30564 35516
rect 30616 35504 30622 35556
rect 45830 35504 45836 35556
rect 45888 35544 45894 35556
rect 48133 35547 48191 35553
rect 48133 35544 48145 35547
rect 45888 35516 48145 35544
rect 45888 35504 45894 35516
rect 48133 35513 48145 35516
rect 48179 35513 48191 35547
rect 48133 35507 48191 35513
rect 29273 35479 29331 35485
rect 29273 35445 29285 35479
rect 29319 35445 29331 35479
rect 29454 35476 29460 35488
rect 29415 35448 29460 35476
rect 29273 35439 29331 35445
rect 29454 35436 29460 35448
rect 29512 35436 29518 35488
rect 33502 35476 33508 35488
rect 33463 35448 33508 35476
rect 33502 35436 33508 35448
rect 33560 35436 33566 35488
rect 46290 35476 46296 35488
rect 46251 35448 46296 35476
rect 46290 35436 46296 35448
rect 46348 35436 46354 35488
rect 46474 35436 46480 35488
rect 46532 35476 46538 35488
rect 46845 35479 46903 35485
rect 46845 35476 46857 35479
rect 46532 35448 46857 35476
rect 46532 35436 46538 35448
rect 46845 35445 46857 35448
rect 46891 35445 46903 35479
rect 46845 35439 46903 35445
rect 1104 35386 48852 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 48852 35386
rect 1104 35312 48852 35334
rect 19334 35232 19340 35284
rect 19392 35272 19398 35284
rect 19429 35275 19487 35281
rect 19429 35272 19441 35275
rect 19392 35244 19441 35272
rect 19392 35232 19398 35244
rect 19429 35241 19441 35244
rect 19475 35241 19487 35275
rect 20990 35272 20996 35284
rect 20951 35244 20996 35272
rect 19429 35235 19487 35241
rect 20990 35232 20996 35244
rect 21048 35232 21054 35284
rect 24673 35275 24731 35281
rect 24673 35241 24685 35275
rect 24719 35272 24731 35275
rect 25038 35272 25044 35284
rect 24719 35244 25044 35272
rect 24719 35241 24731 35244
rect 24673 35235 24731 35241
rect 25038 35232 25044 35244
rect 25096 35232 25102 35284
rect 25498 35272 25504 35284
rect 25459 35244 25504 35272
rect 25498 35232 25504 35244
rect 25556 35232 25562 35284
rect 29454 35232 29460 35284
rect 29512 35272 29518 35284
rect 29549 35275 29607 35281
rect 29549 35272 29561 35275
rect 29512 35244 29561 35272
rect 29512 35232 29518 35244
rect 29549 35241 29561 35244
rect 29595 35241 29607 35275
rect 29549 35235 29607 35241
rect 30282 35232 30288 35284
rect 30340 35272 30346 35284
rect 30561 35275 30619 35281
rect 30561 35272 30573 35275
rect 30340 35244 30573 35272
rect 30340 35232 30346 35244
rect 30561 35241 30573 35244
rect 30607 35241 30619 35275
rect 30561 35235 30619 35241
rect 31941 35275 31999 35281
rect 31941 35241 31953 35275
rect 31987 35272 31999 35275
rect 32214 35272 32220 35284
rect 31987 35244 32220 35272
rect 31987 35241 31999 35244
rect 31941 35235 31999 35241
rect 32214 35232 32220 35244
rect 32272 35232 32278 35284
rect 1762 35164 1768 35216
rect 1820 35204 1826 35216
rect 2590 35204 2596 35216
rect 1820 35176 2596 35204
rect 1820 35164 1826 35176
rect 2590 35164 2596 35176
rect 2648 35164 2654 35216
rect 19610 35164 19616 35216
rect 19668 35204 19674 35216
rect 21821 35207 21879 35213
rect 21821 35204 21833 35207
rect 19668 35176 21833 35204
rect 19668 35164 19674 35176
rect 21821 35173 21833 35176
rect 21867 35173 21879 35207
rect 21821 35167 21879 35173
rect 24210 35164 24216 35216
rect 24268 35204 24274 35216
rect 24268 35176 25452 35204
rect 24268 35164 24274 35176
rect 2041 35139 2099 35145
rect 2041 35105 2053 35139
rect 2087 35136 2099 35139
rect 20070 35136 20076 35148
rect 2087 35108 6914 35136
rect 20031 35108 20076 35136
rect 2087 35105 2099 35108
rect 2041 35099 2099 35105
rect 1762 35028 1768 35080
rect 1820 35068 1826 35080
rect 2685 35071 2743 35077
rect 2685 35068 2697 35071
rect 1820 35040 2697 35068
rect 1820 35028 1826 35040
rect 2685 35037 2697 35040
rect 2731 35037 2743 35071
rect 6886 35068 6914 35108
rect 20070 35096 20076 35108
rect 20128 35096 20134 35148
rect 24486 35136 24492 35148
rect 24447 35108 24492 35136
rect 24486 35096 24492 35108
rect 24544 35096 24550 35148
rect 24302 35068 24308 35080
rect 6886 35040 24308 35068
rect 2685 35031 2743 35037
rect 24302 35028 24308 35040
rect 24360 35028 24366 35080
rect 24670 35068 24676 35080
rect 24631 35040 24676 35068
rect 24670 35028 24676 35040
rect 24728 35028 24734 35080
rect 25424 35077 25452 35176
rect 29362 35164 29368 35216
rect 29420 35204 29426 35216
rect 29420 35176 31754 35204
rect 29420 35164 29426 35176
rect 31110 35136 31116 35148
rect 30576 35108 31116 35136
rect 25409 35071 25467 35077
rect 25409 35037 25421 35071
rect 25455 35037 25467 35071
rect 25409 35031 25467 35037
rect 28718 35028 28724 35080
rect 28776 35068 28782 35080
rect 29549 35071 29607 35077
rect 29549 35068 29561 35071
rect 28776 35040 29561 35068
rect 28776 35028 28782 35040
rect 29549 35037 29561 35040
rect 29595 35037 29607 35071
rect 29549 35031 29607 35037
rect 29733 35071 29791 35077
rect 29733 35037 29745 35071
rect 29779 35068 29791 35071
rect 30466 35068 30472 35080
rect 29779 35040 30472 35068
rect 29779 35037 29791 35040
rect 29733 35031 29791 35037
rect 30466 35028 30472 35040
rect 30524 35028 30530 35080
rect 1854 35000 1860 35012
rect 1815 34972 1860 35000
rect 1854 34960 1860 34972
rect 1912 34960 1918 35012
rect 19518 34960 19524 35012
rect 19576 35000 19582 35012
rect 19797 35003 19855 35009
rect 19797 35000 19809 35003
rect 19576 34972 19809 35000
rect 19576 34960 19582 34972
rect 19797 34969 19809 34972
rect 19843 35000 19855 35003
rect 20898 35000 20904 35012
rect 19843 34972 20208 35000
rect 20859 34972 20904 35000
rect 19843 34969 19855 34972
rect 19797 34963 19855 34969
rect 19889 34935 19947 34941
rect 19889 34901 19901 34935
rect 19935 34932 19947 34935
rect 20070 34932 20076 34944
rect 19935 34904 20076 34932
rect 19935 34901 19947 34904
rect 19889 34895 19947 34901
rect 20070 34892 20076 34904
rect 20128 34892 20134 34944
rect 20180 34932 20208 34972
rect 20898 34960 20904 34972
rect 20956 34960 20962 35012
rect 21637 35003 21695 35009
rect 21637 34969 21649 35003
rect 21683 35000 21695 35003
rect 22646 35000 22652 35012
rect 21683 34972 22652 35000
rect 21683 34969 21695 34972
rect 21637 34963 21695 34969
rect 22646 34960 22652 34972
rect 22704 34960 22710 35012
rect 24118 34960 24124 35012
rect 24176 35000 24182 35012
rect 30576 35009 30604 35108
rect 31110 35096 31116 35108
rect 31168 35096 31174 35148
rect 31726 35136 31754 35176
rect 32217 35139 32275 35145
rect 32217 35136 32229 35139
rect 31726 35108 32229 35136
rect 32217 35105 32229 35108
rect 32263 35136 32275 35139
rect 33502 35136 33508 35148
rect 32263 35108 33508 35136
rect 32263 35105 32275 35108
rect 32217 35099 32275 35105
rect 33502 35096 33508 35108
rect 33560 35096 33566 35148
rect 46290 35136 46296 35148
rect 46251 35108 46296 35136
rect 46290 35096 46296 35108
rect 46348 35096 46354 35148
rect 46474 35136 46480 35148
rect 46435 35108 46480 35136
rect 46474 35096 46480 35108
rect 46532 35096 46538 35148
rect 48130 35136 48136 35148
rect 48091 35108 48136 35136
rect 48130 35096 48136 35108
rect 48188 35096 48194 35148
rect 30742 35028 30748 35080
rect 30800 35028 30806 35080
rect 31570 35028 31576 35080
rect 31628 35068 31634 35080
rect 32030 35068 32036 35080
rect 31628 35040 32036 35068
rect 31628 35028 31634 35040
rect 32030 35028 32036 35040
rect 32088 35068 32094 35080
rect 32125 35071 32183 35077
rect 32125 35068 32137 35071
rect 32088 35040 32137 35068
rect 32088 35028 32094 35040
rect 32125 35037 32137 35040
rect 32171 35037 32183 35071
rect 32125 35031 32183 35037
rect 32309 35071 32367 35077
rect 32309 35037 32321 35071
rect 32355 35037 32367 35071
rect 32309 35031 32367 35037
rect 32401 35071 32459 35077
rect 32401 35037 32413 35071
rect 32447 35068 32459 35071
rect 32674 35068 32680 35080
rect 32447 35040 32680 35068
rect 32447 35037 32459 35040
rect 32401 35031 32459 35037
rect 24397 35003 24455 35009
rect 24397 35000 24409 35003
rect 24176 34972 24409 35000
rect 24176 34960 24182 34972
rect 24397 34969 24409 34972
rect 24443 34969 24455 35003
rect 24397 34963 24455 34969
rect 30377 35003 30435 35009
rect 30377 34969 30389 35003
rect 30423 34969 30435 35003
rect 30576 35003 30635 35009
rect 30576 34972 30589 35003
rect 30377 34963 30435 34969
rect 30577 34969 30589 34972
rect 30623 34969 30635 35003
rect 30760 35000 30788 35028
rect 30577 34963 30635 34969
rect 30668 34972 30788 35000
rect 21266 34932 21272 34944
rect 20180 34904 21272 34932
rect 21266 34892 21272 34904
rect 21324 34892 21330 34944
rect 24854 34932 24860 34944
rect 24815 34904 24860 34932
rect 24854 34892 24860 34904
rect 24912 34892 24918 34944
rect 25590 34892 25596 34944
rect 25648 34932 25654 34944
rect 29917 34935 29975 34941
rect 29917 34932 29929 34935
rect 25648 34904 29929 34932
rect 25648 34892 25654 34904
rect 29917 34901 29929 34904
rect 29963 34901 29975 34935
rect 30392 34932 30420 34963
rect 30668 34932 30696 34972
rect 30834 34960 30840 35012
rect 30892 35000 30898 35012
rect 31662 35000 31668 35012
rect 30892 34972 31668 35000
rect 30892 34960 30898 34972
rect 31662 34960 31668 34972
rect 31720 35000 31726 35012
rect 32324 35000 32352 35031
rect 32674 35028 32680 35040
rect 32732 35028 32738 35080
rect 31720 34972 32352 35000
rect 31720 34960 31726 34972
rect 30392 34904 30696 34932
rect 30745 34935 30803 34941
rect 29917 34895 29975 34901
rect 30745 34901 30757 34935
rect 30791 34932 30803 34935
rect 31202 34932 31208 34944
rect 30791 34904 31208 34932
rect 30791 34901 30803 34904
rect 30745 34895 30803 34901
rect 31202 34892 31208 34904
rect 31260 34892 31266 34944
rect 1104 34842 48852 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 48852 34842
rect 1104 34768 48852 34790
rect 23566 34728 23572 34740
rect 23527 34700 23572 34728
rect 23566 34688 23572 34700
rect 23624 34728 23630 34740
rect 24397 34731 24455 34737
rect 24397 34728 24409 34731
rect 23624 34700 24409 34728
rect 23624 34688 23630 34700
rect 24397 34697 24409 34700
rect 24443 34728 24455 34731
rect 24486 34728 24492 34740
rect 24443 34700 24492 34728
rect 24443 34697 24455 34700
rect 24397 34691 24455 34697
rect 24486 34688 24492 34700
rect 24544 34688 24550 34740
rect 28718 34728 28724 34740
rect 28679 34700 28724 34728
rect 28718 34688 28724 34700
rect 28776 34688 28782 34740
rect 31110 34688 31116 34740
rect 31168 34728 31174 34740
rect 32030 34728 32036 34740
rect 31168 34700 32036 34728
rect 31168 34688 31174 34700
rect 32030 34688 32036 34700
rect 32088 34728 32094 34740
rect 32509 34731 32567 34737
rect 32509 34728 32521 34731
rect 32088 34700 32521 34728
rect 32088 34688 32094 34700
rect 32509 34697 32521 34700
rect 32555 34697 32567 34731
rect 32674 34728 32680 34740
rect 32635 34700 32680 34728
rect 32509 34691 32567 34697
rect 32674 34688 32680 34700
rect 32732 34688 32738 34740
rect 1949 34663 2007 34669
rect 1949 34629 1961 34663
rect 1995 34660 2007 34663
rect 2406 34660 2412 34672
rect 1995 34632 2412 34660
rect 1995 34629 2007 34632
rect 1949 34623 2007 34629
rect 2406 34620 2412 34632
rect 2464 34620 2470 34672
rect 24762 34660 24768 34672
rect 22204 34632 24768 34660
rect 1762 34592 1768 34604
rect 1723 34564 1768 34592
rect 1762 34552 1768 34564
rect 1820 34552 1826 34604
rect 19426 34552 19432 34604
rect 19484 34592 19490 34604
rect 19705 34595 19763 34601
rect 19705 34592 19717 34595
rect 19484 34564 19717 34592
rect 19484 34552 19490 34564
rect 19705 34561 19717 34564
rect 19751 34561 19763 34595
rect 20346 34592 20352 34604
rect 20307 34564 20352 34592
rect 19705 34555 19763 34561
rect 2774 34524 2780 34536
rect 2735 34496 2780 34524
rect 2774 34484 2780 34496
rect 2832 34484 2838 34536
rect 19720 34456 19748 34555
rect 20346 34552 20352 34564
rect 20404 34552 20410 34604
rect 20530 34552 20536 34604
rect 20588 34592 20594 34604
rect 22204 34601 22232 34632
rect 24762 34620 24768 34632
rect 24820 34620 24826 34672
rect 25332 34632 27752 34660
rect 22462 34601 22468 34604
rect 22189 34595 22247 34601
rect 20588 34564 20681 34592
rect 20588 34552 20594 34564
rect 20640 34536 20668 34564
rect 22189 34561 22201 34595
rect 22235 34561 22247 34595
rect 22189 34555 22247 34561
rect 22456 34555 22468 34601
rect 22520 34592 22526 34604
rect 24489 34595 24547 34601
rect 22520 34564 22556 34592
rect 22462 34552 22468 34555
rect 22520 34552 22526 34564
rect 24489 34561 24501 34595
rect 24535 34592 24547 34595
rect 25332 34592 25360 34632
rect 24535 34564 25360 34592
rect 24535 34561 24547 34564
rect 24489 34555 24547 34561
rect 25406 34552 25412 34604
rect 25464 34592 25470 34604
rect 25501 34595 25559 34601
rect 25501 34592 25513 34595
rect 25464 34564 25513 34592
rect 25464 34552 25470 34564
rect 25501 34561 25513 34564
rect 25547 34561 25559 34595
rect 25774 34592 25780 34604
rect 25735 34564 25780 34592
rect 25501 34555 25559 34561
rect 25774 34552 25780 34564
rect 25832 34552 25838 34604
rect 20622 34484 20628 34536
rect 20680 34484 20686 34536
rect 20717 34527 20775 34533
rect 20717 34493 20729 34527
rect 20763 34524 20775 34527
rect 24578 34524 24584 34536
rect 20763 34496 22232 34524
rect 24539 34496 24584 34524
rect 20763 34493 20775 34496
rect 20717 34487 20775 34493
rect 22204 34468 22232 34496
rect 24578 34484 24584 34496
rect 24636 34484 24642 34536
rect 25222 34484 25228 34536
rect 25280 34524 25286 34536
rect 25593 34527 25651 34533
rect 25593 34524 25605 34527
rect 25280 34496 25605 34524
rect 25280 34484 25286 34496
rect 25593 34493 25605 34496
rect 25639 34493 25651 34527
rect 27724 34524 27752 34632
rect 27798 34620 27804 34672
rect 27856 34660 27862 34672
rect 31478 34660 31484 34672
rect 27856 34632 29224 34660
rect 27856 34620 27862 34632
rect 28258 34592 28264 34604
rect 28219 34564 28264 34592
rect 28258 34552 28264 34564
rect 28316 34552 28322 34604
rect 28537 34595 28595 34601
rect 28537 34561 28549 34595
rect 28583 34592 28595 34595
rect 28626 34592 28632 34604
rect 28583 34564 28632 34592
rect 28583 34561 28595 34564
rect 28537 34555 28595 34561
rect 28626 34552 28632 34564
rect 28684 34552 28690 34604
rect 29196 34601 29224 34632
rect 29380 34632 31484 34660
rect 29181 34595 29239 34601
rect 29181 34561 29193 34595
rect 29227 34561 29239 34595
rect 29181 34555 29239 34561
rect 28353 34527 28411 34533
rect 28353 34524 28365 34527
rect 27724 34496 28365 34524
rect 25593 34487 25651 34493
rect 28353 34493 28365 34496
rect 28399 34524 28411 34527
rect 29380 34524 29408 34632
rect 31478 34620 31484 34632
rect 31536 34620 31542 34672
rect 32309 34663 32367 34669
rect 32309 34629 32321 34663
rect 32355 34629 32367 34663
rect 46014 34660 46020 34672
rect 32309 34623 32367 34629
rect 41386 34632 46020 34660
rect 29457 34595 29515 34601
rect 29457 34561 29469 34595
rect 29503 34592 29515 34595
rect 30282 34592 30288 34604
rect 29503 34564 30288 34592
rect 29503 34561 29515 34564
rect 29457 34555 29515 34561
rect 30282 34552 30288 34564
rect 30340 34552 30346 34604
rect 30558 34552 30564 34604
rect 30616 34592 30622 34604
rect 30834 34592 30840 34604
rect 30616 34564 30840 34592
rect 30616 34552 30622 34564
rect 30834 34552 30840 34564
rect 30892 34552 30898 34604
rect 30929 34595 30987 34601
rect 30929 34561 30941 34595
rect 30975 34592 30987 34595
rect 31202 34592 31208 34604
rect 30975 34564 31208 34592
rect 30975 34561 30987 34564
rect 30929 34555 30987 34561
rect 31202 34552 31208 34564
rect 31260 34552 31266 34604
rect 32324 34592 32352 34623
rect 41386 34592 41414 34632
rect 46014 34620 46020 34632
rect 46072 34620 46078 34672
rect 46750 34592 46756 34604
rect 32324 34564 41414 34592
rect 46711 34564 46756 34592
rect 46750 34552 46756 34564
rect 46808 34552 46814 34604
rect 28399 34496 29408 34524
rect 28399 34493 28411 34496
rect 28353 34487 28411 34493
rect 19720 34428 22094 34456
rect 19334 34348 19340 34400
rect 19392 34388 19398 34400
rect 19797 34391 19855 34397
rect 19797 34388 19809 34391
rect 19392 34360 19809 34388
rect 19392 34348 19398 34360
rect 19797 34357 19809 34360
rect 19843 34357 19855 34391
rect 22066 34388 22094 34428
rect 22186 34416 22192 34468
rect 22244 34416 22250 34468
rect 25608 34456 25636 34487
rect 29638 34484 29644 34536
rect 29696 34524 29702 34536
rect 30653 34527 30711 34533
rect 30653 34524 30665 34527
rect 29696 34496 30665 34524
rect 29696 34484 29702 34496
rect 30653 34493 30665 34496
rect 30699 34493 30711 34527
rect 30653 34487 30711 34493
rect 30742 34484 30748 34536
rect 30800 34524 30806 34536
rect 30800 34496 30845 34524
rect 30800 34484 30806 34496
rect 28074 34456 28080 34468
rect 25608 34428 28080 34456
rect 28074 34416 28080 34428
rect 28132 34416 28138 34468
rect 30282 34416 30288 34468
rect 30340 34456 30346 34468
rect 30340 34428 31754 34456
rect 30340 34416 30346 34428
rect 23474 34388 23480 34400
rect 22066 34360 23480 34388
rect 19797 34351 19855 34357
rect 23474 34348 23480 34360
rect 23532 34348 23538 34400
rect 24026 34388 24032 34400
rect 23987 34360 24032 34388
rect 24026 34348 24032 34360
rect 24084 34348 24090 34400
rect 25314 34348 25320 34400
rect 25372 34388 25378 34400
rect 25501 34391 25559 34397
rect 25501 34388 25513 34391
rect 25372 34360 25513 34388
rect 25372 34348 25378 34360
rect 25501 34357 25513 34360
rect 25547 34357 25559 34391
rect 25958 34388 25964 34400
rect 25919 34360 25964 34388
rect 25501 34351 25559 34357
rect 25958 34348 25964 34360
rect 26016 34348 26022 34400
rect 27982 34348 27988 34400
rect 28040 34388 28046 34400
rect 28261 34391 28319 34397
rect 28261 34388 28273 34391
rect 28040 34360 28273 34388
rect 28040 34348 28046 34360
rect 28261 34357 28273 34360
rect 28307 34357 28319 34391
rect 28261 34351 28319 34357
rect 30374 34348 30380 34400
rect 30432 34388 30438 34400
rect 30469 34391 30527 34397
rect 30469 34388 30481 34391
rect 30432 34360 30481 34388
rect 30432 34348 30438 34360
rect 30469 34357 30481 34360
rect 30515 34357 30527 34391
rect 31726 34388 31754 34428
rect 32493 34391 32551 34397
rect 32493 34388 32505 34391
rect 31726 34360 32505 34388
rect 30469 34351 30527 34357
rect 32493 34357 32505 34360
rect 32539 34357 32551 34391
rect 32493 34351 32551 34357
rect 46474 34348 46480 34400
rect 46532 34388 46538 34400
rect 46845 34391 46903 34397
rect 46845 34388 46857 34391
rect 46532 34360 46857 34388
rect 46532 34348 46538 34360
rect 46845 34357 46857 34360
rect 46891 34357 46903 34391
rect 47762 34388 47768 34400
rect 47723 34360 47768 34388
rect 46845 34351 46903 34357
rect 47762 34348 47768 34360
rect 47820 34348 47826 34400
rect 1104 34298 48852 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 48852 34298
rect 1104 34224 48852 34246
rect 20346 34144 20352 34196
rect 20404 34184 20410 34196
rect 20441 34187 20499 34193
rect 20441 34184 20453 34187
rect 20404 34156 20453 34184
rect 20404 34144 20410 34156
rect 20441 34153 20453 34156
rect 20487 34153 20499 34187
rect 20441 34147 20499 34153
rect 22005 34187 22063 34193
rect 22005 34153 22017 34187
rect 22051 34184 22063 34187
rect 22462 34184 22468 34196
rect 22051 34156 22468 34184
rect 22051 34153 22063 34156
rect 22005 34147 22063 34153
rect 22462 34144 22468 34156
rect 22520 34144 22526 34196
rect 24578 34144 24584 34196
rect 24636 34184 24642 34196
rect 24765 34187 24823 34193
rect 24765 34184 24777 34187
rect 24636 34156 24777 34184
rect 24636 34144 24642 34156
rect 24765 34153 24777 34156
rect 24811 34153 24823 34187
rect 24765 34147 24823 34153
rect 25222 34116 25228 34128
rect 20916 34088 25228 34116
rect 19794 34008 19800 34060
rect 19852 34048 19858 34060
rect 20622 34048 20628 34060
rect 19852 34020 20628 34048
rect 19852 34008 19858 34020
rect 20622 34008 20628 34020
rect 20680 34008 20686 34060
rect 20916 34057 20944 34088
rect 25222 34076 25228 34088
rect 25280 34076 25286 34128
rect 25406 34076 25412 34128
rect 25464 34116 25470 34128
rect 47762 34116 47768 34128
rect 25464 34088 27936 34116
rect 25464 34076 25470 34088
rect 20901 34051 20959 34057
rect 20901 34017 20913 34051
rect 20947 34017 20959 34051
rect 20901 34011 20959 34017
rect 21085 34051 21143 34057
rect 21085 34017 21097 34051
rect 21131 34048 21143 34051
rect 21174 34048 21180 34060
rect 21131 34020 21180 34048
rect 21131 34017 21143 34020
rect 21085 34011 21143 34017
rect 21174 34008 21180 34020
rect 21232 34008 21238 34060
rect 23845 34051 23903 34057
rect 23845 34048 23857 34051
rect 22572 34020 23857 34048
rect 19613 33983 19671 33989
rect 19613 33949 19625 33983
rect 19659 33980 19671 33983
rect 20530 33980 20536 33992
rect 19659 33952 20536 33980
rect 19659 33949 19671 33952
rect 19613 33943 19671 33949
rect 20530 33940 20536 33952
rect 20588 33940 20594 33992
rect 22281 33983 22339 33989
rect 22486 33983 22544 33989
rect 22281 33949 22293 33983
rect 22327 33949 22339 33983
rect 22281 33943 22339 33949
rect 22370 33977 22428 33983
rect 22370 33943 22382 33977
rect 22416 33943 22428 33977
rect 22486 33949 22498 33983
rect 22532 33980 22544 33983
rect 22572 33980 22600 34020
rect 23845 34017 23857 34020
rect 23891 34017 23903 34051
rect 23845 34011 23903 34017
rect 24854 34008 24860 34060
rect 24912 34048 24918 34060
rect 24912 34020 25820 34048
rect 24912 34008 24918 34020
rect 22532 33952 22600 33980
rect 22649 33983 22707 33989
rect 22532 33949 22544 33952
rect 22486 33943 22544 33949
rect 22649 33949 22661 33983
rect 22695 33949 22707 33983
rect 22649 33943 22707 33949
rect 23477 33983 23535 33989
rect 23477 33949 23489 33983
rect 23523 33980 23535 33983
rect 24026 33980 24032 33992
rect 23523 33952 24032 33980
rect 23523 33949 23535 33952
rect 23477 33943 23535 33949
rect 19794 33912 19800 33924
rect 19755 33884 19800 33912
rect 19794 33872 19800 33884
rect 19852 33872 19858 33924
rect 20346 33872 20352 33924
rect 20404 33912 20410 33924
rect 20809 33915 20867 33921
rect 20809 33912 20821 33915
rect 20404 33884 20821 33912
rect 20404 33872 20410 33884
rect 20809 33881 20821 33884
rect 20855 33881 20867 33915
rect 20809 33875 20867 33881
rect 22296 33856 22324 33943
rect 22370 33937 22428 33943
rect 22385 33856 22413 33937
rect 22664 33912 22692 33943
rect 24026 33940 24032 33952
rect 24084 33940 24090 33992
rect 24118 33940 24124 33992
rect 24176 33980 24182 33992
rect 25409 33983 25467 33989
rect 24176 33952 24808 33980
rect 24176 33940 24182 33952
rect 22572 33884 22692 33912
rect 23661 33915 23719 33921
rect 22572 33856 22600 33884
rect 23661 33881 23673 33915
rect 23707 33881 23719 33915
rect 23661 33875 23719 33881
rect 1762 33804 1768 33856
rect 1820 33844 1826 33856
rect 1857 33847 1915 33853
rect 1857 33844 1869 33847
rect 1820 33816 1869 33844
rect 1820 33804 1826 33816
rect 1857 33813 1869 33816
rect 1903 33813 1915 33847
rect 1857 33807 1915 33813
rect 19981 33847 20039 33853
rect 19981 33813 19993 33847
rect 20027 33844 20039 33847
rect 20622 33844 20628 33856
rect 20027 33816 20628 33844
rect 20027 33813 20039 33816
rect 19981 33807 20039 33813
rect 20622 33804 20628 33816
rect 20680 33804 20686 33856
rect 22278 33804 22284 33856
rect 22336 33804 22342 33856
rect 22370 33804 22376 33856
rect 22428 33804 22434 33856
rect 22554 33804 22560 33856
rect 22612 33804 22618 33856
rect 23676 33844 23704 33875
rect 24210 33872 24216 33924
rect 24268 33912 24274 33924
rect 24486 33912 24492 33924
rect 24268 33884 24492 33912
rect 24268 33872 24274 33884
rect 24486 33872 24492 33884
rect 24544 33912 24550 33924
rect 24673 33915 24731 33921
rect 24673 33912 24685 33915
rect 24544 33884 24685 33912
rect 24544 33872 24550 33884
rect 24673 33881 24685 33884
rect 24719 33881 24731 33915
rect 24780 33912 24808 33952
rect 25409 33949 25421 33983
rect 25455 33980 25467 33983
rect 25498 33980 25504 33992
rect 25455 33952 25504 33980
rect 25455 33949 25467 33952
rect 25409 33943 25467 33949
rect 25498 33940 25504 33952
rect 25556 33940 25562 33992
rect 25792 33989 25820 34020
rect 25593 33983 25651 33989
rect 25593 33949 25605 33983
rect 25639 33949 25651 33983
rect 25593 33943 25651 33949
rect 25777 33983 25835 33989
rect 25777 33949 25789 33983
rect 25823 33949 25835 33983
rect 25958 33980 25964 33992
rect 25919 33952 25964 33980
rect 25777 33943 25835 33949
rect 25608 33912 25636 33943
rect 25958 33940 25964 33952
rect 26016 33940 26022 33992
rect 27908 33989 27936 34088
rect 46308 34088 47768 34116
rect 28074 34048 28080 34060
rect 28035 34020 28080 34048
rect 28074 34008 28080 34020
rect 28132 34008 28138 34060
rect 29546 34048 29552 34060
rect 29507 34020 29552 34048
rect 29546 34008 29552 34020
rect 29604 34008 29610 34060
rect 32030 34048 32036 34060
rect 31991 34020 32036 34048
rect 32030 34008 32036 34020
rect 32088 34008 32094 34060
rect 46308 34057 46336 34088
rect 47762 34076 47768 34088
rect 47820 34076 47826 34128
rect 46293 34051 46351 34057
rect 46293 34017 46305 34051
rect 46339 34017 46351 34051
rect 46474 34048 46480 34060
rect 46435 34020 46480 34048
rect 46293 34011 46351 34017
rect 46474 34008 46480 34020
rect 46532 34008 46538 34060
rect 48130 34048 48136 34060
rect 48091 34020 48136 34048
rect 48130 34008 48136 34020
rect 48188 34008 48194 34060
rect 26697 33983 26755 33989
rect 26697 33949 26709 33983
rect 26743 33980 26755 33983
rect 27893 33983 27951 33989
rect 26743 33952 27568 33980
rect 26743 33949 26755 33952
rect 26697 33943 26755 33949
rect 26050 33912 26056 33924
rect 24780 33884 25636 33912
rect 25700 33884 26056 33912
rect 24673 33875 24731 33881
rect 23750 33844 23756 33856
rect 23663 33816 23756 33844
rect 23750 33804 23756 33816
rect 23808 33844 23814 33856
rect 25700 33844 25728 33884
rect 26050 33872 26056 33884
rect 26108 33872 26114 33924
rect 26234 33872 26240 33924
rect 26292 33912 26298 33924
rect 26881 33915 26939 33921
rect 26881 33912 26893 33915
rect 26292 33884 26893 33912
rect 26292 33872 26298 33884
rect 26881 33881 26893 33884
rect 26927 33881 26939 33915
rect 26881 33875 26939 33881
rect 23808 33816 25728 33844
rect 25869 33847 25927 33853
rect 23808 33804 23814 33816
rect 25869 33813 25881 33847
rect 25915 33844 25927 33847
rect 25958 33844 25964 33856
rect 25915 33816 25964 33844
rect 25915 33813 25927 33816
rect 25869 33807 25927 33813
rect 25958 33804 25964 33816
rect 26016 33804 26022 33856
rect 27065 33847 27123 33853
rect 27065 33813 27077 33847
rect 27111 33844 27123 33847
rect 27246 33844 27252 33856
rect 27111 33816 27252 33844
rect 27111 33813 27123 33816
rect 27065 33807 27123 33813
rect 27246 33804 27252 33816
rect 27304 33804 27310 33856
rect 27540 33853 27568 33952
rect 27893 33949 27905 33983
rect 27939 33980 27951 33983
rect 28350 33980 28356 33992
rect 27939 33952 28356 33980
rect 27939 33949 27951 33952
rect 27893 33943 27951 33949
rect 28350 33940 28356 33952
rect 28408 33940 28414 33992
rect 29816 33983 29874 33989
rect 29816 33949 29828 33983
rect 29862 33980 29874 33983
rect 30374 33980 30380 33992
rect 29862 33952 30380 33980
rect 29862 33949 29874 33952
rect 29816 33943 29874 33949
rect 30374 33940 30380 33952
rect 30432 33940 30438 33992
rect 31754 33940 31760 33992
rect 31812 33980 31818 33992
rect 31812 33952 31857 33980
rect 31812 33940 31818 33952
rect 27525 33847 27583 33853
rect 27525 33813 27537 33847
rect 27571 33813 27583 33847
rect 27525 33807 27583 33813
rect 27985 33847 28043 33853
rect 27985 33813 27997 33847
rect 28031 33844 28043 33847
rect 28994 33844 29000 33856
rect 28031 33816 29000 33844
rect 28031 33813 28043 33816
rect 27985 33807 28043 33813
rect 28994 33804 29000 33816
rect 29052 33804 29058 33856
rect 30834 33804 30840 33856
rect 30892 33844 30898 33856
rect 30929 33847 30987 33853
rect 30929 33844 30941 33847
rect 30892 33816 30941 33844
rect 30892 33804 30898 33816
rect 30929 33813 30941 33816
rect 30975 33813 30987 33847
rect 30929 33807 30987 33813
rect 1104 33754 48852 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 48852 33754
rect 1104 33680 48852 33702
rect 20530 33640 20536 33652
rect 20491 33612 20536 33640
rect 20530 33600 20536 33612
rect 20588 33600 20594 33652
rect 23293 33643 23351 33649
rect 23293 33609 23305 33643
rect 23339 33640 23351 33643
rect 24118 33640 24124 33652
rect 23339 33612 24124 33640
rect 23339 33609 23351 33612
rect 23293 33603 23351 33609
rect 24118 33600 24124 33612
rect 24176 33600 24182 33652
rect 24762 33600 24768 33652
rect 24820 33640 24826 33652
rect 25685 33643 25743 33649
rect 25685 33640 25697 33643
rect 24820 33612 25697 33640
rect 24820 33600 24826 33612
rect 25685 33609 25697 33612
rect 25731 33609 25743 33643
rect 25685 33603 25743 33609
rect 19334 33572 19340 33584
rect 18064 33544 19340 33572
rect 1762 33504 1768 33516
rect 1723 33476 1768 33504
rect 1762 33464 1768 33476
rect 1820 33464 1826 33516
rect 18064 33513 18092 33544
rect 19334 33532 19340 33544
rect 19392 33532 19398 33584
rect 21821 33575 21879 33581
rect 21821 33572 21833 33575
rect 20079 33544 21833 33572
rect 18049 33507 18107 33513
rect 18049 33473 18061 33507
rect 18095 33473 18107 33507
rect 18049 33467 18107 33473
rect 18316 33507 18374 33513
rect 18316 33473 18328 33507
rect 18362 33504 18374 33507
rect 20079 33504 20107 33544
rect 21821 33541 21833 33544
rect 21867 33541 21879 33575
rect 22554 33572 22560 33584
rect 21821 33535 21879 33541
rect 21928 33544 22560 33572
rect 18362 33476 20107 33504
rect 20901 33507 20959 33513
rect 18362 33473 18374 33476
rect 18316 33467 18374 33473
rect 20901 33473 20913 33507
rect 20947 33504 20959 33507
rect 21082 33504 21088 33516
rect 20947 33476 21088 33504
rect 20947 33473 20959 33476
rect 20901 33467 20959 33473
rect 21082 33464 21088 33476
rect 21140 33464 21146 33516
rect 21634 33464 21640 33516
rect 21692 33504 21698 33516
rect 21928 33504 21956 33544
rect 21692 33476 21956 33504
rect 22097 33507 22155 33513
rect 21692 33464 21698 33476
rect 22097 33473 22109 33507
rect 22143 33473 22155 33507
rect 22097 33467 22155 33473
rect 22189 33507 22247 33513
rect 22189 33473 22201 33507
rect 22235 33473 22247 33507
rect 22189 33467 22247 33473
rect 1946 33436 1952 33448
rect 1907 33408 1952 33436
rect 1946 33396 1952 33408
rect 2004 33396 2010 33448
rect 2774 33436 2780 33448
rect 2735 33408 2780 33436
rect 2774 33396 2780 33408
rect 2832 33396 2838 33448
rect 20993 33439 21051 33445
rect 20993 33405 21005 33439
rect 21039 33405 21051 33439
rect 21174 33436 21180 33448
rect 21135 33408 21180 33436
rect 20993 33399 21051 33405
rect 21008 33368 21036 33399
rect 21174 33396 21180 33408
rect 21232 33396 21238 33448
rect 21910 33396 21916 33448
rect 21968 33436 21974 33448
rect 22112 33436 22140 33467
rect 21968 33408 22140 33436
rect 22217 33436 22245 33467
rect 22278 33464 22284 33516
rect 22336 33504 22342 33516
rect 22480 33513 22508 33544
rect 22554 33532 22560 33544
rect 22612 33572 22618 33584
rect 22612 33544 23060 33572
rect 22612 33532 22618 33544
rect 22465 33507 22523 33513
rect 22336 33476 22381 33504
rect 22336 33464 22342 33476
rect 22465 33473 22477 33507
rect 22511 33473 22523 33507
rect 22922 33504 22928 33516
rect 22883 33476 22928 33504
rect 22465 33467 22523 33473
rect 22922 33464 22928 33476
rect 22980 33464 22986 33516
rect 23032 33504 23060 33544
rect 23474 33532 23480 33584
rect 23532 33572 23538 33584
rect 25593 33575 25651 33581
rect 25593 33572 25605 33575
rect 23532 33544 25605 33572
rect 23532 33532 23538 33544
rect 25593 33541 25605 33544
rect 25639 33541 25651 33575
rect 25700 33572 25728 33603
rect 26050 33600 26056 33652
rect 26108 33640 26114 33652
rect 26237 33643 26295 33649
rect 26237 33640 26249 33643
rect 26108 33612 26249 33640
rect 26108 33600 26114 33612
rect 26237 33609 26249 33612
rect 26283 33609 26295 33643
rect 28350 33640 28356 33652
rect 28311 33612 28356 33640
rect 26237 33603 26295 33609
rect 28350 33600 28356 33612
rect 28408 33600 28414 33652
rect 29546 33600 29552 33652
rect 29604 33640 29610 33652
rect 31113 33643 31171 33649
rect 31113 33640 31125 33643
rect 29604 33612 31125 33640
rect 29604 33600 29610 33612
rect 31113 33609 31125 33612
rect 31159 33609 31171 33643
rect 31113 33603 31171 33609
rect 25700 33544 27016 33572
rect 25593 33535 25651 33541
rect 26988 33516 27016 33544
rect 31754 33532 31760 33584
rect 31812 33572 31818 33584
rect 32309 33575 32367 33581
rect 32309 33572 32321 33575
rect 31812 33544 32321 33572
rect 31812 33532 31818 33544
rect 32309 33541 32321 33544
rect 32355 33541 32367 33575
rect 32309 33535 32367 33541
rect 23934 33504 23940 33516
rect 23032 33476 23940 33504
rect 23934 33464 23940 33476
rect 23992 33464 23998 33516
rect 24210 33464 24216 33516
rect 24268 33504 24274 33516
rect 24673 33507 24731 33513
rect 24673 33504 24685 33507
rect 24268 33476 24685 33504
rect 24268 33464 24274 33476
rect 24673 33473 24685 33476
rect 24719 33473 24731 33507
rect 24673 33467 24731 33473
rect 24765 33507 24823 33513
rect 24765 33473 24777 33507
rect 24811 33504 24823 33507
rect 25406 33504 25412 33516
rect 24811 33476 25412 33504
rect 24811 33473 24823 33476
rect 24765 33467 24823 33473
rect 25406 33464 25412 33476
rect 25464 33464 25470 33516
rect 26418 33504 26424 33516
rect 26379 33476 26424 33504
rect 26418 33464 26424 33476
rect 26476 33464 26482 33516
rect 26970 33504 26976 33516
rect 26883 33476 26976 33504
rect 26970 33464 26976 33476
rect 27028 33464 27034 33516
rect 27062 33464 27068 33516
rect 27120 33504 27126 33516
rect 27229 33507 27287 33513
rect 27229 33504 27241 33507
rect 27120 33476 27241 33504
rect 27120 33464 27126 33476
rect 27229 33473 27241 33476
rect 27275 33473 27287 33507
rect 27229 33467 27287 33473
rect 29641 33507 29699 33513
rect 29641 33473 29653 33507
rect 29687 33504 29699 33507
rect 30558 33504 30564 33516
rect 29687 33476 30564 33504
rect 29687 33473 29699 33476
rect 29641 33467 29699 33473
rect 30558 33464 30564 33476
rect 30616 33464 30622 33516
rect 31018 33504 31024 33516
rect 30979 33476 31024 33504
rect 31018 33464 31024 33476
rect 31076 33464 31082 33516
rect 31938 33464 31944 33516
rect 31996 33504 32002 33516
rect 32125 33507 32183 33513
rect 32125 33504 32137 33507
rect 31996 33476 32137 33504
rect 31996 33464 32002 33476
rect 32125 33473 32137 33476
rect 32171 33473 32183 33507
rect 32125 33467 32183 33473
rect 46014 33464 46020 33516
rect 46072 33504 46078 33516
rect 46477 33507 46535 33513
rect 46477 33504 46489 33507
rect 46072 33476 46489 33504
rect 46072 33464 46078 33476
rect 46477 33473 46489 33476
rect 46523 33473 46535 33507
rect 46477 33467 46535 33473
rect 22370 33436 22376 33448
rect 22217 33408 22376 33436
rect 21968 33396 21974 33408
rect 22370 33396 22376 33408
rect 22428 33396 22434 33448
rect 22554 33396 22560 33448
rect 22612 33436 22618 33448
rect 23017 33439 23075 33445
rect 23017 33436 23029 33439
rect 22612 33408 23029 33436
rect 22612 33396 22618 33408
rect 23017 33405 23029 33408
rect 23063 33405 23075 33439
rect 23017 33399 23075 33405
rect 24578 33396 24584 33448
rect 24636 33436 24642 33448
rect 24857 33439 24915 33445
rect 24857 33436 24869 33439
rect 24636 33408 24869 33436
rect 24636 33396 24642 33408
rect 24857 33405 24869 33408
rect 24903 33405 24915 33439
rect 24857 33399 24915 33405
rect 29365 33439 29423 33445
rect 29365 33405 29377 33439
rect 29411 33405 29423 33439
rect 46198 33436 46204 33448
rect 46159 33408 46204 33436
rect 29365 33399 29423 33405
rect 25314 33368 25320 33380
rect 21008 33340 22048 33368
rect 19429 33303 19487 33309
rect 19429 33269 19441 33303
rect 19475 33300 19487 33303
rect 19886 33300 19892 33312
rect 19475 33272 19892 33300
rect 19475 33269 19487 33272
rect 19429 33263 19487 33269
rect 19886 33260 19892 33272
rect 19944 33260 19950 33312
rect 20438 33260 20444 33312
rect 20496 33300 20502 33312
rect 21358 33300 21364 33312
rect 20496 33272 21364 33300
rect 20496 33260 20502 33272
rect 21358 33260 21364 33272
rect 21416 33260 21422 33312
rect 22020 33300 22048 33340
rect 23032 33340 25320 33368
rect 23032 33300 23060 33340
rect 25314 33328 25320 33340
rect 25372 33328 25378 33380
rect 22020 33272 23060 33300
rect 23109 33303 23167 33309
rect 23109 33269 23121 33303
rect 23155 33300 23167 33303
rect 23290 33300 23296 33312
rect 23155 33272 23296 33300
rect 23155 33269 23167 33272
rect 23109 33263 23167 33269
rect 23290 33260 23296 33272
rect 23348 33260 23354 33312
rect 23566 33260 23572 33312
rect 23624 33300 23630 33312
rect 24305 33303 24363 33309
rect 24305 33300 24317 33303
rect 23624 33272 24317 33300
rect 23624 33260 23630 33272
rect 24305 33269 24317 33272
rect 24351 33269 24363 33303
rect 24305 33263 24363 33269
rect 24394 33260 24400 33312
rect 24452 33300 24458 33312
rect 29380 33300 29408 33399
rect 46198 33396 46204 33408
rect 46256 33396 46262 33448
rect 24452 33272 29408 33300
rect 32493 33303 32551 33309
rect 24452 33260 24458 33272
rect 32493 33269 32505 33303
rect 32539 33300 32551 33303
rect 32858 33300 32864 33312
rect 32539 33272 32864 33300
rect 32539 33269 32551 33272
rect 32493 33263 32551 33269
rect 32858 33260 32864 33272
rect 32916 33260 32922 33312
rect 47762 33300 47768 33312
rect 47723 33272 47768 33300
rect 47762 33260 47768 33272
rect 47820 33260 47826 33312
rect 1104 33210 48852 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 48852 33210
rect 1104 33136 48852 33158
rect 1946 33056 1952 33108
rect 2004 33096 2010 33108
rect 2133 33099 2191 33105
rect 2133 33096 2145 33099
rect 2004 33068 2145 33096
rect 2004 33056 2010 33068
rect 2133 33065 2145 33068
rect 2179 33065 2191 33099
rect 2133 33059 2191 33065
rect 19978 33056 19984 33108
rect 20036 33096 20042 33108
rect 20438 33096 20444 33108
rect 20036 33068 20444 33096
rect 20036 33056 20042 33068
rect 20438 33056 20444 33068
rect 20496 33056 20502 33108
rect 20533 33099 20591 33105
rect 20533 33065 20545 33099
rect 20579 33065 20591 33099
rect 20533 33059 20591 33065
rect 20717 33099 20775 33105
rect 20717 33065 20729 33099
rect 20763 33096 20775 33099
rect 22922 33096 22928 33108
rect 20763 33068 22928 33096
rect 20763 33065 20775 33068
rect 20717 33059 20775 33065
rect 20548 33028 20576 33059
rect 22922 33056 22928 33068
rect 22980 33056 22986 33108
rect 23017 33099 23075 33105
rect 23017 33065 23029 33099
rect 23063 33096 23075 33099
rect 23842 33096 23848 33108
rect 23063 33068 23848 33096
rect 23063 33065 23075 33068
rect 23017 33059 23075 33065
rect 23842 33056 23848 33068
rect 23900 33056 23906 33108
rect 24762 33096 24768 33108
rect 24412 33068 24768 33096
rect 20990 33028 20996 33040
rect 20548 33000 20996 33028
rect 20990 32988 20996 33000
rect 21048 32988 21054 33040
rect 24210 33028 24216 33040
rect 21100 33000 24216 33028
rect 15194 32920 15200 32972
rect 15252 32960 15258 32972
rect 16025 32963 16083 32969
rect 16025 32960 16037 32963
rect 15252 32932 16037 32960
rect 15252 32920 15258 32932
rect 16025 32929 16037 32932
rect 16071 32929 16083 32963
rect 16025 32923 16083 32929
rect 19978 32920 19984 32972
rect 20036 32960 20042 32972
rect 20346 32960 20352 32972
rect 20036 32932 20352 32960
rect 20036 32920 20042 32932
rect 20346 32920 20352 32932
rect 20404 32920 20410 32972
rect 21100 32960 21128 33000
rect 24210 32988 24216 33000
rect 24268 32988 24274 33040
rect 20456 32932 21128 32960
rect 21177 32963 21235 32969
rect 1581 32895 1639 32901
rect 1581 32861 1593 32895
rect 1627 32892 1639 32895
rect 1946 32892 1952 32904
rect 1627 32864 1952 32892
rect 1627 32861 1639 32864
rect 1581 32855 1639 32861
rect 1946 32852 1952 32864
rect 2004 32852 2010 32904
rect 2041 32895 2099 32901
rect 2041 32861 2053 32895
rect 2087 32892 2099 32895
rect 2130 32892 2136 32904
rect 2087 32864 2136 32892
rect 2087 32861 2099 32864
rect 2041 32855 2099 32861
rect 2130 32852 2136 32864
rect 2188 32892 2194 32904
rect 2406 32892 2412 32904
rect 2188 32864 2412 32892
rect 2188 32852 2194 32864
rect 2406 32852 2412 32864
rect 2464 32852 2470 32904
rect 2682 32892 2688 32904
rect 2643 32864 2688 32892
rect 2682 32852 2688 32864
rect 2740 32852 2746 32904
rect 15562 32892 15568 32904
rect 15523 32864 15568 32892
rect 15562 32852 15568 32864
rect 15620 32852 15626 32904
rect 20070 32852 20076 32904
rect 20128 32892 20134 32904
rect 20257 32895 20315 32901
rect 20257 32892 20269 32895
rect 20128 32864 20269 32892
rect 20128 32852 20134 32864
rect 20257 32861 20269 32864
rect 20303 32892 20315 32895
rect 20456 32892 20484 32932
rect 21177 32929 21189 32963
rect 21223 32960 21235 32963
rect 22002 32960 22008 32972
rect 21223 32932 22008 32960
rect 21223 32929 21235 32932
rect 21177 32923 21235 32929
rect 22002 32920 22008 32932
rect 22060 32920 22066 32972
rect 22572 32932 23704 32960
rect 20303 32864 20484 32892
rect 20303 32861 20315 32864
rect 20257 32855 20315 32861
rect 20530 32852 20536 32904
rect 20588 32892 20594 32904
rect 20588 32864 20633 32892
rect 20588 32852 20594 32864
rect 20806 32852 20812 32904
rect 20864 32892 20870 32904
rect 21453 32895 21511 32901
rect 21453 32892 21465 32895
rect 20864 32864 21465 32892
rect 20864 32852 20870 32864
rect 21453 32861 21465 32864
rect 21499 32861 21511 32895
rect 21453 32855 21511 32861
rect 15746 32824 15752 32836
rect 15707 32796 15752 32824
rect 15746 32784 15752 32796
rect 15804 32784 15810 32836
rect 19613 32827 19671 32833
rect 19613 32793 19625 32827
rect 19659 32824 19671 32827
rect 20714 32824 20720 32836
rect 19659 32796 20720 32824
rect 19659 32793 19671 32796
rect 19613 32787 19671 32793
rect 20714 32784 20720 32796
rect 20772 32824 20778 32836
rect 20898 32824 20904 32836
rect 20772 32796 20904 32824
rect 20772 32784 20778 32796
rect 20898 32784 20904 32796
rect 20956 32784 20962 32836
rect 22572 32824 22600 32932
rect 22649 32895 22707 32901
rect 22649 32861 22661 32895
rect 22695 32892 22707 32895
rect 23566 32892 23572 32904
rect 22695 32864 23572 32892
rect 22695 32861 22707 32864
rect 22649 32855 22707 32861
rect 23566 32852 23572 32864
rect 23624 32852 23630 32904
rect 23676 32901 23704 32932
rect 23661 32895 23719 32901
rect 23661 32861 23673 32895
rect 23707 32892 23719 32895
rect 23750 32892 23756 32904
rect 23707 32864 23756 32892
rect 23707 32861 23719 32864
rect 23661 32855 23719 32861
rect 23750 32852 23756 32864
rect 23808 32852 23814 32904
rect 24228 32892 24256 32988
rect 24302 32920 24308 32972
rect 24360 32960 24366 32972
rect 24412 32969 24440 33068
rect 24762 33056 24768 33068
rect 24820 33056 24826 33108
rect 26789 33099 26847 33105
rect 26789 33065 26801 33099
rect 26835 33096 26847 33099
rect 27062 33096 27068 33108
rect 26835 33068 27068 33096
rect 26835 33065 26847 33068
rect 26789 33059 26847 33065
rect 27062 33056 27068 33068
rect 27120 33056 27126 33108
rect 30285 33099 30343 33105
rect 30285 33065 30297 33099
rect 30331 33065 30343 33099
rect 30466 33096 30472 33108
rect 30427 33068 30472 33096
rect 30285 33059 30343 33065
rect 25777 33031 25835 33037
rect 25777 32997 25789 33031
rect 25823 32997 25835 33031
rect 30300 33028 30328 33059
rect 30466 33056 30472 33068
rect 30524 33056 30530 33108
rect 30558 33056 30564 33108
rect 30616 33096 30622 33108
rect 35894 33096 35900 33108
rect 30616 33068 35900 33096
rect 30616 33056 30622 33068
rect 35894 33056 35900 33068
rect 35952 33056 35958 33108
rect 31294 33028 31300 33040
rect 30300 33000 31300 33028
rect 25777 32991 25835 32997
rect 24397 32963 24455 32969
rect 24397 32960 24409 32963
rect 24360 32932 24409 32960
rect 24360 32920 24366 32932
rect 24397 32929 24409 32932
rect 24443 32929 24455 32963
rect 24397 32923 24455 32929
rect 25792 32892 25820 32991
rect 31294 32988 31300 33000
rect 31352 32988 31358 33040
rect 27338 32960 27344 32972
rect 27172 32932 27344 32960
rect 24228 32864 25820 32892
rect 26142 32852 26148 32904
rect 26200 32892 26206 32904
rect 27172 32901 27200 32932
rect 27338 32920 27344 32932
rect 27396 32920 27402 32972
rect 28810 32960 28816 32972
rect 28552 32932 28816 32960
rect 27065 32895 27123 32901
rect 27065 32892 27077 32895
rect 26200 32864 27077 32892
rect 26200 32852 26206 32864
rect 27065 32861 27077 32864
rect 27111 32861 27123 32895
rect 27065 32855 27123 32861
rect 27157 32895 27215 32901
rect 27157 32861 27169 32895
rect 27203 32861 27215 32895
rect 27157 32855 27215 32861
rect 27246 32852 27252 32904
rect 27304 32892 27310 32904
rect 27433 32895 27491 32901
rect 27304 32864 27349 32892
rect 27304 32852 27310 32864
rect 27433 32861 27445 32895
rect 27479 32892 27491 32895
rect 27706 32892 27712 32904
rect 27479 32864 27712 32892
rect 27479 32861 27491 32864
rect 27433 32855 27491 32861
rect 27706 32852 27712 32864
rect 27764 32852 27770 32904
rect 22833 32827 22891 32833
rect 22833 32824 22845 32827
rect 22572 32796 22845 32824
rect 22833 32793 22845 32796
rect 22879 32793 22891 32827
rect 23474 32824 23480 32836
rect 23435 32796 23480 32824
rect 22833 32787 22891 32793
rect 23474 32784 23480 32796
rect 23532 32784 23538 32836
rect 24642 32827 24700 32833
rect 24642 32824 24654 32827
rect 23768 32796 24654 32824
rect 2130 32716 2136 32768
rect 2188 32756 2194 32768
rect 2777 32759 2835 32765
rect 2777 32756 2789 32759
rect 2188 32728 2789 32756
rect 2188 32716 2194 32728
rect 2777 32725 2789 32728
rect 2823 32725 2835 32759
rect 2777 32719 2835 32725
rect 19705 32759 19763 32765
rect 19705 32725 19717 32759
rect 19751 32756 19763 32759
rect 20806 32756 20812 32768
rect 19751 32728 20812 32756
rect 19751 32725 19763 32728
rect 19705 32719 19763 32725
rect 20806 32716 20812 32728
rect 20864 32716 20870 32768
rect 23198 32716 23204 32768
rect 23256 32756 23262 32768
rect 23768 32756 23796 32796
rect 24642 32793 24654 32796
rect 24688 32793 24700 32827
rect 24642 32787 24700 32793
rect 25774 32784 25780 32836
rect 25832 32824 25838 32836
rect 28074 32824 28080 32836
rect 25832 32796 28080 32824
rect 25832 32784 25838 32796
rect 28074 32784 28080 32796
rect 28132 32824 28138 32836
rect 28552 32824 28580 32932
rect 28810 32920 28816 32932
rect 28868 32920 28874 32972
rect 30193 32963 30251 32969
rect 30193 32960 30205 32963
rect 30024 32932 30205 32960
rect 28721 32895 28779 32901
rect 28721 32861 28733 32895
rect 28767 32892 28779 32895
rect 30024 32892 30052 32932
rect 30193 32929 30205 32932
rect 30239 32960 30251 32963
rect 30834 32960 30840 32972
rect 30239 32932 30840 32960
rect 30239 32929 30251 32932
rect 30193 32923 30251 32929
rect 30834 32920 30840 32932
rect 30892 32920 30898 32972
rect 31662 32960 31668 32972
rect 31623 32932 31668 32960
rect 31662 32920 31668 32932
rect 31720 32920 31726 32972
rect 32122 32920 32128 32972
rect 32180 32960 32186 32972
rect 32582 32960 32588 32972
rect 32180 32932 32588 32960
rect 32180 32920 32186 32932
rect 32582 32920 32588 32932
rect 32640 32920 32646 32972
rect 46293 32963 46351 32969
rect 46293 32929 46305 32963
rect 46339 32960 46351 32963
rect 47762 32960 47768 32972
rect 46339 32932 47768 32960
rect 46339 32929 46351 32932
rect 46293 32923 46351 32929
rect 47762 32920 47768 32932
rect 47820 32920 47826 32972
rect 48038 32960 48044 32972
rect 47999 32932 48044 32960
rect 48038 32920 48044 32932
rect 48096 32920 48102 32972
rect 28767 32864 30052 32892
rect 30101 32895 30159 32901
rect 28767 32861 28779 32864
rect 28721 32855 28779 32861
rect 30101 32861 30113 32895
rect 30147 32861 30159 32895
rect 31478 32892 31484 32904
rect 31439 32864 31484 32892
rect 30101 32855 30159 32861
rect 28132 32796 28580 32824
rect 30116 32824 30144 32855
rect 31478 32852 31484 32864
rect 31536 32892 31542 32904
rect 31536 32864 31754 32892
rect 31536 32852 31542 32864
rect 31202 32824 31208 32836
rect 30116 32796 31208 32824
rect 28132 32784 28138 32796
rect 31202 32784 31208 32796
rect 31260 32824 31266 32836
rect 31573 32827 31631 32833
rect 31573 32824 31585 32827
rect 31260 32796 31585 32824
rect 31260 32784 31266 32796
rect 31573 32793 31585 32796
rect 31619 32793 31631 32827
rect 31573 32787 31631 32793
rect 23256 32728 23796 32756
rect 23845 32759 23903 32765
rect 23256 32716 23262 32728
rect 23845 32725 23857 32759
rect 23891 32756 23903 32759
rect 24854 32756 24860 32768
rect 23891 32728 24860 32756
rect 23891 32725 23903 32728
rect 23845 32719 23903 32725
rect 24854 32716 24860 32728
rect 24912 32716 24918 32768
rect 28166 32716 28172 32768
rect 28224 32756 28230 32768
rect 28261 32759 28319 32765
rect 28261 32756 28273 32759
rect 28224 32728 28273 32756
rect 28224 32716 28230 32728
rect 28261 32725 28273 32728
rect 28307 32725 28319 32759
rect 28626 32756 28632 32768
rect 28587 32728 28632 32756
rect 28261 32719 28319 32725
rect 28626 32716 28632 32728
rect 28684 32716 28690 32768
rect 31110 32756 31116 32768
rect 31071 32728 31116 32756
rect 31110 32716 31116 32728
rect 31168 32716 31174 32768
rect 31726 32756 31754 32864
rect 32306 32852 32312 32904
rect 32364 32892 32370 32904
rect 36081 32895 36139 32901
rect 36081 32892 36093 32895
rect 32364 32864 36093 32892
rect 32364 32852 32370 32864
rect 36081 32861 36093 32864
rect 36127 32861 36139 32895
rect 36081 32855 36139 32861
rect 32398 32784 32404 32836
rect 32456 32824 32462 32836
rect 32830 32827 32888 32833
rect 32830 32824 32842 32827
rect 32456 32796 32842 32824
rect 32456 32784 32462 32796
rect 32830 32793 32842 32796
rect 32876 32793 32888 32827
rect 46474 32824 46480 32836
rect 46435 32796 46480 32824
rect 32830 32787 32888 32793
rect 46474 32784 46480 32796
rect 46532 32784 46538 32836
rect 33965 32759 34023 32765
rect 33965 32756 33977 32759
rect 31726 32728 33977 32756
rect 33965 32725 33977 32728
rect 34011 32725 34023 32759
rect 33965 32719 34023 32725
rect 34054 32716 34060 32768
rect 34112 32756 34118 32768
rect 36265 32759 36323 32765
rect 36265 32756 36277 32759
rect 34112 32728 36277 32756
rect 34112 32716 34118 32728
rect 36265 32725 36277 32728
rect 36311 32756 36323 32759
rect 40770 32756 40776 32768
rect 36311 32728 40776 32756
rect 36311 32725 36323 32728
rect 36265 32719 36323 32725
rect 40770 32716 40776 32728
rect 40828 32716 40834 32768
rect 1104 32666 48852 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 48852 32666
rect 1104 32592 48852 32614
rect 15657 32555 15715 32561
rect 15657 32521 15669 32555
rect 15703 32552 15715 32555
rect 15746 32552 15752 32564
rect 15703 32524 15752 32552
rect 15703 32521 15715 32524
rect 15657 32515 15715 32521
rect 15746 32512 15752 32524
rect 15804 32512 15810 32564
rect 19426 32512 19432 32564
rect 19484 32552 19490 32564
rect 19613 32555 19671 32561
rect 19613 32552 19625 32555
rect 19484 32524 19625 32552
rect 19484 32512 19490 32524
rect 19613 32521 19625 32524
rect 19659 32521 19671 32555
rect 23198 32552 23204 32564
rect 23159 32524 23204 32552
rect 19613 32515 19671 32521
rect 23198 32512 23204 32524
rect 23256 32512 23262 32564
rect 23382 32512 23388 32564
rect 23440 32512 23446 32564
rect 23474 32512 23480 32564
rect 23532 32552 23538 32564
rect 24305 32555 24363 32561
rect 24305 32552 24317 32555
rect 23532 32524 24317 32552
rect 23532 32512 23538 32524
rect 24305 32521 24317 32524
rect 24351 32521 24363 32555
rect 24670 32552 24676 32564
rect 24631 32524 24676 32552
rect 24305 32515 24363 32521
rect 24670 32512 24676 32524
rect 24728 32512 24734 32564
rect 24765 32555 24823 32561
rect 24765 32521 24777 32555
rect 24811 32552 24823 32555
rect 28626 32552 28632 32564
rect 24811 32524 28632 32552
rect 24811 32521 24823 32524
rect 24765 32515 24823 32521
rect 28626 32512 28632 32524
rect 28684 32552 28690 32564
rect 28721 32555 28779 32561
rect 28721 32552 28733 32555
rect 28684 32524 28733 32552
rect 28684 32512 28690 32524
rect 28721 32521 28733 32524
rect 28767 32521 28779 32555
rect 28721 32515 28779 32521
rect 28902 32512 28908 32564
rect 28960 32552 28966 32564
rect 30837 32555 30895 32561
rect 28960 32524 30696 32552
rect 28960 32512 28966 32524
rect 2130 32484 2136 32496
rect 2091 32456 2136 32484
rect 2130 32444 2136 32456
rect 2188 32444 2194 32496
rect 19521 32487 19579 32493
rect 15580 32456 18552 32484
rect 1946 32416 1952 32428
rect 1907 32388 1952 32416
rect 1946 32376 1952 32388
rect 2004 32376 2010 32428
rect 12618 32376 12624 32428
rect 12676 32416 12682 32428
rect 15580 32425 15608 32456
rect 15565 32419 15623 32425
rect 15565 32416 15577 32419
rect 12676 32388 15577 32416
rect 12676 32376 12682 32388
rect 15565 32385 15577 32388
rect 15611 32385 15623 32419
rect 18230 32416 18236 32428
rect 18191 32388 18236 32416
rect 15565 32379 15623 32385
rect 18230 32376 18236 32388
rect 18288 32376 18294 32428
rect 18414 32416 18420 32428
rect 18375 32388 18420 32416
rect 18414 32376 18420 32388
rect 18472 32376 18478 32428
rect 18524 32416 18552 32456
rect 19521 32453 19533 32487
rect 19567 32484 19579 32487
rect 21542 32484 21548 32496
rect 19567 32456 21548 32484
rect 19567 32453 19579 32456
rect 19521 32447 19579 32453
rect 21542 32444 21548 32456
rect 21600 32444 21606 32496
rect 22554 32484 22560 32496
rect 22515 32456 22560 32484
rect 22554 32444 22560 32456
rect 22612 32444 22618 32496
rect 22741 32487 22799 32493
rect 22741 32453 22753 32487
rect 22787 32484 22799 32487
rect 22922 32484 22928 32496
rect 22787 32456 22928 32484
rect 22787 32453 22799 32456
rect 22741 32447 22799 32453
rect 22922 32444 22928 32456
rect 22980 32444 22986 32496
rect 20346 32416 20352 32428
rect 18524 32388 20352 32416
rect 20346 32376 20352 32388
rect 20404 32376 20410 32428
rect 20441 32419 20499 32425
rect 20441 32385 20453 32419
rect 20487 32385 20499 32419
rect 20441 32379 20499 32385
rect 20533 32419 20591 32425
rect 20533 32385 20545 32419
rect 20579 32385 20591 32419
rect 20533 32379 20591 32385
rect 2774 32348 2780 32360
rect 2735 32320 2780 32348
rect 2774 32308 2780 32320
rect 2832 32308 2838 32360
rect 20456 32348 20484 32379
rect 12406 32320 20484 32348
rect 20548 32348 20576 32379
rect 20622 32376 20628 32428
rect 20680 32416 20686 32428
rect 20680 32388 20725 32416
rect 20680 32376 20686 32388
rect 20806 32376 20812 32428
rect 20864 32416 20870 32428
rect 21634 32416 21640 32428
rect 20864 32388 21640 32416
rect 20864 32376 20870 32388
rect 21634 32376 21640 32388
rect 21692 32376 21698 32428
rect 21821 32419 21879 32425
rect 21821 32385 21833 32419
rect 21867 32385 21879 32419
rect 21821 32379 21879 32385
rect 21836 32348 21864 32379
rect 22002 32376 22008 32428
rect 22060 32416 22066 32428
rect 23400 32419 23428 32512
rect 24026 32444 24032 32496
rect 24084 32484 24090 32496
rect 30558 32484 30564 32496
rect 24084 32456 30564 32484
rect 24084 32444 24090 32456
rect 30558 32444 30564 32456
rect 30616 32444 30622 32496
rect 30668 32484 30696 32524
rect 30837 32521 30849 32555
rect 30883 32552 30895 32555
rect 31938 32552 31944 32564
rect 30883 32524 31944 32552
rect 30883 32521 30895 32524
rect 30837 32515 30895 32521
rect 31938 32512 31944 32524
rect 31996 32512 32002 32564
rect 32122 32512 32128 32564
rect 32180 32552 32186 32564
rect 32490 32552 32496 32564
rect 32180 32524 32496 32552
rect 32180 32512 32186 32524
rect 32490 32512 32496 32524
rect 32548 32512 32554 32564
rect 32582 32512 32588 32564
rect 32640 32552 32646 32564
rect 33778 32552 33784 32564
rect 32640 32524 33784 32552
rect 32640 32512 32646 32524
rect 33778 32512 33784 32524
rect 33836 32512 33842 32564
rect 33965 32555 34023 32561
rect 33965 32521 33977 32555
rect 34011 32521 34023 32555
rect 36446 32552 36452 32564
rect 36407 32524 36452 32552
rect 33965 32515 34023 32521
rect 32306 32484 32312 32496
rect 30668 32456 32312 32484
rect 32306 32444 32312 32456
rect 32364 32444 32370 32496
rect 33980 32484 34008 32515
rect 36446 32512 36452 32524
rect 36504 32512 36510 32564
rect 39114 32484 39120 32496
rect 32416 32456 34008 32484
rect 39075 32456 39120 32484
rect 23457 32419 23515 32425
rect 23569 32419 23627 32425
rect 22060 32388 22692 32416
rect 23400 32391 23469 32419
rect 22060 32376 22066 32388
rect 22186 32348 22192 32360
rect 20548 32320 20832 32348
rect 21836 32320 22192 32348
rect 1946 32240 1952 32292
rect 2004 32280 2010 32292
rect 12406 32280 12434 32320
rect 2004 32252 12434 32280
rect 2004 32240 2010 32252
rect 18414 32240 18420 32292
rect 18472 32280 18478 32292
rect 20804 32280 20832 32320
rect 22186 32308 22192 32320
rect 22244 32308 22250 32360
rect 22370 32280 22376 32292
rect 18472 32252 20760 32280
rect 20804 32252 22376 32280
rect 18472 32240 18478 32252
rect 15654 32172 15660 32224
rect 15712 32212 15718 32224
rect 16850 32212 16856 32224
rect 15712 32184 16856 32212
rect 15712 32172 15718 32184
rect 16850 32172 16856 32184
rect 16908 32172 16914 32224
rect 17954 32172 17960 32224
rect 18012 32212 18018 32224
rect 18601 32215 18659 32221
rect 18601 32212 18613 32215
rect 18012 32184 18613 32212
rect 18012 32172 18018 32184
rect 18601 32181 18613 32184
rect 18647 32181 18659 32215
rect 18601 32175 18659 32181
rect 19426 32172 19432 32224
rect 19484 32212 19490 32224
rect 19978 32212 19984 32224
rect 19484 32184 19984 32212
rect 19484 32172 19490 32184
rect 19978 32172 19984 32184
rect 20036 32172 20042 32224
rect 20070 32172 20076 32224
rect 20128 32212 20134 32224
rect 20165 32215 20223 32221
rect 20165 32212 20177 32215
rect 20128 32184 20177 32212
rect 20128 32172 20134 32184
rect 20165 32181 20177 32184
rect 20211 32181 20223 32215
rect 20732 32212 20760 32252
rect 22370 32240 22376 32252
rect 22428 32240 22434 32292
rect 22664 32280 22692 32388
rect 23457 32385 23469 32391
rect 23503 32388 23520 32419
rect 23569 32412 23581 32419
rect 23615 32412 23627 32419
rect 23661 32422 23719 32428
rect 23503 32385 23515 32388
rect 23457 32379 23515 32385
rect 23566 32360 23572 32412
rect 23624 32360 23630 32412
rect 23661 32388 23673 32422
rect 23707 32388 23719 32422
rect 23661 32382 23719 32388
rect 23845 32419 23903 32425
rect 23845 32385 23857 32419
rect 23891 32416 23903 32419
rect 23934 32416 23940 32428
rect 23891 32388 23940 32416
rect 23891 32385 23903 32388
rect 23676 32348 23704 32382
rect 23845 32379 23903 32385
rect 23934 32376 23940 32388
rect 23992 32376 23998 32428
rect 24486 32376 24492 32428
rect 24544 32416 24550 32428
rect 25593 32419 25651 32425
rect 25593 32416 25605 32419
rect 24544 32388 25605 32416
rect 24544 32376 24550 32388
rect 25593 32385 25605 32388
rect 25639 32385 25651 32419
rect 26418 32416 26424 32428
rect 25593 32379 25651 32385
rect 25700 32388 26424 32416
rect 23750 32348 23756 32360
rect 23676 32320 23756 32348
rect 23750 32308 23756 32320
rect 23808 32308 23814 32360
rect 24578 32308 24584 32360
rect 24636 32348 24642 32360
rect 24857 32351 24915 32357
rect 24857 32348 24869 32351
rect 24636 32320 24869 32348
rect 24636 32308 24642 32320
rect 24857 32317 24869 32320
rect 24903 32317 24915 32351
rect 24857 32311 24915 32317
rect 25700 32280 25728 32388
rect 26418 32376 26424 32388
rect 26476 32376 26482 32428
rect 26970 32376 26976 32428
rect 27028 32416 27034 32428
rect 27341 32419 27399 32425
rect 27341 32416 27353 32419
rect 27028 32388 27353 32416
rect 27028 32376 27034 32388
rect 27341 32385 27353 32388
rect 27387 32385 27399 32419
rect 27341 32379 27399 32385
rect 27430 32376 27436 32428
rect 27488 32416 27494 32428
rect 27597 32419 27655 32425
rect 27597 32416 27609 32419
rect 27488 32388 27609 32416
rect 27488 32376 27494 32388
rect 27597 32385 27609 32388
rect 27643 32385 27655 32419
rect 27597 32379 27655 32385
rect 27982 32376 27988 32428
rect 28040 32416 28046 32428
rect 31205 32419 31263 32425
rect 31205 32416 31217 32419
rect 28040 32388 31217 32416
rect 28040 32376 28046 32388
rect 31205 32385 31217 32388
rect 31251 32416 31263 32419
rect 32416 32416 32444 32456
rect 39114 32444 39120 32456
rect 39172 32444 39178 32496
rect 32582 32416 32588 32428
rect 31251 32388 32444 32416
rect 32543 32388 32588 32416
rect 31251 32385 31263 32388
rect 31205 32379 31263 32385
rect 32582 32376 32588 32388
rect 32640 32376 32646 32428
rect 32841 32419 32899 32425
rect 32841 32416 32853 32419
rect 32692 32388 32853 32416
rect 28350 32308 28356 32360
rect 28408 32348 28414 32360
rect 28902 32348 28908 32360
rect 28408 32320 28908 32348
rect 28408 32308 28414 32320
rect 28902 32308 28908 32320
rect 28960 32308 28966 32360
rect 31294 32348 31300 32360
rect 31255 32320 31300 32348
rect 31294 32308 31300 32320
rect 31352 32308 31358 32360
rect 31389 32351 31447 32357
rect 31389 32317 31401 32351
rect 31435 32348 31447 32351
rect 31662 32348 31668 32360
rect 31435 32320 31668 32348
rect 31435 32317 31447 32320
rect 31389 32311 31447 32317
rect 26234 32280 26240 32292
rect 22664 32252 25728 32280
rect 26195 32252 26240 32280
rect 26234 32240 26240 32252
rect 26292 32240 26298 32292
rect 28810 32240 28816 32292
rect 28868 32280 28874 32292
rect 31404 32280 31432 32311
rect 31662 32308 31668 32320
rect 31720 32308 31726 32360
rect 32490 32308 32496 32360
rect 32548 32348 32554 32360
rect 32692 32348 32720 32388
rect 32841 32385 32853 32388
rect 32887 32385 32899 32419
rect 36354 32416 36360 32428
rect 36315 32388 36360 32416
rect 32841 32379 32899 32385
rect 36354 32376 36360 32388
rect 36412 32376 36418 32428
rect 46382 32416 46388 32428
rect 46343 32388 46388 32416
rect 46382 32376 46388 32388
rect 46440 32376 46446 32428
rect 32548 32320 32720 32348
rect 37277 32351 37335 32357
rect 32548 32308 32554 32320
rect 37277 32317 37289 32351
rect 37323 32317 37335 32351
rect 37458 32348 37464 32360
rect 37419 32320 37464 32348
rect 37277 32311 37335 32317
rect 28868 32252 31432 32280
rect 28868 32240 28874 32252
rect 21450 32212 21456 32224
rect 20732 32184 21456 32212
rect 20165 32175 20223 32181
rect 21450 32172 21456 32184
rect 21508 32172 21514 32224
rect 21913 32215 21971 32221
rect 21913 32181 21925 32215
rect 21959 32212 21971 32215
rect 22554 32212 22560 32224
rect 21959 32184 22560 32212
rect 21959 32181 21971 32184
rect 21913 32175 21971 32181
rect 22554 32172 22560 32184
rect 22612 32172 22618 32224
rect 22830 32172 22836 32224
rect 22888 32212 22894 32224
rect 23198 32212 23204 32224
rect 22888 32184 23204 32212
rect 22888 32172 22894 32184
rect 23198 32172 23204 32184
rect 23256 32172 23262 32224
rect 23474 32172 23480 32224
rect 23532 32212 23538 32224
rect 24486 32212 24492 32224
rect 23532 32184 24492 32212
rect 23532 32172 23538 32184
rect 24486 32172 24492 32184
rect 24544 32172 24550 32224
rect 25685 32215 25743 32221
rect 25685 32181 25697 32215
rect 25731 32212 25743 32215
rect 25774 32212 25780 32224
rect 25731 32184 25780 32212
rect 25731 32181 25743 32184
rect 25685 32175 25743 32181
rect 25774 32172 25780 32184
rect 25832 32172 25838 32224
rect 26252 32212 26280 32240
rect 28350 32212 28356 32224
rect 26252 32184 28356 32212
rect 28350 32172 28356 32184
rect 28408 32172 28414 32224
rect 32030 32172 32036 32224
rect 32088 32212 32094 32224
rect 37292 32212 37320 32311
rect 37458 32308 37464 32320
rect 37516 32308 37522 32360
rect 46198 32308 46204 32360
rect 46256 32348 46262 32360
rect 46661 32351 46719 32357
rect 46661 32348 46673 32351
rect 46256 32320 46673 32348
rect 46256 32308 46262 32320
rect 46661 32317 46673 32320
rect 46707 32317 46719 32351
rect 46661 32311 46719 32317
rect 32088 32184 37320 32212
rect 32088 32172 32094 32184
rect 1104 32122 48852 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 48852 32122
rect 1104 32048 48852 32070
rect 15562 31968 15568 32020
rect 15620 32008 15626 32020
rect 16669 32011 16727 32017
rect 16669 32008 16681 32011
rect 15620 31980 16681 32008
rect 15620 31968 15626 31980
rect 16669 31977 16681 31980
rect 16715 31977 16727 32011
rect 16669 31971 16727 31977
rect 16850 31968 16856 32020
rect 16908 32008 16914 32020
rect 22186 32008 22192 32020
rect 16908 31980 22192 32008
rect 16908 31968 16914 31980
rect 22186 31968 22192 31980
rect 22244 32008 22250 32020
rect 23014 32008 23020 32020
rect 22244 31980 23020 32008
rect 22244 31968 22250 31980
rect 23014 31968 23020 31980
rect 23072 31968 23078 32020
rect 23934 31968 23940 32020
rect 23992 32008 23998 32020
rect 27065 32011 27123 32017
rect 23992 31980 25084 32008
rect 23992 31968 23998 31980
rect 21174 31940 21180 31952
rect 21135 31912 21180 31940
rect 21174 31900 21180 31912
rect 21232 31900 21238 31952
rect 22370 31940 22376 31952
rect 22283 31912 22376 31940
rect 22370 31900 22376 31912
rect 22428 31940 22434 31952
rect 23566 31940 23572 31952
rect 22428 31912 23572 31940
rect 22428 31900 22434 31912
rect 23566 31900 23572 31912
rect 23624 31940 23630 31952
rect 23624 31912 24808 31940
rect 23624 31900 23630 31912
rect 1581 31875 1639 31881
rect 1581 31841 1593 31875
rect 1627 31872 1639 31875
rect 2774 31872 2780 31884
rect 1627 31844 2780 31872
rect 1627 31841 1639 31844
rect 1581 31835 1639 31841
rect 2774 31832 2780 31844
rect 2832 31832 2838 31884
rect 2866 31832 2872 31884
rect 2924 31872 2930 31884
rect 2924 31844 2969 31872
rect 2924 31832 2930 31844
rect 19334 31832 19340 31884
rect 19392 31832 19398 31884
rect 20806 31832 20812 31884
rect 20864 31872 20870 31884
rect 23290 31872 23296 31884
rect 20864 31844 23296 31872
rect 20864 31832 20870 31844
rect 23290 31832 23296 31844
rect 23348 31832 23354 31884
rect 1397 31807 1455 31813
rect 1397 31773 1409 31807
rect 1443 31773 1455 31807
rect 1397 31767 1455 31773
rect 15289 31807 15347 31813
rect 15289 31773 15301 31807
rect 15335 31804 15347 31807
rect 16574 31804 16580 31816
rect 15335 31776 16580 31804
rect 15335 31773 15347 31776
rect 15289 31767 15347 31773
rect 1412 31736 1440 31767
rect 16574 31764 16580 31776
rect 16632 31804 16638 31816
rect 17129 31807 17187 31813
rect 17129 31804 17141 31807
rect 16632 31776 17141 31804
rect 16632 31764 16638 31776
rect 17129 31773 17141 31776
rect 17175 31804 17187 31807
rect 19352 31804 19380 31832
rect 19797 31807 19855 31813
rect 19797 31804 19809 31807
rect 17175 31776 19809 31804
rect 17175 31773 17187 31776
rect 17129 31767 17187 31773
rect 19797 31773 19809 31776
rect 19843 31804 19855 31807
rect 21818 31804 21824 31816
rect 19843 31776 21824 31804
rect 19843 31773 19855 31776
rect 19797 31767 19855 31773
rect 21818 31764 21824 31776
rect 21876 31764 21882 31816
rect 22189 31807 22247 31813
rect 22189 31773 22201 31807
rect 22235 31804 22247 31807
rect 22278 31804 22284 31816
rect 22235 31776 22284 31804
rect 22235 31773 22247 31776
rect 22189 31767 22247 31773
rect 22278 31764 22284 31776
rect 22336 31764 22342 31816
rect 23474 31764 23480 31816
rect 23532 31804 23538 31816
rect 23532 31776 23577 31804
rect 23532 31764 23538 31776
rect 24118 31764 24124 31816
rect 24176 31804 24182 31816
rect 24780 31813 24808 31912
rect 24673 31807 24731 31813
rect 24673 31804 24685 31807
rect 24176 31776 24685 31804
rect 24176 31764 24182 31776
rect 24673 31773 24685 31776
rect 24719 31773 24731 31807
rect 24673 31767 24731 31773
rect 24765 31807 24823 31813
rect 24765 31773 24777 31807
rect 24811 31773 24823 31807
rect 24765 31767 24823 31773
rect 24854 31764 24860 31816
rect 24912 31804 24918 31816
rect 25056 31813 25084 31980
rect 27065 31977 27077 32011
rect 27111 32008 27123 32011
rect 27430 32008 27436 32020
rect 27111 31980 27436 32008
rect 27111 31977 27123 31980
rect 27065 31971 27123 31977
rect 27430 31968 27436 31980
rect 27488 31968 27494 32020
rect 27706 31968 27712 32020
rect 27764 32008 27770 32020
rect 35713 32011 35771 32017
rect 27764 31980 32812 32008
rect 27764 31968 27770 31980
rect 26605 31943 26663 31949
rect 26605 31940 26617 31943
rect 26160 31912 26617 31940
rect 25041 31807 25099 31813
rect 24912 31776 24957 31804
rect 24912 31764 24918 31776
rect 25041 31773 25053 31807
rect 25087 31773 25099 31807
rect 25041 31767 25099 31773
rect 25222 31764 25228 31816
rect 25280 31804 25286 31816
rect 25685 31807 25743 31813
rect 25280 31776 25636 31804
rect 25280 31764 25286 31776
rect 2038 31736 2044 31748
rect 1412 31708 2044 31736
rect 2038 31696 2044 31708
rect 2096 31696 2102 31748
rect 15556 31739 15614 31745
rect 15556 31705 15568 31739
rect 15602 31736 15614 31739
rect 15654 31736 15660 31748
rect 15602 31708 15660 31736
rect 15602 31705 15614 31708
rect 15556 31699 15614 31705
rect 15654 31696 15660 31708
rect 15712 31696 15718 31748
rect 16850 31696 16856 31748
rect 16908 31736 16914 31748
rect 20070 31745 20076 31748
rect 17374 31739 17432 31745
rect 17374 31736 17386 31739
rect 16908 31708 17386 31736
rect 16908 31696 16914 31708
rect 17374 31705 17386 31708
rect 17420 31705 17432 31739
rect 17374 31699 17432 31705
rect 20064 31699 20076 31745
rect 20128 31736 20134 31748
rect 20128 31708 20164 31736
rect 20070 31696 20076 31699
rect 20128 31696 20134 31708
rect 23014 31696 23020 31748
rect 23072 31736 23078 31748
rect 23293 31739 23351 31745
rect 23293 31736 23305 31739
rect 23072 31708 23305 31736
rect 23072 31696 23078 31708
rect 23293 31705 23305 31708
rect 23339 31705 23351 31739
rect 25608 31736 25636 31776
rect 25685 31773 25697 31807
rect 25731 31804 25743 31807
rect 26160 31804 26188 31912
rect 26605 31909 26617 31912
rect 26651 31940 26663 31943
rect 27338 31940 27344 31952
rect 26651 31912 27344 31940
rect 26651 31909 26663 31912
rect 26605 31903 26663 31909
rect 27338 31900 27344 31912
rect 27396 31940 27402 31952
rect 32030 31940 32036 31952
rect 27396 31912 32036 31940
rect 27396 31900 27402 31912
rect 27338 31804 27344 31816
rect 25731 31776 26188 31804
rect 27299 31776 27344 31804
rect 25731 31773 25743 31776
rect 25685 31767 25743 31773
rect 27338 31764 27344 31776
rect 27396 31764 27402 31816
rect 27448 31813 27476 31912
rect 32030 31900 32036 31912
rect 32088 31900 32094 31952
rect 32398 31940 32404 31952
rect 32359 31912 32404 31940
rect 32398 31900 32404 31912
rect 32456 31900 32462 31952
rect 32784 31940 32812 31980
rect 35713 31977 35725 32011
rect 35759 32008 35771 32011
rect 37458 32008 37464 32020
rect 35759 31980 37464 32008
rect 35759 31977 35771 31980
rect 35713 31971 35771 31977
rect 37458 31968 37464 31980
rect 37516 31968 37522 32020
rect 46474 31968 46480 32020
rect 46532 32008 46538 32020
rect 46753 32011 46811 32017
rect 46753 32008 46765 32011
rect 46532 31980 46765 32008
rect 46532 31968 46538 31980
rect 46753 31977 46765 31980
rect 46799 31977 46811 32011
rect 46753 31971 46811 31977
rect 32524 31912 32720 31940
rect 32784 31912 32884 31940
rect 28537 31875 28595 31881
rect 28537 31872 28549 31875
rect 27540 31844 28549 31872
rect 27540 31813 27568 31844
rect 28537 31841 28549 31844
rect 28583 31841 28595 31875
rect 32048 31872 32076 31900
rect 32524 31872 32552 31912
rect 32048 31844 32552 31872
rect 32692 31872 32720 31912
rect 32856 31872 32884 31912
rect 33226 31872 33232 31884
rect 32692 31844 32809 31872
rect 32856 31844 33232 31872
rect 28537 31835 28595 31841
rect 27433 31807 27491 31813
rect 27433 31773 27445 31807
rect 27479 31773 27491 31807
rect 27433 31767 27491 31773
rect 27525 31807 27583 31813
rect 27525 31773 27537 31807
rect 27571 31773 27583 31807
rect 27706 31804 27712 31816
rect 27667 31776 27712 31804
rect 27525 31767 27583 31773
rect 27706 31764 27712 31776
rect 27764 31764 27770 31816
rect 28166 31804 28172 31816
rect 28127 31776 28172 31804
rect 28166 31764 28172 31776
rect 28224 31764 28230 31816
rect 28350 31804 28356 31816
rect 28311 31776 28356 31804
rect 28350 31764 28356 31776
rect 28408 31764 28414 31816
rect 28460 31776 31064 31804
rect 26421 31739 26479 31745
rect 26421 31736 26433 31739
rect 23293 31699 23351 31705
rect 23400 31708 24624 31736
rect 25608 31708 26433 31736
rect 18506 31668 18512 31680
rect 18467 31640 18512 31668
rect 18506 31628 18512 31640
rect 18564 31628 18570 31680
rect 21726 31628 21732 31680
rect 21784 31668 21790 31680
rect 22186 31668 22192 31680
rect 21784 31640 22192 31668
rect 21784 31628 21790 31640
rect 22186 31628 22192 31640
rect 22244 31668 22250 31680
rect 23400 31668 23428 31708
rect 22244 31640 23428 31668
rect 24397 31671 24455 31677
rect 22244 31628 22250 31640
rect 24397 31637 24409 31671
rect 24443 31668 24455 31671
rect 24486 31668 24492 31680
rect 24443 31640 24492 31668
rect 24443 31637 24455 31640
rect 24397 31631 24455 31637
rect 24486 31628 24492 31640
rect 24544 31628 24550 31680
rect 24596 31668 24624 31708
rect 26421 31705 26433 31708
rect 26467 31736 26479 31739
rect 26602 31736 26608 31748
rect 26467 31708 26608 31736
rect 26467 31705 26479 31708
rect 26421 31699 26479 31705
rect 26602 31696 26608 31708
rect 26660 31696 26666 31748
rect 27246 31696 27252 31748
rect 27304 31736 27310 31748
rect 28460 31736 28488 31776
rect 27304 31708 28488 31736
rect 31036 31736 31064 31776
rect 31110 31764 31116 31816
rect 31168 31804 31174 31816
rect 31573 31807 31631 31813
rect 31573 31804 31585 31807
rect 31168 31776 31585 31804
rect 31168 31764 31174 31776
rect 31573 31773 31585 31776
rect 31619 31773 31631 31807
rect 31573 31767 31631 31773
rect 31754 31764 31760 31816
rect 31812 31804 31818 31816
rect 32677 31807 32735 31813
rect 32781 31810 32809 31844
rect 31812 31776 31857 31804
rect 31812 31764 31818 31776
rect 32677 31773 32689 31807
rect 32723 31773 32735 31807
rect 32677 31767 32735 31773
rect 32766 31804 32824 31810
rect 32766 31770 32778 31804
rect 32812 31770 32824 31804
rect 32122 31736 32128 31748
rect 31036 31708 32128 31736
rect 27304 31696 27310 31708
rect 32122 31696 32128 31708
rect 32180 31696 32186 31748
rect 32692 31736 32720 31767
rect 32766 31764 32824 31770
rect 32861 31807 32919 31813
rect 32861 31773 32873 31807
rect 32907 31804 32919 31807
rect 32950 31804 32956 31816
rect 32907 31776 32956 31804
rect 32907 31773 32919 31776
rect 32861 31767 32919 31773
rect 32950 31764 32956 31776
rect 33008 31764 33014 31816
rect 33060 31813 33088 31844
rect 33226 31832 33232 31844
rect 33284 31872 33290 31884
rect 34054 31872 34060 31884
rect 33284 31844 34060 31872
rect 33284 31832 33290 31844
rect 34054 31832 34060 31844
rect 34112 31832 34118 31884
rect 38562 31872 38568 31884
rect 38523 31844 38568 31872
rect 38562 31832 38568 31844
rect 38620 31832 38626 31884
rect 46566 31832 46572 31884
rect 46624 31872 46630 31884
rect 47581 31875 47639 31881
rect 47581 31872 47593 31875
rect 46624 31844 47593 31872
rect 46624 31832 46630 31844
rect 47581 31841 47593 31844
rect 47627 31841 47639 31875
rect 47581 31835 47639 31841
rect 33045 31807 33103 31813
rect 33045 31773 33057 31807
rect 33091 31773 33103 31807
rect 33594 31804 33600 31816
rect 33555 31776 33600 31804
rect 33045 31767 33103 31773
rect 33594 31764 33600 31776
rect 33652 31764 33658 31816
rect 35621 31807 35679 31813
rect 35621 31773 35633 31807
rect 35667 31804 35679 31807
rect 35894 31804 35900 31816
rect 35667 31776 35900 31804
rect 35667 31773 35679 31776
rect 35621 31767 35679 31773
rect 35894 31764 35900 31776
rect 35952 31764 35958 31816
rect 36265 31807 36323 31813
rect 36265 31773 36277 31807
rect 36311 31804 36323 31807
rect 36354 31804 36360 31816
rect 36311 31776 36360 31804
rect 36311 31773 36323 31776
rect 36265 31767 36323 31773
rect 36354 31764 36360 31776
rect 36412 31764 36418 31816
rect 36541 31807 36599 31813
rect 36541 31773 36553 31807
rect 36587 31804 36599 31807
rect 36630 31804 36636 31816
rect 36587 31776 36636 31804
rect 36587 31773 36599 31776
rect 36541 31767 36599 31773
rect 36630 31764 36636 31776
rect 36688 31764 36694 31816
rect 37182 31804 37188 31816
rect 37143 31776 37188 31804
rect 37182 31764 37188 31776
rect 37240 31764 37246 31816
rect 45462 31764 45468 31816
rect 45520 31804 45526 31816
rect 46661 31807 46719 31813
rect 46661 31804 46673 31807
rect 45520 31776 46673 31804
rect 45520 31764 45526 31776
rect 46661 31773 46673 31776
rect 46707 31773 46719 31807
rect 46661 31767 46719 31773
rect 47305 31807 47363 31813
rect 47305 31773 47317 31807
rect 47351 31804 47363 31807
rect 47394 31804 47400 31816
rect 47351 31776 47400 31804
rect 47351 31773 47363 31776
rect 47305 31767 47363 31773
rect 47394 31764 47400 31776
rect 47452 31764 47458 31816
rect 33778 31736 33784 31748
rect 32692 31708 33088 31736
rect 33739 31708 33784 31736
rect 33060 31680 33088 31708
rect 33778 31696 33784 31708
rect 33836 31696 33842 31748
rect 37366 31736 37372 31748
rect 37327 31708 37372 31736
rect 37366 31696 37372 31708
rect 37424 31696 37430 31748
rect 25777 31671 25835 31677
rect 25777 31668 25789 31671
rect 24596 31640 25789 31668
rect 25777 31637 25789 31640
rect 25823 31637 25835 31671
rect 25777 31631 25835 31637
rect 31941 31671 31999 31677
rect 31941 31637 31953 31671
rect 31987 31668 31999 31671
rect 32950 31668 32956 31680
rect 31987 31640 32956 31668
rect 31987 31637 31999 31640
rect 31941 31631 31999 31637
rect 32950 31628 32956 31640
rect 33008 31628 33014 31680
rect 33042 31628 33048 31680
rect 33100 31628 33106 31680
rect 35802 31628 35808 31680
rect 35860 31668 35866 31680
rect 46198 31668 46204 31680
rect 35860 31640 46204 31668
rect 35860 31628 35866 31640
rect 46198 31628 46204 31640
rect 46256 31628 46262 31680
rect 1104 31578 48852 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 48852 31578
rect 1104 31504 48852 31526
rect 2774 31464 2780 31476
rect 2735 31436 2780 31464
rect 2774 31424 2780 31436
rect 2832 31424 2838 31476
rect 16850 31464 16856 31476
rect 16811 31436 16856 31464
rect 16850 31424 16856 31436
rect 16908 31424 16914 31476
rect 16960 31436 18092 31464
rect 16960 31396 16988 31436
rect 17954 31396 17960 31408
rect 1688 31368 16988 31396
rect 17328 31368 17960 31396
rect 1394 31328 1400 31340
rect 1355 31300 1400 31328
rect 1394 31288 1400 31300
rect 1452 31288 1458 31340
rect 1688 31337 1716 31368
rect 1673 31331 1731 31337
rect 1673 31297 1685 31331
rect 1719 31297 1731 31331
rect 1673 31291 1731 31297
rect 1762 31288 1768 31340
rect 1820 31328 1826 31340
rect 2685 31331 2743 31337
rect 2685 31328 2697 31331
rect 1820 31300 2697 31328
rect 1820 31288 1826 31300
rect 2685 31297 2697 31300
rect 2731 31297 2743 31331
rect 2685 31291 2743 31297
rect 3694 31288 3700 31340
rect 3752 31328 3758 31340
rect 17328 31337 17356 31368
rect 17954 31356 17960 31368
rect 18012 31356 18018 31408
rect 18064 31396 18092 31436
rect 18230 31424 18236 31476
rect 18288 31464 18294 31476
rect 18509 31467 18567 31473
rect 18509 31464 18521 31467
rect 18288 31436 18521 31464
rect 18288 31424 18294 31436
rect 18509 31433 18521 31436
rect 18555 31433 18567 31467
rect 18509 31427 18567 31433
rect 18969 31467 19027 31473
rect 18969 31433 18981 31467
rect 19015 31464 19027 31467
rect 19426 31464 19432 31476
rect 19015 31436 19432 31464
rect 19015 31433 19027 31436
rect 18969 31427 19027 31433
rect 19426 31424 19432 31436
rect 19484 31424 19490 31476
rect 20162 31424 20168 31476
rect 20220 31464 20226 31476
rect 20622 31464 20628 31476
rect 20220 31436 20628 31464
rect 20220 31424 20226 31436
rect 20622 31424 20628 31436
rect 20680 31424 20686 31476
rect 28442 31464 28448 31476
rect 20732 31436 25912 31464
rect 28403 31436 28448 31464
rect 20732 31405 20760 31436
rect 20257 31399 20315 31405
rect 18064 31368 19012 31396
rect 17129 31331 17187 31337
rect 17129 31328 17141 31331
rect 3752 31300 17141 31328
rect 3752 31288 3758 31300
rect 17129 31297 17141 31300
rect 17175 31297 17187 31331
rect 17129 31291 17187 31297
rect 17221 31331 17279 31337
rect 17221 31297 17233 31331
rect 17267 31297 17279 31331
rect 17221 31291 17279 31297
rect 17313 31331 17371 31337
rect 17313 31297 17325 31331
rect 17359 31297 17371 31331
rect 17494 31328 17500 31340
rect 17455 31300 17500 31328
rect 17313 31291 17371 31297
rect 17236 31260 17264 31291
rect 17494 31288 17500 31300
rect 17552 31288 17558 31340
rect 18506 31288 18512 31340
rect 18564 31328 18570 31340
rect 18877 31331 18935 31337
rect 18877 31328 18889 31331
rect 18564 31300 18889 31328
rect 18564 31288 18570 31300
rect 18877 31297 18889 31300
rect 18923 31297 18935 31331
rect 18984 31328 19012 31368
rect 20257 31365 20269 31399
rect 20303 31396 20315 31399
rect 20717 31399 20775 31405
rect 20717 31396 20729 31399
rect 20303 31368 20729 31396
rect 20303 31365 20315 31368
rect 20257 31359 20315 31365
rect 20717 31365 20729 31368
rect 20763 31365 20775 31399
rect 20717 31359 20775 31365
rect 21910 31356 21916 31408
rect 21968 31396 21974 31408
rect 22370 31396 22376 31408
rect 21968 31368 22376 31396
rect 21968 31356 21974 31368
rect 22370 31356 22376 31368
rect 22428 31356 22434 31408
rect 23201 31399 23259 31405
rect 23201 31365 23213 31399
rect 23247 31396 23259 31399
rect 23474 31396 23480 31408
rect 23247 31368 23480 31396
rect 23247 31365 23259 31368
rect 23201 31359 23259 31365
rect 23474 31356 23480 31368
rect 23532 31356 23538 31408
rect 20533 31331 20591 31337
rect 20533 31328 20545 31331
rect 18984 31300 20545 31328
rect 18877 31291 18935 31297
rect 20533 31297 20545 31300
rect 20579 31297 20591 31331
rect 22281 31331 22339 31337
rect 22281 31328 22293 31331
rect 20533 31291 20591 31297
rect 22066 31300 22293 31328
rect 17586 31260 17592 31272
rect 17236 31232 17592 31260
rect 17586 31220 17592 31232
rect 17644 31220 17650 31272
rect 18892 31192 18920 31291
rect 19150 31260 19156 31272
rect 19111 31232 19156 31260
rect 19150 31220 19156 31232
rect 19208 31220 19214 31272
rect 20714 31220 20720 31272
rect 20772 31260 20778 31272
rect 22066 31260 22094 31300
rect 22281 31297 22293 31300
rect 22327 31328 22339 31331
rect 25038 31328 25044 31340
rect 22327 31300 25044 31328
rect 22327 31297 22339 31300
rect 22281 31291 22339 31297
rect 25038 31288 25044 31300
rect 25096 31288 25102 31340
rect 25133 31331 25191 31337
rect 25133 31297 25145 31331
rect 25179 31328 25191 31331
rect 25774 31328 25780 31340
rect 25179 31300 25780 31328
rect 25179 31297 25191 31300
rect 25133 31291 25191 31297
rect 25774 31288 25780 31300
rect 25832 31288 25838 31340
rect 20772 31232 22094 31260
rect 20772 31220 20778 31232
rect 23382 31220 23388 31272
rect 23440 31260 23446 31272
rect 24210 31260 24216 31272
rect 23440 31232 24216 31260
rect 23440 31220 23446 31232
rect 24210 31220 24216 31232
rect 24268 31220 24274 31272
rect 25884 31260 25912 31436
rect 28442 31424 28448 31436
rect 28500 31464 28506 31476
rect 29730 31464 29736 31476
rect 28500 31436 28856 31464
rect 28500 31424 28506 31436
rect 26970 31356 26976 31408
rect 27028 31396 27034 31408
rect 27801 31399 27859 31405
rect 27801 31396 27813 31399
rect 27028 31368 27813 31396
rect 27028 31356 27034 31368
rect 27801 31365 27813 31368
rect 27847 31365 27859 31399
rect 27801 31359 27859 31365
rect 27982 31356 27988 31408
rect 28040 31405 28046 31408
rect 28828 31405 28856 31436
rect 29012 31436 29736 31464
rect 29012 31405 29040 31436
rect 29730 31424 29736 31436
rect 29788 31424 29794 31476
rect 31018 31424 31024 31476
rect 31076 31464 31082 31476
rect 31481 31467 31539 31473
rect 31481 31464 31493 31467
rect 31076 31436 31493 31464
rect 31076 31424 31082 31436
rect 31481 31433 31493 31436
rect 31527 31433 31539 31467
rect 31481 31427 31539 31433
rect 32401 31467 32459 31473
rect 32401 31433 32413 31467
rect 32447 31464 32459 31467
rect 32490 31464 32496 31476
rect 32447 31436 32496 31464
rect 32447 31433 32459 31436
rect 32401 31427 32459 31433
rect 32490 31424 32496 31436
rect 32548 31424 32554 31476
rect 37366 31464 37372 31476
rect 32600 31436 32873 31464
rect 37327 31436 37372 31464
rect 28040 31399 28059 31405
rect 28047 31365 28059 31399
rect 28040 31359 28059 31365
rect 28813 31399 28871 31405
rect 28813 31365 28825 31399
rect 28859 31365 28871 31399
rect 29012 31399 29071 31405
rect 29012 31396 29025 31399
rect 28813 31359 28871 31365
rect 28920 31368 29025 31396
rect 28040 31356 28046 31359
rect 28016 31328 28044 31356
rect 28920 31328 28948 31368
rect 29013 31365 29025 31368
rect 29059 31365 29071 31399
rect 32600 31396 32628 31436
rect 29013 31359 29071 31365
rect 29656 31368 32628 31396
rect 32845 31396 32873 31436
rect 37366 31424 37372 31436
rect 37424 31424 37430 31476
rect 39758 31396 39764 31408
rect 32845 31368 39344 31396
rect 39719 31368 39764 31396
rect 28016 31300 28948 31328
rect 29656 31260 29684 31368
rect 29917 31331 29975 31337
rect 29917 31297 29929 31331
rect 29963 31328 29975 31331
rect 31294 31328 31300 31340
rect 29963 31300 31300 31328
rect 29963 31297 29975 31300
rect 29917 31291 29975 31297
rect 31294 31288 31300 31300
rect 31352 31288 31358 31340
rect 31386 31288 31392 31340
rect 31444 31328 31450 31340
rect 31444 31300 31489 31328
rect 31444 31288 31450 31300
rect 32582 31288 32588 31340
rect 32640 31331 32646 31340
rect 32677 31331 32735 31337
rect 32640 31303 32689 31331
rect 32640 31288 32646 31303
rect 32677 31297 32689 31303
rect 32723 31297 32735 31331
rect 32677 31291 32735 31297
rect 32769 31331 32827 31337
rect 32769 31297 32781 31331
rect 32815 31297 32827 31331
rect 32769 31291 32827 31297
rect 29822 31260 29828 31272
rect 25884 31232 29684 31260
rect 29783 31232 29828 31260
rect 29822 31220 29828 31232
rect 29880 31220 29886 31272
rect 30006 31260 30012 31272
rect 29967 31232 30012 31260
rect 30006 31220 30012 31232
rect 30064 31220 30070 31272
rect 30101 31263 30159 31269
rect 30101 31229 30113 31263
rect 30147 31229 30159 31263
rect 30101 31223 30159 31229
rect 20162 31192 20168 31204
rect 18892 31164 20168 31192
rect 20162 31152 20168 31164
rect 20220 31152 20226 31204
rect 26970 31192 26976 31204
rect 20640 31164 26976 31192
rect 15010 31084 15016 31136
rect 15068 31124 15074 31136
rect 20640 31124 20668 31164
rect 26970 31152 26976 31164
rect 27028 31152 27034 31204
rect 28169 31195 28227 31201
rect 28169 31161 28181 31195
rect 28215 31192 28227 31195
rect 30116 31192 30144 31223
rect 32030 31220 32036 31272
rect 32088 31260 32094 31272
rect 32784 31260 32812 31291
rect 32858 31288 32864 31340
rect 32916 31328 32922 31340
rect 33045 31331 33103 31337
rect 33226 31331 33232 31340
rect 32916 31300 32961 31328
rect 32916 31288 32922 31300
rect 33045 31297 33057 31331
rect 33091 31303 33232 31331
rect 33091 31297 33103 31303
rect 33045 31291 33103 31297
rect 33226 31288 33232 31303
rect 33284 31288 33290 31340
rect 35986 31288 35992 31340
rect 36044 31328 36050 31340
rect 37277 31331 37335 31337
rect 37277 31328 37289 31331
rect 36044 31300 37289 31328
rect 36044 31288 36050 31300
rect 37277 31297 37289 31300
rect 37323 31297 37335 31331
rect 39316 31328 39344 31368
rect 39758 31356 39764 31368
rect 39816 31356 39822 31408
rect 43898 31328 43904 31340
rect 39316 31300 43904 31328
rect 37277 31291 37335 31297
rect 43898 31288 43904 31300
rect 43956 31288 43962 31340
rect 32088 31232 32812 31260
rect 32088 31220 32094 31232
rect 35342 31220 35348 31272
rect 35400 31260 35406 31272
rect 35802 31260 35808 31272
rect 35400 31232 35808 31260
rect 35400 31220 35406 31232
rect 35802 31220 35808 31232
rect 35860 31260 35866 31272
rect 35897 31263 35955 31269
rect 35897 31260 35909 31263
rect 35860 31232 35909 31260
rect 35860 31220 35866 31232
rect 35897 31229 35909 31232
rect 35943 31229 35955 31263
rect 35897 31223 35955 31229
rect 36173 31263 36231 31269
rect 36173 31229 36185 31263
rect 36219 31260 36231 31263
rect 36262 31260 36268 31272
rect 36219 31232 36268 31260
rect 36219 31229 36231 31232
rect 36173 31223 36231 31229
rect 36262 31220 36268 31232
rect 36320 31260 36326 31272
rect 36538 31260 36544 31272
rect 36320 31232 36544 31260
rect 36320 31220 36326 31232
rect 36538 31220 36544 31232
rect 36596 31220 36602 31272
rect 37921 31263 37979 31269
rect 37921 31229 37933 31263
rect 37967 31229 37979 31263
rect 38102 31260 38108 31272
rect 38063 31232 38108 31260
rect 37921 31223 37979 31229
rect 28215 31164 30144 31192
rect 37936 31192 37964 31223
rect 38102 31220 38108 31232
rect 38160 31220 38166 31272
rect 38010 31192 38016 31204
rect 37936 31164 38016 31192
rect 28215 31161 28227 31164
rect 28169 31155 28227 31161
rect 38010 31152 38016 31164
rect 38068 31152 38074 31204
rect 15068 31096 20668 31124
rect 15068 31084 15074 31096
rect 20714 31084 20720 31136
rect 20772 31124 20778 31136
rect 20901 31127 20959 31133
rect 20901 31124 20913 31127
rect 20772 31096 20913 31124
rect 20772 31084 20778 31096
rect 20901 31093 20913 31096
rect 20947 31093 20959 31127
rect 20901 31087 20959 31093
rect 21082 31084 21088 31136
rect 21140 31124 21146 31136
rect 22373 31127 22431 31133
rect 22373 31124 22385 31127
rect 21140 31096 22385 31124
rect 21140 31084 21146 31096
rect 22373 31093 22385 31096
rect 22419 31124 22431 31127
rect 22554 31124 22560 31136
rect 22419 31096 22560 31124
rect 22419 31093 22431 31096
rect 22373 31087 22431 31093
rect 22554 31084 22560 31096
rect 22612 31084 22618 31136
rect 23293 31127 23351 31133
rect 23293 31093 23305 31127
rect 23339 31124 23351 31127
rect 23382 31124 23388 31136
rect 23339 31096 23388 31124
rect 23339 31093 23351 31096
rect 23293 31087 23351 31093
rect 23382 31084 23388 31096
rect 23440 31084 23446 31136
rect 24578 31084 24584 31136
rect 24636 31124 24642 31136
rect 24949 31127 25007 31133
rect 24949 31124 24961 31127
rect 24636 31096 24961 31124
rect 24636 31084 24642 31096
rect 24949 31093 24961 31096
rect 24995 31093 25007 31127
rect 24949 31087 25007 31093
rect 27985 31127 28043 31133
rect 27985 31093 27997 31127
rect 28031 31124 28043 31127
rect 28902 31124 28908 31136
rect 28031 31096 28908 31124
rect 28031 31093 28043 31096
rect 27985 31087 28043 31093
rect 28902 31084 28908 31096
rect 28960 31124 28966 31136
rect 28997 31127 29055 31133
rect 28997 31124 29009 31127
rect 28960 31096 29009 31124
rect 28960 31084 28966 31096
rect 28997 31093 29009 31096
rect 29043 31093 29055 31127
rect 29178 31124 29184 31136
rect 29139 31096 29184 31124
rect 28997 31087 29055 31093
rect 29178 31084 29184 31096
rect 29236 31084 29242 31136
rect 29641 31127 29699 31133
rect 29641 31093 29653 31127
rect 29687 31124 29699 31127
rect 30006 31124 30012 31136
rect 29687 31096 30012 31124
rect 29687 31093 29699 31096
rect 29641 31087 29699 31093
rect 30006 31084 30012 31096
rect 30064 31084 30070 31136
rect 35342 31084 35348 31136
rect 35400 31124 35406 31136
rect 35529 31127 35587 31133
rect 35529 31124 35541 31127
rect 35400 31096 35541 31124
rect 35400 31084 35406 31096
rect 35529 31093 35541 31096
rect 35575 31093 35587 31127
rect 35529 31087 35587 31093
rect 35618 31084 35624 31136
rect 35676 31124 35682 31136
rect 46566 31124 46572 31136
rect 35676 31096 46572 31124
rect 35676 31084 35682 31096
rect 46566 31084 46572 31096
rect 46624 31084 46630 31136
rect 1104 31034 48852 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 48852 31034
rect 1104 30960 48852 30982
rect 2038 30920 2044 30932
rect 1999 30892 2044 30920
rect 2038 30880 2044 30892
rect 2096 30880 2102 30932
rect 17494 30880 17500 30932
rect 17552 30920 17558 30932
rect 20990 30920 20996 30932
rect 17552 30892 20996 30920
rect 17552 30880 17558 30892
rect 20990 30880 20996 30892
rect 21048 30880 21054 30932
rect 21634 30880 21640 30932
rect 21692 30920 21698 30932
rect 27338 30920 27344 30932
rect 21692 30892 27344 30920
rect 21692 30880 21698 30892
rect 27338 30880 27344 30892
rect 27396 30880 27402 30932
rect 28994 30920 29000 30932
rect 28955 30892 29000 30920
rect 28994 30880 29000 30892
rect 29052 30880 29058 30932
rect 31294 30920 31300 30932
rect 31255 30892 31300 30920
rect 31294 30880 31300 30892
rect 31352 30880 31358 30932
rect 38013 30923 38071 30929
rect 38013 30889 38025 30923
rect 38059 30920 38071 30923
rect 38102 30920 38108 30932
rect 38059 30892 38108 30920
rect 38059 30889 38071 30892
rect 38013 30883 38071 30889
rect 38102 30880 38108 30892
rect 38160 30880 38166 30932
rect 17957 30855 18015 30861
rect 17957 30821 17969 30855
rect 18003 30852 18015 30855
rect 18414 30852 18420 30864
rect 18003 30824 18420 30852
rect 18003 30821 18015 30824
rect 17957 30815 18015 30821
rect 18414 30812 18420 30824
rect 18472 30812 18478 30864
rect 21726 30852 21732 30864
rect 20921 30824 21732 30852
rect 16574 30784 16580 30796
rect 16535 30756 16580 30784
rect 16574 30744 16580 30756
rect 16632 30744 16638 30796
rect 17586 30744 17592 30796
rect 17644 30784 17650 30796
rect 20921 30784 20949 30824
rect 21726 30812 21732 30824
rect 21784 30812 21790 30864
rect 22002 30812 22008 30864
rect 22060 30852 22066 30864
rect 22060 30824 22968 30852
rect 22060 30812 22066 30824
rect 17644 30756 20949 30784
rect 17644 30744 17650 30756
rect 19334 30676 19340 30728
rect 19392 30716 19398 30728
rect 19978 30716 19984 30728
rect 19392 30688 19984 30716
rect 19392 30676 19398 30688
rect 19978 30676 19984 30688
rect 20036 30676 20042 30728
rect 20921 30725 20949 30756
rect 21008 30756 21404 30784
rect 21008 30725 21036 30756
rect 20789 30719 20847 30725
rect 20789 30685 20801 30719
rect 20835 30716 20847 30719
rect 20898 30719 20956 30725
rect 20835 30685 20852 30716
rect 20789 30679 20852 30685
rect 20898 30685 20910 30719
rect 20944 30685 20956 30719
rect 20898 30679 20956 30685
rect 20993 30719 21051 30725
rect 20993 30685 21005 30719
rect 21039 30685 21051 30719
rect 20993 30679 21051 30685
rect 16666 30608 16672 30660
rect 16724 30648 16730 30660
rect 16822 30651 16880 30657
rect 16822 30648 16834 30651
rect 16724 30620 16834 30648
rect 16724 30608 16730 30620
rect 16822 30617 16834 30620
rect 16868 30617 16880 30651
rect 16822 30611 16880 30617
rect 18138 30608 18144 30660
rect 18196 30648 18202 30660
rect 19245 30651 19303 30657
rect 19245 30648 19257 30651
rect 18196 30620 19257 30648
rect 18196 30608 18202 30620
rect 19245 30617 19257 30620
rect 19291 30617 19303 30651
rect 19426 30648 19432 30660
rect 19387 30620 19432 30648
rect 19245 30611 19303 30617
rect 19426 30608 19432 30620
rect 19484 30608 19490 30660
rect 17126 30540 17132 30592
rect 17184 30580 17190 30592
rect 19613 30583 19671 30589
rect 19613 30580 19625 30583
rect 17184 30552 19625 30580
rect 17184 30540 17190 30552
rect 19613 30549 19625 30552
rect 19659 30549 19671 30583
rect 19613 30543 19671 30549
rect 20438 30540 20444 30592
rect 20496 30580 20502 30592
rect 20533 30583 20591 30589
rect 20533 30580 20545 30583
rect 20496 30552 20545 30580
rect 20496 30540 20502 30552
rect 20533 30549 20545 30552
rect 20579 30549 20591 30583
rect 20824 30580 20852 30679
rect 21082 30676 21088 30728
rect 21140 30716 21146 30728
rect 21177 30719 21235 30725
rect 21177 30716 21189 30719
rect 21140 30688 21189 30716
rect 21140 30676 21146 30688
rect 21177 30685 21189 30688
rect 21223 30685 21235 30719
rect 21376 30716 21404 30756
rect 21450 30744 21456 30796
rect 21508 30784 21514 30796
rect 22738 30784 22744 30796
rect 21508 30756 21956 30784
rect 21508 30744 21514 30756
rect 21726 30716 21732 30728
rect 21376 30688 21732 30716
rect 21177 30679 21235 30685
rect 21726 30676 21732 30688
rect 21784 30676 21790 30728
rect 21928 30660 21956 30756
rect 22020 30756 22744 30784
rect 22020 30725 22048 30756
rect 22738 30744 22744 30756
rect 22796 30744 22802 30796
rect 22940 30725 22968 30824
rect 28902 30812 28908 30864
rect 28960 30852 28966 30864
rect 29086 30852 29092 30864
rect 28960 30824 29092 30852
rect 28960 30812 28966 30824
rect 29086 30812 29092 30824
rect 29144 30812 29150 30864
rect 24302 30744 24308 30796
rect 24360 30784 24366 30796
rect 24397 30787 24455 30793
rect 24397 30784 24409 30787
rect 24360 30756 24409 30784
rect 24360 30744 24366 30756
rect 24397 30753 24409 30756
rect 24443 30753 24455 30787
rect 24397 30747 24455 30753
rect 27617 30787 27675 30793
rect 27617 30753 27629 30787
rect 27663 30784 27675 30787
rect 27663 30756 27752 30784
rect 27663 30753 27675 30756
rect 27617 30747 27675 30753
rect 22005 30719 22063 30725
rect 22005 30685 22017 30719
rect 22051 30685 22063 30719
rect 22925 30719 22983 30725
rect 22005 30679 22063 30685
rect 22204 30688 22600 30716
rect 21910 30648 21916 30660
rect 21823 30620 21916 30648
rect 21910 30608 21916 30620
rect 21968 30648 21974 30660
rect 22204 30657 22232 30688
rect 22189 30651 22247 30657
rect 22189 30648 22201 30651
rect 21968 30620 22201 30648
rect 21968 30608 21974 30620
rect 22189 30617 22201 30620
rect 22235 30617 22247 30651
rect 22189 30611 22247 30617
rect 22373 30651 22431 30657
rect 22373 30617 22385 30651
rect 22419 30617 22431 30651
rect 22572 30648 22600 30688
rect 22925 30685 22937 30719
rect 22971 30685 22983 30719
rect 22925 30679 22983 30685
rect 24486 30676 24492 30728
rect 24544 30716 24550 30728
rect 24653 30719 24711 30725
rect 24653 30716 24665 30719
rect 24544 30688 24665 30716
rect 24544 30676 24550 30688
rect 24653 30685 24665 30688
rect 24699 30685 24711 30719
rect 24653 30679 24711 30685
rect 27154 30676 27160 30728
rect 27212 30716 27218 30728
rect 27724 30716 27752 30756
rect 29546 30716 29552 30728
rect 27212 30688 27660 30716
rect 27724 30688 29552 30716
rect 27212 30676 27218 30688
rect 23109 30651 23167 30657
rect 23109 30648 23121 30651
rect 22572 30620 23121 30648
rect 22373 30611 22431 30617
rect 23109 30617 23121 30620
rect 23155 30617 23167 30651
rect 23109 30611 23167 30617
rect 22278 30580 22284 30592
rect 20824 30552 22284 30580
rect 20533 30543 20591 30549
rect 22278 30540 22284 30552
rect 22336 30540 22342 30592
rect 22385 30580 22413 30611
rect 23290 30608 23296 30660
rect 23348 30648 23354 30660
rect 24762 30648 24768 30660
rect 23348 30620 24768 30648
rect 23348 30608 23354 30620
rect 24762 30608 24768 30620
rect 24820 30648 24826 30660
rect 27632 30648 27660 30688
rect 29546 30676 29552 30688
rect 29604 30716 29610 30728
rect 29914 30716 29920 30728
rect 29604 30688 29920 30716
rect 29604 30676 29610 30688
rect 29914 30676 29920 30688
rect 29972 30676 29978 30728
rect 30006 30676 30012 30728
rect 30064 30716 30070 30728
rect 30173 30719 30231 30725
rect 30173 30716 30185 30719
rect 30064 30688 30185 30716
rect 30064 30676 30070 30688
rect 30173 30685 30185 30688
rect 30219 30685 30231 30719
rect 30173 30679 30231 30685
rect 35621 30719 35679 30725
rect 35621 30685 35633 30719
rect 35667 30716 35679 30719
rect 36538 30716 36544 30728
rect 35667 30688 36544 30716
rect 35667 30685 35679 30688
rect 35621 30679 35679 30685
rect 36538 30676 36544 30688
rect 36596 30676 36602 30728
rect 36630 30676 36636 30728
rect 36688 30716 36694 30728
rect 37921 30719 37979 30725
rect 37921 30716 37933 30719
rect 36688 30688 37933 30716
rect 36688 30676 36694 30688
rect 37921 30685 37933 30688
rect 37967 30716 37979 30719
rect 45462 30716 45468 30728
rect 37967 30688 45468 30716
rect 37967 30685 37979 30688
rect 37921 30679 37979 30685
rect 45462 30676 45468 30688
rect 45520 30676 45526 30728
rect 27884 30651 27942 30657
rect 24820 30620 25820 30648
rect 27632 30620 27752 30648
rect 24820 30608 24826 30620
rect 22462 30580 22468 30592
rect 22385 30552 22468 30580
rect 22462 30540 22468 30552
rect 22520 30540 22526 30592
rect 22646 30540 22652 30592
rect 22704 30580 22710 30592
rect 23382 30580 23388 30592
rect 22704 30552 23388 30580
rect 22704 30540 22710 30552
rect 23382 30540 23388 30552
rect 23440 30540 23446 30592
rect 25792 30589 25820 30620
rect 25777 30583 25835 30589
rect 25777 30549 25789 30583
rect 25823 30549 25835 30583
rect 27724 30580 27752 30620
rect 27884 30617 27896 30651
rect 27930 30648 27942 30651
rect 28626 30648 28632 30660
rect 27930 30620 28632 30648
rect 27930 30617 27942 30620
rect 27884 30611 27942 30617
rect 28626 30608 28632 30620
rect 28684 30608 28690 30660
rect 35986 30648 35992 30660
rect 35947 30620 35992 30648
rect 35986 30608 35992 30620
rect 36044 30608 36050 30660
rect 36906 30648 36912 30660
rect 36867 30620 36912 30648
rect 36906 30608 36912 30620
rect 36964 30648 36970 30660
rect 46382 30648 46388 30660
rect 36964 30620 46388 30648
rect 36964 30608 36970 30620
rect 46382 30608 46388 30620
rect 46440 30608 46446 30660
rect 36630 30580 36636 30592
rect 27724 30552 36636 30580
rect 25777 30543 25835 30549
rect 36630 30540 36636 30552
rect 36688 30540 36694 30592
rect 1104 30490 48852 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 48852 30490
rect 1104 30416 48852 30438
rect 3418 30336 3424 30388
rect 3476 30376 3482 30388
rect 36906 30376 36912 30388
rect 3476 30348 36912 30376
rect 3476 30336 3482 30348
rect 36906 30336 36912 30348
rect 36964 30336 36970 30388
rect 16666 30308 16672 30320
rect 16627 30280 16672 30308
rect 16666 30268 16672 30280
rect 16724 30268 16730 30320
rect 18601 30311 18659 30317
rect 18601 30277 18613 30311
rect 18647 30308 18659 30311
rect 20530 30308 20536 30320
rect 18647 30280 20536 30308
rect 18647 30277 18659 30280
rect 18601 30271 18659 30277
rect 20530 30268 20536 30280
rect 20588 30268 20594 30320
rect 20806 30308 20812 30320
rect 20732 30280 20812 30308
rect 2133 30243 2191 30249
rect 2133 30209 2145 30243
rect 2179 30240 2191 30243
rect 2406 30240 2412 30252
rect 2179 30212 2412 30240
rect 2179 30209 2191 30212
rect 2133 30203 2191 30209
rect 2406 30200 2412 30212
rect 2464 30200 2470 30252
rect 14826 30200 14832 30252
rect 14884 30240 14890 30252
rect 16945 30243 17003 30249
rect 16945 30240 16957 30243
rect 14884 30212 16957 30240
rect 14884 30200 14890 30212
rect 16945 30209 16957 30212
rect 16991 30209 17003 30243
rect 16945 30203 17003 30209
rect 17034 30243 17092 30249
rect 17034 30209 17046 30243
rect 17080 30209 17092 30243
rect 17034 30203 17092 30209
rect 1854 30132 1860 30184
rect 1912 30172 1918 30184
rect 2222 30172 2228 30184
rect 1912 30144 2228 30172
rect 1912 30132 1918 30144
rect 2222 30132 2228 30144
rect 2280 30132 2286 30184
rect 17049 30116 17077 30203
rect 17126 30200 17132 30252
rect 17184 30249 17190 30252
rect 17184 30240 17192 30249
rect 17313 30243 17371 30249
rect 17184 30212 17229 30240
rect 17184 30203 17192 30212
rect 17313 30209 17325 30243
rect 17359 30240 17371 30243
rect 17494 30240 17500 30252
rect 17359 30212 17500 30240
rect 17359 30209 17371 30212
rect 17313 30203 17371 30209
rect 17184 30200 17190 30203
rect 17494 30200 17500 30212
rect 17552 30200 17558 30252
rect 18414 30200 18420 30252
rect 18472 30240 18478 30252
rect 18509 30243 18567 30249
rect 18509 30240 18521 30243
rect 18472 30212 18521 30240
rect 18472 30200 18478 30212
rect 18509 30209 18521 30212
rect 18555 30209 18567 30243
rect 19702 30240 19708 30252
rect 19663 30212 19708 30240
rect 18509 30203 18567 30209
rect 19702 30200 19708 30212
rect 19760 30200 19766 30252
rect 19797 30243 19855 30249
rect 19797 30209 19809 30243
rect 19843 30240 19855 30243
rect 20732 30240 20760 30280
rect 20806 30268 20812 30280
rect 20864 30268 20870 30320
rect 20993 30311 21051 30317
rect 20993 30277 21005 30311
rect 21039 30308 21051 30311
rect 21174 30308 21180 30320
rect 21039 30280 21180 30308
rect 21039 30277 21051 30280
rect 20993 30271 21051 30277
rect 21174 30268 21180 30280
rect 21232 30268 21238 30320
rect 22278 30268 22284 30320
rect 22336 30308 22342 30320
rect 48133 30311 48191 30317
rect 48133 30308 48145 30311
rect 22336 30280 48145 30308
rect 22336 30268 22342 30280
rect 48133 30277 48145 30280
rect 48179 30277 48191 30311
rect 48133 30271 48191 30277
rect 20898 30240 20904 30252
rect 19843 30212 20760 30240
rect 20859 30212 20904 30240
rect 19843 30209 19855 30212
rect 19797 30203 19855 30209
rect 20898 30200 20904 30212
rect 20956 30200 20962 30252
rect 21821 30243 21879 30249
rect 21821 30240 21833 30243
rect 21100 30212 21833 30240
rect 18785 30175 18843 30181
rect 18785 30141 18797 30175
rect 18831 30141 18843 30175
rect 18785 30135 18843 30141
rect 19981 30175 20039 30181
rect 19981 30141 19993 30175
rect 20027 30172 20039 30175
rect 20027 30144 20208 30172
rect 20027 30141 20039 30144
rect 19981 30135 20039 30141
rect 17034 30104 17040 30116
rect 16947 30076 17040 30104
rect 17034 30064 17040 30076
rect 17092 30104 17098 30116
rect 17586 30104 17592 30116
rect 17092 30076 17592 30104
rect 17092 30064 17098 30076
rect 17586 30064 17592 30076
rect 17644 30064 17650 30116
rect 18138 30104 18144 30116
rect 18099 30076 18144 30104
rect 18138 30064 18144 30076
rect 18196 30064 18202 30116
rect 18800 30104 18828 30135
rect 19150 30104 19156 30116
rect 18800 30076 19156 30104
rect 19150 30064 19156 30076
rect 19208 30104 19214 30116
rect 20180 30104 20208 30144
rect 19208 30076 20208 30104
rect 19208 30064 19214 30076
rect 1394 29996 1400 30048
rect 1452 30036 1458 30048
rect 1673 30039 1731 30045
rect 1673 30036 1685 30039
rect 1452 30008 1685 30036
rect 1452 29996 1458 30008
rect 1673 30005 1685 30008
rect 1719 30005 1731 30039
rect 2222 30036 2228 30048
rect 2183 30008 2228 30036
rect 1673 29999 1731 30005
rect 2222 29996 2228 30008
rect 2280 29996 2286 30048
rect 17770 29996 17776 30048
rect 17828 30036 17834 30048
rect 19337 30039 19395 30045
rect 19337 30036 19349 30039
rect 17828 30008 19349 30036
rect 17828 29996 17834 30008
rect 19337 30005 19349 30008
rect 19383 30005 19395 30039
rect 20180 30036 20208 30076
rect 20533 30107 20591 30113
rect 20533 30073 20545 30107
rect 20579 30104 20591 30107
rect 21100 30104 21128 30212
rect 21821 30209 21833 30212
rect 21867 30209 21879 30243
rect 21821 30203 21879 30209
rect 21910 30200 21916 30252
rect 21968 30240 21974 30252
rect 22005 30243 22063 30249
rect 22005 30240 22017 30243
rect 21968 30212 22017 30240
rect 21968 30200 21974 30212
rect 22005 30209 22017 30212
rect 22051 30209 22063 30243
rect 22005 30203 22063 30209
rect 23201 30243 23259 30249
rect 23201 30209 23213 30243
rect 23247 30240 23259 30243
rect 23934 30240 23940 30252
rect 23247 30212 23940 30240
rect 23247 30209 23259 30212
rect 23201 30203 23259 30209
rect 23934 30200 23940 30212
rect 23992 30200 23998 30252
rect 24578 30200 24584 30252
rect 24636 30240 24642 30252
rect 24673 30243 24731 30249
rect 24673 30240 24685 30243
rect 24636 30212 24685 30240
rect 24636 30200 24642 30212
rect 24673 30209 24685 30212
rect 24719 30209 24731 30243
rect 24854 30240 24860 30252
rect 24815 30212 24860 30240
rect 24673 30203 24731 30209
rect 24854 30200 24860 30212
rect 24912 30200 24918 30252
rect 25590 30240 25596 30252
rect 25551 30212 25596 30240
rect 25590 30200 25596 30212
rect 25648 30200 25654 30252
rect 26418 30200 26424 30252
rect 26476 30240 26482 30252
rect 27430 30240 27436 30252
rect 26476 30212 27436 30240
rect 26476 30200 26482 30212
rect 27430 30200 27436 30212
rect 27488 30200 27494 30252
rect 28902 30240 28908 30252
rect 28863 30212 28908 30240
rect 28902 30200 28908 30212
rect 28960 30200 28966 30252
rect 29089 30243 29147 30249
rect 29089 30209 29101 30243
rect 29135 30240 29147 30243
rect 29178 30240 29184 30252
rect 29135 30212 29184 30240
rect 29135 30209 29147 30212
rect 29089 30203 29147 30209
rect 29178 30200 29184 30212
rect 29236 30200 29242 30252
rect 29914 30240 29920 30252
rect 29875 30212 29920 30240
rect 29914 30200 29920 30212
rect 29972 30200 29978 30252
rect 30006 30200 30012 30252
rect 30064 30240 30070 30252
rect 30173 30243 30231 30249
rect 30173 30240 30185 30243
rect 30064 30212 30185 30240
rect 30064 30200 30070 30212
rect 30173 30209 30185 30212
rect 30219 30209 30231 30243
rect 30173 30203 30231 30209
rect 36538 30200 36544 30252
rect 36596 30240 36602 30252
rect 37277 30243 37335 30249
rect 37277 30240 37289 30243
rect 36596 30212 37289 30240
rect 36596 30200 36602 30212
rect 37277 30209 37289 30212
rect 37323 30209 37335 30243
rect 47946 30240 47952 30252
rect 47907 30212 47952 30240
rect 37277 30203 37335 30209
rect 47946 30200 47952 30212
rect 48004 30200 48010 30252
rect 21177 30175 21235 30181
rect 21177 30141 21189 30175
rect 21223 30141 21235 30175
rect 21177 30135 21235 30141
rect 20579 30076 21128 30104
rect 20579 30073 20591 30076
rect 20533 30067 20591 30073
rect 21192 30036 21220 30135
rect 21726 30132 21732 30184
rect 21784 30172 21790 30184
rect 22189 30175 22247 30181
rect 22189 30172 22201 30175
rect 21784 30144 22201 30172
rect 21784 30132 21790 30144
rect 22189 30141 22201 30144
rect 22235 30141 22247 30175
rect 23290 30172 23296 30184
rect 23251 30144 23296 30172
rect 22189 30135 22247 30141
rect 23290 30132 23296 30144
rect 23348 30132 23354 30184
rect 23382 30132 23388 30184
rect 23440 30172 23446 30184
rect 28626 30172 28632 30184
rect 23440 30144 23485 30172
rect 28587 30144 28632 30172
rect 23440 30132 23446 30144
rect 28626 30132 28632 30144
rect 28684 30132 28690 30184
rect 28813 30175 28871 30181
rect 28813 30141 28825 30175
rect 28859 30141 28871 30175
rect 28813 30135 28871 30141
rect 28997 30175 29055 30181
rect 28997 30141 29009 30175
rect 29043 30172 29055 30175
rect 29362 30172 29368 30184
rect 29043 30144 29368 30172
rect 29043 30141 29055 30144
rect 28997 30135 29055 30141
rect 21542 30064 21548 30116
rect 21600 30104 21606 30116
rect 22002 30104 22008 30116
rect 21600 30076 22008 30104
rect 21600 30064 21606 30076
rect 22002 30064 22008 30076
rect 22060 30104 22066 30116
rect 25777 30107 25835 30113
rect 25777 30104 25789 30107
rect 22060 30076 25789 30104
rect 22060 30064 22066 30076
rect 25777 30073 25789 30076
rect 25823 30073 25835 30107
rect 28828 30104 28856 30135
rect 29362 30132 29368 30144
rect 29420 30132 29426 30184
rect 28828 30076 29040 30104
rect 25777 30067 25835 30073
rect 29012 30048 29040 30076
rect 31202 30064 31208 30116
rect 31260 30104 31266 30116
rect 31297 30107 31355 30113
rect 31297 30104 31309 30107
rect 31260 30076 31309 30104
rect 31260 30064 31266 30076
rect 31297 30073 31309 30076
rect 31343 30073 31355 30107
rect 31297 30067 31355 30073
rect 22646 30036 22652 30048
rect 20180 30008 22652 30036
rect 19337 29999 19395 30005
rect 22646 29996 22652 30008
rect 22704 29996 22710 30048
rect 22738 29996 22744 30048
rect 22796 30036 22802 30048
rect 22833 30039 22891 30045
rect 22833 30036 22845 30039
rect 22796 30008 22845 30036
rect 22796 29996 22802 30008
rect 22833 30005 22845 30008
rect 22879 30005 22891 30039
rect 22833 29999 22891 30005
rect 24946 29996 24952 30048
rect 25004 30036 25010 30048
rect 25041 30039 25099 30045
rect 25041 30036 25053 30039
rect 25004 30008 25053 30036
rect 25004 29996 25010 30008
rect 25041 30005 25053 30008
rect 25087 30005 25099 30039
rect 25041 29999 25099 30005
rect 27338 29996 27344 30048
rect 27396 30036 27402 30048
rect 27525 30039 27583 30045
rect 27525 30036 27537 30039
rect 27396 30008 27537 30036
rect 27396 29996 27402 30008
rect 27525 30005 27537 30008
rect 27571 30036 27583 30039
rect 27982 30036 27988 30048
rect 27571 30008 27988 30036
rect 27571 30005 27583 30008
rect 27525 29999 27583 30005
rect 27982 29996 27988 30008
rect 28040 29996 28046 30048
rect 28994 29996 29000 30048
rect 29052 29996 29058 30048
rect 37458 30036 37464 30048
rect 37419 30008 37464 30036
rect 37458 29996 37464 30008
rect 37516 29996 37522 30048
rect 1104 29946 48852 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 48852 29946
rect 1104 29872 48852 29894
rect 18141 29835 18199 29841
rect 18141 29801 18153 29835
rect 18187 29832 18199 29835
rect 19426 29832 19432 29844
rect 18187 29804 19432 29832
rect 18187 29801 18199 29804
rect 18141 29795 18199 29801
rect 19426 29792 19432 29804
rect 19484 29832 19490 29844
rect 19702 29832 19708 29844
rect 19484 29804 19708 29832
rect 19484 29792 19490 29804
rect 19702 29792 19708 29804
rect 19760 29792 19766 29844
rect 24854 29792 24860 29844
rect 24912 29832 24918 29844
rect 24912 29804 26372 29832
rect 24912 29792 24918 29804
rect 23569 29767 23627 29773
rect 23569 29733 23581 29767
rect 23615 29764 23627 29767
rect 23934 29764 23940 29776
rect 23615 29736 23940 29764
rect 23615 29733 23627 29736
rect 23569 29727 23627 29733
rect 23934 29724 23940 29736
rect 23992 29724 23998 29776
rect 26344 29773 26372 29804
rect 27430 29792 27436 29844
rect 27488 29832 27494 29844
rect 27525 29835 27583 29841
rect 27525 29832 27537 29835
rect 27488 29804 27537 29832
rect 27488 29792 27494 29804
rect 27525 29801 27537 29804
rect 27571 29801 27583 29835
rect 27525 29795 27583 29801
rect 29825 29835 29883 29841
rect 29825 29801 29837 29835
rect 29871 29832 29883 29835
rect 30006 29832 30012 29844
rect 29871 29804 30012 29832
rect 29871 29801 29883 29804
rect 29825 29795 29883 29801
rect 30006 29792 30012 29804
rect 30064 29792 30070 29844
rect 31021 29835 31079 29841
rect 31021 29801 31033 29835
rect 31067 29832 31079 29835
rect 31570 29832 31576 29844
rect 31067 29804 31576 29832
rect 31067 29801 31079 29804
rect 31021 29795 31079 29801
rect 31570 29792 31576 29804
rect 31628 29832 31634 29844
rect 32950 29832 32956 29844
rect 31628 29804 32168 29832
rect 31628 29792 31634 29804
rect 26329 29767 26387 29773
rect 26329 29733 26341 29767
rect 26375 29764 26387 29767
rect 26375 29736 31892 29764
rect 26375 29733 26387 29736
rect 26329 29727 26387 29733
rect 1394 29696 1400 29708
rect 1355 29668 1400 29696
rect 1394 29656 1400 29668
rect 1452 29656 1458 29708
rect 1581 29699 1639 29705
rect 1581 29665 1593 29699
rect 1627 29696 1639 29699
rect 2222 29696 2228 29708
rect 1627 29668 2228 29696
rect 1627 29665 1639 29668
rect 1581 29659 1639 29665
rect 2222 29656 2228 29668
rect 2280 29656 2286 29708
rect 2774 29696 2780 29708
rect 2735 29668 2780 29696
rect 2774 29656 2780 29668
rect 2832 29656 2838 29708
rect 21818 29656 21824 29708
rect 21876 29696 21882 29708
rect 22189 29699 22247 29705
rect 22189 29696 22201 29699
rect 21876 29668 22201 29696
rect 21876 29656 21882 29668
rect 22189 29665 22201 29668
rect 22235 29665 22247 29699
rect 22189 29659 22247 29665
rect 28994 29656 29000 29708
rect 29052 29696 29058 29708
rect 29822 29696 29828 29708
rect 29052 29668 29828 29696
rect 29052 29656 29058 29668
rect 29822 29656 29828 29668
rect 29880 29696 29886 29708
rect 30006 29696 30012 29708
rect 29880 29668 30012 29696
rect 29880 29656 29886 29668
rect 30006 29656 30012 29668
rect 30064 29656 30070 29708
rect 30101 29699 30159 29705
rect 30101 29665 30113 29699
rect 30147 29696 30159 29699
rect 31202 29696 31208 29708
rect 30147 29668 31208 29696
rect 30147 29665 30159 29668
rect 30101 29659 30159 29665
rect 31202 29656 31208 29668
rect 31260 29656 31266 29708
rect 16761 29631 16819 29637
rect 16761 29597 16773 29631
rect 16807 29628 16819 29631
rect 16850 29628 16856 29640
rect 16807 29600 16856 29628
rect 16807 29597 16819 29600
rect 16761 29591 16819 29597
rect 16850 29588 16856 29600
rect 16908 29628 16914 29640
rect 20438 29637 20444 29640
rect 20165 29631 20223 29637
rect 20165 29628 20177 29631
rect 16908 29600 20177 29628
rect 16908 29588 16914 29600
rect 20165 29597 20177 29600
rect 20211 29597 20223 29631
rect 20432 29628 20444 29637
rect 20399 29600 20444 29628
rect 20165 29591 20223 29597
rect 20432 29591 20444 29600
rect 20438 29588 20444 29591
rect 20496 29588 20502 29640
rect 24949 29631 25007 29637
rect 24949 29597 24961 29631
rect 24995 29628 25007 29631
rect 25038 29628 25044 29640
rect 24995 29600 25044 29628
rect 24995 29597 25007 29600
rect 24949 29591 25007 29597
rect 25038 29588 25044 29600
rect 25096 29588 25102 29640
rect 29362 29588 29368 29640
rect 29420 29628 29426 29640
rect 30190 29628 30196 29640
rect 29420 29600 30196 29628
rect 29420 29588 29426 29600
rect 30190 29588 30196 29600
rect 30248 29588 30254 29640
rect 30282 29588 30288 29640
rect 30340 29628 30346 29640
rect 30340 29600 30385 29628
rect 30340 29588 30346 29600
rect 16666 29520 16672 29572
rect 16724 29560 16730 29572
rect 17006 29563 17064 29569
rect 17006 29560 17018 29563
rect 16724 29532 17018 29560
rect 16724 29520 16730 29532
rect 17006 29529 17018 29532
rect 17052 29529 17064 29563
rect 17006 29523 17064 29529
rect 22278 29520 22284 29572
rect 22336 29560 22342 29572
rect 22434 29563 22492 29569
rect 22434 29560 22446 29563
rect 22336 29532 22446 29560
rect 22336 29520 22342 29532
rect 22434 29529 22446 29532
rect 22480 29529 22492 29563
rect 22434 29523 22492 29529
rect 24302 29520 24308 29572
rect 24360 29560 24366 29572
rect 25194 29563 25252 29569
rect 25194 29560 25206 29563
rect 24360 29532 25206 29560
rect 24360 29520 24366 29532
rect 25194 29529 25206 29532
rect 25240 29529 25252 29563
rect 25194 29523 25252 29529
rect 27433 29563 27491 29569
rect 27433 29529 27445 29563
rect 27479 29560 27491 29563
rect 27982 29560 27988 29572
rect 27479 29532 27988 29560
rect 27479 29529 27491 29532
rect 27433 29523 27491 29529
rect 27982 29520 27988 29532
rect 28040 29560 28046 29572
rect 28353 29563 28411 29569
rect 28353 29560 28365 29563
rect 28040 29532 28365 29560
rect 28040 29520 28046 29532
rect 28353 29529 28365 29532
rect 28399 29529 28411 29563
rect 28353 29523 28411 29529
rect 30006 29520 30012 29572
rect 30064 29560 30070 29572
rect 30929 29563 30987 29569
rect 30929 29560 30941 29563
rect 30064 29532 30941 29560
rect 30064 29520 30070 29532
rect 30929 29529 30941 29532
rect 30975 29529 30987 29563
rect 31754 29560 31760 29572
rect 30929 29523 30987 29529
rect 31726 29520 31760 29560
rect 31812 29520 31818 29572
rect 20898 29452 20904 29504
rect 20956 29492 20962 29504
rect 21545 29495 21603 29501
rect 21545 29492 21557 29495
rect 20956 29464 21557 29492
rect 20956 29452 20962 29464
rect 21545 29461 21557 29464
rect 21591 29492 21603 29495
rect 21726 29492 21732 29504
rect 21591 29464 21732 29492
rect 21591 29461 21603 29464
rect 21545 29455 21603 29461
rect 21726 29452 21732 29464
rect 21784 29452 21790 29504
rect 28445 29495 28503 29501
rect 28445 29461 28457 29495
rect 28491 29492 28503 29495
rect 28718 29492 28724 29504
rect 28491 29464 28724 29492
rect 28491 29461 28503 29464
rect 28445 29455 28503 29461
rect 28718 29452 28724 29464
rect 28776 29492 28782 29504
rect 31726 29492 31754 29520
rect 28776 29464 31754 29492
rect 31864 29492 31892 29736
rect 32140 29637 32168 29804
rect 32324 29804 32956 29832
rect 32324 29637 32352 29804
rect 32950 29792 32956 29804
rect 33008 29832 33014 29844
rect 34790 29832 34796 29844
rect 33008 29804 33732 29832
rect 34751 29804 34796 29832
rect 33008 29792 33014 29804
rect 33704 29764 33732 29804
rect 34790 29792 34796 29804
rect 34848 29792 34854 29844
rect 38654 29832 38660 29844
rect 38615 29804 38660 29832
rect 38654 29792 38660 29804
rect 38712 29792 38718 29844
rect 35069 29767 35127 29773
rect 35069 29764 35081 29767
rect 33704 29736 35081 29764
rect 35069 29733 35081 29736
rect 35115 29733 35127 29767
rect 35069 29727 35127 29733
rect 33778 29656 33784 29708
rect 33836 29696 33842 29708
rect 37277 29699 37335 29705
rect 37277 29696 37289 29699
rect 33836 29668 37289 29696
rect 33836 29656 33842 29668
rect 37277 29665 37289 29668
rect 37323 29665 37335 29699
rect 37277 29659 37335 29665
rect 32125 29631 32183 29637
rect 32125 29597 32137 29631
rect 32171 29597 32183 29631
rect 32125 29591 32183 29597
rect 32309 29631 32367 29637
rect 32309 29597 32321 29631
rect 32355 29597 32367 29631
rect 32309 29591 32367 29597
rect 32769 29631 32827 29637
rect 32769 29597 32781 29631
rect 32815 29628 32827 29631
rect 33796 29628 33824 29656
rect 34698 29628 34704 29640
rect 32815 29600 33824 29628
rect 34659 29600 34704 29628
rect 32815 29597 32827 29600
rect 32769 29591 32827 29597
rect 34698 29588 34704 29600
rect 34756 29588 34762 29640
rect 34882 29628 34888 29640
rect 34843 29600 34888 29628
rect 34882 29588 34888 29600
rect 34940 29588 34946 29640
rect 46290 29588 46296 29640
rect 46348 29628 46354 29640
rect 47673 29631 47731 29637
rect 47673 29628 47685 29631
rect 46348 29600 47685 29628
rect 46348 29588 46354 29600
rect 47673 29597 47685 29600
rect 47719 29597 47731 29631
rect 47673 29591 47731 29597
rect 32217 29563 32275 29569
rect 32217 29529 32229 29563
rect 32263 29560 32275 29563
rect 33014 29563 33072 29569
rect 33014 29560 33026 29563
rect 32263 29532 33026 29560
rect 32263 29529 32275 29532
rect 32217 29523 32275 29529
rect 33014 29529 33026 29532
rect 33060 29529 33072 29563
rect 37274 29560 37280 29572
rect 33014 29523 33072 29529
rect 33152 29532 37280 29560
rect 33152 29492 33180 29532
rect 37274 29520 37280 29532
rect 37332 29520 37338 29572
rect 37550 29569 37556 29572
rect 37544 29523 37556 29569
rect 37608 29560 37614 29572
rect 37608 29532 37644 29560
rect 37550 29520 37556 29523
rect 37608 29520 37614 29532
rect 31864 29464 33180 29492
rect 28776 29452 28782 29464
rect 33870 29452 33876 29504
rect 33928 29492 33934 29504
rect 34149 29495 34207 29501
rect 34149 29492 34161 29495
rect 33928 29464 34161 29492
rect 33928 29452 33934 29464
rect 34149 29461 34161 29464
rect 34195 29461 34207 29495
rect 34149 29455 34207 29461
rect 1104 29402 48852 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 48852 29402
rect 1104 29328 48852 29350
rect 16666 29288 16672 29300
rect 16627 29260 16672 29288
rect 16666 29248 16672 29260
rect 16724 29248 16730 29300
rect 22005 29291 22063 29297
rect 22005 29257 22017 29291
rect 22051 29288 22063 29291
rect 22278 29288 22284 29300
rect 22051 29260 22284 29288
rect 22051 29257 22063 29260
rect 22005 29251 22063 29257
rect 22278 29248 22284 29260
rect 22336 29248 22342 29300
rect 24302 29288 24308 29300
rect 24263 29260 24308 29288
rect 24302 29248 24308 29260
rect 24360 29248 24366 29300
rect 28721 29291 28779 29297
rect 28721 29257 28733 29291
rect 28767 29288 28779 29291
rect 28994 29288 29000 29300
rect 28767 29260 29000 29288
rect 28767 29257 28779 29260
rect 28721 29251 28779 29257
rect 28994 29248 29000 29260
rect 29052 29248 29058 29300
rect 29178 29248 29184 29300
rect 29236 29288 29242 29300
rect 29236 29260 29776 29288
rect 29236 29248 29242 29260
rect 18141 29223 18199 29229
rect 18141 29220 18153 29223
rect 17144 29192 18153 29220
rect 17031 29164 17037 29167
rect 8846 29112 8852 29164
rect 8904 29152 8910 29164
rect 16899 29155 16957 29161
rect 16899 29152 16911 29155
rect 8904 29124 16911 29152
rect 8904 29112 8910 29124
rect 16899 29121 16911 29124
rect 16945 29121 16957 29155
rect 16899 29115 16957 29121
rect 17018 29158 17037 29164
rect 17018 29124 17030 29158
rect 17018 29118 17037 29124
rect 17031 29115 17037 29118
rect 17089 29115 17095 29167
rect 17144 29164 17172 29192
rect 18141 29189 18153 29192
rect 18187 29189 18199 29223
rect 18141 29183 18199 29189
rect 22186 29180 22192 29232
rect 22244 29220 22250 29232
rect 22244 29192 22416 29220
rect 22244 29180 22250 29192
rect 17129 29158 17187 29164
rect 17129 29124 17141 29158
rect 17175 29124 17187 29158
rect 17129 29118 17187 29124
rect 17313 29155 17371 29161
rect 17313 29121 17325 29155
rect 17359 29152 17371 29155
rect 17494 29152 17500 29164
rect 17359 29124 17500 29152
rect 17359 29121 17371 29124
rect 17313 29115 17371 29121
rect 17494 29112 17500 29124
rect 17552 29112 17558 29164
rect 17770 29152 17776 29164
rect 17731 29124 17776 29152
rect 17770 29112 17776 29124
rect 17828 29112 17834 29164
rect 17957 29155 18015 29161
rect 17957 29121 17969 29155
rect 18003 29152 18015 29155
rect 19334 29152 19340 29164
rect 18003 29124 19340 29152
rect 18003 29121 18015 29124
rect 17957 29115 18015 29121
rect 19334 29112 19340 29124
rect 19392 29112 19398 29164
rect 22388 29161 22416 29192
rect 22554 29180 22560 29232
rect 22612 29220 22618 29232
rect 29748 29229 29776 29260
rect 29822 29248 29828 29300
rect 29880 29288 29886 29300
rect 29933 29291 29991 29297
rect 29933 29288 29945 29291
rect 29880 29260 29945 29288
rect 29880 29248 29886 29260
rect 29933 29257 29945 29260
rect 29979 29257 29991 29291
rect 29933 29251 29991 29257
rect 30101 29291 30159 29297
rect 30101 29257 30113 29291
rect 30147 29288 30159 29291
rect 30282 29288 30288 29300
rect 30147 29260 30288 29288
rect 30147 29257 30159 29260
rect 30101 29251 30159 29257
rect 30282 29248 30288 29260
rect 30340 29248 30346 29300
rect 31386 29248 31392 29300
rect 31444 29288 31450 29300
rect 32582 29288 32588 29300
rect 31444 29260 32588 29288
rect 31444 29248 31450 29260
rect 32582 29248 32588 29260
rect 32640 29288 32646 29300
rect 32677 29291 32735 29297
rect 32677 29288 32689 29291
rect 32640 29260 32689 29288
rect 32640 29248 32646 29260
rect 32677 29257 32689 29260
rect 32723 29257 32735 29291
rect 32677 29251 32735 29257
rect 46934 29248 46940 29300
rect 46992 29288 46998 29300
rect 47394 29288 47400 29300
rect 46992 29260 47400 29288
rect 46992 29248 46998 29260
rect 47394 29248 47400 29260
rect 47452 29248 47458 29300
rect 27433 29223 27491 29229
rect 22612 29192 22692 29220
rect 22612 29180 22618 29192
rect 22281 29155 22339 29161
rect 22281 29121 22293 29155
rect 22327 29121 22339 29155
rect 22281 29115 22339 29121
rect 22373 29155 22431 29161
rect 22373 29121 22385 29155
rect 22419 29121 22431 29155
rect 22373 29115 22431 29121
rect 3418 28976 3424 29028
rect 3476 29016 3482 29028
rect 15470 29016 15476 29028
rect 3476 28988 15476 29016
rect 3476 28976 3482 28988
rect 15470 28976 15476 28988
rect 15528 28976 15534 29028
rect 22296 29016 22324 29115
rect 22462 29112 22468 29164
rect 22520 29152 22526 29164
rect 22664 29161 22692 29192
rect 27433 29189 27445 29223
rect 27479 29220 27491 29223
rect 29733 29223 29791 29229
rect 27479 29192 29684 29220
rect 27479 29189 27491 29192
rect 27433 29183 27491 29189
rect 22649 29155 22707 29161
rect 22520 29124 22565 29152
rect 22520 29112 22526 29124
rect 22649 29121 22661 29155
rect 22695 29121 22707 29155
rect 22649 29115 22707 29121
rect 23198 29112 23204 29164
rect 23256 29152 23262 29164
rect 24581 29155 24639 29161
rect 24581 29152 24593 29155
rect 23256 29124 24593 29152
rect 23256 29112 23262 29124
rect 24581 29121 24593 29124
rect 24627 29121 24639 29155
rect 24581 29115 24639 29121
rect 24673 29155 24731 29161
rect 24673 29121 24685 29155
rect 24719 29121 24731 29155
rect 24673 29115 24731 29121
rect 23382 29044 23388 29096
rect 23440 29084 23446 29096
rect 24688 29084 24716 29115
rect 24762 29112 24768 29164
rect 24820 29152 24826 29164
rect 24946 29152 24952 29164
rect 24820 29124 24865 29152
rect 24907 29124 24952 29152
rect 24820 29112 24826 29124
rect 24946 29112 24952 29124
rect 25004 29112 25010 29164
rect 28442 29152 28448 29164
rect 28403 29124 28448 29152
rect 28442 29112 28448 29124
rect 28500 29112 28506 29164
rect 28718 29152 28724 29164
rect 28679 29124 28724 29152
rect 28718 29112 28724 29124
rect 28776 29112 28782 29164
rect 29656 29152 29684 29192
rect 29733 29189 29745 29223
rect 29779 29189 29791 29223
rect 34514 29220 34520 29232
rect 29733 29183 29791 29189
rect 33612 29192 34520 29220
rect 30374 29152 30380 29164
rect 29656 29124 30380 29152
rect 30374 29112 30380 29124
rect 30432 29112 30438 29164
rect 33612 29161 33640 29192
rect 34514 29180 34520 29192
rect 34572 29180 34578 29232
rect 34790 29180 34796 29232
rect 34848 29220 34854 29232
rect 35805 29223 35863 29229
rect 35805 29220 35817 29223
rect 34848 29192 35817 29220
rect 34848 29180 34854 29192
rect 35805 29189 35817 29192
rect 35851 29189 35863 29223
rect 35805 29183 35863 29189
rect 36633 29223 36691 29229
rect 36633 29189 36645 29223
rect 36679 29220 36691 29223
rect 37461 29223 37519 29229
rect 37461 29220 37473 29223
rect 36679 29192 37473 29220
rect 36679 29189 36691 29192
rect 36633 29183 36691 29189
rect 37461 29189 37473 29192
rect 37507 29189 37519 29223
rect 37461 29183 37519 29189
rect 32585 29155 32643 29161
rect 32585 29152 32597 29155
rect 31726 29124 32597 29152
rect 23440 29056 24716 29084
rect 23440 29044 23446 29056
rect 22646 29016 22652 29028
rect 22296 28988 22652 29016
rect 22646 28976 22652 28988
rect 22704 28976 22710 29028
rect 24688 29016 24716 29056
rect 25590 29044 25596 29096
rect 25648 29084 25654 29096
rect 27617 29087 27675 29093
rect 27617 29084 27629 29087
rect 25648 29056 27629 29084
rect 25648 29044 25654 29056
rect 27617 29053 27629 29056
rect 27663 29084 27675 29087
rect 31726 29084 31754 29124
rect 32585 29121 32597 29124
rect 32631 29121 32643 29155
rect 32585 29115 32643 29121
rect 33597 29155 33655 29161
rect 33597 29121 33609 29155
rect 33643 29121 33655 29155
rect 33597 29115 33655 29121
rect 33864 29155 33922 29161
rect 33864 29121 33876 29155
rect 33910 29152 33922 29155
rect 35437 29155 35495 29161
rect 35437 29152 35449 29155
rect 33910 29124 35449 29152
rect 33910 29121 33922 29124
rect 33864 29115 33922 29121
rect 35437 29121 35449 29124
rect 35483 29121 35495 29155
rect 35437 29115 35495 29121
rect 35526 29112 35532 29164
rect 35584 29152 35590 29164
rect 35621 29155 35679 29161
rect 35621 29152 35633 29155
rect 35584 29124 35633 29152
rect 35584 29112 35590 29124
rect 35621 29121 35633 29124
rect 35667 29121 35679 29155
rect 35621 29115 35679 29121
rect 35897 29155 35955 29161
rect 35897 29121 35909 29155
rect 35943 29121 35955 29155
rect 35897 29115 35955 29121
rect 36541 29155 36599 29161
rect 36541 29121 36553 29155
rect 36587 29121 36599 29155
rect 37274 29152 37280 29164
rect 37235 29124 37280 29152
rect 36541 29115 36599 29121
rect 27663 29056 31754 29084
rect 27663 29053 27675 29056
rect 27617 29047 27675 29053
rect 34698 29044 34704 29096
rect 34756 29084 34762 29096
rect 35912 29084 35940 29115
rect 34756 29056 35940 29084
rect 36556 29084 36584 29115
rect 37274 29112 37280 29124
rect 37332 29112 37338 29164
rect 46934 29112 46940 29164
rect 46992 29152 46998 29164
rect 47581 29155 47639 29161
rect 47581 29152 47593 29155
rect 46992 29124 47593 29152
rect 46992 29112 46998 29124
rect 47581 29121 47593 29124
rect 47627 29121 47639 29155
rect 47581 29115 47639 29121
rect 37458 29084 37464 29096
rect 36556 29056 37464 29084
rect 34756 29044 34762 29056
rect 37458 29044 37464 29056
rect 37516 29084 37522 29096
rect 38470 29084 38476 29096
rect 37516 29056 38476 29084
rect 37516 29044 37522 29056
rect 38470 29044 38476 29056
rect 38528 29044 38534 29096
rect 39117 29087 39175 29093
rect 39117 29053 39129 29087
rect 39163 29084 39175 29087
rect 39574 29084 39580 29096
rect 39163 29056 39580 29084
rect 39163 29053 39175 29056
rect 39117 29047 39175 29053
rect 39574 29044 39580 29056
rect 39632 29044 39638 29096
rect 28994 29016 29000 29028
rect 24688 28988 29000 29016
rect 28994 28976 29000 28988
rect 29052 29016 29058 29028
rect 29362 29016 29368 29028
rect 29052 28988 29368 29016
rect 29052 28976 29058 28988
rect 29362 28976 29368 28988
rect 29420 28976 29426 29028
rect 34882 29016 34888 29028
rect 34716 28988 34888 29016
rect 2038 28948 2044 28960
rect 1999 28920 2044 28948
rect 2038 28908 2044 28920
rect 2096 28908 2102 28960
rect 29086 28908 29092 28960
rect 29144 28948 29150 28960
rect 29822 28948 29828 28960
rect 29144 28920 29828 28948
rect 29144 28908 29150 28920
rect 29822 28908 29828 28920
rect 29880 28948 29886 28960
rect 29917 28951 29975 28957
rect 29917 28948 29929 28951
rect 29880 28920 29929 28948
rect 29880 28908 29886 28920
rect 29917 28917 29929 28920
rect 29963 28917 29975 28951
rect 29917 28911 29975 28917
rect 34238 28908 34244 28960
rect 34296 28948 34302 28960
rect 34716 28948 34744 28988
rect 34882 28976 34888 28988
rect 34940 28976 34946 29028
rect 46566 28976 46572 29028
rect 46624 29016 46630 29028
rect 47673 29019 47731 29025
rect 47673 29016 47685 29019
rect 46624 28988 47685 29016
rect 46624 28976 46630 28988
rect 47673 28985 47685 28988
rect 47719 28985 47731 29019
rect 47673 28979 47731 28985
rect 34296 28920 34744 28948
rect 34296 28908 34302 28920
rect 34790 28908 34796 28960
rect 34848 28948 34854 28960
rect 34977 28951 35035 28957
rect 34977 28948 34989 28951
rect 34848 28920 34989 28948
rect 34848 28908 34854 28920
rect 34977 28917 34989 28920
rect 35023 28917 35035 28951
rect 34977 28911 35035 28917
rect 1104 28858 48852 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 48852 28858
rect 1104 28784 48852 28806
rect 26418 28744 26424 28756
rect 19260 28716 26424 28744
rect 1397 28611 1455 28617
rect 1397 28577 1409 28611
rect 1443 28608 1455 28611
rect 2038 28608 2044 28620
rect 1443 28580 2044 28608
rect 1443 28577 1455 28580
rect 1397 28571 1455 28577
rect 2038 28568 2044 28580
rect 2096 28568 2102 28620
rect 2774 28608 2780 28620
rect 2735 28580 2780 28608
rect 2774 28568 2780 28580
rect 2832 28568 2838 28620
rect 19260 28549 19288 28716
rect 26418 28704 26424 28716
rect 26476 28704 26482 28756
rect 26602 28704 26608 28756
rect 26660 28744 26666 28756
rect 26881 28747 26939 28753
rect 26881 28744 26893 28747
rect 26660 28716 26893 28744
rect 26660 28704 26666 28716
rect 26881 28713 26893 28716
rect 26927 28713 26939 28747
rect 27982 28744 27988 28756
rect 27943 28716 27988 28744
rect 26881 28707 26939 28713
rect 27982 28704 27988 28716
rect 28040 28704 28046 28756
rect 32214 28744 32220 28756
rect 31680 28716 32220 28744
rect 24670 28636 24676 28688
rect 24728 28676 24734 28688
rect 28905 28679 28963 28685
rect 24728 28648 28764 28676
rect 24728 28636 24734 28648
rect 22830 28568 22836 28620
rect 22888 28608 22894 28620
rect 25774 28608 25780 28620
rect 22888 28580 24808 28608
rect 22888 28568 22894 28580
rect 19245 28543 19303 28549
rect 19245 28509 19257 28543
rect 19291 28509 19303 28543
rect 19245 28503 19303 28509
rect 22002 28500 22008 28552
rect 22060 28540 22066 28552
rect 22189 28543 22247 28549
rect 22189 28540 22201 28543
rect 22060 28512 22201 28540
rect 22060 28500 22066 28512
rect 22189 28509 22201 28512
rect 22235 28509 22247 28543
rect 24670 28540 24676 28552
rect 24631 28512 24676 28540
rect 22189 28503 22247 28509
rect 24670 28500 24676 28512
rect 24728 28500 24734 28552
rect 24780 28549 24808 28580
rect 25516 28580 25780 28608
rect 24765 28543 24823 28549
rect 24765 28509 24777 28543
rect 24811 28509 24823 28543
rect 24765 28503 24823 28509
rect 24854 28500 24860 28552
rect 24912 28540 24918 28552
rect 25041 28543 25099 28549
rect 24912 28512 24957 28540
rect 24912 28500 24918 28512
rect 25041 28509 25053 28543
rect 25087 28540 25099 28543
rect 25222 28540 25228 28552
rect 25087 28512 25228 28540
rect 25087 28509 25099 28512
rect 25041 28503 25099 28509
rect 25222 28500 25228 28512
rect 25280 28500 25286 28552
rect 25516 28549 25544 28580
rect 25774 28568 25780 28580
rect 25832 28568 25838 28620
rect 26418 28568 26424 28620
rect 26476 28608 26482 28620
rect 27154 28608 27160 28620
rect 26476 28580 27160 28608
rect 26476 28568 26482 28580
rect 27154 28568 27160 28580
rect 27212 28568 27218 28620
rect 27617 28611 27675 28617
rect 27617 28577 27629 28611
rect 27663 28608 27675 28611
rect 27663 28580 28580 28608
rect 27663 28577 27675 28580
rect 27617 28571 27675 28577
rect 25501 28543 25559 28549
rect 25501 28509 25513 28543
rect 25547 28509 25559 28543
rect 25501 28503 25559 28509
rect 26326 28500 26332 28552
rect 26384 28540 26390 28552
rect 26789 28543 26847 28549
rect 26789 28540 26801 28543
rect 26384 28512 26801 28540
rect 26384 28500 26390 28512
rect 26789 28509 26801 28512
rect 26835 28509 26847 28543
rect 26789 28503 26847 28509
rect 27065 28543 27123 28549
rect 27065 28509 27077 28543
rect 27111 28540 27123 28543
rect 27632 28540 27660 28571
rect 27111 28512 27660 28540
rect 27801 28543 27859 28549
rect 27111 28509 27123 28512
rect 27065 28503 27123 28509
rect 27801 28509 27813 28543
rect 27847 28509 27859 28543
rect 27801 28503 27859 28509
rect 1581 28475 1639 28481
rect 1581 28441 1593 28475
rect 1627 28472 1639 28475
rect 2314 28472 2320 28484
rect 1627 28444 2320 28472
rect 1627 28441 1639 28444
rect 1581 28435 1639 28441
rect 2314 28432 2320 28444
rect 2372 28432 2378 28484
rect 17310 28432 17316 28484
rect 17368 28472 17374 28484
rect 17681 28475 17739 28481
rect 17681 28472 17693 28475
rect 17368 28444 17693 28472
rect 17368 28432 17374 28444
rect 17681 28441 17693 28444
rect 17727 28441 17739 28475
rect 17681 28435 17739 28441
rect 17865 28475 17923 28481
rect 17865 28441 17877 28475
rect 17911 28472 17923 28475
rect 18322 28472 18328 28484
rect 17911 28444 18328 28472
rect 17911 28441 17923 28444
rect 17865 28435 17923 28441
rect 18322 28432 18328 28444
rect 18380 28432 18386 28484
rect 21174 28432 21180 28484
rect 21232 28472 21238 28484
rect 23382 28472 23388 28484
rect 21232 28444 23388 28472
rect 21232 28432 21238 28444
rect 23382 28432 23388 28444
rect 23440 28432 23446 28484
rect 23477 28475 23535 28481
rect 23477 28441 23489 28475
rect 23523 28472 23535 28475
rect 24578 28472 24584 28484
rect 23523 28444 24584 28472
rect 23523 28441 23535 28444
rect 23477 28435 23535 28441
rect 24578 28432 24584 28444
rect 24636 28472 24642 28484
rect 25685 28475 25743 28481
rect 25685 28472 25697 28475
rect 24636 28444 25697 28472
rect 24636 28432 24642 28444
rect 25685 28441 25697 28444
rect 25731 28441 25743 28475
rect 26804 28472 26832 28503
rect 27430 28472 27436 28484
rect 26804 28444 27436 28472
rect 25685 28435 25743 28441
rect 27430 28432 27436 28444
rect 27488 28472 27494 28484
rect 27816 28472 27844 28503
rect 28552 28484 28580 28580
rect 28736 28549 28764 28648
rect 28905 28645 28917 28679
rect 28951 28676 28963 28679
rect 28994 28676 29000 28688
rect 28951 28648 29000 28676
rect 28951 28645 28963 28648
rect 28905 28639 28963 28645
rect 28994 28636 29000 28648
rect 29052 28636 29058 28688
rect 31680 28549 31708 28716
rect 32214 28704 32220 28716
rect 32272 28744 32278 28756
rect 32272 28716 36492 28744
rect 32272 28704 32278 28716
rect 31754 28636 31760 28688
rect 31812 28676 31818 28688
rect 31812 28648 32904 28676
rect 31812 28636 31818 28648
rect 32876 28549 32904 28648
rect 36464 28617 36492 28716
rect 37458 28636 37464 28688
rect 37516 28676 37522 28688
rect 38749 28679 38807 28685
rect 38749 28676 38761 28679
rect 37516 28648 38761 28676
rect 37516 28636 37522 28648
rect 38749 28645 38761 28648
rect 38795 28645 38807 28679
rect 38749 28639 38807 28645
rect 36449 28611 36507 28617
rect 33888 28580 35296 28608
rect 33888 28552 33916 28580
rect 28721 28543 28779 28549
rect 28721 28509 28733 28543
rect 28767 28509 28779 28543
rect 31680 28543 31756 28549
rect 31680 28512 31710 28543
rect 28721 28503 28779 28509
rect 31698 28509 31710 28512
rect 31744 28509 31756 28543
rect 31698 28503 31756 28509
rect 32125 28543 32183 28549
rect 32125 28509 32137 28543
rect 32171 28509 32183 28543
rect 32125 28503 32183 28509
rect 32217 28543 32275 28549
rect 32217 28509 32229 28543
rect 32263 28509 32275 28543
rect 32217 28503 32275 28509
rect 32861 28543 32919 28549
rect 32861 28509 32873 28543
rect 32907 28509 32919 28543
rect 32861 28503 32919 28509
rect 27488 28444 27844 28472
rect 27488 28432 27494 28444
rect 28534 28432 28540 28484
rect 28592 28472 28598 28484
rect 31846 28472 31852 28484
rect 28592 28444 31852 28472
rect 28592 28432 28598 28444
rect 31846 28432 31852 28444
rect 31904 28472 31910 28484
rect 32140 28472 32168 28503
rect 31904 28444 32168 28472
rect 32232 28472 32260 28503
rect 32950 28500 32956 28552
rect 33008 28540 33014 28552
rect 33045 28543 33103 28549
rect 33045 28540 33057 28543
rect 33008 28512 33057 28540
rect 33008 28500 33014 28512
rect 33045 28509 33057 28512
rect 33091 28509 33103 28543
rect 33870 28540 33876 28552
rect 33831 28512 33876 28540
rect 33045 28503 33103 28509
rect 33870 28500 33876 28512
rect 33928 28500 33934 28552
rect 34057 28543 34115 28549
rect 34057 28509 34069 28543
rect 34103 28509 34115 28543
rect 34057 28503 34115 28509
rect 32674 28472 32680 28484
rect 32232 28444 32680 28472
rect 31904 28432 31910 28444
rect 32674 28432 32680 28444
rect 32732 28472 32738 28484
rect 34072 28472 34100 28503
rect 34146 28500 34152 28552
rect 34204 28540 34210 28552
rect 35268 28549 35296 28580
rect 36449 28577 36461 28611
rect 36495 28577 36507 28611
rect 36449 28571 36507 28577
rect 38289 28611 38347 28617
rect 38289 28577 38301 28611
rect 38335 28608 38347 28611
rect 39298 28608 39304 28620
rect 38335 28580 39304 28608
rect 38335 28577 38347 28580
rect 38289 28571 38347 28577
rect 39298 28568 39304 28580
rect 39356 28568 39362 28620
rect 48130 28608 48136 28620
rect 48091 28580 48136 28608
rect 48130 28568 48136 28580
rect 48188 28568 48194 28620
rect 34701 28543 34759 28549
rect 34701 28540 34713 28543
rect 34204 28512 34713 28540
rect 34204 28500 34210 28512
rect 34701 28509 34713 28512
rect 34747 28509 34759 28543
rect 34701 28503 34759 28509
rect 34885 28543 34943 28549
rect 34885 28509 34897 28543
rect 34931 28509 34943 28543
rect 34885 28503 34943 28509
rect 35253 28543 35311 28549
rect 35253 28509 35265 28543
rect 35299 28509 35311 28543
rect 35253 28503 35311 28509
rect 34790 28472 34796 28484
rect 32732 28444 33824 28472
rect 34072 28444 34796 28472
rect 32732 28432 32738 28444
rect 18049 28407 18107 28413
rect 18049 28373 18061 28407
rect 18095 28404 18107 28407
rect 18690 28404 18696 28416
rect 18095 28376 18696 28404
rect 18095 28373 18107 28376
rect 18049 28367 18107 28373
rect 18690 28364 18696 28376
rect 18748 28364 18754 28416
rect 19334 28404 19340 28416
rect 19295 28376 19340 28404
rect 19334 28364 19340 28376
rect 19392 28364 19398 28416
rect 19978 28364 19984 28416
rect 20036 28404 20042 28416
rect 20346 28404 20352 28416
rect 20036 28376 20352 28404
rect 20036 28364 20042 28376
rect 20346 28364 20352 28376
rect 20404 28364 20410 28416
rect 22278 28404 22284 28416
rect 22239 28376 22284 28404
rect 22278 28364 22284 28376
rect 22336 28364 22342 28416
rect 23569 28407 23627 28413
rect 23569 28373 23581 28407
rect 23615 28404 23627 28407
rect 23658 28404 23664 28416
rect 23615 28376 23664 28404
rect 23615 28373 23627 28376
rect 23569 28367 23627 28373
rect 23658 28364 23664 28376
rect 23716 28364 23722 28416
rect 24394 28404 24400 28416
rect 24355 28376 24400 28404
rect 24394 28364 24400 28376
rect 24452 28364 24458 28416
rect 25222 28364 25228 28416
rect 25280 28404 25286 28416
rect 25869 28407 25927 28413
rect 25869 28404 25881 28407
rect 25280 28376 25881 28404
rect 25280 28364 25286 28376
rect 25869 28373 25881 28376
rect 25915 28373 25927 28407
rect 31570 28404 31576 28416
rect 31531 28376 31576 28404
rect 25869 28367 25927 28373
rect 31570 28364 31576 28376
rect 31628 28364 31634 28416
rect 31757 28407 31815 28413
rect 31757 28373 31769 28407
rect 31803 28404 31815 28407
rect 32953 28407 33011 28413
rect 32953 28404 32965 28407
rect 31803 28376 32965 28404
rect 31803 28373 31815 28376
rect 31757 28367 31815 28373
rect 32953 28373 32965 28376
rect 32999 28373 33011 28407
rect 32953 28367 33011 28373
rect 33594 28364 33600 28416
rect 33652 28404 33658 28416
rect 33689 28407 33747 28413
rect 33689 28404 33701 28407
rect 33652 28376 33701 28404
rect 33652 28364 33658 28376
rect 33689 28373 33701 28376
rect 33735 28373 33747 28407
rect 33796 28404 33824 28444
rect 34790 28432 34796 28444
rect 34848 28472 34854 28484
rect 34900 28472 34928 28503
rect 38654 28500 38660 28552
rect 38712 28540 38718 28552
rect 38933 28543 38991 28549
rect 38933 28540 38945 28543
rect 38712 28512 38945 28540
rect 38712 28500 38718 28512
rect 38933 28509 38945 28512
rect 38979 28509 38991 28543
rect 38933 28503 38991 28509
rect 39022 28500 39028 28552
rect 39080 28540 39086 28552
rect 39080 28512 39125 28540
rect 39080 28500 39086 28512
rect 46106 28500 46112 28552
rect 46164 28540 46170 28552
rect 46293 28543 46351 28549
rect 46293 28540 46305 28543
rect 46164 28512 46305 28540
rect 46164 28500 46170 28512
rect 46293 28509 46305 28512
rect 46339 28509 46351 28543
rect 46293 28503 46351 28509
rect 34848 28444 34928 28472
rect 35161 28475 35219 28481
rect 34848 28432 34854 28444
rect 35161 28441 35173 28475
rect 35207 28441 35219 28475
rect 36630 28472 36636 28484
rect 36591 28444 36636 28472
rect 35161 28435 35219 28441
rect 35176 28404 35204 28435
rect 36630 28432 36636 28444
rect 36688 28432 36694 28484
rect 38749 28475 38807 28481
rect 38749 28441 38761 28475
rect 38795 28472 38807 28475
rect 39850 28472 39856 28484
rect 38795 28444 39856 28472
rect 38795 28441 38807 28444
rect 38749 28435 38807 28441
rect 39850 28432 39856 28444
rect 39908 28432 39914 28484
rect 46474 28472 46480 28484
rect 46435 28444 46480 28472
rect 46474 28432 46480 28444
rect 46532 28432 46538 28484
rect 37366 28404 37372 28416
rect 33796 28376 37372 28404
rect 33689 28367 33747 28373
rect 37366 28364 37372 28376
rect 37424 28364 37430 28416
rect 1104 28314 48852 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 48852 28314
rect 1104 28240 48852 28262
rect 2314 28200 2320 28212
rect 2275 28172 2320 28200
rect 2314 28160 2320 28172
rect 2372 28160 2378 28212
rect 18322 28160 18328 28212
rect 18380 28200 18386 28212
rect 18380 28172 20024 28200
rect 18380 28160 18386 28172
rect 17580 28135 17638 28141
rect 17580 28101 17592 28135
rect 17626 28132 17638 28135
rect 19153 28135 19211 28141
rect 19153 28132 19165 28135
rect 17626 28104 19165 28132
rect 17626 28101 17638 28104
rect 17580 28095 17638 28101
rect 19153 28101 19165 28104
rect 19199 28101 19211 28135
rect 19996 28132 20024 28172
rect 20806 28160 20812 28212
rect 20864 28200 20870 28212
rect 20864 28172 25728 28200
rect 20864 28160 20870 28172
rect 20257 28135 20315 28141
rect 19996 28104 20208 28132
rect 19153 28095 19211 28101
rect 2225 28067 2283 28073
rect 2225 28033 2237 28067
rect 2271 28064 2283 28067
rect 2866 28064 2872 28076
rect 2271 28036 2872 28064
rect 2271 28033 2283 28036
rect 2225 28027 2283 28033
rect 2866 28024 2872 28036
rect 2924 28064 2930 28076
rect 3142 28064 3148 28076
rect 2924 28036 3148 28064
rect 2924 28024 2930 28036
rect 3142 28024 3148 28036
rect 3200 28024 3206 28076
rect 12618 28064 12624 28076
rect 12579 28036 12624 28064
rect 12618 28024 12624 28036
rect 12676 28024 12682 28076
rect 19383 28067 19441 28073
rect 19383 28033 19395 28067
rect 19429 28033 19441 28067
rect 19515 28064 19521 28076
rect 19476 28036 19521 28064
rect 19383 28027 19441 28033
rect 1670 27956 1676 28008
rect 1728 27996 1734 28008
rect 2314 27996 2320 28008
rect 1728 27968 2320 27996
rect 1728 27956 1734 27968
rect 2314 27956 2320 27968
rect 2372 27956 2378 28008
rect 16850 27956 16856 28008
rect 16908 27996 16914 28008
rect 17313 27999 17371 28005
rect 17313 27996 17325 27999
rect 16908 27968 17325 27996
rect 16908 27956 16914 27968
rect 17313 27965 17325 27968
rect 17359 27965 17371 27999
rect 17313 27959 17371 27965
rect 12710 27860 12716 27872
rect 12671 27832 12716 27860
rect 12710 27820 12716 27832
rect 12768 27820 12774 27872
rect 18230 27820 18236 27872
rect 18288 27860 18294 27872
rect 18693 27863 18751 27869
rect 18693 27860 18705 27863
rect 18288 27832 18705 27860
rect 18288 27820 18294 27832
rect 18693 27829 18705 27832
rect 18739 27829 18751 27863
rect 19398 27860 19426 28027
rect 19515 28024 19521 28036
rect 19573 28024 19579 28076
rect 19613 28067 19671 28073
rect 19613 28033 19625 28067
rect 19659 28033 19671 28067
rect 19613 28027 19671 28033
rect 19797 28067 19855 28073
rect 19797 28033 19809 28067
rect 19843 28064 19855 28067
rect 20070 28064 20076 28076
rect 19843 28036 20076 28064
rect 19843 28033 19855 28036
rect 19797 28027 19855 28033
rect 19628 27928 19656 28027
rect 20070 28024 20076 28036
rect 20128 28024 20134 28076
rect 20180 28064 20208 28104
rect 20257 28101 20269 28135
rect 20303 28132 20315 28135
rect 20824 28132 20852 28160
rect 23934 28132 23940 28144
rect 20303 28104 20852 28132
rect 22572 28104 23704 28132
rect 20303 28101 20315 28104
rect 20257 28095 20315 28101
rect 22572 28076 22600 28104
rect 20441 28067 20499 28073
rect 20441 28064 20453 28067
rect 20180 28036 20453 28064
rect 20441 28033 20453 28036
rect 20487 28064 20499 28067
rect 21082 28064 21088 28076
rect 20487 28036 21088 28064
rect 20487 28033 20499 28036
rect 20441 28027 20499 28033
rect 21082 28024 21088 28036
rect 21140 28024 21146 28076
rect 21450 28064 21456 28076
rect 21192 28036 21456 28064
rect 21192 27996 21220 28036
rect 21450 28024 21456 28036
rect 21508 28064 21514 28076
rect 22554 28064 22560 28076
rect 21508 28036 22560 28064
rect 21508 28024 21514 28036
rect 22554 28024 22560 28036
rect 22612 28024 22618 28076
rect 22649 28067 22707 28073
rect 22649 28033 22661 28067
rect 22695 28033 22707 28067
rect 22649 28027 22707 28033
rect 22741 28067 22799 28073
rect 22741 28033 22753 28067
rect 22787 28033 22799 28067
rect 22741 28027 22799 28033
rect 22925 28067 22983 28073
rect 22925 28033 22937 28067
rect 22971 28064 22983 28067
rect 23474 28064 23480 28076
rect 22971 28036 23480 28064
rect 22971 28033 22983 28036
rect 22925 28027 22983 28033
rect 19904 27968 21220 27996
rect 19794 27928 19800 27940
rect 19628 27900 19800 27928
rect 19794 27888 19800 27900
rect 19852 27888 19858 27940
rect 19610 27860 19616 27872
rect 19398 27832 19616 27860
rect 18693 27823 18751 27829
rect 19610 27820 19616 27832
rect 19668 27860 19674 27872
rect 19904 27860 19932 27968
rect 21266 27956 21272 28008
rect 21324 27996 21330 28008
rect 22664 27996 22692 28027
rect 21324 27968 22692 27996
rect 22756 27996 22784 28027
rect 23474 28024 23480 28036
rect 23532 28024 23538 28076
rect 23676 28073 23704 28104
rect 23768 28104 23940 28132
rect 23768 28073 23796 28104
rect 23934 28092 23940 28104
rect 23992 28092 23998 28144
rect 24394 28092 24400 28144
rect 24452 28132 24458 28144
rect 25286 28135 25344 28141
rect 25286 28132 25298 28135
rect 24452 28104 25298 28132
rect 24452 28092 24458 28104
rect 25286 28101 25298 28104
rect 25332 28101 25344 28135
rect 25700 28132 25728 28172
rect 25774 28160 25780 28212
rect 25832 28200 25838 28212
rect 26421 28203 26479 28209
rect 26421 28200 26433 28203
rect 25832 28172 26433 28200
rect 25832 28160 25838 28172
rect 26421 28169 26433 28172
rect 26467 28200 26479 28203
rect 36541 28203 36599 28209
rect 26467 28172 35480 28200
rect 26467 28169 26479 28172
rect 26421 28163 26479 28169
rect 34333 28135 34391 28141
rect 25700 28104 33824 28132
rect 25286 28095 25344 28101
rect 23661 28067 23719 28073
rect 23661 28033 23673 28067
rect 23707 28033 23719 28067
rect 23661 28027 23719 28033
rect 23753 28067 23811 28073
rect 23753 28033 23765 28067
rect 23799 28033 23811 28067
rect 23753 28027 23811 28033
rect 23845 28067 23903 28073
rect 23845 28033 23857 28067
rect 23891 28033 23903 28067
rect 24026 28064 24032 28076
rect 23987 28036 24032 28064
rect 23845 28027 23903 28033
rect 23860 27996 23888 28027
rect 24026 28024 24032 28036
rect 24084 28024 24090 28076
rect 25038 28064 25044 28076
rect 24999 28036 25044 28064
rect 25038 28024 25044 28036
rect 25096 28024 25102 28076
rect 28445 28067 28503 28073
rect 28445 28033 28457 28067
rect 28491 28064 28503 28067
rect 28534 28064 28540 28076
rect 28491 28036 28540 28064
rect 28491 28033 28503 28036
rect 28445 28027 28503 28033
rect 28534 28024 28540 28036
rect 28592 28024 28598 28076
rect 29546 28024 29552 28076
rect 29604 28064 29610 28076
rect 29989 28067 30047 28073
rect 29989 28064 30001 28067
rect 29604 28036 30001 28064
rect 29604 28024 29610 28036
rect 29989 28033 30001 28036
rect 30035 28033 30047 28067
rect 29989 28027 30047 28033
rect 31570 28024 31576 28076
rect 31628 28064 31634 28076
rect 32125 28067 32183 28073
rect 32125 28064 32137 28067
rect 31628 28036 32137 28064
rect 31628 28024 31634 28036
rect 32125 28033 32137 28036
rect 32171 28033 32183 28067
rect 32306 28064 32312 28076
rect 32267 28036 32312 28064
rect 32125 28027 32183 28033
rect 32306 28024 32312 28036
rect 32364 28024 32370 28076
rect 24762 27996 24768 28008
rect 22756 27968 24768 27996
rect 21324 27956 21330 27968
rect 24762 27956 24768 27968
rect 24820 27956 24826 28008
rect 29454 27956 29460 28008
rect 29512 27996 29518 28008
rect 29733 27999 29791 28005
rect 29733 27996 29745 27999
rect 29512 27968 29745 27996
rect 29512 27956 29518 27968
rect 29733 27965 29745 27968
rect 29779 27965 29791 27999
rect 29733 27959 29791 27965
rect 21082 27888 21088 27940
rect 21140 27928 21146 27940
rect 23658 27928 23664 27940
rect 21140 27900 23664 27928
rect 21140 27888 21146 27900
rect 23658 27888 23664 27900
rect 23716 27888 23722 27940
rect 31113 27931 31171 27937
rect 31113 27897 31125 27931
rect 31159 27928 31171 27931
rect 31846 27928 31852 27940
rect 31159 27900 31852 27928
rect 31159 27897 31171 27900
rect 31113 27891 31171 27897
rect 31846 27888 31852 27900
rect 31904 27888 31910 27940
rect 31938 27888 31944 27940
rect 31996 27928 32002 27940
rect 33796 27928 33824 28104
rect 34333 28101 34345 28135
rect 34379 28132 34391 28135
rect 34698 28132 34704 28144
rect 34379 28104 34704 28132
rect 34379 28101 34391 28104
rect 34333 28095 34391 28101
rect 34698 28092 34704 28104
rect 34756 28092 34762 28144
rect 33870 28024 33876 28076
rect 33928 28064 33934 28076
rect 34241 28067 34299 28073
rect 34241 28064 34253 28067
rect 33928 28036 34253 28064
rect 33928 28024 33934 28036
rect 34241 28033 34253 28036
rect 34287 28033 34299 28067
rect 34241 28027 34299 28033
rect 35452 27996 35480 28172
rect 36541 28169 36553 28203
rect 36587 28200 36599 28203
rect 36630 28200 36636 28212
rect 36587 28172 36636 28200
rect 36587 28169 36599 28172
rect 36541 28163 36599 28169
rect 36630 28160 36636 28172
rect 36688 28160 36694 28212
rect 37550 28200 37556 28212
rect 37511 28172 37556 28200
rect 37550 28160 37556 28172
rect 37608 28160 37614 28212
rect 35526 28092 35532 28144
rect 35584 28132 35590 28144
rect 38657 28135 38715 28141
rect 35584 28104 37688 28132
rect 35584 28092 35590 28104
rect 35986 28024 35992 28076
rect 36044 28064 36050 28076
rect 36449 28067 36507 28073
rect 36449 28064 36461 28067
rect 36044 28036 36461 28064
rect 36044 28024 36050 28036
rect 36449 28033 36461 28036
rect 36495 28033 36507 28067
rect 37458 28064 37464 28076
rect 37419 28036 37464 28064
rect 36449 28027 36507 28033
rect 37458 28024 37464 28036
rect 37516 28024 37522 28076
rect 37660 28073 37688 28104
rect 38657 28101 38669 28135
rect 38703 28132 38715 28135
rect 39393 28135 39451 28141
rect 39393 28132 39405 28135
rect 38703 28104 39405 28132
rect 38703 28101 38715 28104
rect 38657 28095 38715 28101
rect 39393 28101 39405 28104
rect 39439 28101 39451 28135
rect 39393 28095 39451 28101
rect 37645 28067 37703 28073
rect 37645 28033 37657 28067
rect 37691 28033 37703 28067
rect 37645 28027 37703 28033
rect 38470 28024 38476 28076
rect 38528 28064 38534 28076
rect 38565 28067 38623 28073
rect 38565 28064 38577 28067
rect 38528 28036 38577 28064
rect 38528 28024 38534 28036
rect 38565 28033 38577 28036
rect 38611 28033 38623 28067
rect 47854 28064 47860 28076
rect 47815 28036 47860 28064
rect 38565 28027 38623 28033
rect 47854 28024 47860 28036
rect 47912 28024 47918 28076
rect 39209 27999 39267 28005
rect 39209 27996 39221 27999
rect 35452 27968 39221 27996
rect 39209 27965 39221 27968
rect 39255 27965 39267 27999
rect 39209 27959 39267 27965
rect 41049 27999 41107 28005
rect 41049 27965 41061 27999
rect 41095 27996 41107 27999
rect 44726 27996 44732 28008
rect 41095 27968 44732 27996
rect 41095 27965 41107 27968
rect 41049 27959 41107 27965
rect 44726 27956 44732 27968
rect 44784 27956 44790 28008
rect 45189 27999 45247 28005
rect 45189 27965 45201 27999
rect 45235 27965 45247 27999
rect 45189 27959 45247 27965
rect 45373 27999 45431 28005
rect 45373 27965 45385 27999
rect 45419 27996 45431 27999
rect 45554 27996 45560 28008
rect 45419 27968 45560 27996
rect 45419 27965 45431 27968
rect 45373 27959 45431 27965
rect 45204 27928 45232 27959
rect 45554 27956 45560 27968
rect 45612 27956 45618 28008
rect 46014 27996 46020 28008
rect 45975 27968 46020 27996
rect 46014 27956 46020 27968
rect 46072 27956 46078 28008
rect 31996 27900 33272 27928
rect 33796 27900 45232 27928
rect 31996 27888 32002 27900
rect 33244 27872 33272 27900
rect 19668 27832 19932 27860
rect 19668 27820 19674 27832
rect 19978 27820 19984 27872
rect 20036 27860 20042 27872
rect 20625 27863 20683 27869
rect 20625 27860 20637 27863
rect 20036 27832 20637 27860
rect 20036 27820 20042 27832
rect 20625 27829 20637 27832
rect 20671 27829 20683 27863
rect 20625 27823 20683 27829
rect 22281 27863 22339 27869
rect 22281 27829 22293 27863
rect 22327 27860 22339 27863
rect 22738 27860 22744 27872
rect 22327 27832 22744 27860
rect 22327 27829 22339 27832
rect 22281 27823 22339 27829
rect 22738 27820 22744 27832
rect 22796 27820 22802 27872
rect 23385 27863 23443 27869
rect 23385 27829 23397 27863
rect 23431 27860 23443 27863
rect 23934 27860 23940 27872
rect 23431 27832 23940 27860
rect 23431 27829 23443 27832
rect 23385 27823 23443 27829
rect 23934 27820 23940 27832
rect 23992 27820 23998 27872
rect 27430 27820 27436 27872
rect 27488 27860 27494 27872
rect 28537 27863 28595 27869
rect 28537 27860 28549 27863
rect 27488 27832 28549 27860
rect 27488 27820 27494 27832
rect 28537 27829 28549 27832
rect 28583 27829 28595 27863
rect 28537 27823 28595 27829
rect 28905 27863 28963 27869
rect 28905 27829 28917 27863
rect 28951 27860 28963 27863
rect 29638 27860 29644 27872
rect 28951 27832 29644 27860
rect 28951 27829 28963 27832
rect 28905 27823 28963 27829
rect 29638 27820 29644 27832
rect 29696 27820 29702 27872
rect 32122 27860 32128 27872
rect 32083 27832 32128 27860
rect 32122 27820 32128 27832
rect 32180 27820 32186 27872
rect 33226 27820 33232 27872
rect 33284 27860 33290 27872
rect 39022 27860 39028 27872
rect 33284 27832 39028 27860
rect 33284 27820 33290 27832
rect 39022 27820 39028 27832
rect 39080 27820 39086 27872
rect 47670 27820 47676 27872
rect 47728 27860 47734 27872
rect 48041 27863 48099 27869
rect 48041 27860 48053 27863
rect 47728 27832 48053 27860
rect 47728 27820 47734 27832
rect 48041 27829 48053 27832
rect 48087 27829 48099 27863
rect 48041 27823 48099 27829
rect 1104 27770 48852 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 48852 27770
rect 1104 27696 48852 27718
rect 19794 27656 19800 27668
rect 19306 27628 19800 27656
rect 7006 27548 7012 27600
rect 7064 27588 7070 27600
rect 15746 27588 15752 27600
rect 7064 27560 15752 27588
rect 7064 27548 7070 27560
rect 15746 27548 15752 27560
rect 15804 27548 15810 27600
rect 17310 27588 17316 27600
rect 17271 27560 17316 27588
rect 17310 27548 17316 27560
rect 17368 27548 17374 27600
rect 18506 27548 18512 27600
rect 18564 27588 18570 27600
rect 19306 27588 19334 27628
rect 19794 27616 19800 27628
rect 19852 27656 19858 27668
rect 19852 27628 21956 27656
rect 19852 27616 19858 27628
rect 20806 27588 20812 27600
rect 18564 27560 19334 27588
rect 20767 27560 20812 27588
rect 18564 27548 18570 27560
rect 20806 27548 20812 27560
rect 20864 27548 20870 27600
rect 21726 27548 21732 27600
rect 21784 27548 21790 27600
rect 2590 27480 2596 27532
rect 2648 27520 2654 27532
rect 2958 27520 2964 27532
rect 2648 27492 2964 27520
rect 2648 27480 2654 27492
rect 2958 27480 2964 27492
rect 3016 27480 3022 27532
rect 18156 27492 19564 27520
rect 1762 27452 1768 27464
rect 1723 27424 1768 27452
rect 1762 27412 1768 27424
rect 1820 27412 1826 27464
rect 2225 27455 2283 27461
rect 2225 27421 2237 27455
rect 2271 27421 2283 27455
rect 3050 27452 3056 27464
rect 3011 27424 3056 27452
rect 2225 27415 2283 27421
rect 2240 27384 2268 27415
rect 3050 27412 3056 27424
rect 3108 27412 3114 27464
rect 15933 27455 15991 27461
rect 15933 27421 15945 27455
rect 15979 27452 15991 27455
rect 18156 27452 18184 27492
rect 18279 27455 18337 27461
rect 18279 27452 18291 27455
rect 15979 27424 16896 27452
rect 18156 27424 18291 27452
rect 15979 27421 15991 27424
rect 15933 27415 15991 27421
rect 16868 27396 16896 27424
rect 18279 27421 18291 27424
rect 18325 27421 18337 27455
rect 18414 27452 18420 27464
rect 18375 27424 18420 27452
rect 18279 27415 18337 27421
rect 18414 27412 18420 27424
rect 18472 27412 18478 27464
rect 18506 27412 18512 27464
rect 18564 27452 18570 27464
rect 18690 27452 18696 27464
rect 18564 27424 18609 27452
rect 18651 27424 18696 27452
rect 18564 27412 18570 27424
rect 18690 27412 18696 27424
rect 18748 27412 18754 27464
rect 19426 27452 19432 27464
rect 19306 27424 19432 27452
rect 2590 27384 2596 27396
rect 2240 27356 2596 27384
rect 2590 27344 2596 27356
rect 2648 27384 2654 27396
rect 12250 27384 12256 27396
rect 2648 27356 12256 27384
rect 2648 27344 2654 27356
rect 12250 27344 12256 27356
rect 12308 27344 12314 27396
rect 16200 27387 16258 27393
rect 16200 27353 16212 27387
rect 16246 27384 16258 27387
rect 16246 27356 16804 27384
rect 16246 27353 16258 27356
rect 16200 27347 16258 27353
rect 1946 27276 1952 27328
rect 2004 27316 2010 27328
rect 2317 27319 2375 27325
rect 2317 27316 2329 27319
rect 2004 27288 2329 27316
rect 2004 27276 2010 27288
rect 2317 27285 2329 27288
rect 2363 27285 2375 27319
rect 2317 27279 2375 27285
rect 8294 27276 8300 27328
rect 8352 27316 8358 27328
rect 16574 27316 16580 27328
rect 8352 27288 16580 27316
rect 8352 27276 8358 27288
rect 16574 27276 16580 27288
rect 16632 27276 16638 27328
rect 16776 27316 16804 27356
rect 16850 27344 16856 27396
rect 16908 27384 16914 27396
rect 19306 27384 19334 27424
rect 19426 27412 19432 27424
rect 19484 27412 19490 27464
rect 19536 27452 19564 27492
rect 21174 27452 21180 27464
rect 19536 27424 21180 27452
rect 21174 27412 21180 27424
rect 21232 27412 21238 27464
rect 21450 27412 21456 27464
rect 21508 27452 21514 27464
rect 21744 27461 21772 27548
rect 21591 27455 21649 27461
rect 21591 27452 21603 27455
rect 21508 27424 21603 27452
rect 21508 27412 21514 27424
rect 21591 27421 21603 27424
rect 21637 27421 21649 27455
rect 21591 27415 21649 27421
rect 21729 27455 21787 27461
rect 21729 27421 21741 27455
rect 21775 27421 21787 27455
rect 21729 27415 21787 27421
rect 21842 27455 21900 27461
rect 21842 27421 21854 27455
rect 21888 27452 21900 27455
rect 21928 27452 21956 27628
rect 24026 27616 24032 27668
rect 24084 27656 24090 27668
rect 24765 27659 24823 27665
rect 24765 27656 24777 27659
rect 24084 27628 24777 27656
rect 24084 27616 24090 27628
rect 24765 27625 24777 27628
rect 24811 27625 24823 27659
rect 29546 27656 29552 27668
rect 29507 27628 29552 27656
rect 24765 27619 24823 27625
rect 29546 27616 29552 27628
rect 29604 27616 29610 27668
rect 32306 27656 32312 27668
rect 31128 27628 32312 27656
rect 25958 27548 25964 27600
rect 26016 27548 26022 27600
rect 26050 27548 26056 27600
rect 26108 27588 26114 27600
rect 31128 27588 31156 27628
rect 32306 27616 32312 27628
rect 32364 27616 32370 27668
rect 33226 27656 33232 27668
rect 33187 27628 33232 27656
rect 33226 27616 33232 27628
rect 33284 27616 33290 27668
rect 36004 27628 36952 27656
rect 26108 27560 26372 27588
rect 26108 27548 26114 27560
rect 22554 27480 22560 27532
rect 22612 27520 22618 27532
rect 23293 27523 23351 27529
rect 23293 27520 23305 27523
rect 22612 27492 23305 27520
rect 22612 27480 22618 27492
rect 23293 27489 23305 27492
rect 23339 27489 23351 27523
rect 25976 27520 26004 27548
rect 25976 27492 26096 27520
rect 23293 27483 23351 27489
rect 21888 27424 21956 27452
rect 22005 27455 22063 27461
rect 21888 27421 21900 27424
rect 21842 27415 21900 27421
rect 22005 27421 22017 27455
rect 22051 27421 22063 27455
rect 22005 27415 22063 27421
rect 23017 27455 23075 27461
rect 23017 27421 23029 27455
rect 23063 27452 23075 27455
rect 24670 27452 24676 27464
rect 23063 27424 24676 27452
rect 23063 27421 23075 27424
rect 23017 27415 23075 27421
rect 19674 27387 19732 27393
rect 19674 27384 19686 27387
rect 16908 27356 19334 27384
rect 19536 27356 19686 27384
rect 16908 27344 16914 27356
rect 18049 27319 18107 27325
rect 18049 27316 18061 27319
rect 16776 27288 18061 27316
rect 18049 27285 18061 27288
rect 18095 27285 18107 27319
rect 18049 27279 18107 27285
rect 19242 27276 19248 27328
rect 19300 27316 19306 27328
rect 19536 27316 19564 27356
rect 19674 27353 19686 27356
rect 19720 27353 19732 27387
rect 19674 27347 19732 27353
rect 21266 27344 21272 27396
rect 21324 27384 21330 27396
rect 22020 27384 22048 27415
rect 24670 27412 24676 27424
rect 24728 27412 24734 27464
rect 26068 27461 26096 27492
rect 25961 27455 26019 27461
rect 25961 27452 25973 27455
rect 25608 27424 25973 27452
rect 21324 27356 22048 27384
rect 24397 27387 24455 27393
rect 21324 27344 21330 27356
rect 24397 27353 24409 27387
rect 24443 27353 24455 27387
rect 24578 27384 24584 27396
rect 24539 27356 24584 27384
rect 24397 27347 24455 27353
rect 19300 27288 19564 27316
rect 21361 27319 21419 27325
rect 19300 27276 19306 27288
rect 21361 27285 21373 27319
rect 21407 27316 21419 27319
rect 21910 27316 21916 27328
rect 21407 27288 21916 27316
rect 21407 27285 21419 27288
rect 21361 27279 21419 27285
rect 21910 27276 21916 27288
rect 21968 27276 21974 27328
rect 24412 27316 24440 27347
rect 24578 27344 24584 27356
rect 24636 27344 24642 27396
rect 25222 27316 25228 27328
rect 24412 27288 25228 27316
rect 25222 27276 25228 27288
rect 25280 27276 25286 27328
rect 25608 27316 25636 27424
rect 25961 27421 25973 27424
rect 26007 27421 26019 27455
rect 25961 27415 26019 27421
rect 26053 27455 26111 27461
rect 26053 27421 26065 27455
rect 26099 27421 26111 27455
rect 26053 27415 26111 27421
rect 26142 27412 26148 27464
rect 26200 27452 26206 27464
rect 26344 27461 26372 27560
rect 29564 27560 31156 27588
rect 29454 27520 29460 27532
rect 28552 27492 29460 27520
rect 26329 27455 26387 27461
rect 26200 27424 26245 27452
rect 26200 27412 26206 27424
rect 26329 27421 26341 27455
rect 26375 27421 26387 27455
rect 26329 27415 26387 27421
rect 26789 27455 26847 27461
rect 26789 27421 26801 27455
rect 26835 27452 26847 27455
rect 28552 27452 28580 27492
rect 29454 27480 29460 27492
rect 29512 27480 29518 27532
rect 26835 27424 28580 27452
rect 28629 27455 28687 27461
rect 26835 27421 26847 27424
rect 26789 27415 26847 27421
rect 28629 27421 28641 27455
rect 28675 27421 28687 27455
rect 28629 27415 28687 27421
rect 25685 27387 25743 27393
rect 25685 27353 25697 27387
rect 25731 27384 25743 27387
rect 27034 27387 27092 27393
rect 27034 27384 27046 27387
rect 25731 27356 27046 27384
rect 25731 27353 25743 27356
rect 25685 27347 25743 27353
rect 27034 27353 27046 27356
rect 27080 27353 27092 27387
rect 27034 27347 27092 27353
rect 27706 27344 27712 27396
rect 27764 27384 27770 27396
rect 28442 27384 28448 27396
rect 27764 27356 28448 27384
rect 27764 27344 27770 27356
rect 28442 27344 28448 27356
rect 28500 27384 28506 27396
rect 28644 27384 28672 27415
rect 28500 27356 28672 27384
rect 28500 27344 28506 27356
rect 28718 27344 28724 27396
rect 28776 27384 28782 27396
rect 29564 27393 29592 27560
rect 32214 27548 32220 27600
rect 32272 27588 32278 27600
rect 32493 27591 32551 27597
rect 32493 27588 32505 27591
rect 32272 27560 32505 27588
rect 32272 27548 32278 27560
rect 32493 27557 32505 27560
rect 32539 27557 32551 27591
rect 32493 27551 32551 27557
rect 32766 27548 32772 27600
rect 32824 27588 32830 27600
rect 36004 27588 36032 27628
rect 32824 27560 36032 27588
rect 36924 27588 36952 27628
rect 45554 27588 45560 27600
rect 36924 27560 39896 27588
rect 45515 27560 45560 27588
rect 32824 27548 32830 27560
rect 39666 27520 39672 27532
rect 32508 27492 36124 27520
rect 29638 27412 29644 27464
rect 29696 27452 29702 27464
rect 29825 27455 29883 27461
rect 29825 27452 29837 27455
rect 29696 27424 29837 27452
rect 29696 27412 29702 27424
rect 29825 27421 29837 27424
rect 29871 27421 29883 27455
rect 29825 27415 29883 27421
rect 30190 27412 30196 27464
rect 30248 27452 30254 27464
rect 31113 27455 31171 27461
rect 31113 27452 31125 27455
rect 30248 27424 31125 27452
rect 30248 27412 30254 27424
rect 31113 27421 31125 27424
rect 31159 27421 31171 27455
rect 31113 27415 31171 27421
rect 31380 27455 31438 27461
rect 31380 27421 31392 27455
rect 31426 27452 31438 27455
rect 32122 27452 32128 27464
rect 31426 27424 32128 27452
rect 31426 27421 31438 27424
rect 31380 27415 31438 27421
rect 32122 27412 32128 27424
rect 32180 27412 32186 27464
rect 29549 27387 29607 27393
rect 29549 27384 29561 27387
rect 28776 27356 29561 27384
rect 28776 27344 28782 27356
rect 28166 27316 28172 27328
rect 25608 27288 28172 27316
rect 28166 27276 28172 27288
rect 28224 27276 28230 27328
rect 28828 27325 28856 27356
rect 29549 27353 29561 27356
rect 29595 27353 29607 27387
rect 29549 27347 29607 27353
rect 29733 27387 29791 27393
rect 29733 27353 29745 27387
rect 29779 27384 29791 27387
rect 31938 27384 31944 27396
rect 29779 27356 31944 27384
rect 29779 27353 29791 27356
rect 29733 27347 29791 27353
rect 31938 27344 31944 27356
rect 31996 27344 32002 27396
rect 28813 27319 28871 27325
rect 28813 27285 28825 27319
rect 28859 27285 28871 27319
rect 28813 27279 28871 27285
rect 28902 27276 28908 27328
rect 28960 27316 28966 27328
rect 32508 27316 32536 27492
rect 32674 27412 32680 27464
rect 32732 27452 32738 27464
rect 33045 27455 33103 27461
rect 33045 27452 33057 27455
rect 32732 27424 33057 27452
rect 32732 27412 32738 27424
rect 33045 27421 33057 27424
rect 33091 27421 33103 27455
rect 33045 27415 33103 27421
rect 35802 27412 35808 27464
rect 35860 27452 35866 27464
rect 35989 27455 36047 27461
rect 35989 27452 36001 27455
rect 35860 27424 36001 27452
rect 35860 27412 35866 27424
rect 35989 27421 36001 27424
rect 36035 27421 36047 27455
rect 36096 27452 36124 27492
rect 37016 27492 39672 27520
rect 37016 27452 37044 27492
rect 39666 27480 39672 27492
rect 39724 27480 39730 27532
rect 39868 27529 39896 27560
rect 45554 27548 45560 27560
rect 45612 27548 45618 27600
rect 39853 27523 39911 27529
rect 39853 27489 39865 27523
rect 39899 27489 39911 27523
rect 46290 27520 46296 27532
rect 46251 27492 46296 27520
rect 39853 27483 39911 27489
rect 46290 27480 46296 27492
rect 46348 27480 46354 27532
rect 46477 27523 46535 27529
rect 46477 27489 46489 27523
rect 46523 27520 46535 27523
rect 46566 27520 46572 27532
rect 46523 27492 46572 27520
rect 46523 27489 46535 27492
rect 46477 27483 46535 27489
rect 46566 27480 46572 27492
rect 46624 27480 46630 27532
rect 48133 27523 48191 27529
rect 48133 27489 48145 27523
rect 48179 27520 48191 27523
rect 48222 27520 48228 27532
rect 48179 27492 48228 27520
rect 48179 27489 48191 27492
rect 48133 27483 48191 27489
rect 48222 27480 48228 27492
rect 48280 27480 48286 27532
rect 36096 27424 37044 27452
rect 35989 27415 36047 27421
rect 37090 27412 37096 27464
rect 37148 27452 37154 27464
rect 37148 27424 37412 27452
rect 37148 27412 37154 27424
rect 32582 27344 32588 27396
rect 32640 27384 32646 27396
rect 33873 27387 33931 27393
rect 33873 27384 33885 27387
rect 32640 27356 33885 27384
rect 32640 27344 32646 27356
rect 33873 27353 33885 27356
rect 33919 27353 33931 27387
rect 34054 27384 34060 27396
rect 34015 27356 34060 27384
rect 33873 27347 33931 27353
rect 34054 27344 34060 27356
rect 34112 27344 34118 27396
rect 35158 27384 35164 27396
rect 35119 27356 35164 27384
rect 35158 27344 35164 27356
rect 35216 27344 35222 27396
rect 35345 27387 35403 27393
rect 35345 27353 35357 27387
rect 35391 27384 35403 27387
rect 35618 27384 35624 27396
rect 35391 27356 35624 27384
rect 35391 27353 35403 27356
rect 35345 27347 35403 27353
rect 35618 27344 35624 27356
rect 35676 27344 35682 27396
rect 36256 27387 36314 27393
rect 36256 27353 36268 27387
rect 36302 27384 36314 27387
rect 37274 27384 37280 27396
rect 36302 27356 37280 27384
rect 36302 27353 36314 27356
rect 36256 27347 36314 27353
rect 37274 27344 37280 27356
rect 37332 27344 37338 27396
rect 35526 27316 35532 27328
rect 28960 27288 32536 27316
rect 35487 27288 35532 27316
rect 28960 27276 28966 27288
rect 35526 27276 35532 27288
rect 35584 27276 35590 27328
rect 37384 27325 37412 27424
rect 38470 27412 38476 27464
rect 38528 27452 38534 27464
rect 39117 27455 39175 27461
rect 39117 27452 39129 27455
rect 38528 27424 39129 27452
rect 38528 27412 38534 27424
rect 39117 27421 39129 27424
rect 39163 27421 39175 27455
rect 45462 27452 45468 27464
rect 45423 27424 45468 27452
rect 39117 27415 39175 27421
rect 45462 27412 45468 27424
rect 45520 27412 45526 27464
rect 39209 27387 39267 27393
rect 39209 27353 39221 27387
rect 39255 27384 39267 27387
rect 40037 27387 40095 27393
rect 40037 27384 40049 27387
rect 39255 27356 40049 27384
rect 39255 27353 39267 27356
rect 39209 27347 39267 27353
rect 40037 27353 40049 27356
rect 40083 27353 40095 27387
rect 41690 27384 41696 27396
rect 41651 27356 41696 27384
rect 40037 27347 40095 27353
rect 41690 27344 41696 27356
rect 41748 27344 41754 27396
rect 37369 27319 37427 27325
rect 37369 27285 37381 27319
rect 37415 27285 37427 27319
rect 37369 27279 37427 27285
rect 37458 27276 37464 27328
rect 37516 27316 37522 27328
rect 48038 27316 48044 27328
rect 37516 27288 48044 27316
rect 37516 27276 37522 27288
rect 48038 27276 48044 27288
rect 48096 27276 48102 27328
rect 1104 27226 48852 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 48852 27226
rect 1104 27152 48852 27174
rect 2130 27072 2136 27124
rect 2188 27112 2194 27124
rect 26142 27112 26148 27124
rect 2188 27084 26004 27112
rect 26103 27084 26148 27112
rect 2188 27072 2194 27084
rect 1946 27044 1952 27056
rect 1907 27016 1952 27044
rect 1946 27004 1952 27016
rect 2004 27004 2010 27056
rect 11977 27047 12035 27053
rect 11977 27013 11989 27047
rect 12023 27044 12035 27047
rect 12710 27044 12716 27056
rect 12023 27016 12716 27044
rect 12023 27013 12035 27016
rect 11977 27007 12035 27013
rect 12710 27004 12716 27016
rect 12768 27004 12774 27056
rect 16574 27004 16580 27056
rect 16632 27044 16638 27056
rect 18417 27047 18475 27053
rect 16632 27016 16804 27044
rect 16632 27004 16638 27016
rect 1762 26976 1768 26988
rect 1723 26948 1768 26976
rect 1762 26936 1768 26948
rect 1820 26936 1826 26988
rect 15746 26976 15752 26988
rect 15659 26948 15752 26976
rect 15746 26936 15752 26948
rect 15804 26976 15810 26988
rect 16114 26976 16120 26988
rect 15804 26948 16120 26976
rect 15804 26936 15810 26948
rect 16114 26936 16120 26948
rect 16172 26936 16178 26988
rect 16669 26979 16727 26985
rect 16669 26945 16681 26979
rect 16715 26945 16727 26979
rect 16776 26976 16804 27016
rect 18417 27013 18429 27047
rect 18463 27044 18475 27047
rect 19334 27044 19340 27056
rect 18463 27016 19340 27044
rect 18463 27013 18475 27016
rect 18417 27007 18475 27013
rect 19334 27004 19340 27016
rect 19392 27004 19398 27056
rect 21082 27044 21088 27056
rect 21043 27016 21088 27044
rect 21082 27004 21088 27016
rect 21140 27004 21146 27056
rect 21266 27044 21272 27056
rect 21227 27016 21272 27044
rect 21266 27004 21272 27016
rect 21324 27004 21330 27056
rect 25038 27044 25044 27056
rect 21836 27016 22508 27044
rect 18230 26976 18236 26988
rect 16776 26948 17632 26976
rect 18191 26948 18236 26976
rect 16669 26939 16727 26945
rect 2774 26908 2780 26920
rect 2735 26880 2780 26908
rect 2774 26868 2780 26880
rect 2832 26868 2838 26920
rect 11790 26908 11796 26920
rect 11751 26880 11796 26908
rect 11790 26868 11796 26880
rect 11848 26868 11854 26920
rect 12253 26911 12311 26917
rect 12253 26877 12265 26911
rect 12299 26877 12311 26911
rect 12253 26871 12311 26877
rect 11054 26800 11060 26852
rect 11112 26840 11118 26852
rect 12268 26840 12296 26871
rect 16574 26868 16580 26920
rect 16632 26908 16638 26920
rect 16684 26908 16712 26939
rect 17034 26908 17040 26920
rect 16632 26880 16712 26908
rect 16995 26880 17040 26908
rect 16632 26868 16638 26880
rect 17034 26868 17040 26880
rect 17092 26868 17098 26920
rect 17604 26908 17632 26948
rect 18230 26936 18236 26948
rect 18288 26936 18294 26988
rect 19886 26936 19892 26988
rect 19944 26976 19950 26988
rect 20346 26976 20352 26988
rect 19944 26948 20352 26976
rect 19944 26936 19950 26948
rect 20346 26936 20352 26948
rect 20404 26936 20410 26988
rect 21836 26985 21864 27016
rect 22480 26988 22508 27016
rect 23860 27016 25044 27044
rect 20901 26979 20959 26985
rect 20901 26945 20913 26979
rect 20947 26945 20959 26979
rect 20901 26939 20959 26945
rect 21821 26979 21879 26985
rect 21821 26945 21833 26979
rect 21867 26945 21879 26979
rect 21821 26939 21879 26945
rect 18693 26911 18751 26917
rect 18693 26908 18705 26911
rect 17604 26880 18705 26908
rect 18693 26877 18705 26880
rect 18739 26877 18751 26911
rect 18693 26871 18751 26877
rect 11112 26812 12296 26840
rect 11112 26800 11118 26812
rect 15838 26772 15844 26784
rect 15799 26744 15844 26772
rect 15838 26732 15844 26744
rect 15896 26732 15902 26784
rect 20916 26772 20944 26939
rect 21910 26936 21916 26988
rect 21968 26976 21974 26988
rect 22077 26979 22135 26985
rect 22077 26976 22089 26979
rect 21968 26948 22089 26976
rect 21968 26936 21974 26948
rect 22077 26945 22089 26948
rect 22123 26945 22135 26979
rect 22077 26939 22135 26945
rect 22462 26936 22468 26988
rect 22520 26976 22526 26988
rect 23860 26985 23888 27016
rect 25038 27004 25044 27016
rect 25096 27004 25102 27056
rect 25976 27044 26004 27084
rect 26142 27072 26148 27084
rect 26200 27072 26206 27124
rect 28166 27072 28172 27124
rect 28224 27112 28230 27124
rect 33778 27112 33784 27124
rect 28224 27084 33784 27112
rect 28224 27072 28230 27084
rect 33778 27072 33784 27084
rect 33836 27072 33842 27124
rect 35618 27072 35624 27124
rect 35676 27112 35682 27124
rect 36998 27112 37004 27124
rect 35676 27084 37004 27112
rect 35676 27072 35682 27084
rect 36998 27072 37004 27084
rect 37056 27072 37062 27124
rect 37274 27112 37280 27124
rect 37235 27084 37280 27112
rect 37274 27072 37280 27084
rect 37332 27072 37338 27124
rect 37458 27072 37464 27124
rect 37516 27072 37522 27124
rect 45830 27112 45836 27124
rect 37844 27084 45836 27112
rect 37844 27073 37872 27084
rect 34514 27044 34520 27056
rect 25976 27016 30052 27044
rect 23845 26979 23903 26985
rect 23845 26976 23857 26979
rect 22520 26948 23857 26976
rect 22520 26936 22526 26948
rect 23845 26945 23857 26948
rect 23891 26945 23903 26979
rect 23845 26939 23903 26945
rect 23934 26936 23940 26988
rect 23992 26976 23998 26988
rect 24101 26979 24159 26985
rect 24101 26976 24113 26979
rect 23992 26948 24113 26976
rect 23992 26936 23998 26948
rect 24101 26945 24113 26948
rect 24147 26945 24159 26979
rect 24101 26939 24159 26945
rect 24670 26936 24676 26988
rect 24728 26976 24734 26988
rect 25869 26979 25927 26985
rect 25869 26976 25881 26979
rect 24728 26948 25881 26976
rect 24728 26936 24734 26948
rect 25869 26945 25881 26948
rect 25915 26945 25927 26979
rect 25869 26939 25927 26945
rect 25958 26936 25964 26988
rect 26016 26976 26022 26988
rect 27154 26976 27160 26988
rect 26016 26948 26061 26976
rect 27115 26948 27160 26976
rect 26016 26936 26022 26948
rect 27154 26936 27160 26948
rect 27212 26936 27218 26988
rect 28074 26976 28080 26988
rect 28035 26948 28080 26976
rect 28074 26936 28080 26948
rect 28132 26936 28138 26988
rect 28442 26976 28448 26988
rect 28403 26948 28448 26976
rect 28442 26936 28448 26948
rect 28500 26976 28506 26988
rect 29362 26976 29368 26988
rect 28500 26948 29368 26976
rect 28500 26936 28506 26948
rect 29362 26936 29368 26948
rect 29420 26936 29426 26988
rect 30024 26985 30052 27016
rect 33244 27016 34520 27044
rect 30009 26979 30067 26985
rect 30009 26945 30021 26979
rect 30055 26945 30067 26979
rect 30009 26939 30067 26945
rect 30101 26979 30159 26985
rect 30101 26945 30113 26979
rect 30147 26945 30159 26979
rect 30101 26939 30159 26945
rect 30193 26979 30251 26985
rect 30193 26945 30205 26979
rect 30239 26976 30251 26979
rect 30282 26976 30288 26988
rect 30239 26948 30288 26976
rect 30239 26945 30251 26948
rect 30193 26939 30251 26945
rect 24854 26868 24860 26920
rect 24912 26908 24918 26920
rect 26145 26911 26203 26917
rect 26145 26908 26157 26911
rect 24912 26880 26157 26908
rect 24912 26868 24918 26880
rect 26145 26877 26157 26880
rect 26191 26877 26203 26911
rect 26145 26871 26203 26877
rect 26234 26868 26240 26920
rect 26292 26908 26298 26920
rect 28902 26908 28908 26920
rect 26292 26880 28908 26908
rect 26292 26868 26298 26880
rect 28902 26868 28908 26880
rect 28960 26868 28966 26920
rect 30116 26908 30144 26939
rect 30282 26936 30288 26948
rect 30340 26936 30346 26988
rect 30377 26979 30435 26985
rect 30377 26945 30389 26979
rect 30423 26976 30435 26979
rect 30466 26976 30472 26988
rect 30423 26948 30472 26976
rect 30423 26945 30435 26948
rect 30377 26939 30435 26945
rect 30466 26936 30472 26948
rect 30524 26936 30530 26988
rect 33244 26985 33272 27016
rect 34514 27004 34520 27016
rect 34572 27044 34578 27056
rect 35802 27044 35808 27056
rect 34572 27016 35808 27044
rect 34572 27004 34578 27016
rect 35802 27004 35808 27016
rect 35860 27004 35866 27056
rect 36078 27004 36084 27056
rect 36136 27044 36142 27056
rect 36136 27016 36492 27044
rect 36136 27004 36142 27016
rect 33229 26979 33287 26985
rect 33229 26945 33241 26979
rect 33275 26945 33287 26979
rect 33229 26939 33287 26945
rect 33496 26979 33554 26985
rect 33496 26945 33508 26979
rect 33542 26976 33554 26979
rect 34698 26976 34704 26988
rect 33542 26948 34704 26976
rect 33542 26945 33554 26948
rect 33496 26939 33554 26945
rect 34698 26936 34704 26948
rect 34756 26936 34762 26988
rect 35253 26979 35311 26985
rect 35253 26945 35265 26979
rect 35299 26945 35311 26979
rect 35253 26939 35311 26945
rect 35437 26979 35495 26985
rect 35437 26945 35449 26979
rect 35483 26976 35495 26979
rect 35526 26976 35532 26988
rect 35483 26948 35532 26976
rect 35483 26945 35495 26948
rect 35437 26939 35495 26945
rect 30742 26908 30748 26920
rect 30116 26880 30748 26908
rect 30742 26868 30748 26880
rect 30800 26868 30806 26920
rect 34514 26868 34520 26920
rect 34572 26908 34578 26920
rect 35158 26908 35164 26920
rect 34572 26880 35164 26908
rect 34572 26868 34578 26880
rect 35158 26868 35164 26880
rect 35216 26908 35222 26920
rect 35268 26908 35296 26939
rect 35526 26936 35532 26948
rect 35584 26936 35590 26988
rect 36262 26936 36268 26988
rect 36320 26985 36326 26988
rect 36464 26985 36492 27016
rect 36814 27004 36820 27056
rect 36872 27044 36878 27056
rect 37476 27044 37504 27072
rect 36872 27016 37504 27044
rect 37568 27045 37872 27073
rect 45830 27072 45836 27084
rect 45888 27072 45894 27124
rect 46474 27072 46480 27124
rect 46532 27112 46538 27124
rect 46569 27115 46627 27121
rect 46569 27112 46581 27115
rect 46532 27084 46581 27112
rect 46532 27072 46538 27084
rect 46569 27081 46581 27084
rect 46615 27081 46627 27115
rect 46569 27075 46627 27081
rect 36872 27004 36878 27016
rect 37568 26985 37596 27045
rect 37642 26985 37700 26991
rect 36320 26979 36369 26985
rect 36320 26945 36323 26979
rect 36357 26945 36369 26979
rect 36320 26939 36369 26945
rect 36449 26979 36507 26985
rect 36449 26945 36461 26979
rect 36495 26945 36507 26979
rect 36449 26939 36507 26945
rect 36562 26979 36620 26985
rect 36562 26945 36574 26979
rect 36608 26945 36620 26979
rect 36562 26939 36620 26945
rect 36725 26979 36783 26985
rect 36725 26945 36737 26979
rect 36771 26945 36783 26979
rect 36725 26939 36783 26945
rect 37553 26979 37611 26985
rect 37553 26945 37565 26979
rect 37599 26945 37611 26979
rect 37642 26951 37654 26985
rect 37688 26951 37700 26985
rect 37642 26945 37700 26951
rect 37737 26979 37795 26985
rect 37737 26945 37749 26979
rect 37783 26945 37795 26979
rect 37918 26976 37924 26988
rect 37879 26948 37924 26976
rect 37553 26939 37611 26945
rect 36320 26936 36326 26939
rect 35216 26880 35296 26908
rect 35621 26911 35679 26917
rect 35216 26868 35222 26880
rect 35621 26877 35633 26911
rect 35667 26908 35679 26911
rect 36577 26908 36605 26939
rect 36740 26908 36768 26939
rect 36814 26908 36820 26920
rect 35667 26880 36605 26908
rect 36727 26880 36820 26908
rect 35667 26877 35679 26880
rect 35621 26871 35679 26877
rect 25222 26840 25228 26852
rect 25135 26812 25228 26840
rect 25222 26800 25228 26812
rect 25280 26840 25286 26852
rect 33226 26840 33232 26852
rect 25280 26812 33232 26840
rect 25280 26800 25286 26812
rect 33226 26800 33232 26812
rect 33284 26800 33290 26852
rect 35342 26840 35348 26852
rect 34348 26812 35348 26840
rect 23201 26775 23259 26781
rect 23201 26772 23213 26775
rect 20916 26744 23213 26772
rect 23201 26741 23213 26744
rect 23247 26772 23259 26775
rect 26234 26772 26240 26784
rect 23247 26744 26240 26772
rect 23247 26741 23259 26744
rect 23201 26735 23259 26741
rect 26234 26732 26240 26744
rect 26292 26732 26298 26784
rect 26694 26732 26700 26784
rect 26752 26772 26758 26784
rect 26973 26775 27031 26781
rect 26973 26772 26985 26775
rect 26752 26744 26985 26772
rect 26752 26732 26758 26744
rect 26973 26741 26985 26744
rect 27019 26741 27031 26775
rect 26973 26735 27031 26741
rect 28074 26732 28080 26784
rect 28132 26772 28138 26784
rect 28718 26772 28724 26784
rect 28132 26744 28724 26772
rect 28132 26732 28138 26744
rect 28718 26732 28724 26744
rect 28776 26732 28782 26784
rect 29730 26772 29736 26784
rect 29691 26744 29736 26772
rect 29730 26732 29736 26744
rect 29788 26732 29794 26784
rect 30466 26732 30472 26784
rect 30524 26772 30530 26784
rect 34348 26772 34376 26812
rect 35342 26800 35348 26812
rect 35400 26840 35406 26852
rect 36740 26840 36768 26880
rect 36814 26868 36820 26880
rect 36872 26908 36878 26920
rect 36998 26908 37004 26920
rect 36872 26880 37004 26908
rect 36872 26868 36878 26880
rect 36998 26868 37004 26880
rect 37056 26868 37062 26920
rect 37458 26868 37464 26920
rect 37516 26908 37522 26920
rect 37657 26908 37685 26945
rect 37737 26939 37795 26945
rect 37516 26880 37685 26908
rect 37752 26908 37780 26939
rect 37918 26936 37924 26948
rect 37976 26936 37982 26988
rect 38470 26936 38476 26988
rect 38528 26976 38534 26988
rect 38565 26979 38623 26985
rect 38565 26976 38577 26979
rect 38528 26948 38577 26976
rect 38528 26936 38534 26948
rect 38565 26945 38577 26948
rect 38611 26945 38623 26979
rect 38565 26939 38623 26945
rect 46382 26936 46388 26988
rect 46440 26976 46446 26988
rect 46477 26979 46535 26985
rect 46477 26976 46489 26979
rect 46440 26948 46489 26976
rect 46440 26936 46446 26948
rect 46477 26945 46489 26948
rect 46523 26945 46535 26979
rect 46477 26939 46535 26945
rect 38102 26908 38108 26920
rect 37752 26880 38108 26908
rect 37516 26868 37522 26880
rect 38102 26868 38108 26880
rect 38160 26868 38166 26920
rect 39209 26911 39267 26917
rect 39209 26877 39221 26911
rect 39255 26877 39267 26911
rect 39390 26908 39396 26920
rect 39351 26880 39396 26908
rect 39209 26871 39267 26877
rect 35400 26812 36768 26840
rect 35400 26800 35406 26812
rect 37734 26800 37740 26852
rect 37792 26840 37798 26852
rect 39224 26840 39252 26871
rect 39390 26868 39396 26880
rect 39448 26868 39454 26920
rect 41049 26911 41107 26917
rect 41049 26877 41061 26911
rect 41095 26908 41107 26911
rect 48498 26908 48504 26920
rect 41095 26880 48504 26908
rect 41095 26877 41107 26880
rect 41049 26871 41107 26877
rect 48498 26868 48504 26880
rect 48556 26868 48562 26920
rect 37792 26812 39252 26840
rect 37792 26800 37798 26812
rect 30524 26744 34376 26772
rect 30524 26732 30530 26744
rect 34422 26732 34428 26784
rect 34480 26772 34486 26784
rect 34609 26775 34667 26781
rect 34609 26772 34621 26775
rect 34480 26744 34621 26772
rect 34480 26732 34486 26744
rect 34609 26741 34621 26744
rect 34655 26741 34667 26775
rect 34609 26735 34667 26741
rect 36081 26775 36139 26781
rect 36081 26741 36093 26775
rect 36127 26772 36139 26775
rect 36446 26772 36452 26784
rect 36127 26744 36452 26772
rect 36127 26741 36139 26744
rect 36081 26735 36139 26741
rect 36446 26732 36452 26744
rect 36504 26732 36510 26784
rect 38657 26775 38715 26781
rect 38657 26741 38669 26775
rect 38703 26772 38715 26775
rect 40034 26772 40040 26784
rect 38703 26744 40040 26772
rect 38703 26741 38715 26744
rect 38657 26735 38715 26741
rect 40034 26732 40040 26744
rect 40092 26732 40098 26784
rect 1104 26682 48852 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 48852 26682
rect 1104 26608 48852 26630
rect 2958 26528 2964 26580
rect 3016 26568 3022 26580
rect 11790 26568 11796 26580
rect 3016 26540 11796 26568
rect 3016 26528 3022 26540
rect 11790 26528 11796 26540
rect 11848 26528 11854 26580
rect 19242 26568 19248 26580
rect 19203 26540 19248 26568
rect 19242 26528 19248 26540
rect 19300 26528 19306 26580
rect 19426 26528 19432 26580
rect 19484 26568 19490 26580
rect 20717 26571 20775 26577
rect 20717 26568 20729 26571
rect 19484 26540 20729 26568
rect 19484 26528 19490 26540
rect 20717 26537 20729 26540
rect 20763 26537 20775 26571
rect 22830 26568 22836 26580
rect 20717 26531 20775 26537
rect 22066 26540 22836 26568
rect 3050 26500 3056 26512
rect 1412 26472 3056 26500
rect 1412 26441 1440 26472
rect 3050 26460 3056 26472
rect 3108 26460 3114 26512
rect 17310 26500 17316 26512
rect 15672 26472 17316 26500
rect 1397 26435 1455 26441
rect 1397 26401 1409 26435
rect 1443 26401 1455 26435
rect 2774 26432 2780 26444
rect 2735 26404 2780 26432
rect 1397 26395 1455 26401
rect 2774 26392 2780 26404
rect 2832 26392 2838 26444
rect 15672 26441 15700 26472
rect 17310 26460 17316 26472
rect 17368 26460 17374 26512
rect 18601 26503 18659 26509
rect 18601 26469 18613 26503
rect 18647 26500 18659 26503
rect 20070 26500 20076 26512
rect 18647 26472 20076 26500
rect 18647 26469 18659 26472
rect 18601 26463 18659 26469
rect 20070 26460 20076 26472
rect 20128 26460 20134 26512
rect 22066 26500 22094 26540
rect 22830 26528 22836 26540
rect 22888 26528 22894 26580
rect 23198 26528 23204 26580
rect 23256 26568 23262 26580
rect 24854 26568 24860 26580
rect 23256 26540 24860 26568
rect 23256 26528 23262 26540
rect 24854 26528 24860 26540
rect 24912 26528 24918 26580
rect 24949 26571 25007 26577
rect 24949 26537 24961 26571
rect 24995 26568 25007 26571
rect 25038 26568 25044 26580
rect 24995 26540 25044 26568
rect 24995 26537 25007 26540
rect 24949 26531 25007 26537
rect 25038 26528 25044 26540
rect 25096 26528 25102 26580
rect 26050 26568 26056 26580
rect 26011 26540 26056 26568
rect 26050 26528 26056 26540
rect 26108 26528 26114 26580
rect 27706 26568 27712 26580
rect 26252 26540 27712 26568
rect 20548 26472 22094 26500
rect 15657 26435 15715 26441
rect 15657 26401 15669 26435
rect 15703 26401 15715 26435
rect 15838 26432 15844 26444
rect 15799 26404 15844 26432
rect 15657 26395 15715 26401
rect 15838 26392 15844 26404
rect 15896 26392 15902 26444
rect 17034 26392 17040 26444
rect 17092 26432 17098 26444
rect 20162 26432 20168 26444
rect 17092 26404 19380 26432
rect 17092 26392 17098 26404
rect 18230 26364 18236 26376
rect 18191 26336 18236 26364
rect 18230 26324 18236 26336
rect 18288 26324 18294 26376
rect 18322 26324 18328 26376
rect 18380 26364 18386 26376
rect 18417 26367 18475 26373
rect 18417 26364 18429 26367
rect 18380 26336 18429 26364
rect 18380 26324 18386 26336
rect 18417 26333 18429 26336
rect 18463 26333 18475 26367
rect 18417 26327 18475 26333
rect 18506 26324 18512 26376
rect 18564 26364 18570 26376
rect 19242 26364 19248 26376
rect 18564 26336 19248 26364
rect 18564 26324 18570 26336
rect 19242 26324 19248 26336
rect 19300 26324 19306 26376
rect 1581 26299 1639 26305
rect 1581 26265 1593 26299
rect 1627 26296 1639 26299
rect 2774 26296 2780 26308
rect 1627 26268 2780 26296
rect 1627 26265 1639 26268
rect 1581 26259 1639 26265
rect 2774 26256 2780 26268
rect 2832 26256 2838 26308
rect 17497 26299 17555 26305
rect 17497 26265 17509 26299
rect 17543 26296 17555 26299
rect 17770 26296 17776 26308
rect 17543 26268 17776 26296
rect 17543 26265 17555 26268
rect 17497 26259 17555 26265
rect 17770 26256 17776 26268
rect 17828 26256 17834 26308
rect 19352 26296 19380 26404
rect 19628 26404 20168 26432
rect 19518 26364 19524 26376
rect 19479 26336 19524 26364
rect 19518 26324 19524 26336
rect 19576 26324 19582 26376
rect 19628 26373 19656 26404
rect 20162 26392 20168 26404
rect 20220 26392 20226 26444
rect 19613 26367 19671 26373
rect 19613 26333 19625 26367
rect 19659 26333 19671 26367
rect 19613 26327 19671 26333
rect 19702 26324 19708 26376
rect 19760 26364 19766 26376
rect 19889 26367 19947 26373
rect 19760 26336 19805 26364
rect 19760 26324 19766 26336
rect 19889 26333 19901 26367
rect 19935 26364 19947 26367
rect 19978 26364 19984 26376
rect 19935 26336 19984 26364
rect 19935 26333 19947 26336
rect 19889 26327 19947 26333
rect 19978 26324 19984 26336
rect 20036 26324 20042 26376
rect 20548 26296 20576 26472
rect 23566 26460 23572 26512
rect 23624 26500 23630 26512
rect 23845 26503 23903 26509
rect 23845 26500 23857 26503
rect 23624 26472 23857 26500
rect 23624 26460 23630 26472
rect 23845 26469 23857 26472
rect 23891 26500 23903 26503
rect 26142 26500 26148 26512
rect 23891 26472 26148 26500
rect 23891 26469 23903 26472
rect 23845 26463 23903 26469
rect 26142 26460 26148 26472
rect 26200 26460 26206 26512
rect 22278 26432 22284 26444
rect 22066 26404 22284 26432
rect 20625 26367 20683 26373
rect 20625 26333 20637 26367
rect 20671 26364 20683 26367
rect 22066 26364 22094 26404
rect 22278 26392 22284 26404
rect 22336 26432 22342 26444
rect 22336 26404 22600 26432
rect 22336 26392 22342 26404
rect 22462 26364 22468 26376
rect 20671 26336 22094 26364
rect 22423 26336 22468 26364
rect 20671 26333 20683 26336
rect 20625 26327 20683 26333
rect 22462 26324 22468 26336
rect 22520 26324 22526 26376
rect 22572 26364 22600 26404
rect 24118 26392 24124 26444
rect 24176 26432 24182 26444
rect 26252 26432 26280 26540
rect 27706 26528 27712 26540
rect 27764 26528 27770 26580
rect 27798 26528 27804 26580
rect 27856 26568 27862 26580
rect 28626 26568 28632 26580
rect 27856 26540 28632 26568
rect 27856 26528 27862 26540
rect 28626 26528 28632 26540
rect 28684 26528 28690 26580
rect 29454 26528 29460 26580
rect 29512 26568 29518 26580
rect 32309 26571 32367 26577
rect 32309 26568 32321 26571
rect 29512 26540 32321 26568
rect 29512 26528 29518 26540
rect 26418 26460 26424 26512
rect 26476 26500 26482 26512
rect 30098 26500 30104 26512
rect 26476 26472 30104 26500
rect 26476 26460 26482 26472
rect 30098 26460 30104 26472
rect 30156 26460 30162 26512
rect 30208 26444 30236 26540
rect 32309 26537 32321 26540
rect 32355 26568 32367 26571
rect 32674 26568 32680 26580
rect 32355 26540 32680 26568
rect 32355 26537 32367 26540
rect 32309 26531 32367 26537
rect 32674 26528 32680 26540
rect 32732 26528 32738 26580
rect 35526 26528 35532 26580
rect 35584 26568 35590 26580
rect 37090 26568 37096 26580
rect 35584 26540 37096 26568
rect 35584 26528 35590 26540
rect 37090 26528 37096 26540
rect 37148 26568 37154 26580
rect 37737 26571 37795 26577
rect 37737 26568 37749 26571
rect 37148 26540 37749 26568
rect 37148 26528 37154 26540
rect 37737 26537 37749 26540
rect 37783 26537 37795 26571
rect 37737 26531 37795 26537
rect 39209 26571 39267 26577
rect 39209 26537 39221 26571
rect 39255 26568 39267 26571
rect 39390 26568 39396 26580
rect 39255 26540 39396 26568
rect 39255 26537 39267 26540
rect 39209 26531 39267 26537
rect 39390 26528 39396 26540
rect 39448 26528 39454 26580
rect 47486 26568 47492 26580
rect 41432 26540 47492 26568
rect 35066 26460 35072 26512
rect 35124 26460 35130 26512
rect 35342 26500 35348 26512
rect 35268 26472 35348 26500
rect 30006 26432 30012 26444
rect 24176 26404 26280 26432
rect 26436 26404 30012 26432
rect 24176 26392 24182 26404
rect 24857 26367 24915 26373
rect 24857 26364 24869 26367
rect 22572 26336 24869 26364
rect 24857 26333 24869 26336
rect 24903 26333 24915 26367
rect 26436 26364 26464 26404
rect 30006 26392 30012 26404
rect 30064 26392 30070 26444
rect 30190 26432 30196 26444
rect 30151 26404 30196 26432
rect 30190 26392 30196 26404
rect 30248 26392 30254 26444
rect 32766 26432 32772 26444
rect 31726 26404 32772 26432
rect 24857 26327 24915 26333
rect 24955 26336 26464 26364
rect 19352 26268 20576 26296
rect 21910 26256 21916 26308
rect 21968 26296 21974 26308
rect 22480 26296 22508 26324
rect 22738 26305 22744 26308
rect 22732 26296 22744 26305
rect 21968 26268 22508 26296
rect 22699 26268 22744 26296
rect 21968 26256 21974 26268
rect 22732 26259 22744 26268
rect 22738 26256 22744 26259
rect 22796 26256 22802 26308
rect 22830 26256 22836 26308
rect 22888 26296 22894 26308
rect 24955 26296 24983 26336
rect 29730 26324 29736 26376
rect 29788 26364 29794 26376
rect 30449 26367 30507 26373
rect 30449 26364 30461 26367
rect 29788 26336 30461 26364
rect 29788 26324 29794 26336
rect 30449 26333 30461 26336
rect 30495 26333 30507 26367
rect 31726 26364 31754 26404
rect 32766 26392 32772 26404
rect 32824 26392 32830 26444
rect 32950 26392 32956 26444
rect 33008 26432 33014 26444
rect 34514 26432 34520 26444
rect 33008 26404 34520 26432
rect 33008 26392 33014 26404
rect 30449 26327 30507 26333
rect 30576 26336 31754 26364
rect 33612 26364 33640 26404
rect 34514 26392 34520 26404
rect 34572 26392 34578 26444
rect 34698 26432 34704 26444
rect 34659 26404 34704 26432
rect 34698 26392 34704 26404
rect 34756 26392 34762 26444
rect 33689 26367 33747 26373
rect 33689 26364 33701 26367
rect 33612 26336 33701 26364
rect 22888 26268 24983 26296
rect 22888 26256 22894 26268
rect 25130 26256 25136 26308
rect 25188 26296 25194 26308
rect 25961 26299 26019 26305
rect 25961 26296 25973 26299
rect 25188 26268 25973 26296
rect 25188 26256 25194 26268
rect 25961 26265 25973 26268
rect 26007 26296 26019 26299
rect 26142 26296 26148 26308
rect 26007 26268 26148 26296
rect 26007 26265 26019 26268
rect 25961 26259 26019 26265
rect 26142 26256 26148 26268
rect 26200 26256 26206 26308
rect 26234 26256 26240 26308
rect 26292 26296 26298 26308
rect 30576 26296 30604 26336
rect 33689 26333 33701 26336
rect 33735 26333 33747 26367
rect 33689 26327 33747 26333
rect 33870 26324 33876 26376
rect 33928 26364 33934 26376
rect 35081 26373 35109 26460
rect 35268 26432 35296 26472
rect 35342 26460 35348 26472
rect 35400 26460 35406 26512
rect 35268 26404 35388 26432
rect 34957 26367 35015 26373
rect 33928 26336 33973 26364
rect 33928 26324 33934 26336
rect 34957 26333 34969 26367
rect 35003 26364 35015 26367
rect 35066 26367 35124 26373
rect 35003 26333 35020 26364
rect 34957 26327 35020 26333
rect 35066 26333 35078 26367
rect 35112 26333 35124 26367
rect 35066 26327 35124 26333
rect 26292 26268 30604 26296
rect 32217 26299 32275 26305
rect 26292 26256 26298 26268
rect 32217 26265 32229 26299
rect 32263 26296 32275 26299
rect 33778 26296 33784 26308
rect 32263 26268 33784 26296
rect 32263 26265 32275 26268
rect 32217 26259 32275 26265
rect 33778 26256 33784 26268
rect 33836 26256 33842 26308
rect 34992 26296 35020 26327
rect 35158 26324 35164 26376
rect 35216 26364 35222 26376
rect 35360 26373 35388 26404
rect 39666 26392 39672 26444
rect 39724 26432 39730 26444
rect 39853 26435 39911 26441
rect 39853 26432 39865 26435
rect 39724 26404 39865 26432
rect 39724 26392 39730 26404
rect 39853 26401 39865 26404
rect 39899 26401 39911 26435
rect 40034 26432 40040 26444
rect 39995 26404 40040 26432
rect 39853 26395 39911 26401
rect 40034 26392 40040 26404
rect 40092 26392 40098 26444
rect 35339 26367 35397 26373
rect 35216 26336 35258 26364
rect 35216 26324 35222 26336
rect 35339 26333 35351 26367
rect 35385 26333 35397 26367
rect 35339 26327 35397 26333
rect 35802 26324 35808 26376
rect 35860 26364 35866 26376
rect 36262 26364 36268 26376
rect 35860 26336 36268 26364
rect 35860 26324 35866 26336
rect 36262 26324 36268 26336
rect 36320 26364 36326 26376
rect 36357 26367 36415 26373
rect 36357 26364 36369 26367
rect 36320 26336 36369 26364
rect 36320 26324 36326 26336
rect 36357 26333 36369 26336
rect 36403 26333 36415 26367
rect 36357 26327 36415 26333
rect 36446 26324 36452 26376
rect 36504 26364 36510 26376
rect 36613 26367 36671 26373
rect 36613 26364 36625 26367
rect 36504 26336 36625 26364
rect 36504 26324 36510 26336
rect 36613 26333 36625 26336
rect 36659 26333 36671 26367
rect 36613 26327 36671 26333
rect 36998 26324 37004 26376
rect 37056 26364 37062 26376
rect 37458 26364 37464 26376
rect 37056 26336 37464 26364
rect 37056 26324 37062 26336
rect 37458 26324 37464 26336
rect 37516 26324 37522 26376
rect 38470 26324 38476 26376
rect 38528 26364 38534 26376
rect 39117 26367 39175 26373
rect 39117 26364 39129 26367
rect 38528 26336 39129 26364
rect 38528 26324 38534 26336
rect 39117 26333 39129 26336
rect 39163 26333 39175 26367
rect 39117 26327 39175 26333
rect 41432 26296 41460 26540
rect 47486 26528 47492 26540
rect 47544 26528 47550 26580
rect 45554 26460 45560 26512
rect 45612 26500 45618 26512
rect 47949 26503 48007 26509
rect 47949 26500 47961 26503
rect 45612 26472 47961 26500
rect 45612 26460 45618 26472
rect 47949 26469 47961 26472
rect 47995 26469 48007 26503
rect 47949 26463 48007 26469
rect 41506 26324 41512 26376
rect 41564 26364 41570 26376
rect 46934 26364 46940 26376
rect 41564 26336 46940 26364
rect 41564 26324 41570 26336
rect 46934 26324 46940 26336
rect 46992 26324 46998 26376
rect 48130 26364 48136 26376
rect 48091 26336 48136 26364
rect 48130 26324 48136 26336
rect 48188 26324 48194 26376
rect 41690 26296 41696 26308
rect 34992 26268 41460 26296
rect 41651 26268 41696 26296
rect 41690 26256 41696 26268
rect 41748 26256 41754 26308
rect 47302 26296 47308 26308
rect 46952 26268 47308 26296
rect 17586 26188 17592 26240
rect 17644 26228 17650 26240
rect 25774 26228 25780 26240
rect 17644 26200 25780 26228
rect 17644 26188 17650 26200
rect 25774 26188 25780 26200
rect 25832 26188 25838 26240
rect 29730 26188 29736 26240
rect 29788 26228 29794 26240
rect 31294 26228 31300 26240
rect 29788 26200 31300 26228
rect 29788 26188 29794 26200
rect 31294 26188 31300 26200
rect 31352 26228 31358 26240
rect 31573 26231 31631 26237
rect 31573 26228 31585 26231
rect 31352 26200 31585 26228
rect 31352 26188 31358 26200
rect 31573 26197 31585 26200
rect 31619 26197 31631 26231
rect 31573 26191 31631 26197
rect 34057 26231 34115 26237
rect 34057 26197 34069 26231
rect 34103 26228 34115 26231
rect 34698 26228 34704 26240
rect 34103 26200 34704 26228
rect 34103 26197 34115 26200
rect 34057 26191 34115 26197
rect 34698 26188 34704 26200
rect 34756 26188 34762 26240
rect 35526 26188 35532 26240
rect 35584 26228 35590 26240
rect 46952 26228 46980 26268
rect 47302 26256 47308 26268
rect 47360 26256 47366 26308
rect 35584 26200 46980 26228
rect 35584 26188 35590 26200
rect 47026 26188 47032 26240
rect 47084 26228 47090 26240
rect 47854 26228 47860 26240
rect 47084 26200 47860 26228
rect 47084 26188 47090 26200
rect 47854 26188 47860 26200
rect 47912 26188 47918 26240
rect 1104 26138 48852 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 48852 26138
rect 1104 26064 48852 26086
rect 2774 26024 2780 26036
rect 2735 25996 2780 26024
rect 2774 25984 2780 25996
rect 2832 25984 2838 26036
rect 11790 25984 11796 26036
rect 11848 26024 11854 26036
rect 47026 26024 47032 26036
rect 11848 25996 47032 26024
rect 11848 25984 11854 25996
rect 47026 25984 47032 25996
rect 47084 25984 47090 26036
rect 5258 25916 5264 25968
rect 5316 25956 5322 25968
rect 23290 25956 23296 25968
rect 5316 25928 23296 25956
rect 5316 25916 5322 25928
rect 23290 25916 23296 25928
rect 23348 25916 23354 25968
rect 23474 25916 23480 25968
rect 23532 25956 23538 25968
rect 23753 25959 23811 25965
rect 23753 25956 23765 25959
rect 23532 25928 23765 25956
rect 23532 25916 23538 25928
rect 23753 25925 23765 25928
rect 23799 25925 23811 25959
rect 29638 25956 29644 25968
rect 29599 25928 29644 25956
rect 23753 25919 23811 25925
rect 29638 25916 29644 25928
rect 29696 25956 29702 25968
rect 30009 25959 30067 25965
rect 29696 25928 29976 25956
rect 29696 25916 29702 25928
rect 1394 25888 1400 25900
rect 1355 25860 1400 25888
rect 1394 25848 1400 25860
rect 1452 25848 1458 25900
rect 2130 25848 2136 25900
rect 2188 25888 2194 25900
rect 2685 25891 2743 25897
rect 2685 25888 2697 25891
rect 2188 25860 2697 25888
rect 2188 25848 2194 25860
rect 2685 25857 2697 25860
rect 2731 25888 2743 25891
rect 15565 25891 15623 25897
rect 2731 25860 6914 25888
rect 2731 25857 2743 25860
rect 2685 25851 2743 25857
rect 1670 25820 1676 25832
rect 1631 25792 1676 25820
rect 1670 25780 1676 25792
rect 1728 25780 1734 25832
rect 6886 25820 6914 25860
rect 15565 25857 15577 25891
rect 15611 25888 15623 25891
rect 15933 25891 15991 25897
rect 15933 25888 15945 25891
rect 15611 25860 15945 25888
rect 15611 25857 15623 25860
rect 15565 25851 15623 25857
rect 15933 25857 15945 25860
rect 15979 25888 15991 25891
rect 16022 25888 16028 25900
rect 15979 25860 16028 25888
rect 15979 25857 15991 25860
rect 15933 25851 15991 25857
rect 16022 25848 16028 25860
rect 16080 25888 16086 25900
rect 16206 25888 16212 25900
rect 16080 25860 16212 25888
rect 16080 25848 16086 25860
rect 16206 25848 16212 25860
rect 16264 25848 16270 25900
rect 16574 25848 16580 25900
rect 16632 25888 16638 25900
rect 16669 25891 16727 25897
rect 16669 25888 16681 25891
rect 16632 25860 16681 25888
rect 16632 25848 16638 25860
rect 16669 25857 16681 25860
rect 16715 25857 16727 25891
rect 20346 25888 20352 25900
rect 20307 25860 20352 25888
rect 16669 25851 16727 25857
rect 20346 25848 20352 25860
rect 20404 25848 20410 25900
rect 20530 25888 20536 25900
rect 20491 25860 20536 25888
rect 20530 25848 20536 25860
rect 20588 25848 20594 25900
rect 23382 25888 23388 25900
rect 23343 25860 23388 25888
rect 23382 25848 23388 25860
rect 23440 25848 23446 25900
rect 23569 25891 23627 25897
rect 23569 25857 23581 25891
rect 23615 25888 23627 25891
rect 24578 25888 24584 25900
rect 23615 25860 24584 25888
rect 23615 25857 23627 25860
rect 23569 25851 23627 25857
rect 24578 25848 24584 25860
rect 24636 25848 24642 25900
rect 24946 25848 24952 25900
rect 25004 25888 25010 25900
rect 29730 25888 29736 25900
rect 25004 25860 29736 25888
rect 25004 25848 25010 25860
rect 29730 25848 29736 25860
rect 29788 25888 29794 25900
rect 29825 25891 29883 25897
rect 29825 25888 29837 25891
rect 29788 25860 29837 25888
rect 29788 25848 29794 25860
rect 29825 25857 29837 25860
rect 29871 25857 29883 25891
rect 29948 25888 29976 25928
rect 30009 25925 30021 25959
rect 30055 25956 30067 25959
rect 30282 25956 30288 25968
rect 30055 25928 30288 25956
rect 30055 25925 30067 25928
rect 30009 25919 30067 25925
rect 30282 25916 30288 25928
rect 30340 25916 30346 25968
rect 30484 25928 30696 25956
rect 30484 25888 30512 25928
rect 29948 25860 30512 25888
rect 30561 25891 30619 25897
rect 29825 25851 29883 25857
rect 30561 25857 30573 25891
rect 30607 25857 30619 25891
rect 30668 25888 30696 25928
rect 30742 25916 30748 25968
rect 30800 25956 30806 25968
rect 30800 25928 30845 25956
rect 30800 25916 30806 25928
rect 34054 25916 34060 25968
rect 34112 25956 34118 25968
rect 34977 25959 35035 25965
rect 34977 25956 34989 25959
rect 34112 25928 34989 25956
rect 34112 25916 34118 25928
rect 34977 25925 34989 25928
rect 35023 25925 35035 25959
rect 34977 25919 35035 25925
rect 35161 25959 35219 25965
rect 35161 25925 35173 25959
rect 35207 25956 35219 25959
rect 35802 25956 35808 25968
rect 35207 25928 35808 25956
rect 35207 25925 35219 25928
rect 35161 25919 35219 25925
rect 35802 25916 35808 25928
rect 35860 25916 35866 25968
rect 36078 25916 36084 25968
rect 36136 25956 36142 25968
rect 36136 25928 36489 25956
rect 36136 25916 36142 25928
rect 32950 25888 32956 25900
rect 30668 25860 32956 25888
rect 30561 25851 30619 25857
rect 17034 25820 17040 25832
rect 6886 25792 17040 25820
rect 17034 25780 17040 25792
rect 17092 25780 17098 25832
rect 17129 25823 17187 25829
rect 17129 25789 17141 25823
rect 17175 25820 17187 25823
rect 30098 25820 30104 25832
rect 17175 25792 30104 25820
rect 17175 25789 17187 25792
rect 17129 25783 17187 25789
rect 2498 25712 2504 25764
rect 2556 25752 2562 25764
rect 17144 25752 17172 25783
rect 30098 25780 30104 25792
rect 30156 25780 30162 25832
rect 30282 25780 30288 25832
rect 30340 25820 30346 25832
rect 30576 25820 30604 25851
rect 32950 25848 32956 25860
rect 33008 25848 33014 25900
rect 33134 25848 33140 25900
rect 33192 25897 33198 25900
rect 33192 25891 33241 25897
rect 33192 25857 33195 25891
rect 33229 25857 33241 25891
rect 33315 25888 33321 25900
rect 33276 25860 33321 25888
rect 33192 25851 33241 25857
rect 33192 25848 33198 25851
rect 33315 25848 33321 25860
rect 33373 25848 33379 25900
rect 33413 25891 33471 25897
rect 33413 25888 33425 25891
rect 33408 25857 33425 25888
rect 33459 25857 33471 25891
rect 33408 25851 33471 25857
rect 33597 25891 33655 25897
rect 33597 25857 33609 25891
rect 33643 25888 33655 25891
rect 33778 25888 33784 25900
rect 33643 25860 33784 25888
rect 33643 25857 33655 25860
rect 33597 25851 33655 25857
rect 30340 25792 30604 25820
rect 30340 25780 30346 25792
rect 32766 25780 32772 25832
rect 32824 25820 32830 25832
rect 33408 25820 33436 25851
rect 33778 25848 33784 25860
rect 33836 25848 33842 25900
rect 36461 25897 36489 25928
rect 36630 25916 36636 25968
rect 36688 25956 36694 25968
rect 45554 25956 45560 25968
rect 36688 25928 45560 25956
rect 36688 25916 36694 25928
rect 45554 25916 45560 25928
rect 45612 25916 45618 25968
rect 36311 25891 36369 25897
rect 36311 25888 36323 25891
rect 36188 25860 36323 25888
rect 32824 25792 33436 25820
rect 32824 25780 32830 25792
rect 34514 25780 34520 25832
rect 34572 25820 34578 25832
rect 35434 25820 35440 25832
rect 34572 25792 35440 25820
rect 34572 25780 34578 25792
rect 35434 25780 35440 25792
rect 35492 25780 35498 25832
rect 36188 25820 36216 25860
rect 36311 25857 36323 25860
rect 36357 25857 36369 25891
rect 36311 25851 36369 25857
rect 36449 25891 36507 25897
rect 36449 25857 36461 25891
rect 36495 25857 36507 25891
rect 36449 25851 36507 25857
rect 36538 25848 36544 25900
rect 36596 25888 36602 25900
rect 36725 25891 36783 25897
rect 36596 25860 36638 25888
rect 36596 25848 36602 25860
rect 36725 25857 36737 25891
rect 36771 25888 36783 25891
rect 36814 25888 36820 25900
rect 36771 25860 36820 25888
rect 36771 25857 36783 25860
rect 36725 25851 36783 25857
rect 36814 25848 36820 25860
rect 36872 25848 36878 25900
rect 36998 25848 37004 25900
rect 37056 25888 37062 25900
rect 42334 25888 42340 25900
rect 37056 25860 42340 25888
rect 37056 25848 37062 25860
rect 42334 25848 42340 25860
rect 42392 25848 42398 25900
rect 36630 25820 36636 25832
rect 36188 25792 36636 25820
rect 36630 25780 36636 25792
rect 36688 25780 36694 25832
rect 36906 25780 36912 25832
rect 36964 25820 36970 25832
rect 45189 25823 45247 25829
rect 45189 25820 45201 25823
rect 36964 25792 45201 25820
rect 36964 25780 36970 25792
rect 45189 25789 45201 25792
rect 45235 25789 45247 25823
rect 45189 25783 45247 25789
rect 45373 25823 45431 25829
rect 45373 25789 45385 25823
rect 45419 25820 45431 25823
rect 45738 25820 45744 25832
rect 45419 25792 45744 25820
rect 45419 25789 45431 25792
rect 45373 25783 45431 25789
rect 45738 25780 45744 25792
rect 45796 25780 45802 25832
rect 46842 25820 46848 25832
rect 46803 25792 46848 25820
rect 46842 25780 46848 25792
rect 46900 25780 46906 25832
rect 47486 25780 47492 25832
rect 47544 25820 47550 25832
rect 47762 25820 47768 25832
rect 47544 25792 47768 25820
rect 47544 25780 47550 25792
rect 47762 25780 47768 25792
rect 47820 25780 47826 25832
rect 17218 25752 17224 25764
rect 2556 25724 17224 25752
rect 2556 25712 2562 25724
rect 17218 25712 17224 25724
rect 17276 25712 17282 25764
rect 21082 25752 21088 25764
rect 17328 25724 21088 25752
rect 15654 25644 15660 25696
rect 15712 25684 15718 25696
rect 16025 25687 16083 25693
rect 16025 25684 16037 25687
rect 15712 25656 16037 25684
rect 15712 25644 15718 25656
rect 16025 25653 16037 25656
rect 16071 25653 16083 25687
rect 16025 25647 16083 25653
rect 16206 25644 16212 25696
rect 16264 25684 16270 25696
rect 17328 25684 17356 25724
rect 21082 25712 21088 25724
rect 21140 25712 21146 25764
rect 28994 25712 29000 25764
rect 29052 25752 29058 25764
rect 30466 25752 30472 25764
rect 29052 25724 30472 25752
rect 29052 25712 29058 25724
rect 30466 25712 30472 25724
rect 30524 25712 30530 25764
rect 16264 25656 17356 25684
rect 20717 25687 20775 25693
rect 16264 25644 16270 25656
rect 20717 25653 20729 25687
rect 20763 25684 20775 25687
rect 24854 25684 24860 25696
rect 20763 25656 24860 25684
rect 20763 25653 20775 25656
rect 20717 25647 20775 25653
rect 24854 25644 24860 25656
rect 24912 25644 24918 25696
rect 25590 25644 25596 25696
rect 25648 25684 25654 25696
rect 29730 25684 29736 25696
rect 25648 25656 29736 25684
rect 25648 25644 25654 25656
rect 29730 25644 29736 25656
rect 29788 25644 29794 25696
rect 32953 25687 33011 25693
rect 32953 25653 32965 25687
rect 32999 25684 33011 25687
rect 33502 25684 33508 25696
rect 32999 25656 33508 25684
rect 32999 25653 33011 25656
rect 32953 25647 33011 25653
rect 33502 25644 33508 25656
rect 33560 25644 33566 25696
rect 34514 25644 34520 25696
rect 34572 25684 34578 25696
rect 34790 25684 34796 25696
rect 34572 25656 34796 25684
rect 34572 25644 34578 25656
rect 34790 25644 34796 25656
rect 34848 25644 34854 25696
rect 36081 25687 36139 25693
rect 36081 25653 36093 25687
rect 36127 25684 36139 25687
rect 36354 25684 36360 25696
rect 36127 25656 36360 25684
rect 36127 25653 36139 25656
rect 36081 25647 36139 25653
rect 36354 25644 36360 25656
rect 36412 25644 36418 25696
rect 47762 25684 47768 25696
rect 47723 25656 47768 25684
rect 47762 25644 47768 25656
rect 47820 25644 47826 25696
rect 1104 25594 48852 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 48852 25594
rect 1104 25520 48852 25542
rect 1670 25440 1676 25492
rect 1728 25480 1734 25492
rect 1728 25452 6914 25480
rect 1728 25440 1734 25452
rect 2498 25372 2504 25424
rect 2556 25412 2562 25424
rect 2866 25412 2872 25424
rect 2556 25384 2872 25412
rect 2556 25372 2562 25384
rect 2866 25372 2872 25384
rect 2924 25372 2930 25424
rect 6886 25344 6914 25452
rect 11882 25440 11888 25492
rect 11940 25480 11946 25492
rect 19981 25483 20039 25489
rect 11940 25452 12434 25480
rect 11940 25440 11946 25452
rect 12406 25412 12434 25452
rect 19981 25449 19993 25483
rect 20027 25480 20039 25483
rect 20162 25480 20168 25492
rect 20027 25452 20168 25480
rect 20027 25449 20039 25452
rect 19981 25443 20039 25449
rect 20162 25440 20168 25452
rect 20220 25440 20226 25492
rect 20714 25480 20720 25492
rect 20675 25452 20720 25480
rect 20714 25440 20720 25452
rect 20772 25480 20778 25492
rect 20898 25480 20904 25492
rect 20772 25452 20904 25480
rect 20772 25440 20778 25452
rect 20898 25440 20904 25452
rect 20956 25440 20962 25492
rect 25590 25480 25596 25492
rect 21008 25452 25596 25480
rect 12406 25384 20944 25412
rect 18782 25344 18788 25356
rect 6886 25316 18788 25344
rect 18782 25304 18788 25316
rect 18840 25344 18846 25356
rect 19889 25347 19947 25353
rect 18840 25316 19748 25344
rect 18840 25304 18846 25316
rect 15105 25279 15163 25285
rect 15105 25245 15117 25279
rect 15151 25276 15163 25279
rect 16574 25276 16580 25288
rect 15151 25248 16580 25276
rect 15151 25245 15163 25248
rect 15105 25239 15163 25245
rect 16574 25236 16580 25248
rect 16632 25236 16638 25288
rect 17586 25276 17592 25288
rect 17547 25248 17592 25276
rect 17586 25236 17592 25248
rect 17644 25236 17650 25288
rect 19720 25285 19748 25316
rect 19889 25313 19901 25347
rect 19935 25344 19947 25347
rect 20070 25344 20076 25356
rect 19935 25316 20076 25344
rect 19935 25313 19947 25316
rect 19889 25307 19947 25313
rect 20070 25304 20076 25316
rect 20128 25344 20134 25356
rect 20622 25344 20628 25356
rect 20128 25316 20628 25344
rect 20128 25304 20134 25316
rect 20622 25304 20628 25316
rect 20680 25304 20686 25356
rect 20806 25344 20812 25356
rect 20767 25316 20812 25344
rect 20806 25304 20812 25316
rect 20864 25304 20870 25356
rect 19705 25279 19763 25285
rect 19705 25245 19717 25279
rect 19751 25245 19763 25279
rect 19705 25239 19763 25245
rect 19794 25236 19800 25288
rect 19852 25276 19858 25288
rect 19981 25279 20039 25285
rect 19981 25276 19993 25279
rect 19852 25248 19993 25276
rect 19852 25236 19858 25248
rect 19981 25245 19993 25248
rect 20027 25245 20039 25279
rect 19981 25239 20039 25245
rect 20088 25248 20852 25276
rect 6822 25168 6828 25220
rect 6880 25208 6886 25220
rect 15841 25211 15899 25217
rect 6880 25168 6914 25208
rect 15841 25177 15853 25211
rect 15887 25208 15899 25211
rect 16022 25208 16028 25220
rect 15887 25180 16028 25208
rect 15887 25177 15899 25180
rect 15841 25171 15899 25177
rect 16022 25168 16028 25180
rect 16080 25168 16086 25220
rect 19334 25168 19340 25220
rect 19392 25208 19398 25220
rect 20088 25208 20116 25248
rect 20714 25208 20720 25220
rect 19392 25180 20116 25208
rect 20675 25180 20720 25208
rect 19392 25168 19398 25180
rect 20714 25168 20720 25180
rect 20772 25168 20778 25220
rect 6886 25140 6914 25168
rect 17402 25140 17408 25152
rect 6886 25112 17408 25140
rect 17402 25100 17408 25112
rect 17460 25100 17466 25152
rect 20165 25143 20223 25149
rect 20165 25109 20177 25143
rect 20211 25140 20223 25143
rect 20254 25140 20260 25152
rect 20211 25112 20260 25140
rect 20211 25109 20223 25112
rect 20165 25103 20223 25109
rect 20254 25100 20260 25112
rect 20312 25100 20318 25152
rect 20824 25140 20852 25248
rect 20916 25208 20944 25384
rect 21008 25285 21036 25452
rect 25590 25440 25596 25452
rect 25648 25440 25654 25492
rect 25774 25440 25780 25492
rect 25832 25480 25838 25492
rect 35526 25480 35532 25492
rect 25832 25452 35532 25480
rect 25832 25440 25838 25452
rect 35526 25440 35532 25452
rect 35584 25440 35590 25492
rect 35802 25480 35808 25492
rect 35763 25452 35808 25480
rect 35802 25440 35808 25452
rect 35860 25440 35866 25492
rect 45738 25480 45744 25492
rect 36004 25452 40632 25480
rect 45699 25452 45744 25480
rect 21082 25372 21088 25424
rect 21140 25412 21146 25424
rect 34514 25412 34520 25424
rect 21140 25384 34520 25412
rect 21140 25372 21146 25384
rect 34514 25372 34520 25384
rect 34572 25372 34578 25424
rect 24486 25304 24492 25356
rect 24544 25344 24550 25356
rect 26418 25344 26424 25356
rect 24544 25316 25452 25344
rect 24544 25304 24550 25316
rect 20993 25279 21051 25285
rect 20993 25245 21005 25279
rect 21039 25245 21051 25279
rect 20993 25239 21051 25245
rect 23290 25236 23296 25288
rect 23348 25276 23354 25288
rect 25424 25285 25452 25316
rect 25516 25316 26424 25344
rect 25516 25285 25544 25316
rect 26418 25304 26424 25316
rect 26476 25304 26482 25356
rect 28994 25344 29000 25356
rect 28955 25316 29000 25344
rect 28994 25304 29000 25316
rect 29052 25304 29058 25356
rect 30006 25304 30012 25356
rect 30064 25344 30070 25356
rect 36004 25344 36032 25452
rect 30064 25316 30788 25344
rect 30064 25304 30070 25316
rect 25317 25279 25375 25285
rect 25317 25276 25329 25279
rect 23348 25248 25329 25276
rect 23348 25236 23354 25248
rect 25317 25245 25329 25248
rect 25363 25245 25375 25279
rect 25317 25239 25375 25245
rect 25409 25279 25467 25285
rect 25409 25245 25421 25279
rect 25455 25245 25467 25279
rect 25409 25239 25467 25245
rect 25501 25279 25559 25285
rect 25501 25245 25513 25279
rect 25547 25245 25559 25279
rect 25501 25239 25559 25245
rect 25682 25236 25688 25288
rect 25740 25276 25746 25288
rect 26050 25276 26056 25288
rect 25740 25248 26056 25276
rect 25740 25236 25746 25248
rect 26050 25236 26056 25248
rect 26108 25236 26114 25288
rect 30331 25279 30389 25285
rect 30331 25276 30343 25279
rect 26252 25273 28856 25276
rect 28920 25273 30343 25276
rect 26252 25248 30343 25273
rect 26252 25208 26280 25248
rect 28828 25245 28948 25248
rect 30331 25245 30343 25248
rect 30377 25245 30389 25279
rect 30466 25276 30472 25288
rect 30427 25248 30472 25276
rect 30331 25239 30389 25245
rect 30466 25236 30472 25248
rect 30524 25236 30530 25288
rect 30760 25285 30788 25316
rect 33428 25316 36032 25344
rect 33428 25285 33456 25316
rect 30582 25279 30640 25285
rect 30582 25245 30594 25279
rect 30628 25276 30640 25279
rect 30739 25279 30797 25285
rect 30628 25248 30696 25276
rect 30628 25245 30640 25248
rect 30582 25239 30640 25245
rect 20916 25180 26280 25208
rect 27614 25168 27620 25220
rect 27672 25208 27678 25220
rect 28077 25211 28135 25217
rect 28077 25208 28089 25211
rect 27672 25180 28089 25208
rect 27672 25168 27678 25180
rect 28077 25177 28089 25180
rect 28123 25208 28135 25211
rect 28813 25211 28871 25217
rect 28813 25208 28825 25211
rect 28123 25180 28825 25208
rect 28123 25177 28135 25180
rect 28077 25171 28135 25177
rect 28813 25177 28825 25180
rect 28859 25177 28871 25211
rect 28813 25171 28871 25177
rect 21177 25143 21235 25149
rect 21177 25140 21189 25143
rect 20824 25112 21189 25140
rect 21177 25109 21189 25112
rect 21223 25109 21235 25143
rect 21177 25103 21235 25109
rect 25041 25143 25099 25149
rect 25041 25109 25053 25143
rect 25087 25140 25099 25143
rect 25590 25140 25596 25152
rect 25087 25112 25596 25140
rect 25087 25109 25099 25112
rect 25041 25103 25099 25109
rect 25590 25100 25596 25112
rect 25648 25100 25654 25152
rect 26234 25100 26240 25152
rect 26292 25140 26298 25152
rect 28169 25143 28227 25149
rect 28169 25140 28181 25143
rect 26292 25112 28181 25140
rect 26292 25100 26298 25112
rect 28169 25109 28181 25112
rect 28215 25140 28227 25143
rect 30006 25140 30012 25152
rect 28215 25112 30012 25140
rect 28215 25109 28227 25112
rect 28169 25103 28227 25109
rect 30006 25100 30012 25112
rect 30064 25100 30070 25152
rect 30101 25143 30159 25149
rect 30101 25109 30113 25143
rect 30147 25140 30159 25143
rect 30466 25140 30472 25152
rect 30147 25112 30472 25140
rect 30147 25109 30159 25112
rect 30101 25103 30159 25109
rect 30466 25100 30472 25112
rect 30524 25100 30530 25152
rect 30668 25140 30696 25248
rect 30739 25245 30751 25279
rect 30785 25245 30797 25279
rect 30739 25239 30797 25245
rect 33413 25279 33471 25285
rect 33413 25245 33425 25279
rect 33459 25245 33471 25279
rect 33413 25239 33471 25245
rect 33505 25279 33563 25285
rect 33505 25245 33517 25279
rect 33551 25245 33563 25279
rect 33505 25239 33563 25245
rect 30834 25168 30840 25220
rect 30892 25208 30898 25220
rect 31205 25211 31263 25217
rect 31205 25208 31217 25211
rect 30892 25180 31217 25208
rect 30892 25168 30898 25180
rect 31205 25177 31217 25180
rect 31251 25177 31263 25211
rect 31386 25208 31392 25220
rect 31347 25180 31392 25208
rect 31205 25171 31263 25177
rect 31386 25168 31392 25180
rect 31444 25168 31450 25220
rect 32122 25168 32128 25220
rect 32180 25208 32186 25220
rect 33318 25208 33324 25220
rect 32180 25180 33324 25208
rect 32180 25168 32186 25180
rect 33318 25168 33324 25180
rect 33376 25208 33382 25220
rect 33520 25208 33548 25239
rect 33594 25236 33600 25288
rect 33652 25276 33658 25288
rect 33652 25248 33697 25276
rect 33652 25236 33658 25248
rect 33778 25236 33784 25288
rect 33836 25276 33842 25288
rect 36262 25276 36268 25288
rect 33836 25248 33881 25276
rect 36223 25248 36268 25276
rect 33836 25236 33842 25248
rect 36262 25236 36268 25248
rect 36320 25236 36326 25288
rect 36354 25236 36360 25288
rect 36412 25276 36418 25288
rect 36521 25279 36579 25285
rect 36521 25276 36533 25279
rect 36412 25248 36533 25276
rect 36412 25236 36418 25248
rect 36521 25245 36533 25248
rect 36567 25245 36579 25279
rect 36521 25239 36579 25245
rect 40313 25279 40371 25285
rect 40313 25245 40325 25279
rect 40359 25276 40371 25279
rect 40494 25276 40500 25288
rect 40359 25248 40500 25276
rect 40359 25245 40371 25248
rect 40313 25239 40371 25245
rect 40494 25236 40500 25248
rect 40552 25236 40558 25288
rect 40604 25276 40632 25452
rect 45738 25440 45744 25452
rect 45796 25440 45802 25492
rect 47026 25440 47032 25492
rect 47084 25480 47090 25492
rect 47121 25483 47179 25489
rect 47121 25480 47133 25483
rect 47084 25452 47133 25480
rect 47084 25440 47090 25452
rect 47121 25449 47133 25452
rect 47167 25480 47179 25483
rect 47854 25480 47860 25492
rect 47167 25452 47532 25480
rect 47815 25452 47860 25480
rect 47167 25449 47179 25452
rect 47121 25443 47179 25449
rect 40678 25372 40684 25424
rect 40736 25412 40742 25424
rect 47394 25412 47400 25424
rect 40736 25384 47400 25412
rect 40736 25372 40742 25384
rect 47394 25372 47400 25384
rect 47452 25372 47458 25424
rect 47504 25353 47532 25452
rect 47854 25440 47860 25452
rect 47912 25440 47918 25492
rect 47489 25347 47547 25353
rect 47489 25313 47501 25347
rect 47535 25313 47547 25347
rect 47489 25307 47547 25313
rect 41598 25276 41604 25288
rect 40604 25248 41604 25276
rect 41598 25236 41604 25248
rect 41656 25236 41662 25288
rect 45649 25279 45707 25285
rect 45649 25245 45661 25279
rect 45695 25276 45707 25279
rect 46198 25276 46204 25288
rect 45695 25248 46204 25276
rect 45695 25245 45707 25248
rect 45649 25239 45707 25245
rect 46198 25236 46204 25248
rect 46256 25236 46262 25288
rect 46382 25236 46388 25288
rect 46440 25276 46446 25288
rect 47857 25279 47915 25285
rect 47857 25276 47869 25279
rect 46440 25248 47869 25276
rect 46440 25236 46446 25248
rect 47857 25245 47869 25248
rect 47903 25245 47915 25279
rect 47857 25239 47915 25245
rect 33376 25180 33548 25208
rect 33376 25168 33382 25180
rect 35434 25168 35440 25220
rect 35492 25208 35498 25220
rect 35621 25211 35679 25217
rect 35492 25180 35537 25208
rect 35492 25168 35498 25180
rect 35621 25177 35633 25211
rect 35667 25177 35679 25211
rect 35621 25171 35679 25177
rect 31573 25143 31631 25149
rect 31573 25140 31585 25143
rect 30668 25112 31585 25140
rect 31573 25109 31585 25112
rect 31619 25109 31631 25143
rect 31573 25103 31631 25109
rect 33137 25143 33195 25149
rect 33137 25109 33149 25143
rect 33183 25140 33195 25143
rect 34790 25140 34796 25152
rect 33183 25112 34796 25140
rect 33183 25109 33195 25112
rect 33137 25103 33195 25109
rect 34790 25100 34796 25112
rect 34848 25100 34854 25152
rect 35636 25140 35664 25171
rect 35802 25168 35808 25220
rect 35860 25208 35866 25220
rect 35860 25180 47716 25208
rect 35860 25168 35866 25180
rect 37274 25140 37280 25152
rect 35636 25112 37280 25140
rect 37274 25100 37280 25112
rect 37332 25100 37338 25152
rect 37642 25140 37648 25152
rect 37603 25112 37648 25140
rect 37642 25100 37648 25112
rect 37700 25100 37706 25152
rect 40126 25140 40132 25152
rect 40087 25112 40132 25140
rect 40126 25100 40132 25112
rect 40184 25100 40190 25152
rect 47688 25149 47716 25180
rect 47673 25143 47731 25149
rect 47673 25109 47685 25143
rect 47719 25109 47731 25143
rect 47673 25103 47731 25109
rect 1104 25050 48852 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 48852 25050
rect 1104 24976 48852 24998
rect 20165 24939 20223 24945
rect 20165 24905 20177 24939
rect 20211 24936 20223 24939
rect 20530 24936 20536 24948
rect 20211 24908 20536 24936
rect 20211 24905 20223 24908
rect 20165 24899 20223 24905
rect 20530 24896 20536 24908
rect 20588 24896 20594 24948
rect 20714 24896 20720 24948
rect 20772 24936 20778 24948
rect 21085 24939 21143 24945
rect 21085 24936 21097 24939
rect 20772 24908 21097 24936
rect 20772 24896 20778 24908
rect 21085 24905 21097 24908
rect 21131 24905 21143 24939
rect 21085 24899 21143 24905
rect 27982 24896 27988 24948
rect 28040 24936 28046 24948
rect 29086 24936 29092 24948
rect 28040 24908 29092 24936
rect 28040 24896 28046 24908
rect 29086 24896 29092 24908
rect 29144 24896 29150 24948
rect 32766 24936 32772 24948
rect 32727 24908 32772 24936
rect 32766 24896 32772 24908
rect 32824 24896 32830 24948
rect 33778 24936 33784 24948
rect 33244 24908 33784 24936
rect 20070 24868 20076 24880
rect 19628 24840 20076 24868
rect 2130 24800 2136 24812
rect 2091 24772 2136 24800
rect 2130 24760 2136 24772
rect 2188 24760 2194 24812
rect 15654 24760 15660 24812
rect 15712 24800 15718 24812
rect 15749 24803 15807 24809
rect 15749 24800 15761 24803
rect 15712 24772 15761 24800
rect 15712 24760 15718 24772
rect 15749 24769 15761 24772
rect 15795 24769 15807 24803
rect 15749 24763 15807 24769
rect 16117 24803 16175 24809
rect 16117 24769 16129 24803
rect 16163 24800 16175 24803
rect 16574 24800 16580 24812
rect 16163 24772 16580 24800
rect 16163 24769 16175 24772
rect 16117 24763 16175 24769
rect 16574 24760 16580 24772
rect 16632 24800 16638 24812
rect 16669 24803 16727 24809
rect 16669 24800 16681 24803
rect 16632 24772 16681 24800
rect 16632 24760 16638 24772
rect 16669 24769 16681 24772
rect 16715 24769 16727 24803
rect 16669 24763 16727 24769
rect 17494 24760 17500 24812
rect 17552 24800 17558 24812
rect 17862 24800 17868 24812
rect 17552 24772 17868 24800
rect 17552 24760 17558 24772
rect 17862 24760 17868 24772
rect 17920 24760 17926 24812
rect 18782 24800 18788 24812
rect 18743 24772 18788 24800
rect 18782 24760 18788 24772
rect 18840 24760 18846 24812
rect 19061 24803 19119 24809
rect 19061 24769 19073 24803
rect 19107 24800 19119 24803
rect 19628 24800 19656 24840
rect 20070 24828 20076 24840
rect 20128 24828 20134 24880
rect 20254 24828 20260 24880
rect 20312 24868 20318 24880
rect 20806 24868 20812 24880
rect 20312 24840 20812 24868
rect 20312 24828 20318 24840
rect 20806 24828 20812 24840
rect 20864 24828 20870 24880
rect 28442 24868 28448 24880
rect 22756 24840 28448 24868
rect 19107 24772 19656 24800
rect 19705 24803 19763 24809
rect 19107 24769 19119 24772
rect 19061 24763 19119 24769
rect 19705 24769 19717 24803
rect 19751 24769 19763 24803
rect 19978 24800 19984 24812
rect 19939 24772 19984 24800
rect 19705 24763 19763 24769
rect 1854 24692 1860 24744
rect 1912 24732 1918 24744
rect 17129 24735 17187 24741
rect 17129 24732 17141 24735
rect 1912 24704 17141 24732
rect 1912 24692 1918 24704
rect 17129 24701 17141 24704
rect 17175 24732 17187 24735
rect 17310 24732 17316 24744
rect 17175 24704 17316 24732
rect 17175 24701 17187 24704
rect 17129 24695 17187 24701
rect 17310 24692 17316 24704
rect 17368 24692 17374 24744
rect 18877 24735 18935 24741
rect 18877 24701 18889 24735
rect 18923 24732 18935 24735
rect 19720 24732 19748 24763
rect 19978 24760 19984 24772
rect 20036 24760 20042 24812
rect 20622 24800 20628 24812
rect 20583 24772 20628 24800
rect 20622 24760 20628 24772
rect 20680 24760 20686 24812
rect 20714 24760 20720 24812
rect 20772 24800 20778 24812
rect 20901 24803 20959 24809
rect 20901 24800 20913 24803
rect 20772 24772 20913 24800
rect 20772 24760 20778 24772
rect 20901 24769 20913 24772
rect 20947 24769 20959 24803
rect 20901 24763 20959 24769
rect 21818 24760 21824 24812
rect 21876 24800 21882 24812
rect 22756 24809 22784 24840
rect 28442 24828 28448 24840
rect 28500 24828 28506 24880
rect 30006 24828 30012 24880
rect 30064 24868 30070 24880
rect 32214 24868 32220 24880
rect 30064 24840 32220 24868
rect 30064 24828 30070 24840
rect 32214 24828 32220 24840
rect 32272 24868 32278 24880
rect 33244 24868 33272 24908
rect 33778 24896 33784 24908
rect 33836 24896 33842 24948
rect 35894 24896 35900 24948
rect 35952 24936 35958 24948
rect 40678 24936 40684 24948
rect 35952 24908 40684 24936
rect 35952 24896 35958 24908
rect 40678 24896 40684 24908
rect 40736 24896 40742 24948
rect 41800 24908 42840 24936
rect 33502 24877 33508 24880
rect 32272 24840 33272 24868
rect 32272 24828 32278 24840
rect 33496 24831 33508 24877
rect 33560 24868 33566 24880
rect 33560 24840 33596 24868
rect 33502 24828 33508 24831
rect 33560 24828 33566 24840
rect 35526 24828 35532 24880
rect 35584 24868 35590 24880
rect 36906 24868 36912 24880
rect 35584 24840 36912 24868
rect 35584 24828 35590 24840
rect 36906 24828 36912 24840
rect 36964 24828 36970 24880
rect 41046 24868 41052 24880
rect 39684 24840 41052 24868
rect 22741 24803 22799 24809
rect 22741 24800 22753 24803
rect 21876 24772 22753 24800
rect 21876 24760 21882 24772
rect 22741 24769 22753 24772
rect 22787 24769 22799 24803
rect 22741 24763 22799 24769
rect 22925 24803 22983 24809
rect 22925 24769 22937 24803
rect 22971 24769 22983 24803
rect 22925 24763 22983 24769
rect 18923 24704 19748 24732
rect 19889 24735 19947 24741
rect 18923 24701 18935 24704
rect 18877 24695 18935 24701
rect 19889 24701 19901 24735
rect 19935 24701 19947 24735
rect 19889 24695 19947 24701
rect 20809 24735 20867 24741
rect 20809 24701 20821 24735
rect 20855 24732 20867 24735
rect 21082 24732 21088 24744
rect 20855 24704 21088 24732
rect 20855 24701 20867 24704
rect 20809 24695 20867 24701
rect 6730 24624 6736 24676
rect 6788 24664 6794 24676
rect 18892 24664 18920 24695
rect 6788 24636 18920 24664
rect 19245 24667 19303 24673
rect 6788 24624 6794 24636
rect 19245 24633 19257 24667
rect 19291 24664 19303 24667
rect 19702 24664 19708 24676
rect 19291 24636 19708 24664
rect 19291 24633 19303 24636
rect 19245 24627 19303 24633
rect 19702 24624 19708 24636
rect 19760 24624 19766 24676
rect 19904 24664 19932 24695
rect 21082 24692 21088 24704
rect 21140 24692 21146 24744
rect 22940 24732 22968 24763
rect 23014 24760 23020 24812
rect 23072 24800 23078 24812
rect 23474 24800 23480 24812
rect 23072 24772 23117 24800
rect 23435 24772 23480 24800
rect 23072 24760 23078 24772
rect 23474 24760 23480 24772
rect 23532 24760 23538 24812
rect 24949 24803 25007 24809
rect 24949 24769 24961 24803
rect 24995 24800 25007 24803
rect 25038 24800 25044 24812
rect 24995 24772 25044 24800
rect 24995 24769 25007 24772
rect 24949 24763 25007 24769
rect 25038 24760 25044 24772
rect 25096 24760 25102 24812
rect 25222 24809 25228 24812
rect 25216 24763 25228 24809
rect 25280 24800 25286 24812
rect 27982 24800 27988 24812
rect 25280 24772 25316 24800
rect 27943 24772 27988 24800
rect 25222 24760 25228 24763
rect 25280 24760 25286 24772
rect 27982 24760 27988 24772
rect 28040 24760 28046 24812
rect 28261 24803 28319 24809
rect 28261 24769 28273 24803
rect 28307 24800 28319 24803
rect 29181 24803 29239 24809
rect 28307 24772 29132 24800
rect 28307 24769 28319 24772
rect 28261 24763 28319 24769
rect 23566 24732 23572 24744
rect 22940 24704 23572 24732
rect 23566 24692 23572 24704
rect 23624 24692 23630 24744
rect 28169 24735 28227 24741
rect 28169 24701 28181 24735
rect 28215 24732 28227 24735
rect 28534 24732 28540 24744
rect 28215 24704 28540 24732
rect 28215 24701 28227 24704
rect 28169 24695 28227 24701
rect 28534 24692 28540 24704
rect 28592 24692 28598 24744
rect 28905 24735 28963 24741
rect 28905 24701 28917 24735
rect 28951 24732 28963 24735
rect 28994 24732 29000 24744
rect 28951 24704 29000 24732
rect 28951 24701 28963 24704
rect 28905 24695 28963 24701
rect 28994 24692 29000 24704
rect 29052 24692 29058 24744
rect 29104 24732 29132 24772
rect 29181 24769 29193 24803
rect 29227 24800 29239 24803
rect 29638 24800 29644 24812
rect 29227 24772 29644 24800
rect 29227 24769 29239 24772
rect 29181 24763 29239 24769
rect 29638 24760 29644 24772
rect 29696 24760 29702 24812
rect 30466 24809 30472 24812
rect 30460 24800 30472 24809
rect 30427 24772 30472 24800
rect 30460 24763 30472 24772
rect 30466 24760 30472 24763
rect 30524 24760 30530 24812
rect 30834 24760 30840 24812
rect 30892 24800 30898 24812
rect 32398 24800 32404 24812
rect 30892 24772 32404 24800
rect 30892 24760 30898 24772
rect 32398 24760 32404 24772
rect 32456 24760 32462 24812
rect 32585 24803 32643 24809
rect 32585 24769 32597 24803
rect 32631 24800 32643 24803
rect 33318 24800 33324 24812
rect 32631 24772 33324 24800
rect 32631 24769 32643 24772
rect 32585 24763 32643 24769
rect 33318 24760 33324 24772
rect 33376 24800 33382 24812
rect 33376 24772 34468 24800
rect 33376 24760 33382 24772
rect 30098 24732 30104 24744
rect 29104 24704 30104 24732
rect 29656 24676 29684 24704
rect 30098 24692 30104 24704
rect 30156 24692 30162 24744
rect 30190 24692 30196 24744
rect 30248 24732 30254 24744
rect 30248 24704 30293 24732
rect 30248 24692 30254 24704
rect 32674 24692 32680 24744
rect 32732 24732 32738 24744
rect 33229 24735 33287 24741
rect 33229 24732 33241 24735
rect 32732 24704 33241 24732
rect 32732 24692 32738 24704
rect 33229 24701 33241 24704
rect 33275 24701 33287 24735
rect 34440 24732 34468 24772
rect 34514 24760 34520 24812
rect 34572 24800 34578 24812
rect 39684 24800 39712 24840
rect 41046 24828 41052 24840
rect 41104 24828 41110 24880
rect 34572 24772 39712 24800
rect 39752 24803 39810 24809
rect 34572 24760 34578 24772
rect 39752 24769 39764 24803
rect 39798 24800 39810 24803
rect 40126 24800 40132 24812
rect 39798 24772 40132 24800
rect 39798 24769 39810 24772
rect 39752 24763 39810 24769
rect 40126 24760 40132 24772
rect 40184 24760 40190 24812
rect 40218 24760 40224 24812
rect 40276 24800 40282 24812
rect 41800 24800 41828 24908
rect 40276 24772 41828 24800
rect 41877 24803 41935 24809
rect 40276 24760 40282 24772
rect 41877 24769 41889 24803
rect 41923 24800 41935 24803
rect 41966 24800 41972 24812
rect 41923 24772 41972 24800
rect 41923 24769 41935 24772
rect 41877 24763 41935 24769
rect 41966 24760 41972 24772
rect 42024 24760 42030 24812
rect 42426 24800 42432 24812
rect 42092 24772 42432 24800
rect 34440 24704 34652 24732
rect 33229 24695 33287 24701
rect 19904 24636 24808 24664
rect 1946 24556 1952 24608
rect 2004 24596 2010 24608
rect 2225 24599 2283 24605
rect 2225 24596 2237 24599
rect 2004 24568 2237 24596
rect 2004 24556 2010 24568
rect 2225 24565 2237 24568
rect 2271 24565 2283 24599
rect 2225 24559 2283 24565
rect 19061 24599 19119 24605
rect 19061 24565 19073 24599
rect 19107 24596 19119 24599
rect 19904 24596 19932 24636
rect 19107 24568 19932 24596
rect 19981 24599 20039 24605
rect 19107 24565 19119 24568
rect 19061 24559 19119 24565
rect 19981 24565 19993 24599
rect 20027 24596 20039 24599
rect 20254 24596 20260 24608
rect 20027 24568 20260 24596
rect 20027 24565 20039 24568
rect 19981 24559 20039 24565
rect 20254 24556 20260 24568
rect 20312 24556 20318 24608
rect 20901 24599 20959 24605
rect 20901 24565 20913 24599
rect 20947 24596 20959 24599
rect 21450 24596 21456 24608
rect 20947 24568 21456 24596
rect 20947 24565 20959 24568
rect 20901 24559 20959 24565
rect 21450 24556 21456 24568
rect 21508 24556 21514 24608
rect 22554 24596 22560 24608
rect 22515 24568 22560 24596
rect 22554 24556 22560 24568
rect 22612 24556 22618 24608
rect 22646 24556 22652 24608
rect 22704 24596 22710 24608
rect 23382 24596 23388 24608
rect 22704 24568 23388 24596
rect 22704 24556 22710 24568
rect 23382 24556 23388 24568
rect 23440 24556 23446 24608
rect 23566 24556 23572 24608
rect 23624 24596 23630 24608
rect 24670 24596 24676 24608
rect 23624 24568 24676 24596
rect 23624 24556 23630 24568
rect 24670 24556 24676 24568
rect 24728 24556 24734 24608
rect 24780 24596 24808 24636
rect 25884 24636 29500 24664
rect 25884 24596 25912 24636
rect 24780 24568 25912 24596
rect 26329 24599 26387 24605
rect 26329 24565 26341 24599
rect 26375 24596 26387 24599
rect 26602 24596 26608 24608
rect 26375 24568 26608 24596
rect 26375 24565 26387 24568
rect 26329 24559 26387 24565
rect 26602 24556 26608 24568
rect 26660 24596 26666 24608
rect 27246 24596 27252 24608
rect 26660 24568 27252 24596
rect 26660 24556 26666 24568
rect 27246 24556 27252 24568
rect 27304 24556 27310 24608
rect 28261 24599 28319 24605
rect 28261 24565 28273 24599
rect 28307 24596 28319 24599
rect 28350 24596 28356 24608
rect 28307 24568 28356 24596
rect 28307 24565 28319 24568
rect 28261 24559 28319 24565
rect 28350 24556 28356 24568
rect 28408 24556 28414 24608
rect 28445 24599 28503 24605
rect 28445 24565 28457 24599
rect 28491 24596 28503 24599
rect 29362 24596 29368 24608
rect 28491 24568 29368 24596
rect 28491 24565 28503 24568
rect 28445 24559 28503 24565
rect 29362 24556 29368 24568
rect 29420 24556 29426 24608
rect 29472 24596 29500 24636
rect 29638 24624 29644 24676
rect 29696 24624 29702 24676
rect 34624 24673 34652 24704
rect 34698 24692 34704 24744
rect 34756 24732 34762 24744
rect 36262 24732 36268 24744
rect 34756 24704 36268 24732
rect 34756 24692 34762 24704
rect 36262 24692 36268 24704
rect 36320 24732 36326 24744
rect 39485 24735 39543 24741
rect 39485 24732 39497 24735
rect 36320 24704 39497 24732
rect 36320 24692 36326 24704
rect 39485 24701 39497 24704
rect 39531 24701 39543 24735
rect 42092 24732 42120 24772
rect 42426 24760 42432 24772
rect 42484 24760 42490 24812
rect 42685 24803 42743 24809
rect 42685 24800 42697 24803
rect 42536 24772 42697 24800
rect 42536 24732 42564 24772
rect 42685 24769 42697 24772
rect 42731 24769 42743 24803
rect 42812 24800 42840 24908
rect 45186 24800 45192 24812
rect 42812 24772 45192 24800
rect 42685 24763 42743 24769
rect 45186 24760 45192 24772
rect 45244 24760 45250 24812
rect 46845 24803 46903 24809
rect 46845 24769 46857 24803
rect 46891 24800 46903 24803
rect 47486 24800 47492 24812
rect 46891 24772 47492 24800
rect 46891 24769 46903 24772
rect 46845 24763 46903 24769
rect 47486 24760 47492 24772
rect 47544 24760 47550 24812
rect 47854 24800 47860 24812
rect 47815 24772 47860 24800
rect 47854 24760 47860 24772
rect 47912 24760 47918 24812
rect 39485 24695 39543 24701
rect 41386 24704 42120 24732
rect 42444 24704 42564 24732
rect 34609 24667 34667 24673
rect 31128 24636 31754 24664
rect 31128 24596 31156 24636
rect 29472 24568 31156 24596
rect 31202 24556 31208 24608
rect 31260 24596 31266 24608
rect 31386 24596 31392 24608
rect 31260 24568 31392 24596
rect 31260 24556 31266 24568
rect 31386 24556 31392 24568
rect 31444 24596 31450 24608
rect 31573 24599 31631 24605
rect 31573 24596 31585 24599
rect 31444 24568 31585 24596
rect 31444 24556 31450 24568
rect 31573 24565 31585 24568
rect 31619 24565 31631 24599
rect 31726 24596 31754 24636
rect 34609 24633 34621 24667
rect 34655 24633 34667 24667
rect 38286 24664 38292 24676
rect 34609 24627 34667 24633
rect 34716 24636 38292 24664
rect 34716 24596 34744 24636
rect 38286 24624 38292 24636
rect 38344 24624 38350 24676
rect 31726 24568 34744 24596
rect 31573 24559 31631 24565
rect 35342 24556 35348 24608
rect 35400 24596 35406 24608
rect 39390 24596 39396 24608
rect 35400 24568 39396 24596
rect 35400 24556 35406 24568
rect 39390 24556 39396 24568
rect 39448 24556 39454 24608
rect 39500 24596 39528 24695
rect 41386 24664 41414 24704
rect 40420 24636 41414 24664
rect 41693 24667 41751 24673
rect 40420 24596 40448 24636
rect 41693 24633 41705 24667
rect 41739 24664 41751 24667
rect 42444 24664 42472 24704
rect 41739 24636 42472 24664
rect 41739 24633 41751 24636
rect 41693 24627 41751 24633
rect 43438 24624 43444 24676
rect 43496 24664 43502 24676
rect 48041 24667 48099 24673
rect 48041 24664 48053 24667
rect 43496 24636 48053 24664
rect 43496 24624 43502 24636
rect 48041 24633 48053 24636
rect 48087 24633 48099 24667
rect 48041 24627 48099 24633
rect 39500 24568 40448 24596
rect 40865 24599 40923 24605
rect 40865 24565 40877 24599
rect 40911 24596 40923 24599
rect 41138 24596 41144 24608
rect 40911 24568 41144 24596
rect 40911 24565 40923 24568
rect 40865 24559 40923 24565
rect 41138 24556 41144 24568
rect 41196 24556 41202 24608
rect 42334 24556 42340 24608
rect 42392 24596 42398 24608
rect 43809 24599 43867 24605
rect 43809 24596 43821 24599
rect 42392 24568 43821 24596
rect 42392 24556 42398 24568
rect 43809 24565 43821 24568
rect 43855 24565 43867 24599
rect 43809 24559 43867 24565
rect 46474 24556 46480 24608
rect 46532 24596 46538 24608
rect 46937 24599 46995 24605
rect 46937 24596 46949 24599
rect 46532 24568 46949 24596
rect 46532 24556 46538 24568
rect 46937 24565 46949 24568
rect 46983 24565 46995 24599
rect 46937 24559 46995 24565
rect 1104 24506 48852 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 48852 24506
rect 1104 24432 48852 24454
rect 2314 24352 2320 24404
rect 2372 24392 2378 24404
rect 19705 24395 19763 24401
rect 19705 24392 19717 24395
rect 2372 24364 19717 24392
rect 2372 24352 2378 24364
rect 19705 24361 19717 24364
rect 19751 24361 19763 24395
rect 19705 24355 19763 24361
rect 20165 24395 20223 24401
rect 20165 24361 20177 24395
rect 20211 24392 20223 24395
rect 20346 24392 20352 24404
rect 20211 24364 20352 24392
rect 20211 24361 20223 24364
rect 20165 24355 20223 24361
rect 19334 24324 19340 24336
rect 16224 24296 19340 24324
rect 1394 24188 1400 24200
rect 1355 24160 1400 24188
rect 1394 24148 1400 24160
rect 1452 24148 1458 24200
rect 1670 24188 1676 24200
rect 1631 24160 1676 24188
rect 1670 24148 1676 24160
rect 1728 24148 1734 24200
rect 1762 24148 1768 24200
rect 1820 24188 1826 24200
rect 2869 24191 2927 24197
rect 2869 24188 2881 24191
rect 1820 24160 2881 24188
rect 1820 24148 1826 24160
rect 2869 24157 2881 24160
rect 2915 24157 2927 24191
rect 15746 24188 15752 24200
rect 15707 24160 15752 24188
rect 2869 24151 2927 24157
rect 15746 24148 15752 24160
rect 15804 24148 15810 24200
rect 16224 24197 16252 24296
rect 19334 24284 19340 24296
rect 19392 24284 19398 24336
rect 19720 24324 19748 24355
rect 20346 24352 20352 24364
rect 20404 24352 20410 24404
rect 20901 24395 20959 24401
rect 20901 24361 20913 24395
rect 20947 24392 20959 24395
rect 20990 24392 20996 24404
rect 20947 24364 20996 24392
rect 20947 24361 20959 24364
rect 20901 24355 20959 24361
rect 20990 24352 20996 24364
rect 21048 24392 21054 24404
rect 21174 24392 21180 24404
rect 21048 24364 21180 24392
rect 21048 24352 21054 24364
rect 21174 24352 21180 24364
rect 21232 24352 21238 24404
rect 21358 24352 21364 24404
rect 21416 24392 21422 24404
rect 27982 24392 27988 24404
rect 21416 24364 27988 24392
rect 21416 24352 21422 24364
rect 27982 24352 27988 24364
rect 28040 24352 28046 24404
rect 28534 24392 28540 24404
rect 28495 24364 28540 24392
rect 28534 24352 28540 24364
rect 28592 24352 28598 24404
rect 29086 24352 29092 24404
rect 29144 24392 29150 24404
rect 29641 24395 29699 24401
rect 29641 24392 29653 24395
rect 29144 24364 29653 24392
rect 29144 24352 29150 24364
rect 29641 24361 29653 24364
rect 29687 24361 29699 24395
rect 29641 24355 29699 24361
rect 36630 24352 36636 24404
rect 36688 24392 36694 24404
rect 38746 24392 38752 24404
rect 36688 24364 38752 24392
rect 36688 24352 36694 24364
rect 38746 24352 38752 24364
rect 38804 24392 38810 24404
rect 38841 24395 38899 24401
rect 38841 24392 38853 24395
rect 38804 24364 38853 24392
rect 38804 24352 38810 24364
rect 38841 24361 38853 24364
rect 38887 24361 38899 24395
rect 38841 24355 38899 24361
rect 40313 24395 40371 24401
rect 40313 24361 40325 24395
rect 40359 24392 40371 24395
rect 41414 24392 41420 24404
rect 40359 24364 41420 24392
rect 40359 24361 40371 24364
rect 40313 24355 40371 24361
rect 41414 24352 41420 24364
rect 41472 24352 41478 24404
rect 41785 24395 41843 24401
rect 41785 24361 41797 24395
rect 41831 24361 41843 24395
rect 41966 24392 41972 24404
rect 41927 24364 41972 24392
rect 41785 24355 41843 24361
rect 20714 24324 20720 24336
rect 19720 24296 20720 24324
rect 20714 24284 20720 24296
rect 20772 24284 20778 24336
rect 23382 24284 23388 24336
rect 23440 24324 23446 24336
rect 25314 24324 25320 24336
rect 23440 24296 25320 24324
rect 23440 24284 23446 24296
rect 25314 24284 25320 24296
rect 25372 24284 25378 24336
rect 27430 24324 27436 24336
rect 27391 24296 27436 24324
rect 27430 24284 27436 24296
rect 27488 24284 27494 24336
rect 28997 24327 29055 24333
rect 28997 24293 29009 24327
rect 29043 24324 29055 24327
rect 29043 24296 29132 24324
rect 29043 24293 29055 24296
rect 28997 24287 29055 24293
rect 16853 24259 16911 24265
rect 16853 24225 16865 24259
rect 16899 24256 16911 24259
rect 17586 24256 17592 24268
rect 16899 24228 17592 24256
rect 16899 24225 16911 24228
rect 16853 24219 16911 24225
rect 17586 24216 17592 24228
rect 17644 24216 17650 24268
rect 17862 24256 17868 24268
rect 17823 24228 17868 24256
rect 17862 24216 17868 24228
rect 17920 24216 17926 24268
rect 19794 24256 19800 24268
rect 19755 24228 19800 24256
rect 19794 24216 19800 24228
rect 19852 24216 19858 24268
rect 19886 24216 19892 24268
rect 19944 24216 19950 24268
rect 20806 24256 20812 24268
rect 20767 24228 20812 24256
rect 20806 24216 20812 24228
rect 20864 24216 20870 24268
rect 21910 24256 21916 24268
rect 21871 24228 21916 24256
rect 21910 24216 21916 24228
rect 21968 24216 21974 24268
rect 27522 24256 27528 24268
rect 27483 24228 27528 24256
rect 27522 24216 27528 24228
rect 27580 24216 27586 24268
rect 28350 24216 28356 24268
rect 28408 24256 28414 24268
rect 28408 24228 28856 24256
rect 28408 24216 28414 24228
rect 16209 24191 16267 24197
rect 16209 24157 16221 24191
rect 16255 24157 16267 24191
rect 16209 24151 16267 24157
rect 16393 24191 16451 24197
rect 16393 24157 16405 24191
rect 16439 24157 16451 24191
rect 16393 24151 16451 24157
rect 16298 24052 16304 24064
rect 16259 24024 16304 24052
rect 16298 24012 16304 24024
rect 16356 24012 16362 24064
rect 16408 24052 16436 24151
rect 19334 24148 19340 24200
rect 19392 24188 19398 24200
rect 19904 24188 19932 24216
rect 19392 24160 19932 24188
rect 19981 24191 20039 24197
rect 19392 24148 19398 24160
rect 19981 24157 19993 24191
rect 20027 24188 20039 24191
rect 20070 24188 20076 24200
rect 20027 24160 20076 24188
rect 20027 24157 20039 24160
rect 19981 24151 20039 24157
rect 20070 24148 20076 24160
rect 20128 24148 20134 24200
rect 20898 24188 20904 24200
rect 20859 24160 20904 24188
rect 20898 24148 20904 24160
rect 20956 24148 20962 24200
rect 21818 24188 21824 24200
rect 21008 24160 21824 24188
rect 17037 24123 17095 24129
rect 17037 24089 17049 24123
rect 17083 24120 17095 24123
rect 18046 24120 18052 24132
rect 17083 24092 18052 24120
rect 17083 24089 17095 24092
rect 17037 24083 17095 24089
rect 18046 24080 18052 24092
rect 18104 24080 18110 24132
rect 19426 24080 19432 24132
rect 19484 24120 19490 24132
rect 19705 24123 19763 24129
rect 19705 24120 19717 24123
rect 19484 24092 19717 24120
rect 19484 24080 19490 24092
rect 19705 24089 19717 24092
rect 19751 24089 19763 24123
rect 20622 24120 20628 24132
rect 20583 24092 20628 24120
rect 19705 24083 19763 24089
rect 20622 24080 20628 24092
rect 20680 24080 20686 24132
rect 16942 24052 16948 24064
rect 16408 24024 16948 24052
rect 16942 24012 16948 24024
rect 17000 24052 17006 24064
rect 21008 24052 21036 24160
rect 21818 24148 21824 24160
rect 21876 24148 21882 24200
rect 22180 24191 22238 24197
rect 22180 24157 22192 24191
rect 22226 24188 22238 24191
rect 22554 24188 22560 24200
rect 22226 24160 22560 24188
rect 22226 24157 22238 24160
rect 22180 24151 22238 24157
rect 22554 24148 22560 24160
rect 22612 24148 22618 24200
rect 24486 24188 24492 24200
rect 24447 24160 24492 24188
rect 24486 24148 24492 24160
rect 24544 24148 24550 24200
rect 24670 24188 24676 24200
rect 24631 24160 24676 24188
rect 24670 24148 24676 24160
rect 24728 24148 24734 24200
rect 25038 24148 25044 24200
rect 25096 24188 25102 24200
rect 25317 24191 25375 24197
rect 25317 24188 25329 24191
rect 25096 24160 25329 24188
rect 25096 24148 25102 24160
rect 25317 24157 25329 24160
rect 25363 24157 25375 24191
rect 27157 24191 27215 24197
rect 27157 24188 27169 24191
rect 25317 24151 25375 24157
rect 25424 24160 27169 24188
rect 25424 24120 25452 24160
rect 27157 24157 27169 24160
rect 27203 24157 27215 24191
rect 27157 24151 27215 24157
rect 27304 24191 27362 24197
rect 27304 24157 27316 24191
rect 27350 24188 27362 24191
rect 28258 24188 28264 24200
rect 27350 24160 28264 24188
rect 27350 24157 27362 24160
rect 27304 24151 27362 24157
rect 28258 24148 28264 24160
rect 28316 24148 28322 24200
rect 28442 24148 28448 24200
rect 28500 24188 28506 24200
rect 28828 24197 28856 24228
rect 28629 24191 28687 24197
rect 28629 24188 28641 24191
rect 28500 24160 28641 24188
rect 28500 24148 28506 24160
rect 28629 24157 28641 24160
rect 28675 24157 28687 24191
rect 28629 24151 28687 24157
rect 28813 24191 28871 24197
rect 28813 24157 28825 24191
rect 28859 24157 28871 24191
rect 29104 24188 29132 24296
rect 30098 24284 30104 24336
rect 30156 24284 30162 24336
rect 32122 24324 32128 24336
rect 32045 24296 32128 24324
rect 29270 24216 29276 24268
rect 29328 24256 29334 24268
rect 29825 24259 29883 24265
rect 29825 24256 29837 24259
rect 29328 24228 29837 24256
rect 29328 24216 29334 24228
rect 29825 24225 29837 24228
rect 29871 24225 29883 24259
rect 30116 24256 30144 24284
rect 29825 24219 29883 24225
rect 30024 24228 30144 24256
rect 30024 24197 30052 24228
rect 30558 24216 30564 24268
rect 30616 24256 30622 24268
rect 32045 24256 32073 24296
rect 32122 24284 32128 24296
rect 32180 24284 32186 24336
rect 35710 24284 35716 24336
rect 35768 24324 35774 24336
rect 40218 24324 40224 24336
rect 35768 24296 40224 24324
rect 35768 24284 35774 24296
rect 40218 24284 40224 24296
rect 40276 24284 40282 24336
rect 40494 24324 40500 24336
rect 40455 24296 40500 24324
rect 40494 24284 40500 24296
rect 40552 24284 40558 24336
rect 40954 24324 40960 24336
rect 40915 24296 40960 24324
rect 40954 24284 40960 24296
rect 41012 24284 41018 24336
rect 41800 24324 41828 24355
rect 41966 24352 41972 24364
rect 42024 24352 42030 24404
rect 42058 24352 42064 24404
rect 42116 24392 42122 24404
rect 42521 24395 42579 24401
rect 42521 24392 42533 24395
rect 42116 24364 42533 24392
rect 42116 24352 42122 24364
rect 42521 24361 42533 24364
rect 42567 24361 42579 24395
rect 48038 24392 48044 24404
rect 42521 24355 42579 24361
rect 43916 24364 48044 24392
rect 43257 24327 43315 24333
rect 43257 24324 43269 24327
rect 41800 24296 43269 24324
rect 43257 24293 43269 24296
rect 43303 24293 43315 24327
rect 43257 24287 43315 24293
rect 43346 24284 43352 24336
rect 43404 24324 43410 24336
rect 43916 24324 43944 24364
rect 48038 24352 48044 24364
rect 48096 24352 48102 24404
rect 47762 24324 47768 24336
rect 43404 24296 43944 24324
rect 46308 24296 47768 24324
rect 43404 24284 43410 24296
rect 30616 24228 32073 24256
rect 30616 24216 30622 24228
rect 32045 24197 32073 24228
rect 32674 24216 32680 24268
rect 32732 24256 32738 24268
rect 32769 24259 32827 24265
rect 32769 24256 32781 24259
rect 32732 24228 32781 24256
rect 32732 24216 32738 24228
rect 32769 24225 32781 24228
rect 32815 24225 32827 24259
rect 34698 24256 34704 24268
rect 34659 24228 34704 24256
rect 32769 24219 32827 24225
rect 34698 24216 34704 24228
rect 34756 24216 34762 24268
rect 40862 24256 40868 24268
rect 35728 24228 40868 24256
rect 28813 24151 28871 24157
rect 29012 24160 29132 24188
rect 30009 24191 30067 24197
rect 25590 24129 25596 24132
rect 25584 24120 25596 24129
rect 21100 24092 25452 24120
rect 25551 24092 25596 24120
rect 21100 24061 21128 24092
rect 25584 24083 25596 24092
rect 25590 24080 25596 24083
rect 25648 24080 25654 24132
rect 27522 24120 27528 24132
rect 26620 24092 27528 24120
rect 17000 24024 21036 24052
rect 21085 24055 21143 24061
rect 17000 24012 17006 24024
rect 21085 24021 21097 24055
rect 21131 24021 21143 24055
rect 21085 24015 21143 24021
rect 23014 24012 23020 24064
rect 23072 24052 23078 24064
rect 23293 24055 23351 24061
rect 23293 24052 23305 24055
rect 23072 24024 23305 24052
rect 23072 24012 23078 24024
rect 23293 24021 23305 24024
rect 23339 24052 23351 24055
rect 24302 24052 24308 24064
rect 23339 24024 24308 24052
rect 23339 24021 23351 24024
rect 23293 24015 23351 24021
rect 24302 24012 24308 24024
rect 24360 24012 24366 24064
rect 24673 24055 24731 24061
rect 24673 24021 24685 24055
rect 24719 24052 24731 24055
rect 25130 24052 25136 24064
rect 24719 24024 25136 24052
rect 24719 24021 24731 24024
rect 24673 24015 24731 24021
rect 25130 24012 25136 24024
rect 25188 24012 25194 24064
rect 25314 24012 25320 24064
rect 25372 24052 25378 24064
rect 26620 24052 26648 24092
rect 27522 24080 27528 24092
rect 27580 24080 27586 24132
rect 28074 24080 28080 24132
rect 28132 24120 28138 24132
rect 28353 24123 28411 24129
rect 28353 24120 28365 24123
rect 28132 24092 28365 24120
rect 28132 24080 28138 24092
rect 28353 24089 28365 24092
rect 28399 24089 28411 24123
rect 28353 24083 28411 24089
rect 25372 24024 26648 24052
rect 26697 24055 26755 24061
rect 25372 24012 25378 24024
rect 26697 24021 26709 24055
rect 26743 24052 26755 24055
rect 26878 24052 26884 24064
rect 26743 24024 26884 24052
rect 26743 24021 26755 24024
rect 26697 24015 26755 24021
rect 26878 24012 26884 24024
rect 26936 24012 26942 24064
rect 27706 24012 27712 24064
rect 27764 24052 27770 24064
rect 27801 24055 27859 24061
rect 27801 24052 27813 24055
rect 27764 24024 27813 24052
rect 27764 24012 27770 24024
rect 27801 24021 27813 24024
rect 27847 24021 27859 24055
rect 29012 24052 29040 24160
rect 30009 24157 30021 24191
rect 30055 24157 30067 24191
rect 30009 24151 30067 24157
rect 31941 24191 31999 24197
rect 31941 24157 31953 24191
rect 31987 24157 31999 24191
rect 31941 24151 31999 24157
rect 32030 24191 32088 24197
rect 32030 24157 32042 24191
rect 32076 24157 32088 24191
rect 32030 24151 32088 24157
rect 32125 24191 32183 24197
rect 32125 24157 32137 24191
rect 32171 24157 32183 24191
rect 32125 24151 32183 24157
rect 29086 24080 29092 24132
rect 29144 24120 29150 24132
rect 29546 24120 29552 24132
rect 29144 24092 29552 24120
rect 29144 24080 29150 24092
rect 29546 24080 29552 24092
rect 29604 24080 29610 24132
rect 30834 24120 30840 24132
rect 30795 24092 30840 24120
rect 30834 24080 30840 24092
rect 30892 24080 30898 24132
rect 30926 24080 30932 24132
rect 30984 24120 30990 24132
rect 31021 24123 31079 24129
rect 31021 24120 31033 24123
rect 30984 24092 31033 24120
rect 30984 24080 30990 24092
rect 31021 24089 31033 24092
rect 31067 24089 31079 24123
rect 31662 24120 31668 24132
rect 31623 24092 31668 24120
rect 31021 24083 31079 24089
rect 31662 24080 31668 24092
rect 31720 24080 31726 24132
rect 31846 24080 31852 24132
rect 31904 24120 31910 24132
rect 31956 24120 31984 24151
rect 31904 24092 31984 24120
rect 31904 24080 31910 24092
rect 29270 24052 29276 24064
rect 29012 24024 29276 24052
rect 27801 24015 27859 24021
rect 29270 24012 29276 24024
rect 29328 24012 29334 24064
rect 30193 24055 30251 24061
rect 30193 24021 30205 24055
rect 30239 24052 30251 24055
rect 30466 24052 30472 24064
rect 30239 24024 30472 24052
rect 30239 24021 30251 24024
rect 30193 24015 30251 24021
rect 30466 24012 30472 24024
rect 30524 24012 30530 24064
rect 31205 24055 31263 24061
rect 31205 24021 31217 24055
rect 31251 24052 31263 24055
rect 32140 24052 32168 24151
rect 32214 24148 32220 24200
rect 32272 24188 32278 24200
rect 32309 24191 32367 24197
rect 32309 24188 32321 24191
rect 32272 24160 32321 24188
rect 32272 24148 32278 24160
rect 32309 24157 32321 24160
rect 32355 24157 32367 24191
rect 32309 24151 32367 24157
rect 34790 24148 34796 24200
rect 34848 24188 34854 24200
rect 34957 24191 35015 24197
rect 34957 24188 34969 24191
rect 34848 24160 34969 24188
rect 34848 24148 34854 24160
rect 34957 24157 34969 24160
rect 35003 24157 35015 24191
rect 34957 24151 35015 24157
rect 35434 24148 35440 24200
rect 35492 24188 35498 24200
rect 35728 24188 35756 24228
rect 40862 24216 40868 24228
rect 40920 24216 40926 24268
rect 41046 24216 41052 24268
rect 41104 24256 41110 24268
rect 42150 24256 42156 24268
rect 41104 24228 42156 24256
rect 41104 24216 41110 24228
rect 42150 24216 42156 24228
rect 42208 24216 42214 24268
rect 46308 24265 46336 24296
rect 47762 24284 47768 24296
rect 47820 24284 47826 24336
rect 46293 24259 46351 24265
rect 42536 24228 43392 24256
rect 35492 24160 35756 24188
rect 37093 24191 37151 24197
rect 35492 24148 35498 24160
rect 37093 24157 37105 24191
rect 37139 24188 37151 24191
rect 37366 24188 37372 24200
rect 37139 24160 37372 24188
rect 37139 24157 37151 24160
rect 37093 24151 37151 24157
rect 37366 24148 37372 24160
rect 37424 24188 37430 24200
rect 37642 24188 37648 24200
rect 37424 24160 37648 24188
rect 37424 24148 37430 24160
rect 37642 24148 37648 24160
rect 37700 24148 37706 24200
rect 38102 24188 38108 24200
rect 38063 24160 38108 24188
rect 38102 24148 38108 24160
rect 38160 24148 38166 24200
rect 38749 24191 38807 24197
rect 38749 24157 38761 24191
rect 38795 24188 38807 24191
rect 39758 24188 39764 24200
rect 38795 24160 39764 24188
rect 38795 24157 38807 24160
rect 38749 24151 38807 24157
rect 39758 24148 39764 24160
rect 39816 24148 39822 24200
rect 39850 24148 39856 24200
rect 39908 24188 39914 24200
rect 39945 24191 40003 24197
rect 39945 24188 39957 24191
rect 39908 24160 39957 24188
rect 39908 24148 39914 24160
rect 39945 24157 39957 24160
rect 39991 24157 40003 24191
rect 41138 24188 41144 24200
rect 41099 24160 41144 24188
rect 39945 24151 40003 24157
rect 41138 24148 41144 24160
rect 41196 24148 41202 24200
rect 42536 24188 42564 24228
rect 43364 24200 43392 24228
rect 46293 24225 46305 24259
rect 46339 24225 46351 24259
rect 46474 24256 46480 24268
rect 46435 24228 46480 24256
rect 46293 24219 46351 24225
rect 46474 24216 46480 24228
rect 46532 24216 46538 24268
rect 48130 24256 48136 24268
rect 48091 24228 48136 24256
rect 48130 24216 48136 24228
rect 48188 24216 48194 24268
rect 42593 24191 42651 24197
rect 42593 24188 42605 24191
rect 42536 24160 42605 24188
rect 42593 24157 42605 24160
rect 42639 24157 42651 24191
rect 42593 24151 42651 24157
rect 42717 24169 42775 24175
rect 42717 24135 42729 24169
rect 42763 24166 42775 24169
rect 42886 24166 42892 24200
rect 42763 24148 42892 24166
rect 42944 24148 42950 24200
rect 43162 24188 43168 24200
rect 43123 24160 43168 24188
rect 43162 24148 43168 24160
rect 43220 24148 43226 24200
rect 43346 24188 43352 24200
rect 43307 24160 43352 24188
rect 43346 24148 43352 24160
rect 43404 24148 43410 24200
rect 43438 24148 43444 24200
rect 43496 24188 43502 24200
rect 43993 24191 44051 24197
rect 43993 24188 44005 24191
rect 43496 24160 44005 24188
rect 43496 24148 43502 24160
rect 43993 24157 44005 24160
rect 44039 24157 44051 24191
rect 43993 24151 44051 24157
rect 42763 24138 42932 24148
rect 42763 24135 42775 24138
rect 32858 24080 32864 24132
rect 32916 24120 32922 24132
rect 33014 24123 33072 24129
rect 33014 24120 33026 24123
rect 32916 24092 33026 24120
rect 32916 24080 32922 24092
rect 33014 24089 33026 24092
rect 33060 24089 33072 24123
rect 33014 24083 33072 24089
rect 38289 24123 38347 24129
rect 38289 24089 38301 24123
rect 38335 24120 38347 24123
rect 40586 24120 40592 24132
rect 38335 24092 40592 24120
rect 38335 24089 38347 24092
rect 38289 24083 38347 24089
rect 40586 24080 40592 24092
rect 40644 24080 40650 24132
rect 41414 24080 41420 24132
rect 41472 24120 41478 24132
rect 41601 24123 41659 24129
rect 41601 24120 41613 24123
rect 41472 24092 41613 24120
rect 41472 24080 41478 24092
rect 41601 24089 41613 24092
rect 41647 24089 41659 24123
rect 41601 24083 41659 24089
rect 42242 24080 42248 24132
rect 42300 24120 42306 24132
rect 42717 24129 42775 24135
rect 42429 24123 42487 24129
rect 42429 24120 42441 24123
rect 42300 24092 42441 24120
rect 42300 24080 42306 24092
rect 42429 24089 42441 24092
rect 42475 24089 42487 24123
rect 47670 24120 47676 24132
rect 42429 24083 42487 24089
rect 43456 24092 47676 24120
rect 31251 24024 32168 24052
rect 34149 24055 34207 24061
rect 31251 24021 31263 24024
rect 31205 24015 31263 24021
rect 34149 24021 34161 24055
rect 34195 24052 34207 24055
rect 34790 24052 34796 24064
rect 34195 24024 34796 24052
rect 34195 24021 34207 24024
rect 34149 24015 34207 24021
rect 34790 24012 34796 24024
rect 34848 24012 34854 24064
rect 36078 24052 36084 24064
rect 36039 24024 36084 24052
rect 36078 24012 36084 24024
rect 36136 24012 36142 24064
rect 37274 24052 37280 24064
rect 37187 24024 37280 24052
rect 37274 24012 37280 24024
rect 37332 24052 37338 24064
rect 37918 24052 37924 24064
rect 37332 24024 37924 24052
rect 37332 24012 37338 24024
rect 37918 24012 37924 24024
rect 37976 24012 37982 24064
rect 38838 24012 38844 24064
rect 38896 24052 38902 24064
rect 39209 24055 39267 24061
rect 39209 24052 39221 24055
rect 38896 24024 39221 24052
rect 38896 24012 38902 24024
rect 39209 24021 39221 24024
rect 39255 24021 39267 24055
rect 39209 24015 39267 24021
rect 39666 24012 39672 24064
rect 39724 24052 39730 24064
rect 40313 24055 40371 24061
rect 40313 24052 40325 24055
rect 39724 24024 40325 24052
rect 39724 24012 39730 24024
rect 40313 24021 40325 24024
rect 40359 24021 40371 24055
rect 40313 24015 40371 24021
rect 41782 24012 41788 24064
rect 41840 24061 41846 24064
rect 41840 24055 41859 24061
rect 41847 24021 41859 24055
rect 41840 24015 41859 24021
rect 41840 24012 41846 24015
rect 43254 24012 43260 24064
rect 43312 24052 43318 24064
rect 43456 24052 43484 24092
rect 47670 24080 47676 24092
rect 47728 24080 47734 24132
rect 43806 24052 43812 24064
rect 43312 24024 43484 24052
rect 43767 24024 43812 24052
rect 43312 24012 43318 24024
rect 43806 24012 43812 24024
rect 43864 24012 43870 24064
rect 1104 23962 48852 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 48852 23962
rect 1104 23888 48852 23910
rect 15562 23808 15568 23860
rect 15620 23848 15626 23860
rect 15620 23820 16068 23848
rect 15620 23808 15626 23820
rect 16040 23792 16068 23820
rect 17310 23808 17316 23860
rect 17368 23848 17374 23860
rect 20898 23848 20904 23860
rect 17368 23820 20904 23848
rect 17368 23808 17374 23820
rect 20898 23808 20904 23820
rect 20956 23808 20962 23860
rect 21082 23848 21088 23860
rect 21043 23820 21088 23848
rect 21082 23808 21088 23820
rect 21140 23808 21146 23860
rect 24949 23851 25007 23857
rect 24949 23817 24961 23851
rect 24995 23848 25007 23851
rect 25222 23848 25228 23860
rect 24995 23820 25228 23848
rect 24995 23817 25007 23820
rect 24949 23811 25007 23817
rect 25222 23808 25228 23820
rect 25280 23808 25286 23860
rect 26234 23848 26240 23860
rect 25608 23820 26240 23848
rect 1946 23780 1952 23792
rect 1907 23752 1952 23780
rect 1946 23740 1952 23752
rect 2004 23740 2010 23792
rect 15930 23780 15936 23792
rect 15891 23752 15936 23780
rect 15930 23740 15936 23752
rect 15988 23740 15994 23792
rect 16022 23740 16028 23792
rect 16080 23780 16086 23792
rect 19705 23783 19763 23789
rect 16080 23752 18368 23780
rect 16080 23740 16086 23752
rect 1762 23712 1768 23724
rect 1723 23684 1768 23712
rect 1762 23672 1768 23684
rect 1820 23672 1826 23724
rect 15654 23712 15660 23724
rect 15567 23684 15660 23712
rect 15654 23672 15660 23684
rect 15712 23672 15718 23724
rect 15746 23672 15752 23724
rect 15804 23712 15810 23724
rect 16945 23715 17003 23721
rect 16945 23712 16957 23715
rect 15804 23684 16957 23712
rect 15804 23672 15810 23684
rect 16945 23681 16957 23684
rect 16991 23681 17003 23715
rect 18340 23712 18368 23752
rect 19705 23749 19717 23783
rect 19751 23780 19763 23783
rect 20346 23780 20352 23792
rect 19751 23752 20352 23780
rect 19751 23749 19763 23752
rect 19705 23743 19763 23749
rect 20346 23740 20352 23752
rect 20404 23740 20410 23792
rect 25130 23740 25136 23792
rect 25188 23780 25194 23792
rect 25188 23752 25452 23780
rect 25188 23740 25194 23752
rect 19886 23712 19892 23724
rect 18340 23684 19892 23712
rect 16945 23675 17003 23681
rect 19886 23672 19892 23684
rect 19944 23672 19950 23724
rect 19981 23715 20039 23721
rect 19981 23681 19993 23715
rect 20027 23681 20039 23715
rect 19981 23675 20039 23681
rect 1486 23604 1492 23656
rect 1544 23644 1550 23656
rect 1946 23644 1952 23656
rect 1544 23616 1952 23644
rect 1544 23604 1550 23616
rect 1946 23604 1952 23616
rect 2004 23604 2010 23656
rect 2774 23644 2780 23656
rect 2735 23616 2780 23644
rect 2774 23604 2780 23616
rect 2832 23604 2838 23656
rect 15672 23644 15700 23672
rect 16482 23644 16488 23656
rect 15672 23616 16488 23644
rect 16482 23604 16488 23616
rect 16540 23604 16546 23656
rect 17126 23644 17132 23656
rect 17087 23616 17132 23644
rect 17126 23604 17132 23616
rect 17184 23604 17190 23656
rect 17494 23644 17500 23656
rect 17455 23616 17500 23644
rect 17494 23604 17500 23616
rect 17552 23604 17558 23656
rect 19334 23604 19340 23656
rect 19392 23644 19398 23656
rect 19392 23616 19656 23644
rect 19392 23604 19398 23616
rect 1670 23536 1676 23588
rect 1728 23576 1734 23588
rect 19426 23576 19432 23588
rect 1728 23548 19432 23576
rect 1728 23536 1734 23548
rect 19426 23536 19432 23548
rect 19484 23536 19490 23588
rect 19628 23576 19656 23616
rect 19702 23604 19708 23656
rect 19760 23644 19766 23656
rect 19797 23647 19855 23653
rect 19797 23644 19809 23647
rect 19760 23616 19809 23644
rect 19760 23604 19766 23616
rect 19797 23613 19809 23616
rect 19843 23613 19855 23647
rect 19996 23644 20024 23675
rect 20254 23672 20260 23724
rect 20312 23712 20318 23724
rect 20625 23715 20683 23721
rect 20625 23712 20637 23715
rect 20312 23684 20637 23712
rect 20312 23672 20318 23684
rect 20625 23681 20637 23684
rect 20671 23681 20683 23715
rect 20625 23675 20683 23681
rect 20714 23672 20720 23724
rect 20772 23712 20778 23724
rect 20809 23715 20867 23721
rect 20809 23712 20821 23715
rect 20772 23684 20821 23712
rect 20772 23672 20778 23684
rect 20809 23681 20821 23684
rect 20855 23681 20867 23715
rect 20809 23675 20867 23681
rect 20901 23715 20959 23721
rect 20901 23681 20913 23715
rect 20947 23712 20959 23715
rect 20990 23712 20996 23724
rect 20947 23684 20996 23712
rect 20947 23681 20959 23684
rect 20901 23675 20959 23681
rect 20990 23672 20996 23684
rect 21048 23672 21054 23724
rect 21910 23672 21916 23724
rect 21968 23712 21974 23724
rect 22373 23715 22431 23721
rect 22373 23712 22385 23715
rect 21968 23684 22385 23712
rect 21968 23672 21974 23684
rect 22373 23681 22385 23684
rect 22419 23681 22431 23715
rect 22373 23675 22431 23681
rect 22640 23715 22698 23721
rect 22640 23681 22652 23715
rect 22686 23712 22698 23715
rect 23198 23712 23204 23724
rect 22686 23684 23204 23712
rect 22686 23681 22698 23684
rect 22640 23675 22698 23681
rect 23198 23672 23204 23684
rect 23256 23672 23262 23724
rect 24302 23712 24308 23724
rect 24263 23684 24308 23712
rect 24302 23672 24308 23684
rect 24360 23672 24366 23724
rect 24489 23715 24547 23721
rect 24489 23681 24501 23715
rect 24535 23712 24547 23715
rect 24670 23712 24676 23724
rect 24535 23684 24676 23712
rect 24535 23681 24547 23684
rect 24489 23675 24547 23681
rect 19797 23607 19855 23613
rect 19904 23616 20024 23644
rect 19904 23576 19932 23616
rect 23474 23604 23480 23656
rect 23532 23644 23538 23656
rect 24504 23644 24532 23675
rect 24670 23672 24676 23684
rect 24728 23672 24734 23724
rect 25222 23712 25228 23724
rect 25183 23684 25228 23712
rect 25222 23672 25228 23684
rect 25280 23672 25286 23724
rect 25424 23721 25452 23752
rect 25608 23721 25636 23820
rect 26234 23808 26240 23820
rect 26292 23808 26298 23860
rect 26418 23848 26424 23860
rect 26379 23820 26424 23848
rect 26418 23808 26424 23820
rect 26476 23808 26482 23860
rect 28074 23808 28080 23860
rect 28132 23848 28138 23860
rect 28994 23848 29000 23860
rect 28132 23820 29000 23848
rect 28132 23808 28138 23820
rect 28994 23808 29000 23820
rect 29052 23808 29058 23860
rect 29089 23851 29147 23857
rect 29089 23817 29101 23851
rect 29135 23848 29147 23851
rect 33137 23851 33195 23857
rect 29135 23820 32996 23848
rect 29135 23817 29147 23820
rect 29089 23811 29147 23817
rect 25774 23740 25780 23792
rect 25832 23780 25838 23792
rect 30006 23780 30012 23792
rect 25832 23752 29040 23780
rect 25832 23740 25838 23752
rect 25314 23715 25372 23721
rect 25314 23681 25326 23715
rect 25360 23681 25372 23715
rect 25424 23715 25488 23721
rect 25424 23684 25442 23715
rect 25314 23675 25372 23681
rect 25430 23681 25442 23684
rect 25476 23681 25488 23715
rect 25430 23675 25488 23681
rect 25593 23715 25651 23721
rect 25593 23681 25605 23715
rect 25639 23681 25651 23715
rect 26050 23712 26056 23724
rect 26011 23684 26056 23712
rect 25593 23675 25651 23681
rect 23532 23616 24532 23644
rect 25323 23644 25351 23675
rect 26050 23672 26056 23684
rect 26108 23672 26114 23724
rect 26237 23715 26295 23721
rect 26237 23681 26249 23715
rect 26283 23712 26295 23715
rect 26878 23712 26884 23724
rect 26283 23684 26884 23712
rect 26283 23681 26295 23684
rect 26237 23675 26295 23681
rect 26878 23672 26884 23684
rect 26936 23672 26942 23724
rect 28166 23712 28172 23724
rect 28127 23684 28172 23712
rect 28166 23672 28172 23684
rect 28224 23672 28230 23724
rect 28534 23712 28540 23724
rect 28495 23684 28540 23712
rect 28534 23672 28540 23684
rect 28592 23672 28598 23724
rect 29012 23712 29040 23752
rect 29288 23752 30012 23780
rect 29288 23712 29316 23752
rect 30006 23740 30012 23752
rect 30064 23740 30070 23792
rect 29012 23684 29316 23712
rect 29362 23672 29368 23724
rect 29420 23712 29426 23724
rect 29420 23684 29465 23712
rect 29420 23672 29426 23684
rect 29546 23672 29552 23724
rect 29604 23712 29610 23724
rect 30116 23712 30144 23820
rect 31662 23740 31668 23792
rect 31720 23780 31726 23792
rect 32858 23780 32864 23792
rect 31720 23752 32864 23780
rect 31720 23740 31726 23752
rect 32858 23740 32864 23752
rect 32916 23740 32922 23792
rect 32968 23780 32996 23820
rect 33137 23817 33149 23851
rect 33183 23848 33195 23851
rect 33594 23848 33600 23860
rect 33183 23820 33600 23848
rect 33183 23817 33195 23820
rect 33137 23811 33195 23817
rect 33594 23808 33600 23820
rect 33652 23808 33658 23860
rect 35802 23848 35808 23860
rect 33704 23820 35808 23848
rect 33704 23780 33732 23820
rect 35802 23808 35808 23820
rect 35860 23808 35866 23860
rect 36633 23851 36691 23857
rect 36633 23817 36645 23851
rect 36679 23848 36691 23851
rect 38838 23848 38844 23860
rect 36679 23820 37504 23848
rect 38799 23820 38844 23848
rect 36679 23817 36691 23820
rect 36633 23811 36691 23817
rect 35710 23780 35716 23792
rect 32968 23752 33732 23780
rect 35623 23752 35716 23780
rect 35710 23740 35716 23752
rect 35768 23780 35774 23792
rect 36078 23780 36084 23792
rect 35768 23752 36084 23780
rect 35768 23740 35774 23752
rect 36078 23740 36084 23752
rect 36136 23740 36142 23792
rect 37274 23740 37280 23792
rect 37332 23780 37338 23792
rect 37476 23789 37504 23820
rect 38838 23808 38844 23820
rect 38896 23808 38902 23860
rect 38933 23851 38991 23857
rect 38933 23817 38945 23851
rect 38979 23848 38991 23851
rect 40129 23851 40187 23857
rect 40129 23848 40141 23851
rect 38979 23820 40141 23848
rect 38979 23817 38991 23820
rect 38933 23811 38991 23817
rect 40129 23817 40141 23820
rect 40175 23817 40187 23851
rect 40129 23811 40187 23817
rect 40862 23808 40868 23860
rect 40920 23848 40926 23860
rect 40957 23851 41015 23857
rect 40957 23848 40969 23851
rect 40920 23820 40969 23848
rect 40920 23808 40926 23820
rect 40957 23817 40969 23820
rect 41003 23817 41015 23851
rect 40957 23811 41015 23817
rect 41386 23820 42472 23848
rect 37476 23783 37551 23789
rect 37332 23752 37377 23780
rect 37476 23752 37505 23783
rect 37332 23740 37338 23752
rect 37493 23749 37505 23752
rect 37539 23780 37551 23783
rect 38378 23780 38384 23792
rect 37539 23752 38384 23780
rect 37539 23749 37551 23752
rect 37493 23743 37551 23749
rect 38378 23740 38384 23752
rect 38436 23740 38442 23792
rect 41386 23780 41414 23820
rect 38488 23752 41414 23780
rect 41601 23783 41659 23789
rect 30282 23712 30288 23724
rect 29604 23684 30144 23712
rect 30243 23684 30288 23712
rect 29604 23672 29610 23684
rect 30282 23672 30288 23684
rect 30340 23672 30346 23724
rect 32398 23672 32404 23724
rect 32456 23712 32462 23724
rect 32769 23715 32827 23721
rect 32456 23710 32720 23712
rect 32769 23710 32781 23715
rect 32456 23684 32781 23710
rect 32456 23672 32462 23684
rect 32692 23682 32781 23684
rect 32769 23681 32781 23682
rect 32815 23681 32827 23715
rect 32769 23675 32827 23681
rect 32953 23715 33011 23721
rect 32953 23681 32965 23715
rect 32999 23712 33011 23715
rect 33042 23712 33048 23724
rect 32999 23684 33048 23712
rect 32999 23681 33011 23684
rect 32953 23675 33011 23681
rect 33042 23672 33048 23684
rect 33100 23672 33106 23724
rect 35897 23715 35955 23721
rect 35897 23681 35909 23715
rect 35943 23712 35955 23715
rect 35986 23712 35992 23724
rect 35943 23684 35992 23712
rect 35943 23681 35955 23684
rect 35897 23675 35955 23681
rect 35986 23672 35992 23684
rect 36044 23712 36050 23724
rect 36357 23715 36415 23721
rect 36357 23712 36369 23715
rect 36044 23684 36369 23712
rect 36044 23672 36050 23684
rect 36357 23681 36369 23684
rect 36403 23681 36415 23715
rect 38488 23712 38516 23752
rect 41601 23749 41613 23783
rect 41647 23780 41659 23783
rect 42334 23780 42340 23792
rect 41647 23752 42340 23780
rect 41647 23749 41659 23752
rect 41601 23743 41659 23749
rect 42334 23740 42340 23752
rect 42392 23740 42398 23792
rect 42444 23780 42472 23820
rect 42518 23808 42524 23860
rect 42576 23848 42582 23860
rect 48041 23851 48099 23857
rect 48041 23848 48053 23851
rect 42576 23820 48053 23848
rect 42576 23808 42582 23820
rect 48041 23817 48053 23820
rect 48087 23817 48099 23851
rect 48041 23811 48099 23817
rect 42978 23780 42984 23792
rect 42444 23752 42984 23780
rect 42978 23740 42984 23752
rect 43036 23740 43042 23792
rect 43156 23783 43214 23789
rect 43156 23749 43168 23783
rect 43202 23780 43214 23783
rect 43806 23780 43812 23792
rect 43202 23752 43812 23780
rect 43202 23749 43214 23752
rect 43156 23743 43214 23749
rect 43806 23740 43812 23752
rect 43864 23740 43870 23792
rect 47946 23780 47952 23792
rect 47907 23752 47952 23780
rect 47946 23740 47952 23752
rect 48004 23740 48010 23792
rect 36357 23675 36415 23681
rect 36464 23684 38516 23712
rect 27154 23644 27160 23656
rect 25323 23616 27160 23644
rect 23532 23604 23538 23616
rect 27154 23604 27160 23616
rect 27212 23604 27218 23656
rect 28074 23644 28080 23656
rect 28035 23616 28080 23644
rect 28074 23604 28080 23616
rect 28132 23604 28138 23656
rect 28994 23644 29000 23656
rect 28184 23616 29000 23644
rect 19628 23548 19932 23576
rect 20165 23579 20223 23585
rect 20165 23545 20177 23579
rect 20211 23576 20223 23579
rect 21450 23576 21456 23588
rect 20211 23548 21456 23576
rect 20211 23545 20223 23548
rect 20165 23539 20223 23545
rect 21450 23536 21456 23548
rect 21508 23536 21514 23588
rect 28184 23576 28212 23616
rect 28994 23604 29000 23616
rect 29052 23604 29058 23656
rect 29086 23604 29092 23656
rect 29144 23644 29150 23656
rect 36464 23644 36492 23684
rect 38562 23672 38568 23724
rect 38620 23712 38626 23724
rect 39666 23712 39672 23724
rect 38620 23684 39252 23712
rect 39627 23684 39672 23712
rect 38620 23672 38626 23684
rect 29144 23616 36492 23644
rect 29144 23604 29150 23616
rect 36538 23604 36544 23656
rect 36596 23644 36602 23656
rect 36633 23647 36691 23653
rect 36633 23644 36645 23647
rect 36596 23616 36645 23644
rect 36596 23604 36602 23616
rect 36633 23613 36645 23616
rect 36679 23613 36691 23647
rect 36633 23607 36691 23613
rect 39022 23604 39028 23656
rect 39080 23644 39086 23656
rect 39224 23644 39252 23684
rect 39666 23672 39672 23684
rect 39724 23672 39730 23724
rect 40402 23712 40408 23724
rect 39776 23684 40408 23712
rect 39776 23644 39804 23684
rect 40402 23672 40408 23684
rect 40460 23672 40466 23724
rect 40586 23712 40592 23724
rect 40547 23684 40592 23712
rect 40586 23672 40592 23684
rect 40644 23672 40650 23724
rect 40773 23715 40831 23721
rect 40773 23681 40785 23715
rect 40819 23681 40831 23715
rect 40773 23675 40831 23681
rect 39080 23616 39125 23644
rect 39224 23616 39804 23644
rect 39080 23604 39086 23616
rect 39850 23604 39856 23656
rect 39908 23644 39914 23656
rect 40788 23644 40816 23675
rect 40862 23672 40868 23724
rect 40920 23712 40926 23724
rect 41417 23715 41475 23721
rect 41417 23712 41429 23715
rect 40920 23684 41429 23712
rect 40920 23672 40926 23684
rect 41417 23681 41429 23684
rect 41463 23681 41475 23715
rect 44450 23712 44456 23724
rect 41417 23675 41475 23681
rect 41708 23684 44456 23712
rect 40954 23644 40960 23656
rect 39908 23616 40960 23644
rect 39908 23604 39914 23616
rect 40954 23604 40960 23616
rect 41012 23604 41018 23656
rect 41506 23604 41512 23656
rect 41564 23644 41570 23656
rect 41708 23644 41736 23684
rect 44450 23672 44456 23684
rect 44508 23672 44514 23724
rect 41564 23616 41736 23644
rect 41564 23604 41570 23616
rect 41782 23604 41788 23656
rect 41840 23644 41846 23656
rect 41840 23616 41885 23644
rect 41840 23604 41846 23616
rect 42426 23604 42432 23656
rect 42484 23644 42490 23656
rect 42889 23647 42947 23653
rect 42889 23644 42901 23647
rect 42484 23616 42901 23644
rect 42484 23604 42490 23616
rect 42889 23613 42901 23616
rect 42935 23613 42947 23647
rect 42889 23607 42947 23613
rect 23308 23548 28212 23576
rect 28721 23579 28779 23585
rect 1486 23468 1492 23520
rect 1544 23508 1550 23520
rect 1854 23508 1860 23520
rect 1544 23480 1860 23508
rect 1544 23468 1550 23480
rect 1854 23468 1860 23480
rect 1912 23468 1918 23520
rect 3510 23468 3516 23520
rect 3568 23508 3574 23520
rect 17862 23508 17868 23520
rect 3568 23480 17868 23508
rect 3568 23468 3574 23480
rect 17862 23468 17868 23480
rect 17920 23468 17926 23520
rect 19886 23508 19892 23520
rect 19847 23480 19892 23508
rect 19886 23468 19892 23480
rect 19944 23468 19950 23520
rect 20070 23468 20076 23520
rect 20128 23508 20134 23520
rect 20901 23511 20959 23517
rect 20901 23508 20913 23511
rect 20128 23480 20913 23508
rect 20128 23468 20134 23480
rect 20901 23477 20913 23480
rect 20947 23508 20959 23511
rect 23308 23508 23336 23548
rect 28721 23545 28733 23579
rect 28767 23576 28779 23579
rect 29730 23576 29736 23588
rect 28767 23548 29408 23576
rect 29691 23548 29736 23576
rect 28767 23545 28779 23548
rect 28721 23539 28779 23545
rect 20947 23480 23336 23508
rect 20947 23477 20959 23480
rect 20901 23471 20959 23477
rect 23750 23468 23756 23520
rect 23808 23508 23814 23520
rect 24394 23508 24400 23520
rect 23808 23480 23853 23508
rect 24355 23480 24400 23508
rect 23808 23468 23814 23480
rect 24394 23468 24400 23480
rect 24452 23468 24458 23520
rect 28442 23508 28448 23520
rect 28403 23480 28448 23508
rect 28442 23468 28448 23480
rect 28500 23468 28506 23520
rect 29380 23517 29408 23548
rect 29730 23536 29736 23548
rect 29788 23536 29794 23588
rect 30006 23536 30012 23588
rect 30064 23576 30070 23588
rect 42794 23576 42800 23588
rect 30064 23548 42800 23576
rect 30064 23536 30070 23548
rect 42794 23536 42800 23548
rect 42852 23536 42858 23588
rect 29365 23511 29423 23517
rect 29365 23477 29377 23511
rect 29411 23477 29423 23511
rect 29365 23471 29423 23477
rect 30098 23468 30104 23520
rect 30156 23508 30162 23520
rect 30377 23511 30435 23517
rect 30377 23508 30389 23511
rect 30156 23480 30389 23508
rect 30156 23468 30162 23480
rect 30377 23477 30389 23480
rect 30423 23508 30435 23511
rect 30558 23508 30564 23520
rect 30423 23480 30564 23508
rect 30423 23477 30435 23480
rect 30377 23471 30435 23477
rect 30558 23468 30564 23480
rect 30616 23468 30622 23520
rect 36446 23508 36452 23520
rect 36407 23480 36452 23508
rect 36446 23468 36452 23480
rect 36504 23468 36510 23520
rect 37458 23508 37464 23520
rect 37419 23480 37464 23508
rect 37458 23468 37464 23480
rect 37516 23468 37522 23520
rect 37642 23508 37648 23520
rect 37603 23480 37648 23508
rect 37642 23468 37648 23480
rect 37700 23468 37706 23520
rect 38470 23508 38476 23520
rect 38431 23480 38476 23508
rect 38470 23468 38476 23480
rect 38528 23468 38534 23520
rect 38746 23468 38752 23520
rect 38804 23508 38810 23520
rect 39666 23508 39672 23520
rect 38804 23480 39672 23508
rect 38804 23468 38810 23480
rect 39666 23468 39672 23480
rect 39724 23468 39730 23520
rect 39945 23511 40003 23517
rect 39945 23477 39957 23511
rect 39991 23508 40003 23511
rect 41138 23508 41144 23520
rect 39991 23480 41144 23508
rect 39991 23477 40003 23480
rect 39945 23471 40003 23477
rect 41138 23468 41144 23480
rect 41196 23468 41202 23520
rect 42904 23508 42932 23607
rect 43898 23604 43904 23656
rect 43956 23644 43962 23656
rect 47486 23644 47492 23656
rect 43956 23616 47492 23644
rect 43956 23604 43962 23616
rect 47486 23604 47492 23616
rect 47544 23604 47550 23656
rect 43990 23536 43996 23588
rect 44048 23576 44054 23588
rect 44269 23579 44327 23585
rect 44269 23576 44281 23579
rect 44048 23548 44281 23576
rect 44048 23536 44054 23548
rect 44269 23545 44281 23548
rect 44315 23545 44327 23579
rect 44269 23539 44327 23545
rect 44174 23508 44180 23520
rect 42904 23480 44180 23508
rect 44174 23468 44180 23480
rect 44232 23468 44238 23520
rect 1104 23418 48852 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 48852 23418
rect 1104 23344 48852 23366
rect 17586 23304 17592 23316
rect 17547 23276 17592 23304
rect 17586 23264 17592 23276
rect 17644 23264 17650 23316
rect 18046 23264 18052 23316
rect 18104 23304 18110 23316
rect 18141 23307 18199 23313
rect 18141 23304 18153 23307
rect 18104 23276 18153 23304
rect 18104 23264 18110 23276
rect 18141 23273 18153 23276
rect 18187 23273 18199 23307
rect 18141 23267 18199 23273
rect 19702 23264 19708 23316
rect 19760 23304 19766 23316
rect 20070 23304 20076 23316
rect 19760 23276 20076 23304
rect 19760 23264 19766 23276
rect 20070 23264 20076 23276
rect 20128 23264 20134 23316
rect 20165 23307 20223 23313
rect 20165 23273 20177 23307
rect 20211 23304 20223 23307
rect 20254 23304 20260 23316
rect 20211 23276 20260 23304
rect 20211 23273 20223 23276
rect 20165 23267 20223 23273
rect 20254 23264 20260 23276
rect 20312 23264 20318 23316
rect 20349 23307 20407 23313
rect 20349 23273 20361 23307
rect 20395 23304 20407 23307
rect 20622 23304 20628 23316
rect 20395 23276 20628 23304
rect 20395 23273 20407 23276
rect 20349 23267 20407 23273
rect 20622 23264 20628 23276
rect 20680 23264 20686 23316
rect 22646 23264 22652 23316
rect 22704 23304 22710 23316
rect 23106 23304 23112 23316
rect 22704 23276 23112 23304
rect 22704 23264 22710 23276
rect 23106 23264 23112 23276
rect 23164 23264 23170 23316
rect 28353 23307 28411 23313
rect 28353 23273 28365 23307
rect 28399 23304 28411 23307
rect 30466 23304 30472 23316
rect 28399 23276 28764 23304
rect 28399 23273 28411 23276
rect 28353 23267 28411 23273
rect 28736 23248 28764 23276
rect 29472 23276 30472 23304
rect 19886 23196 19892 23248
rect 19944 23236 19950 23248
rect 19944 23208 20668 23236
rect 19944 23196 19950 23208
rect 20640 23180 20668 23208
rect 28258 23196 28264 23248
rect 28316 23236 28322 23248
rect 28537 23239 28595 23245
rect 28537 23236 28549 23239
rect 28316 23208 28549 23236
rect 28316 23196 28322 23208
rect 28537 23205 28549 23208
rect 28583 23205 28595 23239
rect 28537 23199 28595 23205
rect 28718 23196 28724 23248
rect 28776 23196 28782 23248
rect 19334 23128 19340 23180
rect 19392 23168 19398 23180
rect 19981 23171 20039 23177
rect 19981 23168 19993 23171
rect 19392 23140 19993 23168
rect 19392 23128 19398 23140
rect 19981 23137 19993 23140
rect 20027 23137 20039 23171
rect 19981 23131 20039 23137
rect 20622 23128 20628 23180
rect 20680 23128 20686 23180
rect 29472 23168 29500 23276
rect 30466 23264 30472 23276
rect 30524 23264 30530 23316
rect 32490 23264 32496 23316
rect 32548 23304 32554 23316
rect 33042 23304 33048 23316
rect 32548 23276 33048 23304
rect 32548 23264 32554 23276
rect 33042 23264 33048 23276
rect 33100 23264 33106 23316
rect 33318 23264 33324 23316
rect 33376 23304 33382 23316
rect 35713 23307 35771 23313
rect 35713 23304 35725 23307
rect 33376 23276 35725 23304
rect 33376 23264 33382 23276
rect 35713 23273 35725 23276
rect 35759 23304 35771 23307
rect 35986 23304 35992 23316
rect 35759 23276 35992 23304
rect 35759 23273 35771 23276
rect 35713 23267 35771 23273
rect 35986 23264 35992 23276
rect 36044 23304 36050 23316
rect 36538 23304 36544 23316
rect 36044 23276 36544 23304
rect 36044 23264 36050 23276
rect 36538 23264 36544 23276
rect 36596 23264 36602 23316
rect 37185 23307 37243 23313
rect 37185 23273 37197 23307
rect 37231 23304 37243 23307
rect 38470 23304 38476 23316
rect 37231 23276 38476 23304
rect 37231 23273 37243 23276
rect 37185 23267 37243 23273
rect 38470 23264 38476 23276
rect 38528 23264 38534 23316
rect 40221 23307 40279 23313
rect 40221 23273 40233 23307
rect 40267 23304 40279 23307
rect 40494 23304 40500 23316
rect 40267 23276 40500 23304
rect 40267 23273 40279 23276
rect 40221 23267 40279 23273
rect 40494 23264 40500 23276
rect 40552 23304 40558 23316
rect 40862 23304 40868 23316
rect 40552 23276 40868 23304
rect 40552 23264 40558 23276
rect 40862 23264 40868 23276
rect 40920 23264 40926 23316
rect 42150 23304 42156 23316
rect 41386 23276 42156 23304
rect 30006 23196 30012 23248
rect 30064 23236 30070 23248
rect 30193 23239 30251 23245
rect 30193 23236 30205 23239
rect 30064 23208 30205 23236
rect 30064 23196 30070 23208
rect 30193 23205 30205 23208
rect 30239 23236 30251 23239
rect 30282 23236 30288 23248
rect 30239 23208 30288 23236
rect 30239 23205 30251 23208
rect 30193 23199 30251 23205
rect 30282 23196 30288 23208
rect 30340 23196 30346 23248
rect 30926 23196 30932 23248
rect 30984 23236 30990 23248
rect 35253 23239 35311 23245
rect 35253 23236 35265 23239
rect 30984 23208 35265 23236
rect 30984 23196 30990 23208
rect 35253 23205 35265 23208
rect 35299 23236 35311 23239
rect 35299 23208 36124 23236
rect 35299 23205 35311 23208
rect 35253 23199 35311 23205
rect 28184 23140 29500 23168
rect 16209 23103 16267 23109
rect 16209 23069 16221 23103
rect 16255 23100 16267 23103
rect 16850 23100 16856 23112
rect 16255 23072 16856 23100
rect 16255 23069 16267 23072
rect 16209 23063 16267 23069
rect 16850 23060 16856 23072
rect 16908 23060 16914 23112
rect 18049 23103 18107 23109
rect 18049 23069 18061 23103
rect 18095 23069 18107 23103
rect 20162 23100 20168 23112
rect 20123 23072 20168 23100
rect 18049 23063 18107 23069
rect 16298 22992 16304 23044
rect 16356 23032 16362 23044
rect 16454 23035 16512 23041
rect 16454 23032 16466 23035
rect 16356 23004 16466 23032
rect 16356 22992 16362 23004
rect 16454 23001 16466 23004
rect 16500 23001 16512 23035
rect 16454 22995 16512 23001
rect 16758 22992 16764 23044
rect 16816 23032 16822 23044
rect 18064 23032 18092 23063
rect 20162 23060 20168 23072
rect 20220 23100 20226 23112
rect 20990 23100 20996 23112
rect 20220 23072 20996 23100
rect 20220 23060 20226 23072
rect 20990 23060 20996 23072
rect 21048 23060 21054 23112
rect 22922 23060 22928 23112
rect 22980 23100 22986 23112
rect 23477 23103 23535 23109
rect 23477 23100 23489 23103
rect 22980 23072 23489 23100
rect 22980 23060 22986 23072
rect 23477 23069 23489 23072
rect 23523 23100 23535 23103
rect 23750 23100 23756 23112
rect 23523 23072 23756 23100
rect 23523 23069 23535 23072
rect 23477 23063 23535 23069
rect 23750 23060 23756 23072
rect 23808 23060 23814 23112
rect 28184 23109 28212 23140
rect 29546 23128 29552 23180
rect 29604 23168 29610 23180
rect 35434 23168 35440 23180
rect 29604 23140 35440 23168
rect 29604 23128 29610 23140
rect 35434 23128 35440 23140
rect 35492 23128 35498 23180
rect 36096 23168 36124 23208
rect 36170 23196 36176 23248
rect 36228 23236 36234 23248
rect 36228 23208 37780 23236
rect 36228 23196 36234 23208
rect 36446 23168 36452 23180
rect 36096 23140 36452 23168
rect 36446 23128 36452 23140
rect 36504 23128 36510 23180
rect 37277 23171 37335 23177
rect 37277 23137 37289 23171
rect 37323 23168 37335 23171
rect 37642 23168 37648 23180
rect 37323 23140 37648 23168
rect 37323 23137 37335 23140
rect 37277 23131 37335 23137
rect 37642 23128 37648 23140
rect 37700 23128 37706 23180
rect 28169 23103 28227 23109
rect 28169 23069 28181 23103
rect 28215 23069 28227 23103
rect 28169 23063 28227 23069
rect 28353 23103 28411 23109
rect 28353 23069 28365 23103
rect 28399 23100 28411 23103
rect 29454 23100 29460 23112
rect 28399 23072 29460 23100
rect 28399 23069 28411 23072
rect 28353 23063 28411 23069
rect 29454 23060 29460 23072
rect 29512 23060 29518 23112
rect 30837 23103 30895 23109
rect 30837 23069 30849 23103
rect 30883 23100 30895 23103
rect 31938 23100 31944 23112
rect 30883 23072 31944 23100
rect 30883 23069 30895 23072
rect 30837 23063 30895 23069
rect 31938 23060 31944 23072
rect 31996 23100 32002 23112
rect 32125 23103 32183 23109
rect 32125 23100 32137 23103
rect 31996 23072 32137 23100
rect 31996 23060 32002 23072
rect 32125 23069 32137 23072
rect 32171 23069 32183 23103
rect 32125 23063 32183 23069
rect 34790 23060 34796 23112
rect 34848 23100 34854 23112
rect 35069 23103 35127 23109
rect 35069 23100 35081 23103
rect 34848 23072 35081 23100
rect 34848 23060 34854 23072
rect 35069 23069 35081 23072
rect 35115 23100 35127 23103
rect 35713 23103 35771 23109
rect 35713 23100 35725 23103
rect 35115 23072 35725 23100
rect 35115 23069 35127 23072
rect 35069 23063 35127 23069
rect 35713 23069 35725 23072
rect 35759 23100 35771 23103
rect 35802 23100 35808 23112
rect 35759 23072 35808 23100
rect 35759 23069 35771 23072
rect 35713 23063 35771 23069
rect 35802 23060 35808 23072
rect 35860 23060 35866 23112
rect 35897 23103 35955 23109
rect 35897 23069 35909 23103
rect 35943 23069 35955 23103
rect 35897 23063 35955 23069
rect 35989 23103 36047 23109
rect 35989 23069 36001 23103
rect 36035 23100 36047 23103
rect 36262 23100 36268 23112
rect 36035 23072 36268 23100
rect 36035 23069 36047 23072
rect 35989 23063 36047 23069
rect 16816 23004 18092 23032
rect 16816 22992 16822 23004
rect 19426 22992 19432 23044
rect 19484 23032 19490 23044
rect 19889 23035 19947 23041
rect 19889 23032 19901 23035
rect 19484 23004 19901 23032
rect 19484 22992 19490 23004
rect 19889 23001 19901 23004
rect 19935 23001 19947 23035
rect 23290 23032 23296 23044
rect 23251 23004 23296 23032
rect 19889 22995 19947 23001
rect 23290 22992 23296 23004
rect 23348 22992 23354 23044
rect 23661 23035 23719 23041
rect 23661 23001 23673 23035
rect 23707 23032 23719 23035
rect 24578 23032 24584 23044
rect 23707 23004 24584 23032
rect 23707 23001 23719 23004
rect 23661 22995 23719 23001
rect 24578 22992 24584 23004
rect 24636 22992 24642 23044
rect 27525 23035 27583 23041
rect 27525 23001 27537 23035
rect 27571 23032 27583 23035
rect 27798 23032 27804 23044
rect 27571 23004 27804 23032
rect 27571 23001 27583 23004
rect 27525 22995 27583 23001
rect 27798 22992 27804 23004
rect 27856 23032 27862 23044
rect 30009 23035 30067 23041
rect 30009 23032 30021 23035
rect 27856 23004 30021 23032
rect 27856 22992 27862 23004
rect 30009 23001 30021 23004
rect 30055 23001 30067 23035
rect 30009 22995 30067 23001
rect 31021 23035 31079 23041
rect 31021 23001 31033 23035
rect 31067 23032 31079 23035
rect 31110 23032 31116 23044
rect 31067 23004 31116 23032
rect 31067 23001 31079 23004
rect 31021 22995 31079 23001
rect 31110 22992 31116 23004
rect 31168 22992 31174 23044
rect 32030 22992 32036 23044
rect 32088 23032 32094 23044
rect 32309 23035 32367 23041
rect 32309 23032 32321 23035
rect 32088 23004 32321 23032
rect 32088 22992 32094 23004
rect 32309 23001 32321 23004
rect 32355 23001 32367 23035
rect 32309 22995 32367 23001
rect 18598 22924 18604 22976
rect 18656 22964 18662 22976
rect 24946 22964 24952 22976
rect 18656 22936 24952 22964
rect 18656 22924 18662 22936
rect 24946 22924 24952 22936
rect 25004 22924 25010 22976
rect 27338 22924 27344 22976
rect 27396 22964 27402 22976
rect 27617 22967 27675 22973
rect 27617 22964 27629 22967
rect 27396 22936 27629 22964
rect 27396 22924 27402 22936
rect 27617 22933 27629 22936
rect 27663 22933 27675 22967
rect 27617 22927 27675 22933
rect 27706 22924 27712 22976
rect 27764 22964 27770 22976
rect 28718 22964 28724 22976
rect 27764 22936 28724 22964
rect 27764 22924 27770 22936
rect 28718 22924 28724 22936
rect 28776 22924 28782 22976
rect 31205 22967 31263 22973
rect 31205 22933 31217 22967
rect 31251 22964 31263 22967
rect 31386 22964 31392 22976
rect 31251 22936 31392 22964
rect 31251 22933 31263 22936
rect 31205 22927 31263 22933
rect 31386 22924 31392 22936
rect 31444 22924 31450 22976
rect 32493 22967 32551 22973
rect 32493 22933 32505 22967
rect 32539 22964 32551 22967
rect 32674 22964 32680 22976
rect 32539 22936 32680 22964
rect 32539 22933 32551 22936
rect 32493 22927 32551 22933
rect 32674 22924 32680 22936
rect 32732 22924 32738 22976
rect 35710 22924 35716 22976
rect 35768 22964 35774 22976
rect 35912 22964 35940 23063
rect 36262 23060 36268 23072
rect 36320 23060 36326 23112
rect 37369 23103 37427 23109
rect 37369 23069 37381 23103
rect 37415 23100 37427 23103
rect 37550 23100 37556 23112
rect 37415 23072 37556 23100
rect 37415 23069 37427 23072
rect 37369 23063 37427 23069
rect 37550 23060 37556 23072
rect 37608 23060 37614 23112
rect 37752 23100 37780 23208
rect 38102 23196 38108 23248
rect 38160 23236 38166 23248
rect 38749 23239 38807 23245
rect 38160 23208 38700 23236
rect 38160 23196 38166 23208
rect 38470 23168 38476 23180
rect 38431 23140 38476 23168
rect 38470 23128 38476 23140
rect 38528 23128 38534 23180
rect 38672 23168 38700 23208
rect 38749 23205 38761 23239
rect 38795 23236 38807 23239
rect 39022 23236 39028 23248
rect 38795 23208 39028 23236
rect 38795 23205 38807 23208
rect 38749 23199 38807 23205
rect 39022 23196 39028 23208
rect 39080 23196 39086 23248
rect 38672 23140 40080 23168
rect 38381 23103 38439 23109
rect 38381 23100 38393 23103
rect 37752 23072 38393 23100
rect 38381 23069 38393 23072
rect 38427 23069 38439 23103
rect 38381 23063 38439 23069
rect 39758 23060 39764 23112
rect 39816 23100 39822 23112
rect 40052 23109 40080 23140
rect 40586 23128 40592 23180
rect 40644 23168 40650 23180
rect 41386 23168 41414 23276
rect 42150 23264 42156 23276
rect 42208 23264 42214 23316
rect 45922 23264 45928 23316
rect 45980 23304 45986 23316
rect 46934 23304 46940 23316
rect 45980 23276 46940 23304
rect 45980 23264 45986 23276
rect 46934 23264 46940 23276
rect 46992 23264 46998 23316
rect 41509 23171 41567 23177
rect 41509 23168 41521 23171
rect 40644 23140 41521 23168
rect 40644 23128 40650 23140
rect 41509 23137 41521 23140
rect 41555 23137 41567 23171
rect 41509 23131 41567 23137
rect 41693 23171 41751 23177
rect 41693 23137 41705 23171
rect 41739 23168 41751 23171
rect 42334 23168 42340 23180
rect 41739 23140 42212 23168
rect 42295 23140 42340 23168
rect 41739 23137 41751 23140
rect 41693 23131 41751 23137
rect 39853 23103 39911 23109
rect 39853 23100 39865 23103
rect 39816 23072 39865 23100
rect 39816 23060 39822 23072
rect 39853 23069 39865 23072
rect 39899 23069 39911 23103
rect 39853 23063 39911 23069
rect 40037 23103 40095 23109
rect 40037 23069 40049 23103
rect 40083 23069 40095 23103
rect 40037 23063 40095 23069
rect 37093 23035 37151 23041
rect 37093 23001 37105 23035
rect 37139 23032 37151 23035
rect 38102 23032 38108 23044
rect 37139 23004 38108 23032
rect 37139 23001 37151 23004
rect 37093 22995 37151 23001
rect 38102 22992 38108 23004
rect 38160 22992 38166 23044
rect 39868 23032 39896 23063
rect 41598 23060 41604 23112
rect 41656 23100 41662 23112
rect 41785 23103 41843 23109
rect 41656 23072 41701 23100
rect 41656 23060 41662 23072
rect 41785 23069 41797 23103
rect 41831 23069 41843 23103
rect 42184 23100 42212 23140
rect 42334 23128 42340 23140
rect 42392 23128 42398 23180
rect 43625 23171 43683 23177
rect 43625 23137 43637 23171
rect 43671 23168 43683 23171
rect 43990 23168 43996 23180
rect 43671 23140 43996 23168
rect 43671 23137 43683 23140
rect 43625 23131 43683 23137
rect 43990 23128 43996 23140
rect 44048 23128 44054 23180
rect 42610 23100 42616 23112
rect 42184 23072 42616 23100
rect 41785 23063 41843 23069
rect 41616 23032 41644 23060
rect 39868 23004 41644 23032
rect 41800 23032 41828 23063
rect 42610 23060 42616 23072
rect 42668 23100 42674 23112
rect 43346 23100 43352 23112
rect 42668 23072 43352 23100
rect 42668 23060 42674 23072
rect 43346 23060 43352 23072
rect 43404 23060 43410 23112
rect 43901 23103 43959 23109
rect 43901 23069 43913 23103
rect 43947 23100 43959 23103
rect 45002 23100 45008 23112
rect 43947 23072 45008 23100
rect 43947 23069 43959 23072
rect 43901 23063 43959 23069
rect 42426 23032 42432 23044
rect 41800 23004 42432 23032
rect 42426 22992 42432 23004
rect 42484 23032 42490 23044
rect 42886 23032 42892 23044
rect 42484 23004 42892 23032
rect 42484 22992 42490 23004
rect 42886 22992 42892 23004
rect 42944 23032 42950 23044
rect 43916 23032 43944 23063
rect 45002 23060 45008 23072
rect 45060 23060 45066 23112
rect 42944 23004 43944 23032
rect 42944 22992 42950 23004
rect 36170 22964 36176 22976
rect 35768 22936 35940 22964
rect 36131 22936 36176 22964
rect 35768 22924 35774 22936
rect 36170 22924 36176 22936
rect 36228 22924 36234 22976
rect 37550 22964 37556 22976
rect 37511 22936 37556 22964
rect 37550 22924 37556 22936
rect 37608 22924 37614 22976
rect 41325 22967 41383 22973
rect 41325 22933 41337 22967
rect 41371 22964 41383 22967
rect 41966 22964 41972 22976
rect 41371 22936 41972 22964
rect 41371 22933 41383 22936
rect 41325 22927 41383 22933
rect 41966 22924 41972 22936
rect 42024 22924 42030 22976
rect 1104 22874 48852 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 48852 22874
rect 1104 22800 48852 22822
rect 16853 22763 16911 22769
rect 16853 22729 16865 22763
rect 16899 22760 16911 22763
rect 17126 22760 17132 22772
rect 16899 22732 17132 22760
rect 16899 22729 16911 22732
rect 16853 22723 16911 22729
rect 17126 22720 17132 22732
rect 17184 22720 17190 22772
rect 18690 22760 18696 22772
rect 17788 22732 18696 22760
rect 2038 22692 2044 22704
rect 1999 22664 2044 22692
rect 2038 22652 2044 22664
rect 2096 22652 2102 22704
rect 17788 22701 17816 22732
rect 18690 22720 18696 22732
rect 18748 22720 18754 22772
rect 20073 22763 20131 22769
rect 20073 22729 20085 22763
rect 20119 22760 20131 22763
rect 20530 22760 20536 22772
rect 20119 22732 20536 22760
rect 20119 22729 20131 22732
rect 20073 22723 20131 22729
rect 20530 22720 20536 22732
rect 20588 22720 20594 22772
rect 23385 22763 23443 22769
rect 23385 22729 23397 22763
rect 23431 22760 23443 22763
rect 24394 22760 24400 22772
rect 23431 22732 24400 22760
rect 23431 22729 23443 22732
rect 23385 22723 23443 22729
rect 24394 22720 24400 22732
rect 24452 22720 24458 22772
rect 27798 22760 27804 22772
rect 27759 22732 27804 22760
rect 27798 22720 27804 22732
rect 27856 22720 27862 22772
rect 32858 22760 32864 22772
rect 31588 22732 32864 22760
rect 17773 22695 17831 22701
rect 17773 22661 17785 22695
rect 17819 22661 17831 22695
rect 18966 22692 18972 22704
rect 17773 22655 17831 22661
rect 18628 22664 18972 22692
rect 18628 22658 18656 22664
rect 18613 22639 18656 22658
rect 18966 22652 18972 22664
rect 19024 22652 19030 22704
rect 23566 22692 23572 22704
rect 20272 22664 23572 22692
rect 1854 22624 1860 22636
rect 1815 22596 1860 22624
rect 1854 22584 1860 22596
rect 1912 22584 1918 22636
rect 3418 22624 3424 22636
rect 3379 22596 3424 22624
rect 3418 22584 3424 22596
rect 3476 22584 3482 22636
rect 15473 22627 15531 22633
rect 15473 22593 15485 22627
rect 15519 22624 15531 22627
rect 16574 22624 16580 22636
rect 15519 22596 16580 22624
rect 15519 22593 15531 22596
rect 15473 22587 15531 22593
rect 16574 22584 16580 22596
rect 16632 22584 16638 22636
rect 16761 22627 16819 22633
rect 16761 22593 16773 22627
rect 16807 22593 16819 22627
rect 16761 22587 16819 22593
rect 17405 22627 17463 22633
rect 17405 22593 17417 22627
rect 17451 22593 17463 22627
rect 17405 22587 17463 22593
rect 17589 22627 17647 22633
rect 17589 22593 17601 22627
rect 17635 22624 17647 22627
rect 18322 22624 18328 22636
rect 17635 22596 18328 22624
rect 17635 22593 17647 22596
rect 17589 22587 17647 22593
rect 13814 22516 13820 22568
rect 13872 22556 13878 22568
rect 15749 22559 15807 22565
rect 15749 22556 15761 22559
rect 13872 22528 15761 22556
rect 13872 22516 13878 22528
rect 15749 22525 15761 22528
rect 15795 22525 15807 22559
rect 15749 22519 15807 22525
rect 15194 22448 15200 22500
rect 15252 22488 15258 22500
rect 16776 22488 16804 22587
rect 17420 22556 17448 22587
rect 18322 22584 18328 22596
rect 18380 22584 18386 22636
rect 18506 22633 18512 22636
rect 18489 22627 18512 22633
rect 18489 22593 18501 22627
rect 18489 22587 18512 22593
rect 18506 22584 18512 22587
rect 18564 22584 18570 22636
rect 18598 22633 18656 22639
rect 18598 22599 18610 22633
rect 18644 22599 18656 22633
rect 18598 22593 18656 22599
rect 18690 22584 18696 22636
rect 18748 22624 18754 22636
rect 18874 22624 18880 22636
rect 18748 22596 18790 22624
rect 18835 22596 18880 22624
rect 18748 22584 18754 22596
rect 18874 22584 18880 22596
rect 18932 22624 18938 22636
rect 19242 22624 19248 22636
rect 18932 22596 19248 22624
rect 18932 22584 18938 22596
rect 19242 22584 19248 22596
rect 19300 22584 19306 22636
rect 19518 22584 19524 22636
rect 19576 22624 19582 22636
rect 19613 22627 19671 22633
rect 19613 22624 19625 22627
rect 19576 22596 19625 22624
rect 19576 22584 19582 22596
rect 19613 22593 19625 22596
rect 19659 22593 19671 22627
rect 19886 22624 19892 22636
rect 19847 22596 19892 22624
rect 19613 22587 19671 22593
rect 19886 22584 19892 22596
rect 19944 22584 19950 22636
rect 18138 22556 18144 22568
rect 17420 22528 18144 22556
rect 18138 22516 18144 22528
rect 18196 22516 18202 22568
rect 19426 22516 19432 22568
rect 19484 22556 19490 22568
rect 19705 22559 19763 22565
rect 19705 22556 19717 22559
rect 19484 22528 19717 22556
rect 19484 22516 19490 22528
rect 19705 22525 19717 22528
rect 19751 22525 19763 22559
rect 19705 22519 19763 22525
rect 15252 22460 16804 22488
rect 15252 22448 15258 22460
rect 18506 22448 18512 22500
rect 18564 22488 18570 22500
rect 20272 22488 20300 22664
rect 23566 22652 23572 22664
rect 23624 22652 23630 22704
rect 24486 22652 24492 22704
rect 24544 22692 24550 22704
rect 25406 22692 25412 22704
rect 24544 22664 25412 22692
rect 24544 22652 24550 22664
rect 23201 22627 23259 22633
rect 23201 22593 23213 22627
rect 23247 22624 23259 22627
rect 23477 22627 23535 22633
rect 23247 22596 23428 22624
rect 23247 22593 23259 22596
rect 23201 22587 23259 22593
rect 23198 22488 23204 22500
rect 18564 22460 20300 22488
rect 23159 22460 23204 22488
rect 18564 22448 18570 22460
rect 23198 22448 23204 22460
rect 23256 22448 23262 22500
rect 23400 22488 23428 22596
rect 23477 22593 23489 22627
rect 23523 22624 23535 22627
rect 23658 22624 23664 22636
rect 23523 22596 23664 22624
rect 23523 22593 23535 22596
rect 23477 22587 23535 22593
rect 23658 22584 23664 22596
rect 23716 22584 23722 22636
rect 24854 22624 24860 22636
rect 24815 22596 24860 22624
rect 24854 22584 24860 22596
rect 24912 22584 24918 22636
rect 24964 22633 24992 22664
rect 25406 22652 25412 22664
rect 25464 22652 25470 22704
rect 27617 22695 27675 22701
rect 27617 22661 27629 22695
rect 27663 22692 27675 22695
rect 28074 22692 28080 22704
rect 27663 22664 28080 22692
rect 27663 22661 27675 22664
rect 27617 22655 27675 22661
rect 28074 22652 28080 22664
rect 28132 22652 28138 22704
rect 31478 22692 31484 22704
rect 28460 22664 28994 22692
rect 24949 22627 25007 22633
rect 24949 22593 24961 22627
rect 24995 22593 25007 22627
rect 24949 22587 25007 22593
rect 25041 22627 25099 22633
rect 25041 22593 25053 22627
rect 25087 22624 25099 22627
rect 25130 22624 25136 22636
rect 25087 22596 25136 22624
rect 25087 22593 25099 22596
rect 25041 22587 25099 22593
rect 25130 22584 25136 22596
rect 25188 22584 25194 22636
rect 25225 22627 25283 22633
rect 25225 22593 25237 22627
rect 25271 22624 25283 22627
rect 25682 22624 25688 22636
rect 25271 22596 25688 22624
rect 25271 22593 25283 22596
rect 25225 22587 25283 22593
rect 25682 22584 25688 22596
rect 25740 22584 25746 22636
rect 27433 22627 27491 22633
rect 27433 22593 27445 22627
rect 27479 22624 27491 22627
rect 27706 22624 27712 22636
rect 27479 22596 27712 22624
rect 27479 22593 27491 22596
rect 27433 22587 27491 22593
rect 27706 22584 27712 22596
rect 27764 22584 27770 22636
rect 28460 22633 28488 22664
rect 28445 22627 28503 22633
rect 28445 22593 28457 22627
rect 28491 22593 28503 22627
rect 28718 22624 28724 22636
rect 28679 22596 28724 22624
rect 28445 22587 28503 22593
rect 28718 22584 28724 22596
rect 28776 22584 28782 22636
rect 28966 22624 28994 22664
rect 31312 22664 31484 22692
rect 29457 22627 29515 22633
rect 29457 22624 29469 22627
rect 28966 22596 29469 22624
rect 29457 22593 29469 22596
rect 29503 22624 29515 22627
rect 29546 22624 29552 22636
rect 29503 22596 29552 22624
rect 29503 22593 29515 22596
rect 29457 22587 29515 22593
rect 29546 22584 29552 22596
rect 29604 22584 29610 22636
rect 30926 22584 30932 22636
rect 30984 22624 30990 22636
rect 31312 22633 31340 22664
rect 31478 22652 31484 22664
rect 31536 22652 31542 22704
rect 31205 22627 31263 22633
rect 31205 22624 31217 22627
rect 30984 22596 31217 22624
rect 30984 22584 30990 22596
rect 31205 22593 31217 22596
rect 31251 22593 31263 22627
rect 31205 22587 31263 22593
rect 31297 22627 31355 22633
rect 31297 22593 31309 22627
rect 31343 22593 31355 22627
rect 31297 22587 31355 22593
rect 31386 22584 31392 22636
rect 31444 22624 31450 22636
rect 31588 22633 31616 22732
rect 32858 22720 32864 22732
rect 32916 22760 32922 22772
rect 33410 22760 33416 22772
rect 32916 22732 33416 22760
rect 32916 22720 32922 22732
rect 33410 22720 33416 22732
rect 33468 22760 33474 22772
rect 33468 22732 34008 22760
rect 33468 22720 33474 22732
rect 31662 22652 31668 22704
rect 31720 22692 31726 22704
rect 33134 22692 33140 22704
rect 31720 22664 33140 22692
rect 31720 22652 31726 22664
rect 31573 22627 31631 22633
rect 31444 22596 31489 22624
rect 31444 22584 31450 22596
rect 31573 22593 31585 22627
rect 31619 22593 31631 22627
rect 32490 22624 32496 22636
rect 32451 22596 32496 22624
rect 31573 22587 31631 22593
rect 32490 22584 32496 22596
rect 32548 22584 32554 22636
rect 32600 22633 32628 22664
rect 33134 22652 33140 22664
rect 33192 22692 33198 22704
rect 33192 22664 33732 22692
rect 33192 22652 33198 22664
rect 32585 22627 32643 22633
rect 32585 22593 32597 22627
rect 32631 22593 32643 22627
rect 32585 22587 32643 22593
rect 32674 22584 32680 22636
rect 32732 22624 32738 22636
rect 32732 22596 32777 22624
rect 32732 22584 32738 22596
rect 32858 22584 32864 22636
rect 32916 22624 32922 22636
rect 32916 22596 32961 22624
rect 32916 22584 32922 22596
rect 33318 22584 33324 22636
rect 33376 22624 33382 22636
rect 33704 22633 33732 22664
rect 33980 22633 34008 22732
rect 37274 22720 37280 22772
rect 37332 22760 37338 22772
rect 40310 22760 40316 22772
rect 37332 22732 40316 22760
rect 37332 22720 37338 22732
rect 38120 22701 38148 22732
rect 40310 22720 40316 22732
rect 40368 22720 40374 22772
rect 40494 22720 40500 22772
rect 40552 22760 40558 22772
rect 40552 22732 40597 22760
rect 40552 22720 40558 22732
rect 44450 22720 44456 22772
rect 44508 22760 44514 22772
rect 48041 22763 48099 22769
rect 48041 22760 48053 22763
rect 44508 22732 48053 22760
rect 44508 22720 44514 22732
rect 48041 22729 48053 22732
rect 48087 22729 48099 22763
rect 48041 22723 48099 22729
rect 38105 22695 38163 22701
rect 38105 22661 38117 22695
rect 38151 22661 38163 22695
rect 38105 22655 38163 22661
rect 40862 22652 40868 22704
rect 40920 22692 40926 22704
rect 40920 22664 41414 22692
rect 40920 22652 40926 22664
rect 33597 22627 33655 22633
rect 33597 22624 33609 22627
rect 33376 22596 33609 22624
rect 33376 22584 33382 22596
rect 33597 22593 33609 22596
rect 33643 22593 33655 22627
rect 33597 22587 33655 22593
rect 33689 22627 33747 22633
rect 33689 22593 33701 22627
rect 33735 22593 33747 22627
rect 33689 22587 33747 22593
rect 33781 22627 33839 22633
rect 33781 22593 33793 22627
rect 33827 22593 33839 22627
rect 33781 22587 33839 22593
rect 33965 22627 34023 22633
rect 33965 22593 33977 22627
rect 34011 22593 34023 22627
rect 35802 22624 35808 22636
rect 35763 22596 35808 22624
rect 33965 22587 34023 22593
rect 23566 22516 23572 22568
rect 23624 22556 23630 22568
rect 28905 22559 28963 22565
rect 28905 22556 28917 22559
rect 23624 22528 28917 22556
rect 23624 22516 23630 22528
rect 28905 22525 28917 22528
rect 28951 22556 28963 22559
rect 28951 22528 31754 22556
rect 28951 22525 28963 22528
rect 28905 22519 28963 22525
rect 28626 22488 28632 22500
rect 23400 22460 28632 22488
rect 28626 22448 28632 22460
rect 28684 22448 28690 22500
rect 31726 22488 31754 22528
rect 32398 22516 32404 22568
rect 32456 22556 32462 22568
rect 33796 22556 33824 22587
rect 35802 22584 35808 22596
rect 35860 22584 35866 22636
rect 35986 22624 35992 22636
rect 35947 22596 35992 22624
rect 35986 22584 35992 22596
rect 36044 22584 36050 22636
rect 36170 22584 36176 22636
rect 36228 22624 36234 22636
rect 36814 22624 36820 22636
rect 36228 22596 36820 22624
rect 36228 22584 36234 22596
rect 36814 22584 36820 22596
rect 36872 22624 36878 22636
rect 37277 22627 37335 22633
rect 37277 22624 37289 22627
rect 36872 22596 37289 22624
rect 36872 22584 36878 22596
rect 37277 22593 37289 22596
rect 37323 22593 37335 22627
rect 37277 22587 37335 22593
rect 38289 22627 38347 22633
rect 38289 22593 38301 22627
rect 38335 22593 38347 22627
rect 38289 22587 38347 22593
rect 32456 22528 33824 22556
rect 32456 22516 32462 22528
rect 37090 22516 37096 22568
rect 37148 22556 37154 22568
rect 37369 22559 37427 22565
rect 37369 22556 37381 22559
rect 37148 22528 37381 22556
rect 37148 22516 37154 22528
rect 37369 22525 37381 22528
rect 37415 22525 37427 22559
rect 38304 22556 38332 22587
rect 38378 22584 38384 22636
rect 38436 22624 38442 22636
rect 40405 22627 40463 22633
rect 38436 22596 38481 22624
rect 38436 22584 38442 22596
rect 40405 22593 40417 22627
rect 40451 22593 40463 22627
rect 41386 22624 41414 22664
rect 41598 22652 41604 22704
rect 41656 22692 41662 22704
rect 42429 22695 42487 22701
rect 42429 22692 42441 22695
rect 41656 22664 42441 22692
rect 41656 22652 41662 22664
rect 42429 22661 42441 22664
rect 42475 22661 42487 22695
rect 42429 22655 42487 22661
rect 41785 22627 41843 22633
rect 41785 22624 41797 22627
rect 41386 22596 41797 22624
rect 40405 22587 40463 22593
rect 41785 22593 41797 22596
rect 41831 22624 41843 22627
rect 42705 22627 42763 22633
rect 42705 22624 42717 22627
rect 41831 22596 42717 22624
rect 41831 22593 41843 22596
rect 41785 22587 41843 22593
rect 42705 22593 42717 22596
rect 42751 22624 42763 22627
rect 43070 22624 43076 22636
rect 42751 22596 43076 22624
rect 42751 22593 42763 22596
rect 42705 22587 42763 22593
rect 37369 22519 37427 22525
rect 37936 22528 38332 22556
rect 32122 22488 32128 22500
rect 31726 22460 32128 22488
rect 32122 22448 32128 22460
rect 32180 22448 32186 22500
rect 32490 22448 32496 22500
rect 32548 22488 32554 22500
rect 36078 22488 36084 22500
rect 32548 22460 36084 22488
rect 32548 22448 32554 22460
rect 3510 22420 3516 22432
rect 3471 22392 3516 22420
rect 3510 22380 3516 22392
rect 3568 22380 3574 22432
rect 18230 22420 18236 22432
rect 18191 22392 18236 22420
rect 18230 22380 18236 22392
rect 18288 22380 18294 22432
rect 19334 22380 19340 22432
rect 19392 22420 19398 22432
rect 19613 22423 19671 22429
rect 19613 22420 19625 22423
rect 19392 22392 19625 22420
rect 19392 22380 19398 22392
rect 19613 22389 19625 22392
rect 19659 22389 19671 22423
rect 19613 22383 19671 22389
rect 20070 22380 20076 22432
rect 20128 22420 20134 22432
rect 20530 22420 20536 22432
rect 20128 22392 20536 22420
rect 20128 22380 20134 22392
rect 20530 22380 20536 22392
rect 20588 22380 20594 22432
rect 24581 22423 24639 22429
rect 24581 22389 24593 22423
rect 24627 22420 24639 22423
rect 24946 22420 24952 22432
rect 24627 22392 24952 22420
rect 24627 22389 24639 22392
rect 24581 22383 24639 22389
rect 24946 22380 24952 22392
rect 25004 22380 25010 22432
rect 28074 22380 28080 22432
rect 28132 22420 28138 22432
rect 28350 22420 28356 22432
rect 28132 22392 28356 22420
rect 28132 22380 28138 22392
rect 28350 22380 28356 22392
rect 28408 22420 28414 22432
rect 29549 22423 29607 22429
rect 29549 22420 29561 22423
rect 28408 22392 29561 22420
rect 28408 22380 28414 22392
rect 29549 22389 29561 22392
rect 29595 22389 29607 22423
rect 30926 22420 30932 22432
rect 30887 22392 30932 22420
rect 29549 22383 29607 22389
rect 30926 22380 30932 22392
rect 30984 22380 30990 22432
rect 32214 22420 32220 22432
rect 32175 22392 32220 22420
rect 32214 22380 32220 22392
rect 32272 22380 32278 22432
rect 33318 22420 33324 22432
rect 33279 22392 33324 22420
rect 33318 22380 33324 22392
rect 33376 22380 33382 22432
rect 35912 22429 35940 22460
rect 36078 22448 36084 22460
rect 36136 22448 36142 22500
rect 37458 22488 37464 22500
rect 36188 22460 37464 22488
rect 36188 22432 36216 22460
rect 37458 22448 37464 22460
rect 37516 22488 37522 22500
rect 37936 22488 37964 22528
rect 38470 22516 38476 22568
rect 38528 22556 38534 22568
rect 40420 22556 40448 22587
rect 43070 22584 43076 22596
rect 43128 22584 43134 22636
rect 44082 22584 44088 22636
rect 44140 22624 44146 22636
rect 45281 22627 45339 22633
rect 45281 22624 45293 22627
rect 44140 22596 45293 22624
rect 44140 22584 44146 22596
rect 45281 22593 45293 22596
rect 45327 22593 45339 22627
rect 45281 22587 45339 22593
rect 45465 22627 45523 22633
rect 45465 22593 45477 22627
rect 45511 22624 45523 22627
rect 46842 22624 46848 22636
rect 45511 22596 46848 22624
rect 45511 22593 45523 22596
rect 45465 22587 45523 22593
rect 46842 22584 46848 22596
rect 46900 22584 46906 22636
rect 47946 22624 47952 22636
rect 47907 22596 47952 22624
rect 47946 22584 47952 22596
rect 48004 22584 48010 22636
rect 38528 22528 41000 22556
rect 38528 22516 38534 22528
rect 38102 22488 38108 22500
rect 37516 22460 37964 22488
rect 38063 22460 38108 22488
rect 37516 22448 37522 22460
rect 38102 22448 38108 22460
rect 38160 22448 38166 22500
rect 40129 22491 40187 22497
rect 40129 22457 40141 22491
rect 40175 22488 40187 22491
rect 40862 22488 40868 22500
rect 40175 22460 40868 22488
rect 40175 22457 40187 22460
rect 40129 22451 40187 22457
rect 40862 22448 40868 22460
rect 40920 22448 40926 22500
rect 40972 22488 41000 22528
rect 41322 22516 41328 22568
rect 41380 22556 41386 22568
rect 41509 22559 41567 22565
rect 41509 22556 41521 22559
rect 41380 22528 41521 22556
rect 41380 22516 41386 22528
rect 41509 22525 41521 22528
rect 41555 22525 41567 22559
rect 41509 22519 41567 22525
rect 41601 22559 41659 22565
rect 41601 22525 41613 22559
rect 41647 22525 41659 22559
rect 41601 22519 41659 22525
rect 41693 22559 41751 22565
rect 41693 22525 41705 22559
rect 41739 22556 41751 22559
rect 42426 22556 42432 22568
rect 41739 22528 42432 22556
rect 41739 22525 41751 22528
rect 41693 22519 41751 22525
rect 41616 22488 41644 22519
rect 42426 22516 42432 22528
rect 42484 22516 42490 22568
rect 42610 22556 42616 22568
rect 42571 22528 42616 22556
rect 42610 22516 42616 22528
rect 42668 22516 42674 22568
rect 42334 22488 42340 22500
rect 40972 22460 42340 22488
rect 42334 22448 42340 22460
rect 42392 22448 42398 22500
rect 35897 22423 35955 22429
rect 35897 22389 35909 22423
rect 35943 22389 35955 22423
rect 36170 22420 36176 22432
rect 36131 22392 36176 22420
rect 35897 22383 35955 22389
rect 36170 22380 36176 22392
rect 36228 22380 36234 22432
rect 37366 22420 37372 22432
rect 37327 22392 37372 22420
rect 37366 22380 37372 22392
rect 37424 22380 37430 22432
rect 37642 22420 37648 22432
rect 37603 22392 37648 22420
rect 37642 22380 37648 22392
rect 37700 22380 37706 22432
rect 40678 22420 40684 22432
rect 40639 22392 40684 22420
rect 40678 22380 40684 22392
rect 40736 22380 40742 22432
rect 40954 22380 40960 22432
rect 41012 22420 41018 22432
rect 41325 22423 41383 22429
rect 41325 22420 41337 22423
rect 41012 22392 41337 22420
rect 41012 22380 41018 22392
rect 41325 22389 41337 22392
rect 41371 22389 41383 22423
rect 42426 22420 42432 22432
rect 42387 22392 42432 22420
rect 41325 22383 41383 22389
rect 42426 22380 42432 22392
rect 42484 22380 42490 22432
rect 42518 22380 42524 22432
rect 42576 22420 42582 22432
rect 42889 22423 42947 22429
rect 42889 22420 42901 22423
rect 42576 22392 42901 22420
rect 42576 22380 42582 22392
rect 42889 22389 42901 22392
rect 42935 22389 42947 22423
rect 42889 22383 42947 22389
rect 45462 22380 45468 22432
rect 45520 22420 45526 22432
rect 45649 22423 45707 22429
rect 45649 22420 45661 22423
rect 45520 22392 45661 22420
rect 45520 22380 45526 22392
rect 45649 22389 45661 22392
rect 45695 22389 45707 22423
rect 45649 22383 45707 22389
rect 1104 22330 48852 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 48852 22330
rect 1104 22256 48852 22278
rect 18506 22216 18512 22228
rect 14108 22188 18512 22216
rect 2866 22040 2872 22092
rect 2924 22080 2930 22092
rect 14108 22089 14136 22188
rect 18506 22176 18512 22188
rect 18564 22176 18570 22228
rect 25038 22216 25044 22228
rect 24688 22188 25044 22216
rect 18233 22151 18291 22157
rect 18233 22117 18245 22151
rect 18279 22148 18291 22151
rect 18322 22148 18328 22160
rect 18279 22120 18328 22148
rect 18279 22117 18291 22120
rect 18233 22111 18291 22117
rect 18322 22108 18328 22120
rect 18380 22108 18386 22160
rect 4249 22083 4307 22089
rect 4249 22080 4261 22083
rect 2924 22052 4261 22080
rect 2924 22040 2930 22052
rect 4249 22049 4261 22052
rect 4295 22049 4307 22083
rect 4249 22043 4307 22049
rect 14093 22083 14151 22089
rect 14093 22049 14105 22083
rect 14139 22049 14151 22083
rect 15470 22080 15476 22092
rect 15431 22052 15476 22080
rect 14093 22043 14151 22049
rect 15470 22040 15476 22052
rect 15528 22040 15534 22092
rect 18138 22040 18144 22092
rect 18196 22080 18202 22092
rect 18414 22080 18420 22092
rect 18196 22052 18420 22080
rect 18196 22040 18202 22052
rect 18414 22040 18420 22052
rect 18472 22080 18478 22092
rect 21818 22080 21824 22092
rect 18472 22052 19288 22080
rect 18472 22040 18478 22052
rect 3053 22015 3111 22021
rect 3053 21981 3065 22015
rect 3099 22012 3111 22015
rect 3418 22012 3424 22024
rect 3099 21984 3424 22012
rect 3099 21981 3111 21984
rect 3053 21975 3111 21981
rect 3418 21972 3424 21984
rect 3476 21972 3482 22024
rect 3786 22012 3792 22024
rect 3747 21984 3792 22012
rect 3786 21972 3792 21984
rect 3844 21972 3850 22024
rect 16850 22012 16856 22024
rect 16763 21984 16856 22012
rect 16850 21972 16856 21984
rect 16908 22012 16914 22024
rect 17402 22012 17408 22024
rect 16908 21984 17408 22012
rect 16908 21972 16914 21984
rect 17402 21972 17408 21984
rect 17460 21972 17466 22024
rect 18230 22012 18236 22024
rect 18156 21984 18236 22012
rect 3145 21947 3203 21953
rect 3145 21913 3157 21947
rect 3191 21944 3203 21947
rect 3973 21947 4031 21953
rect 3973 21944 3985 21947
rect 3191 21916 3985 21944
rect 3191 21913 3203 21916
rect 3145 21907 3203 21913
rect 3973 21913 3985 21916
rect 4019 21913 4031 21947
rect 3973 21907 4031 21913
rect 13906 21904 13912 21956
rect 13964 21944 13970 21956
rect 14277 21947 14335 21953
rect 14277 21944 14289 21947
rect 13964 21916 14289 21944
rect 13964 21904 13970 21916
rect 14277 21913 14289 21916
rect 14323 21913 14335 21947
rect 14277 21907 14335 21913
rect 17120 21947 17178 21953
rect 17120 21913 17132 21947
rect 17166 21944 17178 21947
rect 18156 21944 18184 21984
rect 18230 21972 18236 21984
rect 18288 21972 18294 22024
rect 19260 22021 19288 22052
rect 19352 22052 21824 22080
rect 19245 22015 19303 22021
rect 19245 21981 19257 22015
rect 19291 21981 19303 22015
rect 19245 21975 19303 21981
rect 17166 21916 18184 21944
rect 17166 21913 17178 21916
rect 17120 21907 17178 21913
rect 18690 21904 18696 21956
rect 18748 21944 18754 21956
rect 19352 21944 19380 22052
rect 21818 22040 21824 22052
rect 21876 22080 21882 22092
rect 22094 22080 22100 22092
rect 21876 22052 22100 22080
rect 21876 22040 21882 22052
rect 22094 22040 22100 22052
rect 22152 22040 22158 22092
rect 24688 22089 24716 22188
rect 25038 22176 25044 22188
rect 25096 22176 25102 22228
rect 25406 22176 25412 22228
rect 25464 22216 25470 22228
rect 27338 22216 27344 22228
rect 25464 22188 27344 22216
rect 25464 22176 25470 22188
rect 27338 22176 27344 22188
rect 27396 22176 27402 22228
rect 30650 22176 30656 22228
rect 30708 22216 30714 22228
rect 32030 22216 32036 22228
rect 30708 22188 32036 22216
rect 30708 22176 30714 22188
rect 32030 22176 32036 22188
rect 32088 22216 32094 22228
rect 34057 22219 34115 22225
rect 34057 22216 34069 22219
rect 32088 22188 34069 22216
rect 32088 22176 32094 22188
rect 34057 22185 34069 22188
rect 34103 22185 34115 22219
rect 34057 22179 34115 22185
rect 40497 22219 40555 22225
rect 40497 22185 40509 22219
rect 40543 22216 40555 22219
rect 41322 22216 41328 22228
rect 40543 22188 41328 22216
rect 40543 22185 40555 22188
rect 40497 22179 40555 22185
rect 41322 22176 41328 22188
rect 41380 22176 41386 22228
rect 42058 22216 42064 22228
rect 42019 22188 42064 22216
rect 42058 22176 42064 22188
rect 42116 22176 42122 22228
rect 42168 22188 46934 22216
rect 30374 22108 30380 22160
rect 30432 22148 30438 22160
rect 31570 22148 31576 22160
rect 30432 22120 31576 22148
rect 30432 22108 30438 22120
rect 31570 22108 31576 22120
rect 31628 22148 31634 22160
rect 31757 22151 31815 22157
rect 31757 22148 31769 22151
rect 31628 22120 31769 22148
rect 31628 22108 31634 22120
rect 31757 22117 31769 22120
rect 31803 22117 31815 22151
rect 41141 22151 41199 22157
rect 41141 22148 41153 22151
rect 31757 22111 31815 22117
rect 40604 22120 41153 22148
rect 24673 22083 24731 22089
rect 24673 22049 24685 22083
rect 24719 22049 24731 22083
rect 24673 22043 24731 22049
rect 25682 22040 25688 22092
rect 25740 22080 25746 22092
rect 28445 22083 28503 22089
rect 25740 22052 27660 22080
rect 25740 22040 25746 22052
rect 27203 22015 27261 22021
rect 27203 21981 27215 22015
rect 27249 21981 27261 22015
rect 27338 22012 27344 22024
rect 27299 21984 27344 22012
rect 27203 21975 27261 21981
rect 18748 21916 19380 21944
rect 19429 21947 19487 21953
rect 18748 21904 18754 21916
rect 19429 21913 19441 21947
rect 19475 21944 19487 21947
rect 20530 21944 20536 21956
rect 19475 21916 20536 21944
rect 19475 21913 19487 21916
rect 19429 21907 19487 21913
rect 18506 21836 18512 21888
rect 18564 21876 18570 21888
rect 19444 21876 19472 21907
rect 20530 21904 20536 21916
rect 20588 21904 20594 21956
rect 20714 21904 20720 21956
rect 20772 21944 20778 21956
rect 23566 21944 23572 21956
rect 20772 21916 23572 21944
rect 20772 21904 20778 21916
rect 23566 21904 23572 21916
rect 23624 21904 23630 21956
rect 24946 21953 24952 21956
rect 24940 21944 24952 21953
rect 24907 21916 24952 21944
rect 24940 21907 24952 21916
rect 24946 21904 24952 21907
rect 25004 21904 25010 21956
rect 27218 21944 27246 21975
rect 27338 21972 27344 21984
rect 27396 21972 27402 22024
rect 27433 22015 27491 22021
rect 27433 21981 27445 22015
rect 27479 22012 27491 22015
rect 27522 22012 27528 22024
rect 27479 21984 27528 22012
rect 27479 21981 27491 21984
rect 27433 21975 27491 21981
rect 27522 21972 27528 21984
rect 27580 21972 27586 22024
rect 27632 22021 27660 22052
rect 28445 22049 28457 22083
rect 28491 22080 28503 22083
rect 28810 22080 28816 22092
rect 28491 22052 28816 22080
rect 28491 22049 28503 22052
rect 28445 22043 28503 22049
rect 28810 22040 28816 22052
rect 28868 22040 28874 22092
rect 36814 22080 36820 22092
rect 36775 22052 36820 22080
rect 36814 22040 36820 22052
rect 36872 22040 36878 22092
rect 37182 22040 37188 22092
rect 37240 22080 37246 22092
rect 40604 22080 40632 22120
rect 41141 22117 41153 22120
rect 41187 22117 41199 22151
rect 41141 22111 41199 22117
rect 42168 22080 42196 22188
rect 42245 22151 42303 22157
rect 42245 22117 42257 22151
rect 42291 22148 42303 22151
rect 43438 22148 43444 22160
rect 42291 22120 43444 22148
rect 42291 22117 42303 22120
rect 42245 22111 42303 22117
rect 43438 22108 43444 22120
rect 43496 22108 43502 22160
rect 37240 22052 40632 22080
rect 41248 22052 42196 22080
rect 37240 22040 37246 22052
rect 27617 22015 27675 22021
rect 27617 21981 27629 22015
rect 27663 21981 27675 22015
rect 28166 22012 28172 22024
rect 28127 21984 28172 22012
rect 27617 21975 27675 21981
rect 28166 21972 28172 21984
rect 28224 21972 28230 22024
rect 28258 21972 28264 22024
rect 28316 22012 28322 22024
rect 31018 22012 31024 22024
rect 28316 21984 31024 22012
rect 28316 21972 28322 21984
rect 31018 21972 31024 21984
rect 31076 22012 31082 22024
rect 32582 22012 32588 22024
rect 31076 21984 32588 22012
rect 31076 21972 31082 21984
rect 32582 21972 32588 21984
rect 32640 21972 32646 22024
rect 32677 22015 32735 22021
rect 32677 21981 32689 22015
rect 32723 22012 32735 22015
rect 34698 22012 34704 22024
rect 32723 21984 34704 22012
rect 32723 21981 32735 21984
rect 32677 21975 32735 21981
rect 34698 21972 34704 21984
rect 34756 21972 34762 22024
rect 36170 22012 36176 22024
rect 36131 21984 36176 22012
rect 36170 21972 36176 21984
rect 36228 21972 36234 22024
rect 36262 21972 36268 22024
rect 36320 22012 36326 22024
rect 36357 22015 36415 22021
rect 36357 22012 36369 22015
rect 36320 21984 36369 22012
rect 36320 21972 36326 21984
rect 36357 21981 36369 21984
rect 36403 21981 36415 22015
rect 36357 21975 36415 21981
rect 37093 22015 37151 22021
rect 37093 21981 37105 22015
rect 37139 22012 37151 22015
rect 37826 22012 37832 22024
rect 37139 21984 37832 22012
rect 37139 21981 37151 21984
rect 37093 21975 37151 21981
rect 37826 21972 37832 21984
rect 37884 21972 37890 22024
rect 40405 22015 40463 22021
rect 40405 21981 40417 22015
rect 40451 22012 40463 22015
rect 40494 22012 40500 22024
rect 40451 21984 40500 22012
rect 40451 21981 40463 21984
rect 40405 21975 40463 21981
rect 40494 21972 40500 21984
rect 40552 21972 40558 22024
rect 41138 22012 41144 22024
rect 41099 21984 41144 22012
rect 41138 21972 41144 21984
rect 41196 21972 41202 22024
rect 30466 21944 30472 21956
rect 27218 21916 29500 21944
rect 30427 21916 30472 21944
rect 18564 21848 19472 21876
rect 19613 21879 19671 21885
rect 18564 21836 18570 21848
rect 19613 21845 19625 21879
rect 19659 21876 19671 21879
rect 19978 21876 19984 21888
rect 19659 21848 19984 21876
rect 19659 21845 19671 21848
rect 19613 21839 19671 21845
rect 19978 21836 19984 21848
rect 20036 21836 20042 21888
rect 25682 21836 25688 21888
rect 25740 21876 25746 21888
rect 26053 21879 26111 21885
rect 26053 21876 26065 21879
rect 25740 21848 26065 21876
rect 25740 21836 25746 21848
rect 26053 21845 26065 21848
rect 26099 21845 26111 21879
rect 26053 21839 26111 21845
rect 26973 21879 27031 21885
rect 26973 21845 26985 21879
rect 27019 21876 27031 21879
rect 27430 21876 27436 21888
rect 27019 21848 27436 21876
rect 27019 21845 27031 21848
rect 26973 21839 27031 21845
rect 27430 21836 27436 21848
rect 27488 21836 27494 21888
rect 28166 21836 28172 21888
rect 28224 21876 28230 21888
rect 28994 21876 29000 21888
rect 28224 21848 29000 21876
rect 28224 21836 28230 21848
rect 28994 21836 29000 21848
rect 29052 21836 29058 21888
rect 29472 21876 29500 21916
rect 30466 21904 30472 21916
rect 30524 21904 30530 21956
rect 32214 21904 32220 21956
rect 32272 21944 32278 21956
rect 32922 21947 32980 21953
rect 32922 21944 32934 21947
rect 32272 21916 32934 21944
rect 32272 21904 32278 21916
rect 32922 21913 32934 21916
rect 32968 21913 32980 21947
rect 41248 21944 41276 22052
rect 44174 22040 44180 22092
rect 44232 22080 44238 22092
rect 45097 22083 45155 22089
rect 45097 22080 45109 22083
rect 44232 22052 45109 22080
rect 44232 22040 44238 22052
rect 45097 22049 45109 22052
rect 45143 22049 45155 22083
rect 45097 22043 45155 22049
rect 41325 22015 41383 22021
rect 41325 21981 41337 22015
rect 41371 22012 41383 22015
rect 42518 22012 42524 22024
rect 41371 21984 42524 22012
rect 41371 21981 41383 21984
rect 41325 21975 41383 21981
rect 42518 21972 42524 21984
rect 42576 21972 42582 22024
rect 42610 21972 42616 22024
rect 42668 22012 42674 22024
rect 43211 22015 43269 22021
rect 43211 22012 43223 22015
rect 42668 21984 43223 22012
rect 42668 21972 42674 21984
rect 43211 21981 43223 21984
rect 43257 21981 43269 22015
rect 43346 22012 43352 22024
rect 43307 21984 43352 22012
rect 43211 21975 43269 21981
rect 43346 21972 43352 21984
rect 43404 21972 43410 22024
rect 43438 21972 43444 22024
rect 43496 22021 43502 22024
rect 43496 22012 43504 22021
rect 43625 22015 43683 22021
rect 43496 21984 43541 22012
rect 43496 21975 43504 21984
rect 43625 21981 43637 22015
rect 43671 21981 43683 22015
rect 46906 22012 46934 22188
rect 48133 22015 48191 22021
rect 48133 22012 48145 22015
rect 46906 21984 48145 22012
rect 43625 21975 43683 21981
rect 48133 21981 48145 21984
rect 48179 21981 48191 22015
rect 48133 21975 48191 21981
rect 43496 21972 43502 21975
rect 32922 21907 32980 21913
rect 36188 21916 41276 21944
rect 36188 21876 36216 21916
rect 41414 21904 41420 21956
rect 41472 21944 41478 21956
rect 41782 21944 41788 21956
rect 41472 21916 41788 21944
rect 41472 21904 41478 21916
rect 41782 21904 41788 21916
rect 41840 21944 41846 21956
rect 41877 21947 41935 21953
rect 41877 21944 41889 21947
rect 41840 21916 41889 21944
rect 41840 21904 41846 21916
rect 41877 21913 41889 21916
rect 41923 21913 41935 21947
rect 41877 21907 41935 21913
rect 41966 21904 41972 21956
rect 42024 21944 42030 21956
rect 42077 21947 42135 21953
rect 42077 21944 42089 21947
rect 42024 21916 42089 21944
rect 42024 21904 42030 21916
rect 42077 21913 42089 21916
rect 42123 21913 42135 21947
rect 42077 21907 42135 21913
rect 42426 21904 42432 21956
rect 42484 21944 42490 21956
rect 43640 21944 43668 21975
rect 42484 21916 43668 21944
rect 42484 21904 42490 21916
rect 44450 21904 44456 21956
rect 44508 21944 44514 21956
rect 45342 21947 45400 21953
rect 45342 21944 45354 21947
rect 44508 21916 45354 21944
rect 44508 21904 44514 21916
rect 45342 21913 45354 21916
rect 45388 21913 45400 21947
rect 47946 21944 47952 21956
rect 47907 21916 47952 21944
rect 45342 21907 45400 21913
rect 47946 21904 47952 21916
rect 48004 21904 48010 21956
rect 36354 21876 36360 21888
rect 29472 21848 36216 21876
rect 36315 21848 36360 21876
rect 36354 21836 36360 21848
rect 36412 21836 36418 21888
rect 42981 21879 43039 21885
rect 42981 21845 42993 21879
rect 43027 21876 43039 21879
rect 43622 21876 43628 21888
rect 43027 21848 43628 21876
rect 43027 21845 43039 21848
rect 42981 21839 43039 21845
rect 43622 21836 43628 21848
rect 43680 21836 43686 21888
rect 46106 21836 46112 21888
rect 46164 21876 46170 21888
rect 46474 21876 46480 21888
rect 46164 21848 46480 21876
rect 46164 21836 46170 21848
rect 46474 21836 46480 21848
rect 46532 21836 46538 21888
rect 1104 21786 48852 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 48852 21786
rect 1104 21712 48852 21734
rect 3786 21632 3792 21684
rect 3844 21672 3850 21684
rect 13722 21672 13728 21684
rect 3844 21644 13728 21672
rect 3844 21632 3850 21644
rect 13722 21632 13728 21644
rect 13780 21632 13786 21684
rect 13906 21672 13912 21684
rect 13867 21644 13912 21672
rect 13906 21632 13912 21644
rect 13964 21632 13970 21684
rect 24946 21672 24952 21684
rect 14476 21644 24952 21672
rect 3510 21604 3516 21616
rect 3471 21576 3516 21604
rect 3510 21564 3516 21576
rect 3568 21564 3574 21616
rect 14476 21604 14504 21644
rect 24946 21632 24952 21644
rect 25004 21632 25010 21684
rect 30650 21672 30656 21684
rect 25056 21644 30656 21672
rect 16574 21604 16580 21616
rect 5092 21576 14504 21604
rect 14936 21576 16580 21604
rect 2498 21496 2504 21548
rect 2556 21496 2562 21548
rect 2516 21332 2544 21496
rect 3329 21471 3387 21477
rect 3329 21437 3341 21471
rect 3375 21468 3387 21471
rect 5092 21468 5120 21576
rect 14936 21548 14964 21576
rect 16574 21564 16580 21576
rect 16632 21604 16638 21616
rect 17037 21607 17095 21613
rect 17037 21604 17049 21607
rect 16632 21576 17049 21604
rect 16632 21564 16638 21576
rect 17037 21573 17049 21576
rect 17083 21573 17095 21607
rect 17037 21567 17095 21573
rect 18322 21564 18328 21616
rect 18380 21604 18386 21616
rect 18690 21604 18696 21616
rect 18380 21576 18696 21604
rect 18380 21564 18386 21576
rect 18690 21564 18696 21576
rect 18748 21564 18754 21616
rect 19334 21564 19340 21616
rect 19392 21604 19398 21616
rect 19490 21607 19548 21613
rect 19490 21604 19502 21607
rect 19392 21576 19502 21604
rect 19392 21564 19398 21576
rect 19490 21573 19502 21576
rect 19536 21573 19548 21607
rect 25056 21604 25084 21644
rect 30650 21632 30656 21644
rect 30708 21632 30714 21684
rect 30742 21632 30748 21684
rect 30800 21672 30806 21684
rect 31110 21672 31116 21684
rect 30800 21644 31116 21672
rect 30800 21632 30806 21644
rect 31110 21632 31116 21644
rect 31168 21672 31174 21684
rect 31481 21675 31539 21681
rect 31481 21672 31493 21675
rect 31168 21644 31493 21672
rect 31168 21632 31174 21644
rect 31481 21641 31493 21644
rect 31527 21641 31539 21675
rect 31481 21635 31539 21641
rect 33042 21632 33048 21684
rect 33100 21672 33106 21684
rect 36170 21672 36176 21684
rect 33100 21644 36176 21672
rect 33100 21632 33106 21644
rect 36170 21632 36176 21644
rect 36228 21632 36234 21684
rect 36354 21632 36360 21684
rect 36412 21672 36418 21684
rect 37855 21675 37913 21681
rect 37855 21672 37867 21675
rect 36412 21644 37867 21672
rect 36412 21632 36418 21644
rect 37855 21641 37867 21644
rect 37901 21672 37913 21675
rect 37901 21644 38792 21672
rect 37901 21641 37913 21644
rect 37855 21635 37913 21641
rect 30190 21604 30196 21616
rect 19490 21567 19548 21573
rect 23124 21576 25084 21604
rect 27356 21576 30196 21604
rect 13814 21536 13820 21548
rect 13775 21508 13820 21536
rect 13814 21496 13820 21508
rect 13872 21496 13878 21548
rect 14918 21536 14924 21548
rect 14831 21508 14924 21536
rect 14918 21496 14924 21508
rect 14976 21496 14982 21548
rect 17402 21496 17408 21548
rect 17460 21536 17466 21548
rect 19245 21539 19303 21545
rect 19245 21536 19257 21539
rect 17460 21508 19257 21536
rect 17460 21496 17466 21508
rect 19245 21505 19257 21508
rect 19291 21505 19303 21539
rect 21634 21536 21640 21548
rect 19245 21499 19303 21505
rect 19352 21508 21640 21536
rect 3375 21440 5120 21468
rect 3375 21437 3387 21440
rect 3329 21431 3387 21437
rect 5166 21428 5172 21480
rect 5224 21468 5230 21480
rect 5224 21440 5269 21468
rect 5224 21428 5230 21440
rect 15470 21428 15476 21480
rect 15528 21468 15534 21480
rect 15933 21471 15991 21477
rect 15933 21468 15945 21471
rect 15528 21440 15945 21468
rect 15528 21428 15534 21440
rect 15933 21437 15945 21440
rect 15979 21468 15991 21471
rect 19352 21468 19380 21508
rect 21634 21496 21640 21508
rect 21692 21496 21698 21548
rect 21726 21496 21732 21548
rect 21784 21536 21790 21548
rect 21821 21539 21879 21545
rect 21821 21536 21833 21539
rect 21784 21508 21833 21536
rect 21784 21496 21790 21508
rect 21821 21505 21833 21508
rect 21867 21505 21879 21539
rect 21821 21499 21879 21505
rect 21910 21496 21916 21548
rect 21968 21536 21974 21548
rect 22077 21539 22135 21545
rect 22077 21536 22089 21539
rect 21968 21508 22089 21536
rect 21968 21496 21974 21508
rect 22077 21505 22089 21508
rect 22123 21505 22135 21539
rect 22077 21499 22135 21505
rect 15979 21440 19380 21468
rect 15979 21437 15991 21440
rect 15933 21431 15991 21437
rect 13722 21360 13728 21412
rect 13780 21400 13786 21412
rect 13780 21372 18460 21400
rect 13780 21360 13786 21372
rect 18322 21332 18328 21344
rect 2516 21304 18328 21332
rect 18322 21292 18328 21304
rect 18380 21292 18386 21344
rect 18432 21332 18460 21372
rect 20530 21360 20536 21412
rect 20588 21400 20594 21412
rect 20625 21403 20683 21409
rect 20625 21400 20637 21403
rect 20588 21372 20637 21400
rect 20588 21360 20594 21372
rect 20625 21369 20637 21372
rect 20671 21369 20683 21403
rect 20625 21363 20683 21369
rect 23124 21332 23152 21576
rect 23566 21496 23572 21548
rect 23624 21536 23630 21548
rect 23845 21539 23903 21545
rect 23845 21536 23857 21539
rect 23624 21508 23857 21536
rect 23624 21496 23630 21508
rect 23845 21505 23857 21508
rect 23891 21505 23903 21539
rect 24029 21539 24087 21545
rect 24029 21536 24041 21539
rect 23845 21499 23903 21505
rect 23952 21508 24041 21536
rect 23952 21468 23980 21508
rect 24029 21505 24041 21508
rect 24075 21505 24087 21539
rect 24029 21499 24087 21505
rect 24118 21496 24124 21548
rect 24176 21536 24182 21548
rect 25038 21536 25044 21548
rect 24176 21508 24221 21536
rect 24999 21508 25044 21536
rect 24176 21496 24182 21508
rect 25038 21496 25044 21508
rect 25096 21496 25102 21548
rect 25314 21545 25320 21548
rect 25308 21499 25320 21545
rect 25372 21536 25378 21548
rect 27356 21545 27384 21576
rect 27341 21539 27399 21545
rect 25372 21508 25408 21536
rect 25314 21496 25320 21499
rect 25372 21496 25378 21508
rect 27341 21505 27353 21539
rect 27387 21505 27399 21539
rect 27341 21499 27399 21505
rect 27430 21496 27436 21548
rect 27488 21536 27494 21548
rect 27597 21539 27655 21545
rect 27597 21536 27609 21539
rect 27488 21508 27609 21536
rect 27488 21496 27494 21508
rect 27597 21505 27609 21508
rect 27643 21505 27655 21539
rect 27597 21499 27655 21505
rect 28534 21496 28540 21548
rect 28592 21536 28598 21548
rect 28718 21536 28724 21548
rect 28592 21508 28724 21536
rect 28592 21496 28598 21508
rect 28718 21496 28724 21508
rect 28776 21536 28782 21548
rect 29181 21539 29239 21545
rect 29181 21536 29193 21539
rect 28776 21508 29193 21536
rect 28776 21496 28782 21508
rect 29181 21505 29193 21508
rect 29227 21505 29239 21539
rect 29181 21499 29239 21505
rect 29365 21539 29423 21545
rect 29365 21505 29377 21539
rect 29411 21536 29423 21539
rect 29546 21536 29552 21548
rect 29411 21508 29552 21536
rect 29411 21505 29423 21508
rect 29365 21499 29423 21505
rect 29546 21496 29552 21508
rect 29604 21496 29610 21548
rect 30116 21545 30144 21576
rect 30190 21564 30196 21576
rect 30248 21564 30254 21616
rect 30368 21607 30426 21613
rect 30368 21573 30380 21607
rect 30414 21604 30426 21607
rect 30926 21604 30932 21616
rect 30414 21576 30932 21604
rect 30414 21573 30426 21576
rect 30368 21567 30426 21573
rect 30926 21564 30932 21576
rect 30984 21564 30990 21616
rect 32769 21607 32827 21613
rect 32048 21576 32444 21604
rect 30101 21539 30159 21545
rect 30101 21505 30113 21539
rect 30147 21505 30159 21539
rect 32048 21536 32076 21576
rect 30101 21499 30159 21505
rect 30208 21508 32076 21536
rect 30208 21468 30236 21508
rect 32122 21496 32128 21548
rect 32180 21536 32186 21548
rect 32309 21539 32367 21545
rect 32309 21536 32321 21539
rect 32180 21508 32321 21536
rect 32180 21496 32186 21508
rect 32309 21505 32321 21508
rect 32355 21505 32367 21539
rect 32416 21536 32444 21576
rect 32769 21573 32781 21607
rect 32815 21604 32827 21607
rect 34118 21607 34176 21613
rect 34118 21604 34130 21607
rect 32815 21576 34130 21604
rect 32815 21573 32827 21576
rect 32769 21567 32827 21573
rect 34118 21573 34130 21576
rect 34164 21573 34176 21607
rect 34118 21567 34176 21573
rect 37645 21607 37703 21613
rect 37645 21573 37657 21607
rect 37691 21604 37703 21607
rect 38286 21604 38292 21616
rect 37691 21576 38292 21604
rect 37691 21573 37703 21576
rect 37645 21567 37703 21573
rect 38286 21564 38292 21576
rect 38344 21564 38350 21616
rect 38657 21607 38715 21613
rect 38657 21604 38669 21607
rect 38396 21576 38669 21604
rect 32999 21539 33057 21545
rect 32999 21536 33011 21539
rect 32416 21508 33011 21536
rect 32309 21499 32367 21505
rect 32999 21505 33011 21508
rect 33045 21505 33057 21539
rect 33134 21536 33140 21548
rect 33095 21508 33140 21536
rect 32999 21499 33057 21505
rect 33134 21496 33140 21508
rect 33192 21496 33198 21548
rect 33226 21496 33232 21548
rect 33284 21536 33290 21548
rect 33284 21508 33329 21536
rect 33284 21496 33290 21508
rect 33410 21496 33416 21548
rect 33468 21536 33474 21548
rect 33468 21508 33513 21536
rect 33468 21496 33474 21508
rect 37826 21496 37832 21548
rect 37884 21536 37890 21548
rect 38396 21536 38424 21576
rect 38657 21573 38669 21576
rect 38703 21573 38715 21607
rect 38657 21567 38715 21573
rect 38764 21567 38792 21644
rect 40770 21632 40776 21684
rect 40828 21672 40834 21684
rect 42426 21672 42432 21684
rect 40828 21644 42432 21672
rect 40828 21632 40834 21644
rect 42426 21632 42432 21644
rect 42484 21632 42490 21684
rect 46842 21672 46848 21684
rect 46803 21644 46848 21672
rect 46842 21632 46848 21644
rect 46900 21632 46906 21684
rect 40957 21607 41015 21613
rect 40957 21573 40969 21607
rect 41003 21604 41015 21607
rect 41322 21604 41328 21616
rect 41003 21576 41328 21604
rect 41003 21573 41015 21576
rect 40957 21567 41015 21573
rect 38758 21561 38816 21567
rect 41322 21564 41328 21576
rect 41380 21564 41386 21616
rect 43548 21576 45508 21604
rect 37884 21508 38424 21536
rect 38473 21539 38531 21545
rect 37884 21496 37890 21508
rect 38473 21505 38485 21539
rect 38519 21505 38531 21539
rect 38758 21527 38770 21561
rect 38804 21527 38816 21561
rect 40862 21536 40868 21548
rect 38758 21521 38816 21527
rect 38473 21499 38531 21505
rect 38856 21508 40868 21536
rect 23860 21440 23980 21468
rect 28966 21440 30236 21468
rect 23860 21412 23888 21440
rect 23842 21360 23848 21412
rect 23900 21360 23906 21412
rect 18432 21304 23152 21332
rect 23201 21335 23259 21341
rect 23201 21301 23213 21335
rect 23247 21332 23259 21335
rect 23290 21332 23296 21344
rect 23247 21304 23296 21332
rect 23247 21301 23259 21304
rect 23201 21295 23259 21301
rect 23290 21292 23296 21304
rect 23348 21292 23354 21344
rect 23474 21292 23480 21344
rect 23532 21332 23538 21344
rect 23661 21335 23719 21341
rect 23661 21332 23673 21335
rect 23532 21304 23673 21332
rect 23532 21292 23538 21304
rect 23661 21301 23673 21304
rect 23707 21301 23719 21335
rect 23661 21295 23719 21301
rect 26234 21292 26240 21344
rect 26292 21332 26298 21344
rect 26421 21335 26479 21341
rect 26421 21332 26433 21335
rect 26292 21304 26433 21332
rect 26292 21292 26298 21304
rect 26421 21301 26433 21304
rect 26467 21301 26479 21335
rect 26421 21295 26479 21301
rect 27154 21292 27160 21344
rect 27212 21332 27218 21344
rect 28721 21335 28779 21341
rect 28721 21332 28733 21335
rect 27212 21304 28733 21332
rect 27212 21292 27218 21304
rect 28721 21301 28733 21304
rect 28767 21332 28779 21335
rect 28966 21332 28994 21440
rect 32766 21428 32772 21480
rect 32824 21468 32830 21480
rect 33873 21471 33931 21477
rect 33873 21468 33885 21471
rect 32824 21440 33885 21468
rect 32824 21428 32830 21440
rect 33873 21437 33885 21440
rect 33919 21437 33931 21471
rect 38010 21468 38016 21480
rect 33873 21431 33931 21437
rect 35268 21440 38016 21468
rect 35268 21409 35296 21440
rect 38010 21428 38016 21440
rect 38068 21428 38074 21480
rect 38488 21468 38516 21499
rect 38856 21468 38884 21508
rect 40862 21496 40868 21508
rect 40920 21496 40926 21548
rect 38488 21440 38884 21468
rect 40218 21428 40224 21480
rect 40276 21468 40282 21480
rect 43548 21477 43576 21576
rect 43622 21496 43628 21548
rect 43680 21536 43686 21548
rect 45480 21545 45508 21576
rect 45738 21545 45744 21548
rect 43789 21539 43847 21545
rect 43789 21536 43801 21539
rect 43680 21508 43801 21536
rect 43680 21496 43686 21508
rect 43789 21505 43801 21508
rect 43835 21505 43847 21539
rect 43789 21499 43847 21505
rect 45465 21539 45523 21545
rect 45465 21505 45477 21539
rect 45511 21505 45523 21539
rect 45465 21499 45523 21505
rect 45732 21499 45744 21545
rect 45796 21536 45802 21548
rect 45796 21508 45832 21536
rect 45738 21496 45744 21499
rect 45796 21496 45802 21508
rect 43533 21471 43591 21477
rect 43533 21468 43545 21471
rect 40276 21440 43545 21468
rect 40276 21428 40282 21440
rect 43533 21437 43545 21440
rect 43579 21437 43591 21471
rect 43533 21431 43591 21437
rect 35253 21403 35311 21409
rect 35253 21369 35265 21403
rect 35299 21400 35311 21403
rect 35342 21400 35348 21412
rect 35299 21372 35348 21400
rect 35299 21369 35311 21372
rect 35253 21363 35311 21369
rect 35342 21360 35348 21372
rect 35400 21360 35406 21412
rect 37734 21360 37740 21412
rect 37792 21400 37798 21412
rect 38473 21403 38531 21409
rect 38473 21400 38485 21403
rect 37792 21372 38485 21400
rect 37792 21360 37798 21372
rect 38473 21369 38485 21372
rect 38519 21369 38531 21403
rect 38473 21363 38531 21369
rect 40589 21403 40647 21409
rect 40589 21369 40601 21403
rect 40635 21400 40647 21403
rect 40678 21400 40684 21412
rect 40635 21372 40684 21400
rect 40635 21369 40647 21372
rect 40589 21363 40647 21369
rect 40678 21360 40684 21372
rect 40736 21360 40742 21412
rect 29546 21332 29552 21344
rect 28767 21304 28994 21332
rect 29507 21304 29552 21332
rect 28767 21301 28779 21304
rect 28721 21295 28779 21301
rect 29546 21292 29552 21304
rect 29604 21292 29610 21344
rect 31938 21292 31944 21344
rect 31996 21332 32002 21344
rect 32125 21335 32183 21341
rect 32125 21332 32137 21335
rect 31996 21304 32137 21332
rect 31996 21292 32002 21304
rect 32125 21301 32137 21304
rect 32171 21332 32183 21335
rect 34790 21332 34796 21344
rect 32171 21304 34796 21332
rect 32171 21301 32183 21304
rect 32125 21295 32183 21301
rect 34790 21292 34796 21304
rect 34848 21292 34854 21344
rect 37274 21292 37280 21344
rect 37332 21332 37338 21344
rect 37826 21332 37832 21344
rect 37332 21304 37832 21332
rect 37332 21292 37338 21304
rect 37826 21292 37832 21304
rect 37884 21292 37890 21344
rect 38010 21332 38016 21344
rect 37971 21304 38016 21332
rect 38010 21292 38016 21304
rect 38068 21292 38074 21344
rect 38930 21292 38936 21344
rect 38988 21332 38994 21344
rect 40402 21332 40408 21344
rect 38988 21304 40408 21332
rect 38988 21292 38994 21304
rect 40402 21292 40408 21304
rect 40460 21292 40466 21344
rect 40954 21332 40960 21344
rect 40915 21304 40960 21332
rect 40954 21292 40960 21304
rect 41012 21292 41018 21344
rect 41141 21335 41199 21341
rect 41141 21301 41153 21335
rect 41187 21332 41199 21335
rect 41874 21332 41880 21344
rect 41187 21304 41880 21332
rect 41187 21301 41199 21304
rect 41141 21295 41199 21301
rect 41874 21292 41880 21304
rect 41932 21292 41938 21344
rect 44910 21332 44916 21344
rect 44871 21304 44916 21332
rect 44910 21292 44916 21304
rect 44968 21292 44974 21344
rect 47762 21332 47768 21344
rect 47723 21304 47768 21332
rect 47762 21292 47768 21304
rect 47820 21292 47826 21344
rect 1104 21242 48852 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 48852 21242
rect 1104 21168 48852 21190
rect 19245 21131 19303 21137
rect 19245 21097 19257 21131
rect 19291 21128 19303 21131
rect 19334 21128 19340 21140
rect 19291 21100 19340 21128
rect 19291 21097 19303 21100
rect 19245 21091 19303 21097
rect 19334 21088 19340 21100
rect 19392 21088 19398 21140
rect 21177 21131 21235 21137
rect 21177 21128 21189 21131
rect 19444 21100 21189 21128
rect 15654 21020 15660 21072
rect 15712 21060 15718 21072
rect 18046 21060 18052 21072
rect 15712 21032 18052 21060
rect 15712 21020 15718 21032
rect 18046 21020 18052 21032
rect 18104 21020 18110 21072
rect 18874 21020 18880 21072
rect 18932 21060 18938 21072
rect 19444 21060 19472 21100
rect 21177 21097 21189 21100
rect 21223 21097 21235 21131
rect 21910 21128 21916 21140
rect 21871 21100 21916 21128
rect 21177 21091 21235 21097
rect 21910 21088 21916 21100
rect 21968 21088 21974 21140
rect 33042 21128 33048 21140
rect 22066 21100 33048 21128
rect 22066 21060 22094 21100
rect 33042 21088 33048 21100
rect 33100 21088 33106 21140
rect 33134 21088 33140 21140
rect 33192 21128 33198 21140
rect 35069 21131 35127 21137
rect 35069 21128 35081 21131
rect 33192 21100 35081 21128
rect 33192 21088 33198 21100
rect 35069 21097 35081 21100
rect 35115 21097 35127 21131
rect 35069 21091 35127 21097
rect 37550 21088 37556 21140
rect 37608 21128 37614 21140
rect 37645 21131 37703 21137
rect 37645 21128 37657 21131
rect 37608 21100 37657 21128
rect 37608 21088 37614 21100
rect 37645 21097 37657 21100
rect 37691 21097 37703 21131
rect 37645 21091 37703 21097
rect 37734 21088 37740 21140
rect 37792 21128 37798 21140
rect 37792 21100 37837 21128
rect 37792 21088 37798 21100
rect 38286 21088 38292 21140
rect 38344 21128 38350 21140
rect 40126 21128 40132 21140
rect 38344 21100 40132 21128
rect 38344 21088 38350 21100
rect 40126 21088 40132 21100
rect 40184 21128 40190 21140
rect 41233 21131 41291 21137
rect 41233 21128 41245 21131
rect 40184 21100 41245 21128
rect 40184 21088 40190 21100
rect 41233 21097 41245 21100
rect 41279 21097 41291 21131
rect 41233 21091 41291 21097
rect 43438 21088 43444 21140
rect 43496 21128 43502 21140
rect 44453 21131 44511 21137
rect 44453 21128 44465 21131
rect 43496 21100 44465 21128
rect 43496 21088 43502 21100
rect 44453 21097 44465 21100
rect 44499 21097 44511 21131
rect 44453 21091 44511 21097
rect 45005 21131 45063 21137
rect 45005 21097 45017 21131
rect 45051 21128 45063 21131
rect 45738 21128 45744 21140
rect 45051 21100 45744 21128
rect 45051 21097 45063 21100
rect 45005 21091 45063 21097
rect 45738 21088 45744 21100
rect 45796 21088 45802 21140
rect 18932 21032 19472 21060
rect 19536 21032 22094 21060
rect 22833 21063 22891 21069
rect 18932 21020 18938 21032
rect 3418 20952 3424 21004
rect 3476 20992 3482 21004
rect 16577 20995 16635 21001
rect 16577 20992 16589 20995
rect 3476 20964 16589 20992
rect 3476 20952 3482 20964
rect 16577 20961 16589 20964
rect 16623 20961 16635 20995
rect 16577 20955 16635 20961
rect 14918 20924 14924 20936
rect 14879 20896 14924 20924
rect 14918 20884 14924 20896
rect 14976 20884 14982 20936
rect 16025 20927 16083 20933
rect 16025 20893 16037 20927
rect 16071 20893 16083 20927
rect 16025 20887 16083 20893
rect 15473 20859 15531 20865
rect 15473 20856 15485 20859
rect 12406 20828 15485 20856
rect 2406 20748 2412 20800
rect 2464 20788 2470 20800
rect 12406 20788 12434 20828
rect 15473 20825 15485 20828
rect 15519 20856 15531 20859
rect 15654 20856 15660 20868
rect 15519 20828 15660 20856
rect 15519 20825 15531 20828
rect 15473 20819 15531 20825
rect 15654 20816 15660 20828
rect 15712 20816 15718 20868
rect 2464 20760 12434 20788
rect 16040 20788 16068 20887
rect 17402 20884 17408 20936
rect 17460 20924 17466 20936
rect 19536 20933 19564 21032
rect 22833 21029 22845 21063
rect 22879 21029 22891 21063
rect 22833 21023 22891 21029
rect 25041 21063 25099 21069
rect 25041 21029 25053 21063
rect 25087 21060 25099 21063
rect 25314 21060 25320 21072
rect 25087 21032 25320 21060
rect 25087 21029 25099 21032
rect 25041 21023 25099 21029
rect 19978 20992 19984 21004
rect 19720 20964 19984 20992
rect 19720 20933 19748 20964
rect 19978 20952 19984 20964
rect 20036 20952 20042 21004
rect 18509 20927 18567 20933
rect 18509 20924 18521 20927
rect 17460 20896 18521 20924
rect 17460 20884 17466 20896
rect 18509 20893 18521 20896
rect 18555 20893 18567 20927
rect 18509 20887 18567 20893
rect 19521 20927 19579 20933
rect 19521 20893 19533 20927
rect 19567 20893 19579 20927
rect 19521 20887 19579 20893
rect 19613 20927 19671 20933
rect 19613 20893 19625 20927
rect 19659 20893 19671 20927
rect 19613 20887 19671 20893
rect 19705 20927 19763 20933
rect 19705 20893 19717 20927
rect 19751 20893 19763 20927
rect 19705 20887 19763 20893
rect 19889 20927 19947 20933
rect 19889 20893 19901 20927
rect 19935 20924 19947 20927
rect 20530 20924 20536 20936
rect 19935 20896 20536 20924
rect 19935 20893 19947 20896
rect 19889 20887 19947 20893
rect 16206 20856 16212 20868
rect 16167 20828 16212 20856
rect 16206 20816 16212 20828
rect 16264 20816 16270 20868
rect 18322 20856 18328 20868
rect 18283 20828 18328 20856
rect 18322 20816 18328 20828
rect 18380 20816 18386 20868
rect 18966 20816 18972 20868
rect 19024 20856 19030 20868
rect 19628 20856 19656 20887
rect 20530 20884 20536 20896
rect 20588 20884 20594 20936
rect 22094 20884 22100 20936
rect 22152 20924 22158 20936
rect 22278 20924 22284 20936
rect 22152 20896 22197 20924
rect 22239 20896 22284 20924
rect 22152 20884 22158 20896
rect 22278 20884 22284 20896
rect 22336 20884 22342 20936
rect 22373 20927 22431 20933
rect 22373 20893 22385 20927
rect 22419 20893 22431 20927
rect 22848 20924 22876 21023
rect 25314 21020 25320 21032
rect 25372 21020 25378 21072
rect 27154 21060 27160 21072
rect 25424 21032 27160 21060
rect 23382 20992 23388 21004
rect 23343 20964 23388 20992
rect 23382 20952 23388 20964
rect 23440 20952 23446 21004
rect 23566 20952 23572 21004
rect 23624 20992 23630 21004
rect 24118 20992 24124 21004
rect 23624 20964 24124 20992
rect 23624 20952 23630 20964
rect 24118 20952 24124 20964
rect 24176 20952 24182 21004
rect 25424 20992 25452 21032
rect 27154 21020 27160 21032
rect 27212 21020 27218 21072
rect 27341 21063 27399 21069
rect 27341 21029 27353 21063
rect 27387 21060 27399 21063
rect 27522 21060 27528 21072
rect 27387 21032 27528 21060
rect 27387 21029 27399 21032
rect 27341 21023 27399 21029
rect 27522 21020 27528 21032
rect 27580 21020 27586 21072
rect 36170 21020 36176 21072
rect 36228 21060 36234 21072
rect 37918 21060 37924 21072
rect 36228 21032 37924 21060
rect 36228 21020 36234 21032
rect 37918 21020 37924 21032
rect 37976 21020 37982 21072
rect 43346 21060 43352 21072
rect 42904 21032 43352 21060
rect 26513 20995 26571 21001
rect 26513 20992 26525 20995
rect 24780 20964 25452 20992
rect 25516 20964 26525 20992
rect 24397 20927 24455 20933
rect 24397 20924 24409 20927
rect 22848 20896 24409 20924
rect 22373 20887 22431 20893
rect 24397 20893 24409 20896
rect 24443 20893 24455 20927
rect 24397 20887 24455 20893
rect 19024 20828 19656 20856
rect 21085 20859 21143 20865
rect 19024 20816 19030 20828
rect 21085 20825 21097 20859
rect 21131 20856 21143 20859
rect 22388 20856 22416 20887
rect 23014 20856 23020 20868
rect 21131 20828 22094 20856
rect 22388 20828 23020 20856
rect 21131 20825 21143 20828
rect 21085 20819 21143 20825
rect 17402 20788 17408 20800
rect 16040 20760 17408 20788
rect 2464 20748 2470 20760
rect 17402 20748 17408 20760
rect 17460 20748 17466 20800
rect 18690 20788 18696 20800
rect 18651 20760 18696 20788
rect 18690 20748 18696 20760
rect 18748 20748 18754 20800
rect 22066 20788 22094 20828
rect 23014 20816 23020 20828
rect 23072 20856 23078 20868
rect 23290 20856 23296 20868
rect 23072 20828 23296 20856
rect 23072 20816 23078 20828
rect 23290 20816 23296 20828
rect 23348 20816 23354 20868
rect 23842 20856 23848 20868
rect 23492 20828 23848 20856
rect 23106 20788 23112 20800
rect 22066 20760 23112 20788
rect 23106 20748 23112 20760
rect 23164 20748 23170 20800
rect 23201 20791 23259 20797
rect 23201 20757 23213 20791
rect 23247 20788 23259 20791
rect 23492 20788 23520 20828
rect 23842 20816 23848 20828
rect 23900 20856 23906 20868
rect 24780 20856 24808 20964
rect 24854 20884 24860 20936
rect 24912 20924 24918 20936
rect 25271 20927 25329 20933
rect 25271 20924 25283 20927
rect 24912 20896 25283 20924
rect 24912 20884 24918 20896
rect 25271 20893 25283 20896
rect 25317 20893 25329 20927
rect 25406 20924 25412 20936
rect 25367 20896 25412 20924
rect 25271 20887 25329 20893
rect 25406 20884 25412 20896
rect 25464 20884 25470 20936
rect 25516 20933 25544 20964
rect 26513 20961 26525 20964
rect 26559 20961 26571 20995
rect 26513 20955 26571 20961
rect 25501 20927 25559 20933
rect 25501 20893 25513 20927
rect 25547 20893 25559 20927
rect 25501 20887 25559 20893
rect 25590 20884 25596 20936
rect 25648 20924 25654 20936
rect 25685 20927 25743 20933
rect 25685 20924 25697 20927
rect 25648 20896 25697 20924
rect 25648 20884 25654 20896
rect 25685 20893 25697 20896
rect 25731 20893 25743 20927
rect 26142 20924 26148 20936
rect 26055 20896 26148 20924
rect 25685 20887 25743 20893
rect 26142 20884 26148 20896
rect 26200 20924 26206 20936
rect 26418 20924 26424 20936
rect 26200 20896 26424 20924
rect 26200 20884 26206 20896
rect 26418 20884 26424 20896
rect 26476 20924 26482 20936
rect 27172 20933 27200 21020
rect 31754 20992 31760 21004
rect 30668 20964 31760 20992
rect 26973 20927 27031 20933
rect 26973 20924 26985 20927
rect 26476 20896 26985 20924
rect 26476 20884 26482 20896
rect 26973 20893 26985 20896
rect 27019 20893 27031 20927
rect 26973 20887 27031 20893
rect 27157 20927 27215 20933
rect 27157 20893 27169 20927
rect 27203 20893 27215 20927
rect 28350 20924 28356 20936
rect 28311 20896 28356 20924
rect 27157 20887 27215 20893
rect 28350 20884 28356 20896
rect 28408 20884 28414 20936
rect 28534 20924 28540 20936
rect 28495 20896 28540 20924
rect 28534 20884 28540 20896
rect 28592 20884 28598 20936
rect 29549 20927 29607 20933
rect 29549 20893 29561 20927
rect 29595 20924 29607 20927
rect 30668 20924 30696 20964
rect 31754 20952 31760 20964
rect 31812 20992 31818 21004
rect 32766 20992 32772 21004
rect 31812 20964 32772 20992
rect 31812 20952 31818 20964
rect 32766 20952 32772 20964
rect 32824 20952 32830 21004
rect 36262 20992 36268 21004
rect 34624 20964 36268 20992
rect 29595 20896 30696 20924
rect 29595 20893 29607 20896
rect 29549 20887 29607 20893
rect 31294 20884 31300 20936
rect 31352 20924 31358 20936
rect 31389 20927 31447 20933
rect 31389 20924 31401 20927
rect 31352 20896 31401 20924
rect 31352 20884 31358 20896
rect 31389 20893 31401 20896
rect 31435 20893 31447 20927
rect 31662 20924 31668 20936
rect 31623 20896 31668 20924
rect 31389 20887 31447 20893
rect 31662 20884 31668 20896
rect 31720 20884 31726 20936
rect 33036 20927 33094 20933
rect 33036 20893 33048 20927
rect 33082 20924 33094 20927
rect 33318 20924 33324 20936
rect 33082 20896 33324 20924
rect 33082 20893 33094 20896
rect 33036 20887 33094 20893
rect 33318 20884 33324 20896
rect 33376 20884 33382 20936
rect 23900 20828 24808 20856
rect 23900 20816 23906 20828
rect 26234 20816 26240 20868
rect 26292 20856 26298 20868
rect 26329 20859 26387 20865
rect 26329 20856 26341 20859
rect 26292 20828 26341 20856
rect 26292 20816 26298 20828
rect 26329 20825 26341 20828
rect 26375 20825 26387 20859
rect 29805 20859 29863 20865
rect 26329 20819 26387 20825
rect 28460 20828 29776 20856
rect 23247 20760 23520 20788
rect 23247 20757 23259 20760
rect 23201 20751 23259 20757
rect 23566 20748 23572 20800
rect 23624 20788 23630 20800
rect 24489 20791 24547 20797
rect 24489 20788 24501 20791
rect 23624 20760 24501 20788
rect 23624 20748 23630 20760
rect 24489 20757 24501 20760
rect 24535 20757 24547 20791
rect 24489 20751 24547 20757
rect 24946 20748 24952 20800
rect 25004 20788 25010 20800
rect 28460 20788 28488 20828
rect 25004 20760 28488 20788
rect 28537 20791 28595 20797
rect 25004 20748 25010 20760
rect 28537 20757 28549 20791
rect 28583 20788 28595 20791
rect 28994 20788 29000 20800
rect 28583 20760 29000 20788
rect 28583 20757 28595 20760
rect 28537 20751 28595 20757
rect 28994 20748 29000 20760
rect 29052 20748 29058 20800
rect 29748 20788 29776 20828
rect 29805 20825 29817 20859
rect 29851 20856 29863 20859
rect 29914 20856 29920 20868
rect 29851 20828 29920 20856
rect 29851 20825 29863 20828
rect 29805 20819 29863 20825
rect 29914 20816 29920 20828
rect 29972 20816 29978 20868
rect 30374 20816 30380 20868
rect 30432 20856 30438 20868
rect 31202 20856 31208 20868
rect 30432 20828 31208 20856
rect 30432 20816 30438 20828
rect 31202 20816 31208 20828
rect 31260 20856 31266 20868
rect 34624 20856 34652 20964
rect 36262 20952 36268 20964
rect 36320 20952 36326 21004
rect 37829 20995 37887 21001
rect 37829 20961 37841 20995
rect 37875 20992 37887 20995
rect 38010 20992 38016 21004
rect 37875 20964 38016 20992
rect 37875 20961 37887 20964
rect 37829 20955 37887 20961
rect 38010 20952 38016 20964
rect 38068 20952 38074 21004
rect 42904 21001 42932 21032
rect 43346 21020 43352 21032
rect 43404 21060 43410 21072
rect 45370 21060 45376 21072
rect 43404 21032 45376 21060
rect 43404 21020 43410 21032
rect 45370 21020 45376 21032
rect 45428 21020 45434 21072
rect 45462 21020 45468 21072
rect 45520 21060 45526 21072
rect 45520 21020 45554 21060
rect 42613 20995 42671 21001
rect 42613 20992 42625 20995
rect 41386 20964 42625 20992
rect 34701 20927 34759 20933
rect 34701 20893 34713 20927
rect 34747 20924 34759 20927
rect 34790 20924 34796 20936
rect 34747 20896 34796 20924
rect 34747 20893 34759 20896
rect 34701 20887 34759 20893
rect 34790 20884 34796 20896
rect 34848 20884 34854 20936
rect 34885 20927 34943 20933
rect 34885 20893 34897 20927
rect 34931 20924 34943 20927
rect 35342 20924 35348 20936
rect 34931 20896 35348 20924
rect 34931 20893 34943 20896
rect 34885 20887 34943 20893
rect 35342 20884 35348 20896
rect 35400 20884 35406 20936
rect 38102 20924 38108 20936
rect 38063 20896 38108 20924
rect 38102 20884 38108 20896
rect 38160 20884 38166 20936
rect 39853 20927 39911 20933
rect 39853 20893 39865 20927
rect 39899 20924 39911 20927
rect 39899 20896 40264 20924
rect 39899 20893 39911 20896
rect 39853 20887 39911 20893
rect 40236 20868 40264 20896
rect 40402 20884 40408 20936
rect 40460 20924 40466 20936
rect 41386 20924 41414 20964
rect 42613 20961 42625 20964
rect 42659 20961 42671 20995
rect 42613 20955 42671 20961
rect 42889 20995 42947 21001
rect 42889 20961 42901 20995
rect 42935 20961 42947 20995
rect 42889 20955 42947 20961
rect 45002 20952 45008 21004
rect 45060 20992 45066 21004
rect 45060 20964 45278 20992
rect 45060 20952 45066 20964
rect 41874 20924 41880 20936
rect 40460 20896 41414 20924
rect 41835 20896 41880 20924
rect 40460 20884 40466 20896
rect 41874 20884 41880 20896
rect 41932 20884 41938 20936
rect 44082 20924 44088 20936
rect 44043 20896 44088 20924
rect 44082 20884 44088 20896
rect 44140 20884 44146 20936
rect 45250 20933 45278 20964
rect 45526 20933 45554 21020
rect 46293 20995 46351 21001
rect 46293 20961 46305 20995
rect 46339 20992 46351 20995
rect 46842 20992 46848 21004
rect 46339 20964 46848 20992
rect 46339 20961 46351 20964
rect 46293 20955 46351 20961
rect 46842 20952 46848 20964
rect 46900 20952 46906 21004
rect 46934 20952 46940 21004
rect 46992 20992 46998 21004
rect 46992 20964 47037 20992
rect 46992 20952 46998 20964
rect 45235 20927 45293 20933
rect 45367 20930 45373 20933
rect 45235 20893 45247 20927
rect 45281 20893 45293 20927
rect 45235 20887 45293 20893
rect 45354 20924 45373 20930
rect 45354 20890 45366 20924
rect 45354 20884 45373 20890
rect 45367 20881 45373 20884
rect 45425 20881 45431 20933
rect 45486 20927 45554 20933
rect 45486 20893 45498 20927
rect 45532 20896 45554 20927
rect 45532 20893 45544 20896
rect 45486 20887 45544 20893
rect 45646 20884 45652 20936
rect 45704 20924 45710 20936
rect 45704 20896 45749 20924
rect 45704 20884 45710 20896
rect 31260 20828 34652 20856
rect 40120 20859 40178 20865
rect 31260 20816 31266 20828
rect 40120 20825 40132 20859
rect 40166 20825 40178 20859
rect 40120 20819 40178 20825
rect 30742 20788 30748 20800
rect 29748 20760 30748 20788
rect 30742 20748 30748 20760
rect 30800 20748 30806 20800
rect 30926 20788 30932 20800
rect 30887 20760 30932 20788
rect 30926 20748 30932 20760
rect 30984 20748 30990 20800
rect 33134 20748 33140 20800
rect 33192 20788 33198 20800
rect 34149 20791 34207 20797
rect 34149 20788 34161 20791
rect 33192 20760 34161 20788
rect 33192 20748 33198 20760
rect 34149 20757 34161 20760
rect 34195 20757 34207 20791
rect 37366 20788 37372 20800
rect 37327 20760 37372 20788
rect 34149 20751 34207 20757
rect 37366 20748 37372 20760
rect 37424 20748 37430 20800
rect 38010 20788 38016 20800
rect 37971 20760 38016 20788
rect 38010 20748 38016 20760
rect 38068 20748 38074 20800
rect 40144 20788 40172 20819
rect 40218 20816 40224 20868
rect 40276 20816 40282 20868
rect 44269 20859 44327 20865
rect 40788 20828 41414 20856
rect 40788 20788 40816 20828
rect 40144 20760 40816 20788
rect 41386 20788 41414 20828
rect 44269 20825 44281 20859
rect 44315 20856 44327 20859
rect 44910 20856 44916 20868
rect 44315 20828 44916 20856
rect 44315 20825 44327 20828
rect 44269 20819 44327 20825
rect 44910 20816 44916 20828
rect 44968 20816 44974 20868
rect 46477 20859 46535 20865
rect 46477 20825 46489 20859
rect 46523 20856 46535 20859
rect 47670 20856 47676 20868
rect 46523 20828 47676 20856
rect 46523 20825 46535 20828
rect 46477 20819 46535 20825
rect 47670 20816 47676 20828
rect 47728 20816 47734 20868
rect 41693 20791 41751 20797
rect 41693 20788 41705 20791
rect 41386 20760 41705 20788
rect 41693 20757 41705 20760
rect 41739 20757 41751 20791
rect 41693 20751 41751 20757
rect 1104 20698 48852 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 48852 20698
rect 1104 20624 48852 20646
rect 14829 20587 14887 20593
rect 6886 20556 14688 20584
rect 2130 20340 2136 20392
rect 2188 20380 2194 20392
rect 6886 20380 6914 20556
rect 11716 20488 13768 20516
rect 11716 20457 11744 20488
rect 11701 20451 11759 20457
rect 11701 20417 11713 20451
rect 11747 20417 11759 20451
rect 11701 20411 11759 20417
rect 11882 20380 11888 20392
rect 2188 20352 6914 20380
rect 11843 20352 11888 20380
rect 2188 20340 2194 20352
rect 11882 20340 11888 20352
rect 11940 20340 11946 20392
rect 12161 20383 12219 20389
rect 12161 20349 12173 20383
rect 12207 20349 12219 20383
rect 12161 20343 12219 20349
rect 2774 20272 2780 20324
rect 2832 20312 2838 20324
rect 5166 20312 5172 20324
rect 2832 20284 5172 20312
rect 2832 20272 2838 20284
rect 5166 20272 5172 20284
rect 5224 20272 5230 20324
rect 14 20204 20 20256
rect 72 20244 78 20256
rect 12176 20244 12204 20343
rect 72 20216 12204 20244
rect 13740 20244 13768 20488
rect 14660 20380 14688 20556
rect 14829 20553 14841 20587
rect 14875 20584 14887 20587
rect 16206 20584 16212 20596
rect 14875 20556 16212 20584
rect 14875 20553 14887 20556
rect 14829 20547 14887 20553
rect 16206 20544 16212 20556
rect 16264 20544 16270 20596
rect 16574 20544 16580 20596
rect 16632 20584 16638 20596
rect 16853 20587 16911 20593
rect 16853 20584 16865 20587
rect 16632 20556 16865 20584
rect 16632 20544 16638 20556
rect 16853 20553 16865 20556
rect 16899 20553 16911 20587
rect 18782 20584 18788 20596
rect 16853 20547 16911 20553
rect 18156 20556 18788 20584
rect 14737 20451 14795 20457
rect 14737 20417 14749 20451
rect 14783 20448 14795 20451
rect 15194 20448 15200 20460
rect 14783 20420 15200 20448
rect 14783 20417 14795 20420
rect 14737 20411 14795 20417
rect 15194 20408 15200 20420
rect 15252 20408 15258 20460
rect 15473 20451 15531 20457
rect 15473 20417 15485 20451
rect 15519 20448 15531 20451
rect 16574 20448 16580 20460
rect 15519 20420 16580 20448
rect 15519 20417 15531 20420
rect 15473 20411 15531 20417
rect 16574 20408 16580 20420
rect 16632 20408 16638 20460
rect 16666 20408 16672 20460
rect 16724 20448 16730 20460
rect 16724 20420 16769 20448
rect 16724 20408 16730 20420
rect 15930 20380 15936 20392
rect 14660 20352 15936 20380
rect 15930 20340 15936 20352
rect 15988 20380 15994 20392
rect 16758 20380 16764 20392
rect 15988 20352 16764 20380
rect 15988 20340 15994 20352
rect 16758 20340 16764 20352
rect 16816 20340 16822 20392
rect 18156 20380 18184 20556
rect 18782 20544 18788 20556
rect 18840 20584 18846 20596
rect 18966 20584 18972 20596
rect 18840 20556 18972 20584
rect 18840 20544 18846 20556
rect 18966 20544 18972 20556
rect 19024 20584 19030 20596
rect 19383 20587 19441 20593
rect 19383 20584 19395 20587
rect 19024 20556 19395 20584
rect 19024 20544 19030 20556
rect 19383 20553 19395 20556
rect 19429 20553 19441 20587
rect 19383 20547 19441 20553
rect 22094 20544 22100 20596
rect 22152 20584 22158 20596
rect 22741 20587 22799 20593
rect 22741 20584 22753 20587
rect 22152 20556 22753 20584
rect 22152 20544 22158 20556
rect 22741 20553 22753 20556
rect 22787 20553 22799 20587
rect 22741 20547 22799 20553
rect 24213 20587 24271 20593
rect 24213 20553 24225 20587
rect 24259 20553 24271 20587
rect 24213 20547 24271 20553
rect 22554 20516 22560 20528
rect 18248 20488 22560 20516
rect 18248 20457 18276 20488
rect 22554 20476 22560 20488
rect 22612 20476 22618 20528
rect 24228 20516 24256 20547
rect 25130 20544 25136 20596
rect 25188 20584 25194 20596
rect 25225 20587 25283 20593
rect 25225 20584 25237 20587
rect 25188 20556 25237 20584
rect 25188 20544 25194 20556
rect 25225 20553 25237 20556
rect 25271 20553 25283 20587
rect 25225 20547 25283 20553
rect 25314 20544 25320 20596
rect 25372 20584 25378 20596
rect 28813 20587 28871 20593
rect 28813 20584 28825 20587
rect 25372 20556 28825 20584
rect 25372 20544 25378 20556
rect 28813 20553 28825 20556
rect 28859 20584 28871 20587
rect 29730 20584 29736 20596
rect 28859 20556 29736 20584
rect 28859 20553 28871 20556
rect 28813 20547 28871 20553
rect 29730 20544 29736 20556
rect 29788 20544 29794 20596
rect 29914 20584 29920 20596
rect 29875 20556 29920 20584
rect 29914 20544 29920 20556
rect 29972 20544 29978 20596
rect 31662 20584 31668 20596
rect 30300 20556 31668 20584
rect 23124 20488 24256 20516
rect 24857 20519 24915 20525
rect 18213 20451 18276 20457
rect 18213 20417 18225 20451
rect 18259 20420 18276 20451
rect 18306 20451 18364 20457
rect 18259 20417 18271 20420
rect 18213 20411 18271 20417
rect 18306 20417 18318 20451
rect 18352 20417 18364 20451
rect 18306 20411 18364 20417
rect 18417 20451 18475 20457
rect 18417 20417 18429 20451
rect 18463 20417 18475 20451
rect 18417 20414 18475 20417
rect 18601 20451 18659 20457
rect 18601 20417 18613 20451
rect 18647 20448 18659 20451
rect 18874 20448 18880 20460
rect 18647 20420 18880 20448
rect 18647 20417 18659 20420
rect 18417 20411 18532 20414
rect 18601 20411 18659 20417
rect 18321 20380 18349 20411
rect 18432 20386 18532 20411
rect 18874 20408 18880 20420
rect 18932 20448 18938 20460
rect 23017 20451 23075 20457
rect 18932 20420 19334 20448
rect 18932 20408 18938 20420
rect 18156 20352 18349 20380
rect 18504 20380 18532 20386
rect 18690 20380 18696 20392
rect 18504 20352 18696 20380
rect 18690 20340 18696 20352
rect 18748 20340 18754 20392
rect 18966 20340 18972 20392
rect 19024 20380 19030 20392
rect 19153 20383 19211 20389
rect 19153 20380 19165 20383
rect 19024 20352 19165 20380
rect 19024 20340 19030 20352
rect 19153 20349 19165 20352
rect 19199 20349 19211 20383
rect 19153 20343 19211 20349
rect 13814 20272 13820 20324
rect 13872 20312 13878 20324
rect 19306 20312 19334 20420
rect 23017 20417 23029 20451
rect 23063 20448 23075 20451
rect 23124 20448 23152 20488
rect 24857 20485 24869 20519
rect 24903 20516 24915 20519
rect 26142 20516 26148 20528
rect 24903 20488 26148 20516
rect 24903 20485 24915 20488
rect 24857 20479 24915 20485
rect 26142 20476 26148 20488
rect 26200 20476 26206 20528
rect 29454 20516 29460 20528
rect 26252 20488 29460 20516
rect 23063 20420 23152 20448
rect 23201 20451 23259 20457
rect 23063 20417 23075 20420
rect 23017 20411 23075 20417
rect 23201 20417 23213 20451
rect 23247 20448 23259 20451
rect 23474 20448 23480 20460
rect 23247 20420 23480 20448
rect 23247 20417 23259 20420
rect 23201 20411 23259 20417
rect 23474 20408 23480 20420
rect 23532 20408 23538 20460
rect 23566 20408 23572 20460
rect 23624 20448 23630 20460
rect 23753 20451 23811 20457
rect 23753 20448 23765 20451
rect 23624 20420 23765 20448
rect 23624 20408 23630 20420
rect 23753 20417 23765 20420
rect 23799 20417 23811 20451
rect 23753 20411 23811 20417
rect 24029 20451 24087 20457
rect 24029 20417 24041 20451
rect 24075 20448 24087 20451
rect 24946 20448 24952 20460
rect 24075 20420 24952 20448
rect 24075 20417 24087 20420
rect 24029 20411 24087 20417
rect 24946 20408 24952 20420
rect 25004 20408 25010 20460
rect 25041 20451 25099 20457
rect 25041 20417 25053 20451
rect 25087 20448 25099 20451
rect 25130 20448 25136 20460
rect 25087 20420 25136 20448
rect 25087 20417 25099 20420
rect 25041 20411 25099 20417
rect 25130 20408 25136 20420
rect 25188 20448 25194 20460
rect 25682 20448 25688 20460
rect 25188 20420 25688 20448
rect 25188 20408 25194 20420
rect 25682 20408 25688 20420
rect 25740 20448 25746 20460
rect 26252 20448 26280 20488
rect 29454 20476 29460 20488
rect 29512 20476 29518 20528
rect 30300 20463 30328 20556
rect 31662 20544 31668 20556
rect 31720 20544 31726 20596
rect 35618 20544 35624 20596
rect 35676 20584 35682 20596
rect 36725 20587 36783 20593
rect 35676 20556 36676 20584
rect 35676 20544 35682 20556
rect 31481 20519 31539 20525
rect 31481 20485 31493 20519
rect 31527 20516 31539 20519
rect 32309 20519 32367 20525
rect 32309 20516 32321 20519
rect 31527 20488 32321 20516
rect 31527 20485 31539 20488
rect 31481 20479 31539 20485
rect 32309 20485 32321 20488
rect 32355 20485 32367 20519
rect 32309 20479 32367 20485
rect 36265 20519 36323 20525
rect 36265 20485 36277 20519
rect 36311 20516 36323 20519
rect 36648 20516 36676 20556
rect 36725 20553 36737 20587
rect 36771 20584 36783 20587
rect 38010 20584 38016 20596
rect 36771 20556 38016 20584
rect 36771 20553 36783 20556
rect 36725 20547 36783 20553
rect 38010 20544 38016 20556
rect 38068 20544 38074 20596
rect 43257 20587 43315 20593
rect 43257 20553 43269 20587
rect 43303 20584 43315 20587
rect 44082 20584 44088 20596
rect 43303 20556 44088 20584
rect 43303 20553 43315 20556
rect 43257 20547 43315 20553
rect 44082 20544 44088 20556
rect 44140 20544 44146 20596
rect 44450 20584 44456 20596
rect 44411 20556 44456 20584
rect 44450 20544 44456 20556
rect 44508 20544 44514 20596
rect 47670 20584 47676 20596
rect 47631 20556 47676 20584
rect 47670 20544 47676 20556
rect 47728 20544 47734 20596
rect 38028 20516 38056 20544
rect 40126 20516 40132 20528
rect 36311 20488 36492 20516
rect 36648 20488 37504 20516
rect 38028 20488 38516 20516
rect 40087 20488 40132 20516
rect 36311 20485 36323 20488
rect 36265 20479 36323 20485
rect 25740 20420 26280 20448
rect 28629 20451 28687 20457
rect 25740 20408 25746 20420
rect 28629 20417 28641 20451
rect 28675 20448 28687 20451
rect 29546 20448 29552 20460
rect 28675 20420 29552 20448
rect 28675 20417 28687 20420
rect 28629 20411 28687 20417
rect 29546 20408 29552 20420
rect 29604 20408 29610 20460
rect 30190 20448 30196 20460
rect 30151 20420 30196 20448
rect 30190 20408 30196 20420
rect 30248 20408 30254 20460
rect 30282 20457 30340 20463
rect 30282 20423 30294 20457
rect 30328 20423 30340 20457
rect 30282 20417 30340 20423
rect 30374 20408 30380 20460
rect 30432 20448 30438 20460
rect 30432 20420 30477 20448
rect 30432 20408 30438 20420
rect 30558 20408 30564 20460
rect 30616 20448 30622 20460
rect 31389 20451 31447 20457
rect 30616 20420 30661 20448
rect 30616 20408 30622 20420
rect 31389 20417 31401 20451
rect 31435 20417 31447 20451
rect 31389 20411 31447 20417
rect 22922 20380 22928 20392
rect 22883 20352 22928 20380
rect 22922 20340 22928 20352
rect 22980 20340 22986 20392
rect 23106 20340 23112 20392
rect 23164 20380 23170 20392
rect 23164 20352 23209 20380
rect 23164 20340 23170 20352
rect 23290 20340 23296 20392
rect 23348 20380 23354 20392
rect 23845 20383 23903 20389
rect 23845 20380 23857 20383
rect 23348 20352 23857 20380
rect 23348 20340 23354 20352
rect 23845 20349 23857 20352
rect 23891 20349 23903 20383
rect 31404 20380 31432 20411
rect 23845 20343 23903 20349
rect 23952 20352 31432 20380
rect 32125 20383 32183 20389
rect 20530 20312 20536 20324
rect 13872 20284 18092 20312
rect 19306 20284 20536 20312
rect 13872 20272 13878 20284
rect 17586 20244 17592 20256
rect 13740 20216 17592 20244
rect 72 20204 78 20216
rect 17586 20204 17592 20216
rect 17644 20204 17650 20256
rect 17954 20244 17960 20256
rect 17915 20216 17960 20244
rect 17954 20204 17960 20216
rect 18012 20204 18018 20256
rect 18064 20244 18092 20284
rect 20530 20272 20536 20284
rect 20588 20312 20594 20324
rect 21910 20312 21916 20324
rect 20588 20284 21916 20312
rect 20588 20272 20594 20284
rect 21910 20272 21916 20284
rect 21968 20272 21974 20324
rect 23952 20312 23980 20352
rect 32125 20349 32137 20383
rect 32171 20380 32183 20383
rect 33134 20380 33140 20392
rect 32171 20352 33140 20380
rect 32171 20349 32183 20352
rect 32125 20343 32183 20349
rect 33134 20340 33140 20352
rect 33192 20340 33198 20392
rect 33962 20380 33968 20392
rect 33923 20352 33968 20380
rect 33962 20340 33968 20352
rect 34020 20340 34026 20392
rect 36170 20340 36176 20392
rect 36228 20380 36234 20392
rect 36357 20383 36415 20389
rect 36357 20380 36369 20383
rect 36228 20352 36369 20380
rect 36228 20340 36234 20352
rect 36357 20349 36369 20352
rect 36403 20349 36415 20383
rect 36464 20380 36492 20488
rect 36538 20408 36544 20460
rect 36596 20448 36602 20460
rect 37476 20457 37504 20488
rect 38488 20457 38516 20488
rect 40126 20476 40132 20488
rect 40184 20476 40190 20528
rect 40313 20519 40371 20525
rect 40313 20485 40325 20519
rect 40359 20516 40371 20519
rect 40862 20516 40868 20528
rect 40359 20488 40868 20516
rect 40359 20485 40371 20488
rect 40313 20479 40371 20485
rect 40862 20476 40868 20488
rect 40920 20476 40926 20528
rect 45925 20519 45983 20525
rect 45925 20516 45937 20519
rect 45020 20488 45937 20516
rect 37461 20451 37519 20457
rect 36596 20420 36641 20448
rect 36596 20408 36602 20420
rect 37461 20417 37473 20451
rect 37507 20417 37519 20451
rect 37461 20411 37519 20417
rect 38289 20451 38347 20457
rect 38289 20417 38301 20451
rect 38335 20417 38347 20451
rect 38289 20411 38347 20417
rect 38473 20451 38531 20457
rect 38473 20417 38485 20451
rect 38519 20417 38531 20451
rect 38473 20411 38531 20417
rect 40773 20451 40831 20457
rect 40773 20417 40785 20451
rect 40819 20448 40831 20451
rect 41322 20448 41328 20460
rect 40819 20420 41328 20448
rect 40819 20417 40831 20420
rect 40773 20411 40831 20417
rect 37274 20380 37280 20392
rect 36464 20352 37280 20380
rect 36357 20343 36415 20349
rect 37274 20340 37280 20352
rect 37332 20340 37338 20392
rect 37553 20383 37611 20389
rect 37553 20349 37565 20383
rect 37599 20349 37611 20383
rect 37553 20343 37611 20349
rect 37829 20383 37887 20389
rect 37829 20349 37841 20383
rect 37875 20380 37887 20383
rect 38102 20380 38108 20392
rect 37875 20352 38108 20380
rect 37875 20349 37887 20352
rect 37829 20343 37887 20349
rect 22020 20284 23980 20312
rect 22020 20244 22048 20284
rect 24486 20272 24492 20324
rect 24544 20312 24550 20324
rect 29270 20312 29276 20324
rect 24544 20284 29276 20312
rect 24544 20272 24550 20284
rect 29270 20272 29276 20284
rect 29328 20312 29334 20324
rect 30558 20312 30564 20324
rect 29328 20284 30564 20312
rect 29328 20272 29334 20284
rect 30558 20272 30564 20284
rect 30616 20272 30622 20324
rect 31478 20272 31484 20324
rect 31536 20312 31542 20324
rect 36538 20312 36544 20324
rect 31536 20284 36544 20312
rect 31536 20272 31542 20284
rect 36538 20272 36544 20284
rect 36596 20272 36602 20324
rect 37568 20312 37596 20343
rect 38102 20340 38108 20352
rect 38160 20380 38166 20392
rect 38304 20380 38332 20411
rect 41322 20408 41328 20420
rect 41380 20408 41386 20460
rect 42150 20408 42156 20460
rect 42208 20448 42214 20460
rect 42702 20448 42708 20460
rect 42208 20420 42708 20448
rect 42208 20408 42214 20420
rect 42702 20408 42708 20420
rect 42760 20448 42766 20460
rect 43441 20451 43499 20457
rect 43441 20448 43453 20451
rect 42760 20420 43453 20448
rect 42760 20408 42766 20420
rect 43441 20417 43453 20420
rect 43487 20417 43499 20451
rect 43441 20411 43499 20417
rect 44729 20451 44787 20457
rect 44729 20417 44741 20451
rect 44775 20417 44787 20451
rect 44729 20411 44787 20417
rect 44818 20451 44876 20457
rect 44818 20417 44830 20451
rect 44864 20417 44876 20451
rect 44818 20411 44876 20417
rect 44913 20451 44971 20457
rect 44913 20417 44925 20451
rect 44959 20432 44971 20451
rect 45020 20432 45048 20488
rect 45925 20485 45937 20488
rect 45971 20485 45983 20519
rect 45925 20479 45983 20485
rect 44959 20417 45048 20432
rect 44913 20411 45048 20417
rect 45097 20451 45155 20457
rect 45097 20417 45109 20451
rect 45143 20417 45155 20451
rect 45097 20411 45155 20417
rect 38160 20352 38332 20380
rect 41049 20383 41107 20389
rect 38160 20340 38166 20352
rect 41049 20349 41061 20383
rect 41095 20380 41107 20383
rect 41782 20380 41788 20392
rect 41095 20352 41788 20380
rect 41095 20349 41107 20352
rect 41049 20343 41107 20349
rect 41782 20340 41788 20352
rect 41840 20340 41846 20392
rect 44744 20380 44772 20411
rect 43180 20352 44772 20380
rect 40494 20312 40500 20324
rect 37568 20284 40500 20312
rect 40494 20272 40500 20284
rect 40552 20312 40558 20324
rect 40954 20312 40960 20324
rect 40552 20284 40960 20312
rect 40552 20272 40558 20284
rect 40954 20272 40960 20284
rect 41012 20272 41018 20324
rect 43180 20256 43208 20352
rect 44827 20312 44855 20411
rect 44928 20404 45048 20411
rect 45112 20380 45140 20411
rect 45186 20408 45192 20460
rect 45244 20448 45250 20460
rect 45557 20451 45615 20457
rect 45557 20448 45569 20451
rect 45244 20420 45569 20448
rect 45244 20408 45250 20420
rect 45557 20417 45569 20420
rect 45603 20417 45615 20451
rect 45557 20411 45615 20417
rect 45741 20451 45799 20457
rect 45741 20417 45753 20451
rect 45787 20448 45799 20451
rect 46474 20448 46480 20460
rect 45787 20420 46480 20448
rect 45787 20417 45799 20420
rect 45741 20411 45799 20417
rect 46474 20408 46480 20420
rect 46532 20408 46538 20460
rect 46842 20448 46848 20460
rect 46803 20420 46848 20448
rect 46842 20408 46848 20420
rect 46900 20408 46906 20460
rect 47302 20408 47308 20460
rect 47360 20448 47366 20460
rect 47581 20451 47639 20457
rect 47581 20448 47593 20451
rect 47360 20420 47593 20448
rect 47360 20408 47366 20420
rect 47581 20417 47593 20420
rect 47627 20417 47639 20451
rect 47581 20411 47639 20417
rect 45646 20380 45652 20392
rect 45112 20352 45652 20380
rect 45646 20340 45652 20352
rect 45704 20340 45710 20392
rect 45370 20312 45376 20324
rect 44827 20284 45376 20312
rect 45370 20272 45376 20284
rect 45428 20272 45434 20324
rect 18064 20216 22048 20244
rect 22094 20204 22100 20256
rect 22152 20244 22158 20256
rect 23753 20247 23811 20253
rect 23753 20244 23765 20247
rect 22152 20216 23765 20244
rect 22152 20204 22158 20216
rect 23753 20213 23765 20216
rect 23799 20213 23811 20247
rect 23753 20207 23811 20213
rect 24302 20204 24308 20256
rect 24360 20244 24366 20256
rect 27338 20244 27344 20256
rect 24360 20216 27344 20244
rect 24360 20204 24366 20216
rect 27338 20204 27344 20216
rect 27396 20204 27402 20256
rect 29730 20204 29736 20256
rect 29788 20244 29794 20256
rect 31294 20244 31300 20256
rect 29788 20216 31300 20244
rect 29788 20204 29794 20216
rect 31294 20204 31300 20216
rect 31352 20204 31358 20256
rect 34146 20204 34152 20256
rect 34204 20244 34210 20256
rect 36265 20247 36323 20253
rect 36265 20244 36277 20247
rect 34204 20216 36277 20244
rect 34204 20204 34210 20216
rect 36265 20213 36277 20216
rect 36311 20244 36323 20247
rect 37090 20244 37096 20256
rect 36311 20216 37096 20244
rect 36311 20213 36323 20216
rect 36265 20207 36323 20213
rect 37090 20204 37096 20216
rect 37148 20244 37154 20256
rect 37458 20244 37464 20256
rect 37148 20216 37464 20244
rect 37148 20204 37154 20216
rect 37458 20204 37464 20216
rect 37516 20204 37522 20256
rect 38289 20247 38347 20253
rect 38289 20213 38301 20247
rect 38335 20244 38347 20247
rect 38378 20244 38384 20256
rect 38335 20216 38384 20244
rect 38335 20213 38347 20216
rect 38289 20207 38347 20213
rect 38378 20204 38384 20216
rect 38436 20204 38442 20256
rect 40862 20204 40868 20256
rect 40920 20244 40926 20256
rect 43162 20244 43168 20256
rect 40920 20216 43168 20244
rect 40920 20204 40926 20216
rect 43162 20204 43168 20216
rect 43220 20204 43226 20256
rect 46937 20247 46995 20253
rect 46937 20213 46949 20247
rect 46983 20244 46995 20247
rect 47026 20244 47032 20256
rect 46983 20216 47032 20244
rect 46983 20213 46995 20216
rect 46937 20207 46995 20213
rect 47026 20204 47032 20216
rect 47084 20204 47090 20256
rect 1104 20154 48852 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 48852 20154
rect 1104 20080 48852 20102
rect 11882 20040 11888 20052
rect 11843 20012 11888 20040
rect 11882 20000 11888 20012
rect 11940 20000 11946 20052
rect 17129 20043 17187 20049
rect 17129 20009 17141 20043
rect 17175 20040 17187 20043
rect 17402 20040 17408 20052
rect 17175 20012 17408 20040
rect 17175 20009 17187 20012
rect 17129 20003 17187 20009
rect 17402 20000 17408 20012
rect 17460 20000 17466 20052
rect 17586 20000 17592 20052
rect 17644 20040 17650 20052
rect 21910 20040 21916 20052
rect 17644 20012 21916 20040
rect 17644 20000 17650 20012
rect 21910 20000 21916 20012
rect 21968 20000 21974 20052
rect 22554 20040 22560 20052
rect 22066 20012 22560 20040
rect 17218 19932 17224 19984
rect 17276 19972 17282 19984
rect 18230 19972 18236 19984
rect 17276 19944 18236 19972
rect 17276 19932 17282 19944
rect 18230 19932 18236 19944
rect 18288 19972 18294 19984
rect 18506 19972 18512 19984
rect 18288 19944 18512 19972
rect 18288 19932 18294 19944
rect 18506 19932 18512 19944
rect 18564 19972 18570 19984
rect 19245 19975 19303 19981
rect 19245 19972 19257 19975
rect 18564 19944 19257 19972
rect 18564 19932 18570 19944
rect 19245 19941 19257 19944
rect 19291 19941 19303 19975
rect 19245 19935 19303 19941
rect 21726 19932 21732 19984
rect 21784 19972 21790 19984
rect 22066 19972 22094 20012
rect 22554 20000 22560 20012
rect 22612 20000 22618 20052
rect 22738 20000 22744 20052
rect 22796 20040 22802 20052
rect 22833 20043 22891 20049
rect 22833 20040 22845 20043
rect 22796 20012 22845 20040
rect 22796 20000 22802 20012
rect 22833 20009 22845 20012
rect 22879 20040 22891 20043
rect 23290 20040 23296 20052
rect 22879 20012 23296 20040
rect 22879 20009 22891 20012
rect 22833 20003 22891 20009
rect 23290 20000 23296 20012
rect 23348 20000 23354 20052
rect 23382 20000 23388 20052
rect 23440 20040 23446 20052
rect 25777 20043 25835 20049
rect 25777 20040 25789 20043
rect 23440 20012 25789 20040
rect 23440 20000 23446 20012
rect 25777 20009 25789 20012
rect 25823 20009 25835 20043
rect 25777 20003 25835 20009
rect 26418 20000 26424 20052
rect 26476 20040 26482 20052
rect 28629 20043 28687 20049
rect 28629 20040 28641 20043
rect 26476 20012 28641 20040
rect 26476 20000 26482 20012
rect 28629 20009 28641 20012
rect 28675 20040 28687 20043
rect 29086 20040 29092 20052
rect 28675 20012 29092 20040
rect 28675 20009 28687 20012
rect 28629 20003 28687 20009
rect 29086 20000 29092 20012
rect 29144 20000 29150 20052
rect 30374 20000 30380 20052
rect 30432 20040 30438 20052
rect 30469 20043 30527 20049
rect 30469 20040 30481 20043
rect 30432 20012 30481 20040
rect 30432 20000 30438 20012
rect 30469 20009 30481 20012
rect 30515 20009 30527 20043
rect 30469 20003 30527 20009
rect 32309 20043 32367 20049
rect 32309 20009 32321 20043
rect 32355 20040 32367 20043
rect 32398 20040 32404 20052
rect 32355 20012 32404 20040
rect 32355 20009 32367 20012
rect 32309 20003 32367 20009
rect 32398 20000 32404 20012
rect 32456 20000 32462 20052
rect 37642 20000 37648 20052
rect 37700 20040 37706 20052
rect 38197 20043 38255 20049
rect 38197 20040 38209 20043
rect 37700 20012 38209 20040
rect 37700 20000 37706 20012
rect 38197 20009 38209 20012
rect 38243 20040 38255 20043
rect 39390 20040 39396 20052
rect 38243 20012 39396 20040
rect 38243 20009 38255 20012
rect 38197 20003 38255 20009
rect 39390 20000 39396 20012
rect 39448 20000 39454 20052
rect 40402 20000 40408 20052
rect 40460 20040 40466 20052
rect 40773 20043 40831 20049
rect 40773 20040 40785 20043
rect 40460 20012 40785 20040
rect 40460 20000 40466 20012
rect 40773 20009 40785 20012
rect 40819 20009 40831 20043
rect 40773 20003 40831 20009
rect 41138 20000 41144 20052
rect 41196 20040 41202 20052
rect 41233 20043 41291 20049
rect 41233 20040 41245 20043
rect 41196 20012 41245 20040
rect 41196 20000 41202 20012
rect 41233 20009 41245 20012
rect 41279 20009 41291 20043
rect 41233 20003 41291 20009
rect 21784 19944 22094 19972
rect 21784 19932 21790 19944
rect 22186 19932 22192 19984
rect 22244 19972 22250 19984
rect 46842 19972 46848 19984
rect 22244 19944 46848 19972
rect 22244 19932 22250 19944
rect 46842 19932 46848 19944
rect 46900 19932 46906 19984
rect 18782 19904 18788 19916
rect 18321 19876 18788 19904
rect 10778 19796 10784 19848
rect 10836 19836 10842 19848
rect 11793 19839 11851 19845
rect 11793 19836 11805 19839
rect 10836 19808 11805 19836
rect 10836 19796 10842 19808
rect 11793 19805 11805 19808
rect 11839 19836 11851 19839
rect 13814 19836 13820 19848
rect 11839 19808 13820 19836
rect 11839 19805 11851 19808
rect 11793 19799 11851 19805
rect 13814 19796 13820 19808
rect 13872 19796 13878 19848
rect 15746 19836 15752 19848
rect 15707 19808 15752 19836
rect 15746 19796 15752 19808
rect 15804 19796 15810 19848
rect 16016 19839 16074 19845
rect 16016 19805 16028 19839
rect 16062 19836 16074 19839
rect 17954 19836 17960 19848
rect 16062 19808 17960 19836
rect 16062 19805 16074 19808
rect 16016 19799 16074 19805
rect 17954 19796 17960 19808
rect 18012 19796 18018 19848
rect 18321 19845 18349 19876
rect 18782 19864 18788 19876
rect 18840 19864 18846 19916
rect 19334 19864 19340 19916
rect 19392 19904 19398 19916
rect 20625 19907 20683 19913
rect 20625 19904 20637 19907
rect 19392 19876 20637 19904
rect 19392 19864 19398 19876
rect 20625 19873 20637 19876
rect 20671 19873 20683 19907
rect 22695 19907 22753 19913
rect 22695 19904 22707 19907
rect 20625 19867 20683 19873
rect 22388 19876 22707 19904
rect 18213 19839 18271 19845
rect 18213 19805 18225 19839
rect 18259 19805 18271 19839
rect 18213 19799 18271 19805
rect 18306 19839 18364 19845
rect 18306 19805 18318 19839
rect 18352 19805 18364 19839
rect 18306 19799 18364 19805
rect 17957 19703 18015 19709
rect 17957 19669 17969 19703
rect 18003 19700 18015 19703
rect 18046 19700 18052 19712
rect 18003 19672 18052 19700
rect 18003 19669 18015 19672
rect 17957 19663 18015 19669
rect 18046 19660 18052 19672
rect 18104 19660 18110 19712
rect 18228 19700 18256 19799
rect 18414 19796 18420 19848
rect 18472 19845 18478 19848
rect 18472 19836 18480 19845
rect 18601 19839 18659 19845
rect 18472 19808 18517 19836
rect 18472 19799 18480 19808
rect 18601 19805 18613 19839
rect 18647 19836 18659 19839
rect 18874 19836 18880 19848
rect 18647 19808 18880 19836
rect 18647 19805 18659 19808
rect 18601 19799 18659 19805
rect 18472 19796 18478 19799
rect 18874 19796 18880 19808
rect 18932 19796 18938 19848
rect 19150 19796 19156 19848
rect 19208 19836 19214 19848
rect 19429 19839 19487 19845
rect 19429 19836 19441 19839
rect 19208 19808 19441 19836
rect 19208 19796 19214 19808
rect 19429 19805 19441 19808
rect 19475 19836 19487 19839
rect 20714 19836 20720 19848
rect 19475 19808 20720 19836
rect 19475 19805 19487 19808
rect 19429 19799 19487 19805
rect 20714 19796 20720 19808
rect 20772 19796 20778 19848
rect 22094 19796 22100 19848
rect 22152 19836 22158 19848
rect 22388 19836 22416 19876
rect 22695 19873 22707 19876
rect 22741 19873 22753 19907
rect 22695 19867 22753 19873
rect 26602 19864 26608 19916
rect 26660 19904 26666 19916
rect 37093 19907 37151 19913
rect 26660 19876 26705 19904
rect 26660 19864 26666 19876
rect 37093 19873 37105 19907
rect 37139 19904 37151 19907
rect 37274 19904 37280 19916
rect 37139 19876 37280 19904
rect 37139 19873 37151 19876
rect 37093 19867 37151 19873
rect 37274 19864 37280 19876
rect 37332 19864 37338 19916
rect 37369 19907 37427 19913
rect 37369 19873 37381 19907
rect 37415 19904 37427 19907
rect 38746 19904 38752 19916
rect 37415 19876 38752 19904
rect 37415 19873 37427 19876
rect 37369 19867 37427 19873
rect 38746 19864 38752 19876
rect 38804 19864 38810 19916
rect 40862 19904 40868 19916
rect 40823 19876 40868 19904
rect 40862 19864 40868 19876
rect 40920 19864 40926 19916
rect 45094 19904 45100 19916
rect 40972 19876 45100 19904
rect 22152 19808 22416 19836
rect 22557 19839 22615 19845
rect 22152 19796 22158 19808
rect 22557 19805 22569 19839
rect 22603 19805 22615 19839
rect 22557 19799 22615 19805
rect 20892 19771 20950 19777
rect 20892 19737 20904 19771
rect 20938 19768 20950 19771
rect 21910 19768 21916 19780
rect 20938 19740 21916 19768
rect 20938 19737 20950 19740
rect 20892 19731 20950 19737
rect 21910 19728 21916 19740
rect 21968 19728 21974 19780
rect 22370 19728 22376 19780
rect 22428 19768 22434 19780
rect 22572 19768 22600 19799
rect 22830 19796 22836 19848
rect 22888 19836 22894 19848
rect 23017 19839 23075 19845
rect 23017 19836 23029 19839
rect 22888 19808 23029 19836
rect 22888 19796 22894 19808
rect 23017 19805 23029 19808
rect 23063 19805 23075 19839
rect 23017 19799 23075 19805
rect 25593 19839 25651 19845
rect 25593 19805 25605 19839
rect 25639 19836 25651 19839
rect 26142 19836 26148 19848
rect 25639 19808 26148 19836
rect 25639 19805 25651 19808
rect 25593 19799 25651 19805
rect 26142 19796 26148 19808
rect 26200 19796 26206 19848
rect 26329 19839 26387 19845
rect 26329 19805 26341 19839
rect 26375 19805 26387 19839
rect 26329 19799 26387 19805
rect 26421 19839 26479 19845
rect 26421 19805 26433 19839
rect 26467 19805 26479 19839
rect 26421 19799 26479 19805
rect 30101 19839 30159 19845
rect 30101 19805 30113 19839
rect 30147 19836 30159 19839
rect 31938 19836 31944 19848
rect 30147 19808 31944 19836
rect 30147 19805 30159 19808
rect 30101 19799 30159 19805
rect 25774 19768 25780 19780
rect 22428 19740 25780 19768
rect 22428 19728 22434 19740
rect 25774 19728 25780 19740
rect 25832 19768 25838 19780
rect 26344 19768 26372 19799
rect 25832 19740 26372 19768
rect 26436 19768 26464 19799
rect 31938 19796 31944 19808
rect 31996 19796 32002 19848
rect 32125 19839 32183 19845
rect 32125 19805 32137 19839
rect 32171 19836 32183 19839
rect 33134 19836 33140 19848
rect 32171 19808 33140 19836
rect 32171 19805 32183 19808
rect 32125 19799 32183 19805
rect 33134 19796 33140 19808
rect 33192 19796 33198 19848
rect 36170 19796 36176 19848
rect 36228 19836 36234 19848
rect 36998 19836 37004 19848
rect 36228 19808 37004 19836
rect 36228 19796 36234 19808
rect 36998 19796 37004 19808
rect 37056 19796 37062 19848
rect 38470 19796 38476 19848
rect 38528 19836 38534 19848
rect 40972 19836 41000 19876
rect 45094 19864 45100 19876
rect 45152 19864 45158 19916
rect 46293 19907 46351 19913
rect 46293 19873 46305 19907
rect 46339 19904 46351 19907
rect 47762 19904 47768 19916
rect 46339 19876 47768 19904
rect 46339 19873 46351 19876
rect 46293 19867 46351 19873
rect 47762 19864 47768 19876
rect 47820 19864 47826 19916
rect 38528 19808 41000 19836
rect 38528 19796 38534 19808
rect 41046 19796 41052 19848
rect 41104 19836 41110 19848
rect 48130 19836 48136 19848
rect 41104 19808 41149 19836
rect 48091 19808 48136 19836
rect 41104 19796 41110 19808
rect 48130 19796 48136 19808
rect 48188 19796 48194 19848
rect 26786 19768 26792 19780
rect 26436 19740 26792 19768
rect 25832 19728 25838 19740
rect 26786 19728 26792 19740
rect 26844 19728 26850 19780
rect 28258 19728 28264 19780
rect 28316 19768 28322 19780
rect 28537 19771 28595 19777
rect 28537 19768 28549 19771
rect 28316 19740 28549 19768
rect 28316 19728 28322 19740
rect 28537 19737 28549 19740
rect 28583 19737 28595 19771
rect 28537 19731 28595 19737
rect 28718 19728 28724 19780
rect 28776 19768 28782 19780
rect 30285 19771 30343 19777
rect 30285 19768 30297 19771
rect 28776 19740 30297 19768
rect 28776 19728 28782 19740
rect 30285 19737 30297 19740
rect 30331 19768 30343 19771
rect 30926 19768 30932 19780
rect 30331 19740 30932 19768
rect 30331 19737 30343 19740
rect 30285 19731 30343 19737
rect 30926 19728 30932 19740
rect 30984 19728 30990 19780
rect 31018 19728 31024 19780
rect 31076 19768 31082 19780
rect 31205 19771 31263 19777
rect 31076 19740 31121 19768
rect 31076 19728 31082 19740
rect 31205 19737 31217 19771
rect 31251 19768 31263 19771
rect 33410 19768 33416 19780
rect 31251 19740 33416 19768
rect 31251 19737 31263 19740
rect 31205 19731 31263 19737
rect 33410 19728 33416 19740
rect 33468 19768 33474 19780
rect 34054 19768 34060 19780
rect 33468 19740 34060 19768
rect 33468 19728 33474 19740
rect 34054 19728 34060 19740
rect 34112 19728 34118 19780
rect 38010 19768 38016 19780
rect 37971 19740 38016 19768
rect 38010 19728 38016 19740
rect 38068 19728 38074 19780
rect 38194 19728 38200 19780
rect 38252 19777 38258 19780
rect 38252 19771 38271 19777
rect 38259 19737 38271 19771
rect 38252 19731 38271 19737
rect 38252 19728 38258 19731
rect 38562 19728 38568 19780
rect 38620 19768 38626 19780
rect 38654 19768 38660 19780
rect 38620 19740 38660 19768
rect 38620 19728 38626 19740
rect 38654 19728 38660 19740
rect 38712 19728 38718 19780
rect 40770 19768 40776 19780
rect 40731 19740 40776 19768
rect 40770 19728 40776 19740
rect 40828 19728 40834 19780
rect 40954 19728 40960 19780
rect 41012 19768 41018 19780
rect 41693 19771 41751 19777
rect 41693 19768 41705 19771
rect 41012 19740 41705 19768
rect 41012 19728 41018 19740
rect 41693 19737 41705 19740
rect 41739 19737 41751 19771
rect 41874 19768 41880 19780
rect 41835 19740 41880 19768
rect 41693 19731 41751 19737
rect 41874 19728 41880 19740
rect 41932 19728 41938 19780
rect 44082 19728 44088 19780
rect 44140 19768 44146 19780
rect 45097 19771 45155 19777
rect 45097 19768 45109 19771
rect 44140 19740 45109 19768
rect 44140 19728 44146 19740
rect 45097 19737 45109 19740
rect 45143 19768 45155 19771
rect 45186 19768 45192 19780
rect 45143 19740 45192 19768
rect 45143 19737 45155 19740
rect 45097 19731 45155 19737
rect 45186 19728 45192 19740
rect 45244 19728 45250 19780
rect 45281 19771 45339 19777
rect 45281 19737 45293 19771
rect 45327 19768 45339 19771
rect 46290 19768 46296 19780
rect 45327 19740 46296 19768
rect 45327 19737 45339 19740
rect 45281 19731 45339 19737
rect 46290 19728 46296 19740
rect 46348 19728 46354 19780
rect 46477 19771 46535 19777
rect 46477 19737 46489 19771
rect 46523 19768 46535 19771
rect 46934 19768 46940 19780
rect 46523 19740 46940 19768
rect 46523 19737 46535 19740
rect 46477 19731 46535 19737
rect 46934 19728 46940 19740
rect 46992 19728 46998 19780
rect 18598 19700 18604 19712
rect 18228 19672 18604 19700
rect 18598 19660 18604 19672
rect 18656 19660 18662 19712
rect 18966 19660 18972 19712
rect 19024 19700 19030 19712
rect 21726 19700 21732 19712
rect 19024 19672 21732 19700
rect 19024 19660 19030 19672
rect 21726 19660 21732 19672
rect 21784 19660 21790 19712
rect 22005 19703 22063 19709
rect 22005 19669 22017 19703
rect 22051 19700 22063 19703
rect 22830 19700 22836 19712
rect 22051 19672 22836 19700
rect 22051 19669 22063 19672
rect 22005 19663 22063 19669
rect 22830 19660 22836 19672
rect 22888 19660 22894 19712
rect 23017 19703 23075 19709
rect 23017 19669 23029 19703
rect 23063 19700 23075 19703
rect 23106 19700 23112 19712
rect 23063 19672 23112 19700
rect 23063 19669 23075 19672
rect 23017 19663 23075 19669
rect 23106 19660 23112 19672
rect 23164 19660 23170 19712
rect 23198 19660 23204 19712
rect 23256 19700 23262 19712
rect 26418 19700 26424 19712
rect 23256 19672 26424 19700
rect 23256 19660 23262 19672
rect 26418 19660 26424 19672
rect 26476 19660 26482 19712
rect 26605 19703 26663 19709
rect 26605 19669 26617 19703
rect 26651 19700 26663 19703
rect 27154 19700 27160 19712
rect 26651 19672 27160 19700
rect 26651 19669 26663 19672
rect 26605 19663 26663 19669
rect 27154 19660 27160 19672
rect 27212 19660 27218 19712
rect 27338 19660 27344 19712
rect 27396 19700 27402 19712
rect 35618 19700 35624 19712
rect 27396 19672 35624 19700
rect 27396 19660 27402 19672
rect 35618 19660 35624 19672
rect 35676 19660 35682 19712
rect 38381 19703 38439 19709
rect 38381 19669 38393 19703
rect 38427 19700 38439 19703
rect 38470 19700 38476 19712
rect 38427 19672 38476 19700
rect 38427 19669 38439 19672
rect 38381 19663 38439 19669
rect 38470 19660 38476 19672
rect 38528 19660 38534 19712
rect 39114 19660 39120 19712
rect 39172 19700 39178 19712
rect 40862 19700 40868 19712
rect 39172 19672 40868 19700
rect 39172 19660 39178 19672
rect 40862 19660 40868 19672
rect 40920 19660 40926 19712
rect 41414 19660 41420 19712
rect 41472 19700 41478 19712
rect 42061 19703 42119 19709
rect 42061 19700 42073 19703
rect 41472 19672 42073 19700
rect 41472 19660 41478 19672
rect 42061 19669 42073 19672
rect 42107 19669 42119 19703
rect 45462 19700 45468 19712
rect 45423 19672 45468 19700
rect 42061 19663 42119 19669
rect 45462 19660 45468 19672
rect 45520 19660 45526 19712
rect 1104 19610 48852 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 48852 19610
rect 1104 19536 48852 19558
rect 18690 19496 18696 19508
rect 18294 19468 18696 19496
rect 17129 19431 17187 19437
rect 17129 19397 17141 19431
rect 17175 19428 17187 19431
rect 17218 19428 17224 19440
rect 17175 19400 17224 19428
rect 17175 19397 17187 19400
rect 17129 19391 17187 19397
rect 17218 19388 17224 19400
rect 17276 19388 17282 19440
rect 2225 19363 2283 19369
rect 2225 19329 2237 19363
rect 2271 19360 2283 19363
rect 2406 19360 2412 19372
rect 2271 19332 2412 19360
rect 2271 19329 2283 19332
rect 2225 19323 2283 19329
rect 2406 19320 2412 19332
rect 2464 19360 2470 19372
rect 12342 19360 12348 19372
rect 2464 19332 12348 19360
rect 2464 19320 2470 19332
rect 12342 19320 12348 19332
rect 12400 19320 12406 19372
rect 17313 19363 17371 19369
rect 17313 19329 17325 19363
rect 17359 19360 17371 19363
rect 17402 19360 17408 19372
rect 17359 19332 17408 19360
rect 17359 19329 17371 19332
rect 17313 19323 17371 19329
rect 17402 19320 17408 19332
rect 17460 19320 17466 19372
rect 17954 19320 17960 19372
rect 18012 19360 18018 19372
rect 18294 19369 18322 19468
rect 18690 19456 18696 19468
rect 18748 19456 18754 19508
rect 22281 19499 22339 19505
rect 22281 19465 22293 19499
rect 22327 19496 22339 19499
rect 22922 19496 22928 19508
rect 22327 19468 22928 19496
rect 22327 19465 22339 19468
rect 22281 19459 22339 19465
rect 22922 19456 22928 19468
rect 22980 19456 22986 19508
rect 26602 19456 26608 19508
rect 26660 19496 26666 19508
rect 27071 19499 27129 19505
rect 27071 19496 27083 19499
rect 26660 19468 27083 19496
rect 26660 19456 26666 19468
rect 27071 19465 27083 19468
rect 27117 19465 27129 19499
rect 29270 19496 29276 19508
rect 29231 19468 29276 19496
rect 27071 19459 27129 19465
rect 29270 19456 29276 19468
rect 29328 19456 29334 19508
rect 29454 19456 29460 19508
rect 29512 19496 29518 19508
rect 33410 19496 33416 19508
rect 29512 19468 33416 19496
rect 29512 19456 29518 19468
rect 33410 19456 33416 19468
rect 33468 19456 33474 19508
rect 38194 19456 38200 19508
rect 38252 19496 38258 19508
rect 39215 19499 39273 19505
rect 39215 19496 39227 19499
rect 38252 19468 39227 19496
rect 38252 19456 38258 19468
rect 39215 19465 39227 19468
rect 39261 19465 39273 19499
rect 39215 19459 39273 19465
rect 39301 19499 39359 19505
rect 39301 19465 39313 19499
rect 39347 19496 39359 19499
rect 39390 19496 39396 19508
rect 39347 19468 39396 19496
rect 39347 19465 39359 19468
rect 39301 19459 39359 19465
rect 39390 19456 39396 19468
rect 39448 19456 39454 19508
rect 40770 19456 40776 19508
rect 40828 19496 40834 19508
rect 41874 19496 41880 19508
rect 40828 19468 41880 19496
rect 40828 19456 40834 19468
rect 41874 19456 41880 19468
rect 41932 19456 41938 19508
rect 46934 19496 46940 19508
rect 46895 19468 46940 19496
rect 46934 19456 46940 19468
rect 46992 19456 46998 19508
rect 18782 19388 18788 19440
rect 18840 19428 18846 19440
rect 34146 19428 34152 19440
rect 18840 19400 34152 19428
rect 18840 19388 18846 19400
rect 34146 19388 34152 19400
rect 34204 19388 34210 19440
rect 34425 19431 34483 19437
rect 34425 19397 34437 19431
rect 34471 19428 34483 19431
rect 35894 19428 35900 19440
rect 34471 19400 35900 19428
rect 34471 19397 34483 19400
rect 34425 19391 34483 19397
rect 35894 19388 35900 19400
rect 35952 19388 35958 19440
rect 37553 19431 37611 19437
rect 37553 19397 37565 19431
rect 37599 19428 37611 19431
rect 38102 19428 38108 19440
rect 37599 19400 38108 19428
rect 37599 19397 37611 19400
rect 37553 19391 37611 19397
rect 38102 19388 38108 19400
rect 38160 19428 38166 19440
rect 40788 19428 40816 19456
rect 38160 19400 39436 19428
rect 38160 19388 38166 19400
rect 18187 19363 18245 19369
rect 18187 19360 18199 19363
rect 18012 19332 18199 19360
rect 18012 19320 18018 19332
rect 18187 19329 18199 19332
rect 18233 19329 18245 19363
rect 18294 19363 18364 19369
rect 18294 19332 18318 19363
rect 18187 19323 18245 19329
rect 18306 19329 18318 19332
rect 18352 19329 18364 19363
rect 18306 19323 18364 19329
rect 18422 19363 18480 19369
rect 18422 19329 18434 19363
rect 18468 19329 18480 19363
rect 18422 19323 18480 19329
rect 18613 19363 18671 19369
rect 18613 19329 18625 19363
rect 18659 19360 18671 19363
rect 18874 19360 18880 19372
rect 18659 19332 18880 19360
rect 18659 19329 18671 19332
rect 18613 19323 18671 19329
rect 17497 19295 17555 19301
rect 17497 19261 17509 19295
rect 17543 19292 17555 19295
rect 18432 19292 18460 19323
rect 18874 19320 18880 19332
rect 18932 19320 18938 19372
rect 19978 19360 19984 19372
rect 19939 19332 19984 19360
rect 19978 19320 19984 19332
rect 20036 19320 20042 19372
rect 21821 19363 21879 19369
rect 21821 19329 21833 19363
rect 21867 19360 21879 19363
rect 22281 19363 22339 19369
rect 21867 19332 22094 19360
rect 21867 19329 21879 19332
rect 21821 19323 21879 19329
rect 17543 19264 18460 19292
rect 22066 19292 22094 19332
rect 22281 19329 22293 19363
rect 22327 19360 22339 19363
rect 22554 19360 22560 19372
rect 22327 19332 22560 19360
rect 22327 19329 22339 19332
rect 22281 19323 22339 19329
rect 22554 19320 22560 19332
rect 22612 19320 22618 19372
rect 23109 19363 23167 19369
rect 23109 19329 23121 19363
rect 23155 19360 23167 19363
rect 23474 19360 23480 19372
rect 23155 19332 23480 19360
rect 23155 19329 23167 19332
rect 23109 19323 23167 19329
rect 23474 19320 23480 19332
rect 23532 19360 23538 19372
rect 25130 19360 25136 19372
rect 23532 19332 25136 19360
rect 23532 19320 23538 19332
rect 25130 19320 25136 19332
rect 25188 19320 25194 19372
rect 25501 19363 25559 19369
rect 25501 19329 25513 19363
rect 25547 19360 25559 19363
rect 26234 19360 26240 19372
rect 25547 19332 26240 19360
rect 25547 19329 25559 19332
rect 25501 19323 25559 19329
rect 26234 19320 26240 19332
rect 26292 19360 26298 19372
rect 26418 19360 26424 19372
rect 26292 19332 26424 19360
rect 26292 19320 26298 19332
rect 26418 19320 26424 19332
rect 26476 19320 26482 19372
rect 26970 19360 26976 19372
rect 26931 19332 26976 19360
rect 26970 19320 26976 19332
rect 27028 19320 27034 19372
rect 27062 19320 27068 19372
rect 27120 19360 27126 19372
rect 27157 19363 27215 19369
rect 27157 19360 27169 19363
rect 27120 19332 27169 19360
rect 27120 19320 27126 19332
rect 27157 19329 27169 19332
rect 27203 19329 27215 19363
rect 27157 19323 27215 19329
rect 27249 19363 27307 19369
rect 27249 19329 27261 19363
rect 27295 19360 27307 19363
rect 27295 19332 27329 19360
rect 27295 19329 27307 19332
rect 27249 19323 27307 19329
rect 22370 19292 22376 19304
rect 22066 19264 22376 19292
rect 17543 19261 17555 19264
rect 17497 19255 17555 19261
rect 22370 19252 22376 19264
rect 22428 19252 22434 19304
rect 22830 19252 22836 19304
rect 22888 19292 22894 19304
rect 23201 19295 23259 19301
rect 23201 19292 23213 19295
rect 22888 19264 23213 19292
rect 22888 19252 22894 19264
rect 23201 19261 23213 19264
rect 23247 19261 23259 19295
rect 23382 19292 23388 19304
rect 23343 19264 23388 19292
rect 23201 19255 23259 19261
rect 23382 19252 23388 19264
rect 23440 19252 23446 19304
rect 25590 19292 25596 19304
rect 25551 19264 25596 19292
rect 25590 19252 25596 19264
rect 25648 19252 25654 19304
rect 25777 19295 25835 19301
rect 25777 19261 25789 19295
rect 25823 19292 25835 19295
rect 26142 19292 26148 19304
rect 25823 19264 26148 19292
rect 25823 19261 25835 19264
rect 25777 19255 25835 19261
rect 26142 19252 26148 19264
rect 26200 19252 26206 19304
rect 26786 19252 26792 19304
rect 26844 19292 26850 19304
rect 27264 19292 27292 19323
rect 29086 19320 29092 19372
rect 29144 19360 29150 19372
rect 29181 19363 29239 19369
rect 29181 19360 29193 19363
rect 29144 19332 29193 19360
rect 29144 19320 29150 19332
rect 29181 19329 29193 19332
rect 29227 19360 29239 19363
rect 30837 19363 30895 19369
rect 30837 19360 30849 19363
rect 29227 19332 30849 19360
rect 29227 19329 29239 19332
rect 29181 19323 29239 19329
rect 30837 19329 30849 19332
rect 30883 19360 30895 19363
rect 31018 19360 31024 19372
rect 30883 19332 31024 19360
rect 30883 19329 30895 19332
rect 30837 19323 30895 19329
rect 31018 19320 31024 19332
rect 31076 19320 31082 19372
rect 33410 19360 33416 19372
rect 33371 19332 33416 19360
rect 33410 19320 33416 19332
rect 33468 19320 33474 19372
rect 33505 19363 33563 19369
rect 33505 19329 33517 19363
rect 33551 19329 33563 19363
rect 33505 19323 33563 19329
rect 26844 19264 27292 19292
rect 26844 19252 26850 19264
rect 33520 19236 33548 19323
rect 33594 19320 33600 19372
rect 33652 19360 33658 19372
rect 33781 19363 33839 19369
rect 33652 19332 33697 19360
rect 33652 19320 33658 19332
rect 33781 19329 33793 19363
rect 33827 19360 33839 19363
rect 34054 19360 34060 19372
rect 33827 19332 34060 19360
rect 33827 19329 33839 19332
rect 33781 19323 33839 19329
rect 34054 19320 34060 19332
rect 34112 19320 34118 19372
rect 34241 19363 34299 19369
rect 34241 19329 34253 19363
rect 34287 19329 34299 19363
rect 34241 19323 34299 19329
rect 33870 19252 33876 19304
rect 33928 19292 33934 19304
rect 34256 19292 34284 19323
rect 36998 19320 37004 19372
rect 37056 19360 37062 19372
rect 37277 19363 37335 19369
rect 37277 19360 37289 19363
rect 37056 19332 37289 19360
rect 37056 19320 37062 19332
rect 37277 19329 37289 19332
rect 37323 19329 37335 19363
rect 38194 19360 38200 19372
rect 38155 19332 38200 19360
rect 37277 19323 37335 19329
rect 38194 19320 38200 19332
rect 38252 19320 38258 19372
rect 38378 19360 38384 19372
rect 38339 19332 38384 19360
rect 38378 19320 38384 19332
rect 38436 19320 38442 19372
rect 38473 19363 38531 19369
rect 38473 19329 38485 19363
rect 38519 19360 38531 19363
rect 39022 19360 39028 19372
rect 38519 19332 39028 19360
rect 38519 19329 38531 19332
rect 38473 19323 38531 19329
rect 39022 19320 39028 19332
rect 39080 19320 39086 19372
rect 39114 19320 39120 19372
rect 39172 19360 39178 19372
rect 39408 19369 39436 19400
rect 40328 19400 40816 19428
rect 40328 19369 40356 19400
rect 41322 19388 41328 19440
rect 41380 19428 41386 19440
rect 41417 19431 41475 19437
rect 41417 19428 41429 19431
rect 41380 19400 41429 19428
rect 41380 19388 41386 19400
rect 41417 19397 41429 19400
rect 41463 19397 41475 19431
rect 41417 19391 41475 19397
rect 39393 19363 39451 19369
rect 39172 19332 39217 19360
rect 39172 19320 39178 19332
rect 39393 19329 39405 19363
rect 39439 19329 39451 19363
rect 39393 19323 39451 19329
rect 40313 19363 40371 19369
rect 40313 19329 40325 19363
rect 40359 19329 40371 19363
rect 40313 19323 40371 19329
rect 40405 19363 40463 19369
rect 40405 19329 40417 19363
rect 40451 19360 40463 19363
rect 40678 19360 40684 19372
rect 40451 19332 40684 19360
rect 40451 19329 40463 19332
rect 40405 19323 40463 19329
rect 40678 19320 40684 19332
rect 40736 19360 40742 19372
rect 40954 19360 40960 19372
rect 40736 19332 40960 19360
rect 40736 19320 40742 19332
rect 40954 19320 40960 19332
rect 41012 19320 41018 19372
rect 41598 19320 41604 19372
rect 41656 19360 41662 19372
rect 42613 19363 42671 19369
rect 42613 19360 42625 19363
rect 41656 19332 42625 19360
rect 41656 19320 41662 19332
rect 42613 19329 42625 19332
rect 42659 19329 42671 19363
rect 42613 19323 42671 19329
rect 43162 19320 43168 19372
rect 43220 19360 43226 19372
rect 44818 19369 44824 19372
rect 43349 19363 43407 19369
rect 43349 19360 43361 19363
rect 43220 19332 43361 19360
rect 43220 19320 43226 19332
rect 43349 19329 43361 19332
rect 43395 19329 43407 19363
rect 43349 19323 43407 19329
rect 44812 19323 44824 19369
rect 44876 19360 44882 19372
rect 44876 19332 44912 19360
rect 44818 19320 44824 19323
rect 44876 19320 44882 19332
rect 45094 19320 45100 19372
rect 45152 19360 45158 19372
rect 46845 19363 46903 19369
rect 46845 19360 46857 19363
rect 45152 19332 46857 19360
rect 45152 19320 45158 19332
rect 46845 19329 46857 19332
rect 46891 19329 46903 19363
rect 47946 19360 47952 19372
rect 47907 19332 47952 19360
rect 46845 19323 46903 19329
rect 47946 19320 47952 19332
rect 48004 19320 48010 19372
rect 33928 19264 34284 19292
rect 33928 19252 33934 19264
rect 37458 19252 37464 19304
rect 37516 19292 37522 19304
rect 37553 19295 37611 19301
rect 37553 19292 37565 19295
rect 37516 19264 37565 19292
rect 37516 19252 37522 19264
rect 37553 19261 37565 19264
rect 37599 19261 37611 19295
rect 37553 19255 37611 19261
rect 38654 19252 38660 19304
rect 38712 19292 38718 19304
rect 43073 19295 43131 19301
rect 43073 19292 43085 19295
rect 38712 19264 43085 19292
rect 38712 19252 38718 19264
rect 43073 19261 43085 19264
rect 43119 19292 43131 19295
rect 43806 19292 43812 19304
rect 43119 19264 43812 19292
rect 43119 19261 43131 19264
rect 43073 19255 43131 19261
rect 43806 19252 43812 19264
rect 43864 19252 43870 19304
rect 44542 19292 44548 19304
rect 44503 19264 44548 19292
rect 44542 19252 44548 19264
rect 44600 19252 44606 19304
rect 22094 19184 22100 19236
rect 22152 19224 22158 19236
rect 22738 19224 22744 19236
rect 22152 19196 22744 19224
rect 22152 19184 22158 19196
rect 22738 19184 22744 19196
rect 22796 19184 22802 19236
rect 33502 19184 33508 19236
rect 33560 19184 33566 19236
rect 37274 19184 37280 19236
rect 37332 19224 37338 19236
rect 37369 19227 37427 19233
rect 37369 19224 37381 19227
rect 37332 19196 37381 19224
rect 37332 19184 37338 19196
rect 37369 19193 37381 19196
rect 37415 19193 37427 19227
rect 37369 19187 37427 19193
rect 40589 19227 40647 19233
rect 40589 19193 40601 19227
rect 40635 19224 40647 19227
rect 41049 19227 41107 19233
rect 41049 19224 41061 19227
rect 40635 19196 41061 19224
rect 40635 19193 40647 19196
rect 40589 19187 40647 19193
rect 41049 19193 41061 19196
rect 41095 19224 41107 19227
rect 41138 19224 41144 19236
rect 41095 19196 41144 19224
rect 41095 19193 41107 19196
rect 41049 19187 41107 19193
rect 41138 19184 41144 19196
rect 41196 19184 41202 19236
rect 41598 19224 41604 19236
rect 41559 19196 41604 19224
rect 41598 19184 41604 19196
rect 41656 19184 41662 19236
rect 1394 19116 1400 19168
rect 1452 19156 1458 19168
rect 1765 19159 1823 19165
rect 1765 19156 1777 19159
rect 1452 19128 1777 19156
rect 1452 19116 1458 19128
rect 1765 19125 1777 19128
rect 1811 19125 1823 19159
rect 2314 19156 2320 19168
rect 2275 19128 2320 19156
rect 1765 19119 1823 19125
rect 2314 19116 2320 19128
rect 2372 19116 2378 19168
rect 17954 19156 17960 19168
rect 17915 19128 17960 19156
rect 17954 19116 17960 19128
rect 18012 19116 18018 19168
rect 19610 19116 19616 19168
rect 19668 19156 19674 19168
rect 19797 19159 19855 19165
rect 19797 19156 19809 19159
rect 19668 19128 19809 19156
rect 19668 19116 19674 19128
rect 19797 19125 19809 19128
rect 19843 19125 19855 19159
rect 19797 19119 19855 19125
rect 21959 19159 22017 19165
rect 21959 19125 21971 19159
rect 22005 19156 22017 19159
rect 22186 19156 22192 19168
rect 22005 19128 22192 19156
rect 22005 19125 22017 19128
rect 21959 19119 22017 19125
rect 22186 19116 22192 19128
rect 22244 19116 22250 19168
rect 25133 19159 25191 19165
rect 25133 19125 25145 19159
rect 25179 19156 25191 19159
rect 25682 19156 25688 19168
rect 25179 19128 25688 19156
rect 25179 19125 25191 19128
rect 25133 19119 25191 19125
rect 25682 19116 25688 19128
rect 25740 19116 25746 19168
rect 30929 19159 30987 19165
rect 30929 19125 30941 19159
rect 30975 19156 30987 19159
rect 31662 19156 31668 19168
rect 30975 19128 31668 19156
rect 30975 19125 30987 19128
rect 30929 19119 30987 19125
rect 31662 19116 31668 19128
rect 31720 19116 31726 19168
rect 33134 19156 33140 19168
rect 33095 19128 33140 19156
rect 33134 19116 33140 19128
rect 33192 19116 33198 19168
rect 33778 19116 33784 19168
rect 33836 19156 33842 19168
rect 34609 19159 34667 19165
rect 34609 19156 34621 19159
rect 33836 19128 34621 19156
rect 33836 19116 33842 19128
rect 34609 19125 34621 19128
rect 34655 19125 34667 19159
rect 38470 19156 38476 19168
rect 38431 19128 38476 19156
rect 34609 19119 34667 19125
rect 38470 19116 38476 19128
rect 38528 19116 38534 19168
rect 38654 19156 38660 19168
rect 38615 19128 38660 19156
rect 38654 19116 38660 19128
rect 38712 19116 38718 19168
rect 41414 19116 41420 19168
rect 41472 19156 41478 19168
rect 42426 19156 42432 19168
rect 41472 19128 41517 19156
rect 42387 19128 42432 19156
rect 41472 19116 41478 19128
rect 42426 19116 42432 19128
rect 42484 19116 42490 19168
rect 45922 19156 45928 19168
rect 45883 19128 45928 19156
rect 45922 19116 45928 19128
rect 45980 19116 45986 19168
rect 48038 19156 48044 19168
rect 47999 19128 48044 19156
rect 48038 19116 48044 19128
rect 48096 19116 48102 19168
rect 1104 19066 48852 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 48852 19066
rect 1104 18992 48852 19014
rect 18414 18912 18420 18964
rect 18472 18952 18478 18964
rect 18509 18955 18567 18961
rect 18509 18952 18521 18955
rect 18472 18924 18521 18952
rect 18472 18912 18478 18924
rect 18509 18921 18521 18924
rect 18555 18921 18567 18955
rect 18509 18915 18567 18921
rect 22554 18912 22560 18964
rect 22612 18952 22618 18964
rect 24118 18952 24124 18964
rect 22612 18924 24124 18952
rect 22612 18912 22618 18924
rect 24118 18912 24124 18924
rect 24176 18912 24182 18964
rect 25547 18955 25605 18961
rect 25547 18921 25559 18955
rect 25593 18952 25605 18955
rect 25774 18952 25780 18964
rect 25593 18924 25780 18952
rect 25593 18921 25605 18924
rect 25547 18915 25605 18921
rect 25774 18912 25780 18924
rect 25832 18912 25838 18964
rect 32306 18912 32312 18964
rect 32364 18952 32370 18964
rect 32401 18955 32459 18961
rect 32401 18952 32413 18955
rect 32364 18924 32413 18952
rect 32364 18912 32370 18924
rect 32401 18921 32413 18924
rect 32447 18921 32459 18955
rect 32401 18915 32459 18921
rect 32968 18924 34008 18952
rect 22186 18844 22192 18896
rect 22244 18884 22250 18896
rect 22281 18887 22339 18893
rect 22281 18884 22293 18887
rect 22244 18856 22293 18884
rect 22244 18844 22250 18856
rect 22281 18853 22293 18856
rect 22327 18884 22339 18887
rect 25038 18884 25044 18896
rect 22327 18856 25044 18884
rect 22327 18853 22339 18856
rect 22281 18847 22339 18853
rect 25038 18844 25044 18856
rect 25096 18884 25102 18896
rect 26973 18887 27031 18893
rect 26973 18884 26985 18887
rect 25096 18856 26985 18884
rect 25096 18844 25102 18856
rect 26973 18853 26985 18856
rect 27019 18853 27031 18887
rect 26973 18847 27031 18853
rect 1394 18816 1400 18828
rect 1355 18788 1400 18816
rect 1394 18776 1400 18788
rect 1452 18776 1458 18828
rect 1581 18819 1639 18825
rect 1581 18785 1593 18819
rect 1627 18816 1639 18819
rect 2314 18816 2320 18828
rect 1627 18788 2320 18816
rect 1627 18785 1639 18788
rect 1581 18779 1639 18785
rect 2314 18776 2320 18788
rect 2372 18776 2378 18828
rect 2774 18816 2780 18828
rect 2735 18788 2780 18816
rect 2774 18776 2780 18788
rect 2832 18776 2838 18828
rect 22370 18816 22376 18828
rect 22331 18788 22376 18816
rect 22370 18776 22376 18788
rect 22428 18776 22434 18828
rect 23106 18816 23112 18828
rect 23067 18788 23112 18816
rect 23106 18776 23112 18788
rect 23164 18776 23170 18828
rect 31021 18819 31079 18825
rect 31021 18816 31033 18819
rect 24596 18788 25728 18816
rect 15746 18708 15752 18760
rect 15804 18748 15810 18760
rect 16301 18751 16359 18757
rect 16301 18748 16313 18751
rect 15804 18720 16313 18748
rect 15804 18708 15810 18720
rect 16301 18717 16313 18720
rect 16347 18748 16359 18751
rect 19334 18748 19340 18760
rect 16347 18720 19340 18748
rect 16347 18717 16359 18720
rect 16301 18711 16359 18717
rect 19334 18708 19340 18720
rect 19392 18708 19398 18760
rect 19610 18757 19616 18760
rect 19604 18748 19616 18757
rect 19571 18720 19616 18748
rect 19604 18711 19616 18720
rect 19610 18708 19616 18711
rect 19668 18708 19674 18760
rect 22094 18708 22100 18760
rect 22152 18748 22158 18760
rect 22152 18720 22197 18748
rect 22152 18708 22158 18720
rect 22738 18708 22744 18760
rect 22796 18748 22802 18760
rect 22833 18751 22891 18757
rect 22833 18748 22845 18751
rect 22796 18720 22845 18748
rect 22796 18708 22802 18720
rect 22833 18717 22845 18720
rect 22879 18717 22891 18751
rect 22833 18711 22891 18717
rect 23017 18751 23075 18757
rect 23017 18717 23029 18751
rect 23063 18717 23075 18751
rect 23017 18711 23075 18717
rect 23201 18751 23259 18757
rect 23201 18717 23213 18751
rect 23247 18717 23259 18751
rect 23201 18711 23259 18717
rect 23385 18751 23443 18757
rect 23385 18717 23397 18751
rect 23431 18748 23443 18751
rect 23474 18748 23480 18760
rect 23431 18720 23480 18748
rect 23431 18717 23443 18720
rect 23385 18711 23443 18717
rect 16568 18683 16626 18689
rect 16568 18649 16580 18683
rect 16614 18680 16626 18683
rect 17954 18680 17960 18692
rect 16614 18652 17960 18680
rect 16614 18649 16626 18652
rect 16568 18643 16626 18649
rect 17954 18640 17960 18652
rect 18012 18640 18018 18692
rect 18141 18683 18199 18689
rect 18141 18649 18153 18683
rect 18187 18680 18199 18683
rect 18230 18680 18236 18692
rect 18187 18652 18236 18680
rect 18187 18649 18199 18652
rect 18141 18643 18199 18649
rect 18230 18640 18236 18652
rect 18288 18640 18294 18692
rect 18325 18683 18383 18689
rect 18325 18649 18337 18683
rect 18371 18649 18383 18683
rect 18325 18643 18383 18649
rect 16666 18572 16672 18624
rect 16724 18612 16730 18624
rect 17402 18612 17408 18624
rect 16724 18584 17408 18612
rect 16724 18572 16730 18584
rect 17402 18572 17408 18584
rect 17460 18612 17466 18624
rect 17681 18615 17739 18621
rect 17681 18612 17693 18615
rect 17460 18584 17693 18612
rect 17460 18572 17466 18584
rect 17681 18581 17693 18584
rect 17727 18581 17739 18615
rect 17681 18575 17739 18581
rect 17862 18572 17868 18624
rect 17920 18612 17926 18624
rect 18340 18612 18368 18643
rect 19886 18640 19892 18692
rect 19944 18680 19950 18692
rect 21082 18680 21088 18692
rect 19944 18652 21088 18680
rect 19944 18640 19950 18652
rect 21082 18640 21088 18652
rect 21140 18640 21146 18692
rect 21913 18683 21971 18689
rect 21913 18649 21925 18683
rect 21959 18680 21971 18683
rect 23032 18680 23060 18711
rect 21959 18652 23060 18680
rect 23216 18680 23244 18711
rect 23474 18708 23480 18720
rect 23532 18708 23538 18760
rect 24596 18757 24624 18788
rect 25700 18760 25728 18788
rect 29656 18788 31033 18816
rect 24581 18751 24639 18757
rect 24581 18717 24593 18751
rect 24627 18717 24639 18751
rect 24762 18748 24768 18760
rect 24723 18720 24768 18748
rect 24581 18711 24639 18717
rect 24762 18708 24768 18720
rect 24820 18708 24826 18760
rect 24857 18751 24915 18757
rect 24857 18717 24869 18751
rect 24903 18748 24915 18751
rect 24946 18748 24952 18760
rect 24903 18720 24952 18748
rect 24903 18717 24915 18720
rect 24857 18711 24915 18717
rect 24946 18708 24952 18720
rect 25004 18748 25010 18760
rect 25314 18748 25320 18760
rect 25004 18720 25320 18748
rect 25004 18708 25010 18720
rect 25314 18708 25320 18720
rect 25372 18708 25378 18760
rect 25682 18708 25688 18760
rect 25740 18748 25746 18760
rect 26605 18751 26663 18757
rect 26605 18748 26617 18751
rect 25740 18720 26617 18748
rect 25740 18708 25746 18720
rect 26605 18717 26617 18720
rect 26651 18717 26663 18751
rect 26605 18711 26663 18717
rect 27433 18751 27491 18757
rect 27433 18717 27445 18751
rect 27479 18748 27491 18751
rect 29656 18748 29684 18788
rect 31021 18785 31033 18788
rect 31067 18785 31079 18819
rect 31021 18779 31079 18785
rect 27479 18720 29684 18748
rect 27479 18717 27491 18720
rect 27433 18711 27491 18717
rect 29730 18708 29736 18760
rect 29788 18748 29794 18760
rect 30009 18751 30067 18757
rect 29788 18720 29833 18748
rect 29788 18708 29794 18720
rect 30009 18717 30021 18751
rect 30055 18748 30067 18751
rect 30834 18748 30840 18760
rect 30055 18720 30840 18748
rect 30055 18717 30067 18720
rect 30009 18711 30067 18717
rect 30834 18708 30840 18720
rect 30892 18708 30898 18760
rect 31036 18748 31064 18779
rect 31754 18748 31760 18760
rect 31036 18720 31760 18748
rect 31754 18708 31760 18720
rect 31812 18708 31818 18760
rect 23842 18680 23848 18692
rect 23216 18652 23848 18680
rect 21959 18649 21971 18652
rect 21913 18643 21971 18649
rect 23842 18640 23848 18652
rect 23900 18640 23906 18692
rect 26786 18680 26792 18692
rect 26747 18652 26792 18680
rect 26786 18640 26792 18652
rect 26844 18640 26850 18692
rect 27700 18683 27758 18689
rect 27700 18649 27712 18683
rect 27746 18680 27758 18683
rect 27890 18680 27896 18692
rect 27746 18652 27896 18680
rect 27746 18649 27758 18652
rect 27700 18643 27758 18649
rect 27890 18640 27896 18652
rect 27948 18640 27954 18692
rect 28350 18640 28356 18692
rect 28408 18680 28414 18692
rect 28408 18652 28948 18680
rect 28408 18640 28414 18652
rect 17920 18584 18368 18612
rect 17920 18572 17926 18584
rect 20622 18572 20628 18624
rect 20680 18612 20686 18624
rect 20717 18615 20775 18621
rect 20717 18612 20729 18615
rect 20680 18584 20729 18612
rect 20680 18572 20686 18584
rect 20717 18581 20729 18584
rect 20763 18581 20775 18615
rect 20717 18575 20775 18581
rect 22186 18572 22192 18624
rect 22244 18612 22250 18624
rect 23569 18615 23627 18621
rect 23569 18612 23581 18615
rect 22244 18584 23581 18612
rect 22244 18572 22250 18584
rect 23569 18581 23581 18584
rect 23615 18581 23627 18615
rect 23569 18575 23627 18581
rect 24397 18615 24455 18621
rect 24397 18581 24409 18615
rect 24443 18612 24455 18615
rect 25406 18612 25412 18624
rect 24443 18584 25412 18612
rect 24443 18581 24455 18584
rect 24397 18575 24455 18581
rect 25406 18572 25412 18584
rect 25464 18572 25470 18624
rect 27430 18572 27436 18624
rect 27488 18612 27494 18624
rect 28813 18615 28871 18621
rect 28813 18612 28825 18615
rect 27488 18584 28825 18612
rect 27488 18572 27494 18584
rect 28813 18581 28825 18584
rect 28859 18581 28871 18615
rect 28920 18612 28948 18652
rect 28994 18640 29000 18692
rect 29052 18680 29058 18692
rect 29748 18680 29776 18708
rect 29052 18652 29776 18680
rect 29052 18640 29058 18652
rect 30926 18640 30932 18692
rect 30984 18680 30990 18692
rect 31266 18683 31324 18689
rect 31266 18680 31278 18683
rect 30984 18652 31278 18680
rect 30984 18640 30990 18652
rect 31266 18649 31278 18652
rect 31312 18649 31324 18683
rect 31266 18643 31324 18649
rect 31662 18640 31668 18692
rect 31720 18680 31726 18692
rect 32968 18680 32996 18924
rect 33502 18844 33508 18896
rect 33560 18844 33566 18896
rect 33042 18776 33048 18828
rect 33100 18816 33106 18828
rect 33520 18816 33548 18844
rect 33100 18788 33732 18816
rect 33100 18776 33106 18788
rect 33502 18708 33508 18760
rect 33560 18748 33566 18760
rect 33704 18757 33732 18788
rect 33597 18751 33655 18757
rect 33597 18748 33609 18751
rect 33560 18720 33609 18748
rect 33560 18708 33566 18720
rect 33597 18717 33609 18720
rect 33643 18717 33655 18751
rect 33597 18711 33655 18717
rect 33689 18751 33747 18757
rect 33689 18717 33701 18751
rect 33735 18717 33747 18751
rect 33689 18711 33747 18717
rect 33778 18708 33784 18760
rect 33836 18748 33842 18760
rect 33980 18757 34008 18924
rect 35894 18912 35900 18964
rect 35952 18952 35958 18964
rect 36081 18955 36139 18961
rect 36081 18952 36093 18955
rect 35952 18924 36093 18952
rect 35952 18912 35958 18924
rect 36081 18921 36093 18924
rect 36127 18921 36139 18955
rect 36081 18915 36139 18921
rect 37366 18912 37372 18964
rect 37424 18952 37430 18964
rect 37829 18955 37887 18961
rect 37829 18952 37841 18955
rect 37424 18924 37841 18952
rect 37424 18912 37430 18924
rect 37829 18921 37841 18924
rect 37875 18921 37887 18955
rect 37829 18915 37887 18921
rect 39022 18912 39028 18964
rect 39080 18952 39086 18964
rect 39117 18955 39175 18961
rect 39117 18952 39129 18955
rect 39080 18924 39129 18952
rect 39080 18912 39086 18924
rect 39117 18921 39129 18924
rect 39163 18921 39175 18955
rect 39117 18915 39175 18921
rect 40405 18955 40463 18961
rect 40405 18921 40417 18955
rect 40451 18952 40463 18955
rect 40770 18952 40776 18964
rect 40451 18924 40776 18952
rect 40451 18921 40463 18924
rect 40405 18915 40463 18921
rect 40770 18912 40776 18924
rect 40828 18912 40834 18964
rect 41417 18955 41475 18961
rect 41417 18921 41429 18955
rect 41463 18952 41475 18955
rect 41506 18952 41512 18964
rect 41463 18924 41512 18952
rect 41463 18921 41475 18924
rect 41417 18915 41475 18921
rect 41506 18912 41512 18924
rect 41564 18912 41570 18964
rect 37461 18887 37519 18893
rect 37461 18853 37473 18887
rect 37507 18884 37519 18887
rect 40589 18887 40647 18893
rect 37507 18856 40540 18884
rect 37507 18853 37519 18856
rect 37461 18847 37519 18853
rect 38746 18816 38752 18828
rect 38707 18788 38752 18816
rect 38746 18776 38752 18788
rect 38804 18776 38810 18828
rect 40512 18816 40540 18856
rect 40589 18853 40601 18887
rect 40635 18884 40647 18887
rect 41046 18884 41052 18896
rect 40635 18856 41052 18884
rect 40635 18853 40647 18856
rect 40589 18847 40647 18853
rect 41046 18844 41052 18856
rect 41104 18844 41110 18896
rect 45370 18844 45376 18896
rect 45428 18844 45434 18896
rect 45462 18844 45468 18896
rect 45520 18844 45526 18896
rect 46106 18844 46112 18896
rect 46164 18884 46170 18896
rect 46164 18856 47164 18884
rect 46164 18844 46170 18856
rect 40770 18816 40776 18828
rect 40512 18788 40776 18816
rect 40770 18776 40776 18788
rect 40828 18776 40834 18828
rect 41230 18776 41236 18828
rect 41288 18816 41294 18828
rect 41288 18788 42104 18816
rect 41288 18776 41294 18788
rect 33965 18751 34023 18757
rect 33836 18720 33881 18748
rect 33836 18708 33842 18720
rect 33965 18717 33977 18751
rect 34011 18748 34023 18751
rect 34054 18748 34060 18760
rect 34011 18720 34060 18748
rect 34011 18717 34023 18720
rect 33965 18711 34023 18717
rect 34054 18708 34060 18720
rect 34112 18708 34118 18760
rect 34701 18751 34759 18757
rect 34701 18717 34713 18751
rect 34747 18748 34759 18751
rect 35986 18748 35992 18760
rect 34747 18720 35992 18748
rect 34747 18717 34759 18720
rect 34701 18711 34759 18717
rect 35986 18708 35992 18720
rect 36044 18708 36050 18760
rect 37737 18751 37795 18757
rect 37737 18717 37749 18751
rect 37783 18717 37795 18751
rect 37918 18748 37924 18760
rect 37879 18720 37924 18748
rect 37737 18711 37795 18717
rect 31720 18652 32996 18680
rect 33321 18683 33379 18689
rect 31720 18640 31726 18652
rect 33321 18649 33333 18683
rect 33367 18680 33379 18683
rect 34946 18683 35004 18689
rect 34946 18680 34958 18683
rect 33367 18652 34958 18680
rect 33367 18649 33379 18652
rect 33321 18643 33379 18649
rect 34946 18649 34958 18652
rect 34992 18649 35004 18683
rect 37752 18680 37780 18711
rect 37918 18708 37924 18720
rect 37976 18708 37982 18760
rect 38010 18708 38016 18760
rect 38068 18748 38074 18760
rect 38197 18751 38255 18757
rect 38068 18720 38113 18748
rect 38068 18708 38074 18720
rect 38197 18717 38209 18751
rect 38243 18748 38255 18751
rect 38654 18748 38660 18760
rect 38243 18720 38660 18748
rect 38243 18717 38255 18720
rect 38197 18711 38255 18717
rect 38654 18708 38660 18720
rect 38712 18708 38718 18760
rect 42076 18757 42104 18788
rect 43070 18776 43076 18828
rect 43128 18816 43134 18828
rect 43128 18788 44680 18816
rect 43128 18776 43134 18788
rect 38841 18751 38899 18757
rect 38841 18717 38853 18751
rect 38887 18748 38899 18751
rect 42061 18751 42119 18757
rect 38887 18720 40356 18748
rect 38887 18717 38899 18720
rect 38841 18711 38899 18717
rect 40218 18680 40224 18692
rect 34946 18643 35004 18649
rect 36004 18652 37780 18680
rect 40179 18652 40224 18680
rect 36004 18612 36032 18652
rect 40218 18640 40224 18652
rect 40276 18640 40282 18692
rect 40328 18680 40356 18720
rect 42061 18717 42073 18751
rect 42107 18748 42119 18751
rect 44542 18748 44548 18760
rect 42107 18720 44548 18748
rect 42107 18717 42119 18720
rect 42061 18711 42119 18717
rect 44542 18708 44548 18720
rect 44600 18708 44606 18760
rect 44652 18748 44680 18788
rect 45388 18757 45416 18844
rect 45480 18757 45508 18844
rect 46477 18819 46535 18825
rect 46477 18785 46489 18819
rect 46523 18816 46535 18819
rect 47026 18816 47032 18828
rect 46523 18788 47032 18816
rect 46523 18785 46535 18788
rect 46477 18779 46535 18785
rect 47026 18776 47032 18788
rect 47084 18776 47090 18828
rect 47136 18825 47164 18856
rect 47121 18819 47179 18825
rect 47121 18785 47133 18819
rect 47167 18785 47179 18819
rect 47121 18779 47179 18785
rect 45235 18751 45293 18757
rect 45235 18748 45247 18751
rect 44652 18720 45247 18748
rect 45235 18717 45247 18720
rect 45281 18717 45293 18751
rect 45235 18711 45293 18717
rect 45370 18751 45428 18757
rect 45370 18717 45382 18751
rect 45416 18717 45428 18751
rect 45370 18711 45428 18717
rect 45465 18751 45523 18757
rect 45465 18717 45477 18751
rect 45511 18717 45523 18751
rect 45646 18748 45652 18760
rect 45607 18720 45652 18748
rect 45465 18711 45523 18717
rect 45646 18708 45652 18720
rect 45704 18708 45710 18760
rect 45738 18708 45744 18760
rect 45796 18748 45802 18760
rect 46293 18751 46351 18757
rect 46293 18748 46305 18751
rect 45796 18720 46305 18748
rect 45796 18708 45802 18720
rect 46293 18717 46305 18720
rect 46339 18717 46351 18751
rect 46293 18711 46351 18717
rect 42328 18683 42386 18689
rect 40328 18652 42288 18680
rect 28920 18584 36032 18612
rect 40431 18615 40489 18621
rect 28813 18575 28871 18581
rect 40431 18581 40443 18615
rect 40477 18612 40489 18615
rect 40678 18612 40684 18624
rect 40477 18584 40684 18612
rect 40477 18581 40489 18584
rect 40431 18575 40489 18581
rect 40678 18572 40684 18584
rect 40736 18572 40742 18624
rect 40770 18572 40776 18624
rect 40828 18612 40834 18624
rect 41322 18612 41328 18624
rect 40828 18584 41328 18612
rect 40828 18572 40834 18584
rect 41322 18572 41328 18584
rect 41380 18612 41386 18624
rect 41417 18615 41475 18621
rect 41417 18612 41429 18615
rect 41380 18584 41429 18612
rect 41380 18572 41386 18584
rect 41417 18581 41429 18584
rect 41463 18581 41475 18615
rect 41417 18575 41475 18581
rect 41601 18615 41659 18621
rect 41601 18581 41613 18615
rect 41647 18612 41659 18615
rect 42150 18612 42156 18624
rect 41647 18584 42156 18612
rect 41647 18581 41659 18584
rect 41601 18575 41659 18581
rect 42150 18572 42156 18584
rect 42208 18572 42214 18624
rect 42260 18612 42288 18652
rect 42328 18649 42340 18683
rect 42374 18680 42386 18683
rect 42426 18680 42432 18692
rect 42374 18652 42432 18680
rect 42374 18649 42386 18652
rect 42328 18643 42386 18649
rect 42426 18640 42432 18652
rect 42484 18640 42490 18692
rect 44082 18680 44088 18692
rect 44043 18652 44088 18680
rect 44082 18640 44088 18652
rect 44140 18640 44146 18692
rect 44269 18683 44327 18689
rect 44269 18649 44281 18683
rect 44315 18680 44327 18683
rect 45922 18680 45928 18692
rect 44315 18652 45928 18680
rect 44315 18649 44327 18652
rect 44269 18643 44327 18649
rect 45922 18640 45928 18652
rect 45980 18640 45986 18692
rect 43254 18612 43260 18624
rect 42260 18584 43260 18612
rect 43254 18572 43260 18584
rect 43312 18612 43318 18624
rect 43441 18615 43499 18621
rect 43441 18612 43453 18615
rect 43312 18584 43453 18612
rect 43312 18572 43318 18584
rect 43441 18581 43453 18584
rect 43487 18581 43499 18615
rect 44450 18612 44456 18624
rect 44411 18584 44456 18612
rect 43441 18575 43499 18581
rect 44450 18572 44456 18584
rect 44508 18572 44514 18624
rect 45002 18612 45008 18624
rect 44963 18584 45008 18612
rect 45002 18572 45008 18584
rect 45060 18572 45066 18624
rect 1104 18522 48852 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 48852 18522
rect 1104 18448 48852 18470
rect 15746 18408 15752 18420
rect 15304 18380 15752 18408
rect 15304 18349 15332 18380
rect 15746 18368 15752 18380
rect 15804 18368 15810 18420
rect 19978 18368 19984 18420
rect 20036 18408 20042 18420
rect 20257 18411 20315 18417
rect 20257 18408 20269 18411
rect 20036 18380 20269 18408
rect 20036 18368 20042 18380
rect 20257 18377 20269 18380
rect 20303 18377 20315 18411
rect 20257 18371 20315 18377
rect 21910 18368 21916 18420
rect 21968 18408 21974 18420
rect 22005 18411 22063 18417
rect 22005 18408 22017 18411
rect 21968 18380 22017 18408
rect 21968 18368 21974 18380
rect 22005 18377 22017 18380
rect 22051 18377 22063 18411
rect 22005 18371 22063 18377
rect 22373 18411 22431 18417
rect 22373 18377 22385 18411
rect 22419 18408 22431 18411
rect 22830 18408 22836 18420
rect 22419 18380 22836 18408
rect 22419 18377 22431 18380
rect 22373 18371 22431 18377
rect 22830 18368 22836 18380
rect 22888 18368 22894 18420
rect 23014 18368 23020 18420
rect 23072 18408 23078 18420
rect 23072 18380 23152 18408
rect 23072 18368 23078 18380
rect 15289 18343 15347 18349
rect 15289 18309 15301 18343
rect 15335 18309 15347 18343
rect 15289 18303 15347 18309
rect 15378 18300 15384 18352
rect 15436 18340 15442 18352
rect 17028 18343 17086 18349
rect 15436 18312 15481 18340
rect 15436 18300 15442 18312
rect 17028 18309 17040 18343
rect 17074 18340 17086 18343
rect 18046 18340 18052 18352
rect 17074 18312 18052 18340
rect 17074 18309 17086 18312
rect 17028 18303 17086 18309
rect 18046 18300 18052 18312
rect 18104 18300 18110 18352
rect 20717 18343 20775 18349
rect 20717 18309 20729 18343
rect 20763 18340 20775 18343
rect 22848 18340 22876 18368
rect 22925 18343 22983 18349
rect 22925 18340 22937 18343
rect 20763 18312 22784 18340
rect 22848 18312 22937 18340
rect 20763 18309 20775 18312
rect 20717 18303 20775 18309
rect 1946 18232 1952 18284
rect 2004 18272 2010 18284
rect 2041 18275 2099 18281
rect 2041 18272 2053 18275
rect 2004 18244 2053 18272
rect 2004 18232 2010 18244
rect 2041 18241 2053 18244
rect 2087 18241 2099 18275
rect 20622 18272 20628 18284
rect 20535 18244 20628 18272
rect 2041 18235 2099 18241
rect 20622 18232 20628 18244
rect 20680 18272 20686 18284
rect 20680 18244 22094 18272
rect 20680 18232 20686 18244
rect 15565 18207 15623 18213
rect 15565 18173 15577 18207
rect 15611 18173 15623 18207
rect 15565 18167 15623 18173
rect 16761 18207 16819 18213
rect 16761 18173 16773 18207
rect 16807 18173 16819 18207
rect 16761 18167 16819 18173
rect 20901 18207 20959 18213
rect 20901 18173 20913 18207
rect 20947 18204 20959 18207
rect 20990 18204 20996 18216
rect 20947 18176 20996 18204
rect 20947 18173 20959 18176
rect 20901 18167 20959 18173
rect 3418 18096 3424 18148
rect 3476 18136 3482 18148
rect 15580 18136 15608 18167
rect 3476 18108 15608 18136
rect 3476 18096 3482 18108
rect 1578 18028 1584 18080
rect 1636 18068 1642 18080
rect 2133 18071 2191 18077
rect 2133 18068 2145 18071
rect 1636 18040 2145 18068
rect 1636 18028 1642 18040
rect 2133 18037 2145 18040
rect 2179 18037 2191 18071
rect 2866 18068 2872 18080
rect 2827 18040 2872 18068
rect 2133 18031 2191 18037
rect 2866 18028 2872 18040
rect 2924 18028 2930 18080
rect 16776 18068 16804 18167
rect 20990 18164 20996 18176
rect 21048 18164 21054 18216
rect 17862 18096 17868 18148
rect 17920 18136 17926 18148
rect 18141 18139 18199 18145
rect 18141 18136 18153 18139
rect 17920 18108 18153 18136
rect 17920 18096 17926 18108
rect 18141 18105 18153 18108
rect 18187 18105 18199 18139
rect 22066 18136 22094 18244
rect 22186 18232 22192 18284
rect 22244 18272 22250 18284
rect 22465 18275 22523 18281
rect 22244 18244 22289 18272
rect 22244 18232 22250 18244
rect 22465 18241 22477 18275
rect 22511 18272 22523 18275
rect 22554 18272 22560 18284
rect 22511 18244 22560 18272
rect 22511 18241 22523 18244
rect 22465 18235 22523 18241
rect 22554 18232 22560 18244
rect 22612 18232 22618 18284
rect 22756 18204 22784 18312
rect 22925 18309 22937 18312
rect 22971 18309 22983 18343
rect 22925 18303 22983 18309
rect 23124 18281 23152 18380
rect 24762 18368 24768 18420
rect 24820 18408 24826 18420
rect 25685 18411 25743 18417
rect 25685 18408 25697 18411
rect 24820 18380 25697 18408
rect 24820 18368 24826 18380
rect 25685 18377 25697 18380
rect 25731 18408 25743 18411
rect 26786 18408 26792 18420
rect 25731 18380 26792 18408
rect 25731 18377 25743 18380
rect 25685 18371 25743 18377
rect 26786 18368 26792 18380
rect 26844 18368 26850 18420
rect 27890 18408 27896 18420
rect 27851 18380 27896 18408
rect 27890 18368 27896 18380
rect 27948 18368 27954 18420
rect 28258 18368 28264 18420
rect 28316 18408 28322 18420
rect 28537 18411 28595 18417
rect 28537 18408 28549 18411
rect 28316 18380 28549 18408
rect 28316 18368 28322 18380
rect 28537 18377 28549 18380
rect 28583 18377 28595 18411
rect 30926 18408 30932 18420
rect 30887 18380 30932 18408
rect 28537 18371 28595 18377
rect 30926 18368 30932 18380
rect 30984 18368 30990 18420
rect 37918 18368 37924 18420
rect 37976 18408 37982 18420
rect 38657 18411 38715 18417
rect 38657 18408 38669 18411
rect 37976 18380 38669 18408
rect 37976 18368 37982 18380
rect 38657 18377 38669 18380
rect 38703 18377 38715 18411
rect 41506 18408 41512 18420
rect 41467 18380 41512 18408
rect 38657 18371 38715 18377
rect 41506 18368 41512 18380
rect 41564 18368 41570 18420
rect 43806 18408 43812 18420
rect 43767 18380 43812 18408
rect 43806 18368 43812 18380
rect 43864 18368 43870 18420
rect 46290 18368 46296 18420
rect 46348 18408 46354 18420
rect 46477 18411 46535 18417
rect 46477 18408 46489 18411
rect 46348 18380 46489 18408
rect 46348 18368 46354 18380
rect 46477 18377 46489 18380
rect 46523 18377 46535 18411
rect 46477 18371 46535 18377
rect 25590 18340 25596 18352
rect 23216 18312 25596 18340
rect 23216 18284 23244 18312
rect 25590 18300 25596 18312
rect 25648 18300 25654 18352
rect 26418 18300 26424 18352
rect 26476 18340 26482 18352
rect 32493 18343 32551 18349
rect 32493 18340 32505 18343
rect 26476 18312 31248 18340
rect 26476 18300 26482 18312
rect 23109 18275 23167 18281
rect 23109 18241 23121 18275
rect 23155 18241 23167 18275
rect 23109 18235 23167 18241
rect 23198 18232 23204 18284
rect 23256 18272 23262 18284
rect 23256 18244 23349 18272
rect 23256 18232 23262 18244
rect 23382 18232 23388 18284
rect 23440 18272 23446 18284
rect 23845 18275 23903 18281
rect 23845 18272 23857 18275
rect 23440 18244 23857 18272
rect 23440 18232 23446 18244
rect 23845 18241 23857 18244
rect 23891 18241 23903 18275
rect 23845 18235 23903 18241
rect 24949 18275 25007 18281
rect 24949 18241 24961 18275
rect 24995 18272 25007 18275
rect 25314 18272 25320 18284
rect 24995 18244 25320 18272
rect 24995 18241 25007 18244
rect 24949 18235 25007 18241
rect 25314 18232 25320 18244
rect 25372 18232 25378 18284
rect 26053 18275 26111 18281
rect 26053 18241 26065 18275
rect 26099 18272 26111 18275
rect 26602 18272 26608 18284
rect 26099 18244 26608 18272
rect 26099 18241 26111 18244
rect 26053 18235 26111 18241
rect 26602 18232 26608 18244
rect 26660 18232 26666 18284
rect 27154 18272 27160 18284
rect 27115 18244 27160 18272
rect 27154 18232 27160 18244
rect 27212 18232 27218 18284
rect 27338 18272 27344 18284
rect 27299 18244 27344 18272
rect 27338 18232 27344 18244
rect 27396 18232 27402 18284
rect 27525 18275 27583 18281
rect 27525 18241 27537 18275
rect 27571 18272 27583 18275
rect 27614 18272 27620 18284
rect 27571 18244 27620 18272
rect 27571 18241 27583 18244
rect 27525 18235 27583 18241
rect 27614 18232 27620 18244
rect 27672 18232 27678 18284
rect 27709 18275 27767 18281
rect 27709 18241 27721 18275
rect 27755 18241 27767 18275
rect 28350 18272 28356 18284
rect 28311 18244 28356 18272
rect 27709 18235 27767 18241
rect 25130 18204 25136 18216
rect 22756 18176 25136 18204
rect 25130 18164 25136 18176
rect 25188 18164 25194 18216
rect 25225 18207 25283 18213
rect 25225 18173 25237 18207
rect 25271 18204 25283 18207
rect 25774 18204 25780 18216
rect 25271 18176 25780 18204
rect 25271 18173 25283 18176
rect 25225 18167 25283 18173
rect 25774 18164 25780 18176
rect 25832 18164 25838 18216
rect 26145 18207 26203 18213
rect 26145 18173 26157 18207
rect 26191 18173 26203 18207
rect 26145 18167 26203 18173
rect 23014 18136 23020 18148
rect 22066 18108 23020 18136
rect 18141 18099 18199 18105
rect 23014 18096 23020 18108
rect 23072 18096 23078 18148
rect 26160 18136 26188 18167
rect 26234 18164 26240 18216
rect 26292 18204 26298 18216
rect 27430 18204 27436 18216
rect 26292 18176 26337 18204
rect 27343 18176 27436 18204
rect 26292 18164 26298 18176
rect 27430 18164 27436 18176
rect 27488 18164 27494 18216
rect 27448 18136 27476 18164
rect 23124 18108 27476 18136
rect 27724 18136 27752 18235
rect 28350 18232 28356 18244
rect 28408 18232 28414 18284
rect 30006 18272 30012 18284
rect 29967 18244 30012 18272
rect 30006 18232 30012 18244
rect 30064 18232 30070 18284
rect 31220 18281 31248 18312
rect 31404 18312 32505 18340
rect 31404 18281 31432 18312
rect 32493 18309 32505 18312
rect 32539 18309 32551 18343
rect 32493 18303 32551 18309
rect 33134 18300 33140 18352
rect 33192 18340 33198 18352
rect 34210 18343 34268 18349
rect 34210 18340 34222 18343
rect 33192 18312 34222 18340
rect 33192 18300 33198 18312
rect 34210 18309 34222 18312
rect 34256 18309 34268 18343
rect 41138 18340 41144 18352
rect 41099 18312 41144 18340
rect 34210 18303 34268 18309
rect 41138 18300 41144 18312
rect 41196 18300 41202 18352
rect 45002 18300 45008 18352
rect 45060 18340 45066 18352
rect 45342 18343 45400 18349
rect 45342 18340 45354 18343
rect 45060 18312 45354 18340
rect 45060 18300 45066 18312
rect 45342 18309 45354 18312
rect 45388 18309 45400 18343
rect 45342 18303 45400 18309
rect 31205 18275 31263 18281
rect 31205 18241 31217 18275
rect 31251 18241 31263 18275
rect 31205 18235 31263 18241
rect 31297 18275 31355 18281
rect 31297 18241 31309 18275
rect 31343 18241 31355 18275
rect 31297 18235 31355 18241
rect 31389 18275 31447 18281
rect 31389 18241 31401 18275
rect 31435 18241 31447 18275
rect 31389 18235 31447 18241
rect 31573 18275 31631 18281
rect 31573 18241 31585 18275
rect 31619 18272 31631 18275
rect 31662 18272 31668 18284
rect 31619 18244 31668 18272
rect 31619 18241 31631 18244
rect 31573 18235 31631 18241
rect 29362 18164 29368 18216
rect 29420 18204 29426 18216
rect 29825 18207 29883 18213
rect 29825 18204 29837 18207
rect 29420 18176 29837 18204
rect 29420 18164 29426 18176
rect 29825 18173 29837 18176
rect 29871 18173 29883 18207
rect 31312 18204 31340 18235
rect 31662 18232 31668 18244
rect 31720 18232 31726 18284
rect 31754 18232 31760 18284
rect 31812 18272 31818 18284
rect 31812 18244 32076 18272
rect 31812 18232 31818 18244
rect 31846 18204 31852 18216
rect 31312 18176 31852 18204
rect 29825 18167 29883 18173
rect 31846 18164 31852 18176
rect 31904 18164 31910 18216
rect 32048 18204 32076 18244
rect 32122 18232 32128 18284
rect 32180 18272 32186 18284
rect 32306 18272 32312 18284
rect 32180 18244 32225 18272
rect 32267 18244 32312 18272
rect 32180 18232 32186 18244
rect 32306 18232 32312 18244
rect 32364 18232 32370 18284
rect 36538 18232 36544 18284
rect 36596 18272 36602 18284
rect 37461 18275 37519 18281
rect 37461 18272 37473 18275
rect 36596 18244 37473 18272
rect 36596 18232 36602 18244
rect 37461 18241 37473 18244
rect 37507 18241 37519 18275
rect 37918 18272 37924 18284
rect 37831 18244 37924 18272
rect 37461 18235 37519 18241
rect 32858 18204 32864 18216
rect 32048 18176 32864 18204
rect 32858 18164 32864 18176
rect 32916 18204 32922 18216
rect 33965 18207 34023 18213
rect 33965 18204 33977 18207
rect 32916 18176 33977 18204
rect 32916 18164 32922 18176
rect 33965 18173 33977 18176
rect 34011 18173 34023 18207
rect 33965 18167 34023 18173
rect 37553 18207 37611 18213
rect 37553 18173 37565 18207
rect 37599 18204 37611 18207
rect 37642 18204 37648 18216
rect 37599 18176 37648 18204
rect 37599 18173 37611 18176
rect 37553 18167 37611 18173
rect 37642 18164 37648 18176
rect 37700 18164 37706 18216
rect 37844 18213 37872 18244
rect 37918 18232 37924 18244
rect 37976 18272 37982 18284
rect 38473 18275 38531 18281
rect 38473 18272 38485 18275
rect 37976 18244 38485 18272
rect 37976 18232 37982 18244
rect 38473 18241 38485 18244
rect 38519 18241 38531 18275
rect 38473 18235 38531 18241
rect 40218 18232 40224 18284
rect 40276 18272 40282 18284
rect 40862 18272 40868 18284
rect 40276 18244 40868 18272
rect 40276 18232 40282 18244
rect 40862 18232 40868 18244
rect 40920 18272 40926 18284
rect 41325 18275 41383 18281
rect 41325 18272 41337 18275
rect 40920 18244 41337 18272
rect 40920 18232 40926 18244
rect 41325 18241 41337 18244
rect 41371 18241 41383 18275
rect 41325 18235 41383 18241
rect 41966 18232 41972 18284
rect 42024 18272 42030 18284
rect 42685 18275 42743 18281
rect 42685 18272 42697 18275
rect 42024 18244 42697 18272
rect 42024 18232 42030 18244
rect 42685 18241 42697 18244
rect 42731 18241 42743 18275
rect 42685 18235 42743 18241
rect 44542 18232 44548 18284
rect 44600 18272 44606 18284
rect 45097 18275 45155 18281
rect 45097 18272 45109 18275
rect 44600 18244 45109 18272
rect 44600 18232 44606 18244
rect 45097 18241 45109 18244
rect 45143 18241 45155 18275
rect 45097 18235 45155 18241
rect 47302 18232 47308 18284
rect 47360 18272 47366 18284
rect 47581 18275 47639 18281
rect 47581 18272 47593 18275
rect 47360 18244 47593 18272
rect 47360 18232 47366 18244
rect 47581 18241 47593 18244
rect 47627 18241 47639 18275
rect 47581 18235 47639 18241
rect 37829 18207 37887 18213
rect 37829 18173 37841 18207
rect 37875 18173 37887 18207
rect 38286 18204 38292 18216
rect 38247 18176 38292 18204
rect 37829 18167 37887 18173
rect 38286 18164 38292 18176
rect 38344 18164 38350 18216
rect 40126 18164 40132 18216
rect 40184 18204 40190 18216
rect 41230 18204 41236 18216
rect 40184 18176 41236 18204
rect 40184 18164 40190 18176
rect 41230 18164 41236 18176
rect 41288 18204 41294 18216
rect 42429 18207 42487 18213
rect 42429 18204 42441 18207
rect 41288 18176 42441 18204
rect 41288 18164 41294 18176
rect 42429 18173 42441 18176
rect 42475 18173 42487 18207
rect 42429 18167 42487 18173
rect 33502 18136 33508 18148
rect 27724 18108 33508 18136
rect 18874 18068 18880 18080
rect 16776 18040 18880 18068
rect 18874 18028 18880 18040
rect 18932 18028 18938 18080
rect 23124 18077 23152 18108
rect 23109 18071 23167 18077
rect 23109 18037 23121 18071
rect 23155 18037 23167 18071
rect 23109 18031 23167 18037
rect 23198 18028 23204 18080
rect 23256 18068 23262 18080
rect 23385 18071 23443 18077
rect 23385 18068 23397 18071
rect 23256 18040 23397 18068
rect 23256 18028 23262 18040
rect 23385 18037 23397 18040
rect 23431 18037 23443 18071
rect 23385 18031 23443 18037
rect 24029 18071 24087 18077
rect 24029 18037 24041 18071
rect 24075 18068 24087 18071
rect 24210 18068 24216 18080
rect 24075 18040 24216 18068
rect 24075 18037 24087 18040
rect 24029 18031 24087 18037
rect 24210 18028 24216 18040
rect 24268 18028 24274 18080
rect 25038 18068 25044 18080
rect 24999 18040 25044 18068
rect 25038 18028 25044 18040
rect 25096 18028 25102 18080
rect 25133 18071 25191 18077
rect 25133 18037 25145 18071
rect 25179 18068 25191 18071
rect 25498 18068 25504 18080
rect 25179 18040 25504 18068
rect 25179 18037 25191 18040
rect 25133 18031 25191 18037
rect 25498 18028 25504 18040
rect 25556 18028 25562 18080
rect 26602 18028 26608 18080
rect 26660 18068 26666 18080
rect 26878 18068 26884 18080
rect 26660 18040 26884 18068
rect 26660 18028 26666 18040
rect 26878 18028 26884 18040
rect 26936 18068 26942 18080
rect 27724 18068 27752 18108
rect 33502 18096 33508 18108
rect 33560 18096 33566 18148
rect 26936 18040 27752 18068
rect 26936 18028 26942 18040
rect 29270 18028 29276 18080
rect 29328 18068 29334 18080
rect 29822 18068 29828 18080
rect 29328 18040 29828 18068
rect 29328 18028 29334 18040
rect 29822 18028 29828 18040
rect 29880 18028 29886 18080
rect 30193 18071 30251 18077
rect 30193 18037 30205 18071
rect 30239 18068 30251 18071
rect 30282 18068 30288 18080
rect 30239 18040 30288 18068
rect 30239 18037 30251 18040
rect 30193 18031 30251 18037
rect 30282 18028 30288 18040
rect 30340 18028 30346 18080
rect 35342 18068 35348 18080
rect 35255 18040 35348 18068
rect 35342 18028 35348 18040
rect 35400 18068 35406 18080
rect 45738 18068 45744 18080
rect 35400 18040 45744 18068
rect 35400 18028 35406 18040
rect 45738 18028 45744 18040
rect 45796 18028 45802 18080
rect 47670 18068 47676 18080
rect 47631 18040 47676 18068
rect 47670 18028 47676 18040
rect 47728 18028 47734 18080
rect 1104 17978 48852 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 48852 17978
rect 1104 17904 48852 17926
rect 15378 17824 15384 17876
rect 15436 17864 15442 17876
rect 15841 17867 15899 17873
rect 15841 17864 15853 17867
rect 15436 17836 15853 17864
rect 15436 17824 15442 17836
rect 15841 17833 15853 17836
rect 15887 17833 15899 17867
rect 15841 17827 15899 17833
rect 16114 17824 16120 17876
rect 16172 17864 16178 17876
rect 23385 17867 23443 17873
rect 16172 17836 23336 17864
rect 16172 17824 16178 17836
rect 2866 17796 2872 17808
rect 1412 17768 2872 17796
rect 1412 17737 1440 17768
rect 2866 17756 2872 17768
rect 2924 17756 2930 17808
rect 19981 17799 20039 17805
rect 19981 17765 19993 17799
rect 20027 17796 20039 17799
rect 20806 17796 20812 17808
rect 20027 17768 20812 17796
rect 20027 17765 20039 17768
rect 19981 17759 20039 17765
rect 20806 17756 20812 17768
rect 20864 17756 20870 17808
rect 1397 17731 1455 17737
rect 1397 17697 1409 17731
rect 1443 17697 1455 17731
rect 1578 17728 1584 17740
rect 1539 17700 1584 17728
rect 1397 17691 1455 17697
rect 1578 17688 1584 17700
rect 1636 17688 1642 17740
rect 2774 17728 2780 17740
rect 2735 17700 2780 17728
rect 2774 17688 2780 17700
rect 2832 17688 2838 17740
rect 20625 17731 20683 17737
rect 20625 17697 20637 17731
rect 20671 17728 20683 17731
rect 20990 17728 20996 17740
rect 20671 17700 20996 17728
rect 20671 17697 20683 17700
rect 20625 17691 20683 17697
rect 20990 17688 20996 17700
rect 21048 17728 21054 17740
rect 22554 17728 22560 17740
rect 21048 17700 22560 17728
rect 21048 17688 21054 17700
rect 22554 17688 22560 17700
rect 22612 17688 22618 17740
rect 23308 17728 23336 17836
rect 23385 17833 23397 17867
rect 23431 17833 23443 17867
rect 23658 17864 23664 17876
rect 23619 17836 23664 17864
rect 23385 17827 23443 17833
rect 23400 17796 23428 17827
rect 23658 17824 23664 17836
rect 23716 17824 23722 17876
rect 25130 17824 25136 17876
rect 25188 17864 25194 17876
rect 25225 17867 25283 17873
rect 25225 17864 25237 17867
rect 25188 17836 25237 17864
rect 25188 17824 25194 17836
rect 25225 17833 25237 17836
rect 25271 17833 25283 17867
rect 25225 17827 25283 17833
rect 25685 17867 25743 17873
rect 25685 17833 25697 17867
rect 25731 17864 25743 17867
rect 26234 17864 26240 17876
rect 25731 17836 26240 17864
rect 25731 17833 25743 17836
rect 25685 17827 25743 17833
rect 26234 17824 26240 17836
rect 26292 17864 26298 17876
rect 28258 17864 28264 17876
rect 26292 17836 28264 17864
rect 26292 17824 26298 17836
rect 28258 17824 28264 17836
rect 28316 17824 28322 17876
rect 28905 17867 28963 17873
rect 28905 17833 28917 17867
rect 28951 17864 28963 17867
rect 29270 17864 29276 17876
rect 28951 17836 29276 17864
rect 28951 17833 28963 17836
rect 28905 17827 28963 17833
rect 29270 17824 29276 17836
rect 29328 17824 29334 17876
rect 29546 17824 29552 17876
rect 29604 17864 29610 17876
rect 31754 17864 31760 17876
rect 29604 17836 31760 17864
rect 29604 17824 29610 17836
rect 31754 17824 31760 17836
rect 31812 17824 31818 17876
rect 32858 17864 32864 17876
rect 32819 17836 32864 17864
rect 32858 17824 32864 17836
rect 32916 17824 32922 17876
rect 33594 17824 33600 17876
rect 33652 17864 33658 17876
rect 34149 17867 34207 17873
rect 34149 17864 34161 17867
rect 33652 17836 34161 17864
rect 33652 17824 33658 17836
rect 34149 17833 34161 17836
rect 34195 17833 34207 17867
rect 34149 17827 34207 17833
rect 37921 17867 37979 17873
rect 37921 17833 37933 17867
rect 37967 17864 37979 17867
rect 38010 17864 38016 17876
rect 37967 17836 38016 17864
rect 37967 17833 37979 17836
rect 37921 17827 37979 17833
rect 38010 17824 38016 17836
rect 38068 17824 38074 17876
rect 41966 17864 41972 17876
rect 41927 17836 41972 17864
rect 41966 17824 41972 17836
rect 42024 17824 42030 17876
rect 44818 17824 44824 17876
rect 44876 17864 44882 17876
rect 45005 17867 45063 17873
rect 45005 17864 45017 17867
rect 44876 17836 45017 17864
rect 44876 17824 44882 17836
rect 45005 17833 45017 17836
rect 45051 17833 45063 17867
rect 45005 17827 45063 17833
rect 23566 17796 23572 17808
rect 23400 17768 23572 17796
rect 23566 17756 23572 17768
rect 23624 17756 23630 17808
rect 23676 17768 25820 17796
rect 23676 17728 23704 17768
rect 23308 17700 23704 17728
rect 25792 17728 25820 17768
rect 26050 17756 26056 17808
rect 26108 17796 26114 17808
rect 27617 17799 27675 17805
rect 27617 17796 27629 17799
rect 26108 17768 27629 17796
rect 26108 17756 26114 17768
rect 27617 17765 27629 17768
rect 27663 17796 27675 17799
rect 29454 17796 29460 17808
rect 27663 17768 29460 17796
rect 27663 17765 27675 17768
rect 27617 17759 27675 17765
rect 29454 17756 29460 17768
rect 29512 17756 29518 17808
rect 39390 17756 39396 17808
rect 39448 17796 39454 17808
rect 45646 17796 45652 17808
rect 39448 17768 45652 17796
rect 39448 17756 39454 17768
rect 45646 17756 45652 17768
rect 45704 17756 45710 17808
rect 31389 17731 31447 17737
rect 25792 17700 29684 17728
rect 15749 17663 15807 17669
rect 15749 17629 15761 17663
rect 15795 17660 15807 17663
rect 15838 17660 15844 17672
rect 15795 17632 15844 17660
rect 15795 17629 15807 17632
rect 15749 17623 15807 17629
rect 15838 17620 15844 17632
rect 15896 17620 15902 17672
rect 20346 17620 20352 17672
rect 20404 17620 20410 17672
rect 23198 17660 23204 17672
rect 22480 17632 23060 17660
rect 23159 17632 23204 17660
rect 16574 17552 16580 17604
rect 16632 17592 16638 17604
rect 17497 17595 17555 17601
rect 17497 17592 17509 17595
rect 16632 17564 17509 17592
rect 16632 17552 16638 17564
rect 17497 17561 17509 17564
rect 17543 17561 17555 17595
rect 17497 17555 17555 17561
rect 17865 17595 17923 17601
rect 17865 17561 17877 17595
rect 17911 17592 17923 17595
rect 17954 17592 17960 17604
rect 17911 17564 17960 17592
rect 17911 17561 17923 17564
rect 17865 17555 17923 17561
rect 17954 17552 17960 17564
rect 18012 17552 18018 17604
rect 20364 17592 20392 17620
rect 20622 17592 20628 17604
rect 20364 17564 20628 17592
rect 20622 17552 20628 17564
rect 20680 17552 20686 17604
rect 22480 17592 22508 17632
rect 22066 17564 22508 17592
rect 20346 17524 20352 17536
rect 20307 17496 20352 17524
rect 20346 17484 20352 17496
rect 20404 17484 20410 17536
rect 20441 17527 20499 17533
rect 20441 17493 20453 17527
rect 20487 17524 20499 17527
rect 22066 17524 22094 17564
rect 22554 17552 22560 17604
rect 22612 17592 22618 17604
rect 22741 17595 22799 17601
rect 22612 17564 22657 17592
rect 22612 17552 22618 17564
rect 22741 17561 22753 17595
rect 22787 17592 22799 17595
rect 22830 17592 22836 17604
rect 22787 17564 22836 17592
rect 22787 17561 22799 17564
rect 22741 17555 22799 17561
rect 22830 17552 22836 17564
rect 22888 17552 22894 17604
rect 23032 17592 23060 17632
rect 23198 17620 23204 17632
rect 23256 17620 23262 17672
rect 23290 17620 23296 17672
rect 23348 17660 23354 17672
rect 23385 17663 23443 17669
rect 23385 17660 23397 17663
rect 23348 17632 23397 17660
rect 23348 17620 23354 17632
rect 23385 17629 23397 17632
rect 23431 17629 23443 17663
rect 23385 17623 23443 17629
rect 23477 17663 23535 17669
rect 23477 17629 23489 17663
rect 23523 17660 23535 17663
rect 24210 17660 24216 17672
rect 23523 17632 24216 17660
rect 23523 17629 23535 17632
rect 23477 17623 23535 17629
rect 24210 17620 24216 17632
rect 24268 17620 24274 17672
rect 25406 17660 25412 17672
rect 25367 17632 25412 17660
rect 25406 17620 25412 17632
rect 25464 17620 25470 17672
rect 25498 17620 25504 17672
rect 25556 17660 25562 17672
rect 25777 17663 25835 17669
rect 25556 17632 25601 17660
rect 25556 17620 25562 17632
rect 25777 17629 25789 17663
rect 25823 17629 25835 17663
rect 25777 17623 25835 17629
rect 25682 17592 25688 17604
rect 23032 17564 25688 17592
rect 25682 17552 25688 17564
rect 25740 17552 25746 17604
rect 25792 17592 25820 17623
rect 25958 17620 25964 17672
rect 26016 17660 26022 17672
rect 26329 17663 26387 17669
rect 26329 17660 26341 17663
rect 26016 17632 26341 17660
rect 26016 17620 26022 17632
rect 26329 17629 26341 17632
rect 26375 17629 26387 17663
rect 26329 17623 26387 17629
rect 27433 17663 27491 17669
rect 27433 17629 27445 17663
rect 27479 17660 27491 17663
rect 27890 17660 27896 17672
rect 27479 17632 27896 17660
rect 27479 17629 27491 17632
rect 27433 17623 27491 17629
rect 27890 17620 27896 17632
rect 27948 17620 27954 17672
rect 28350 17620 28356 17672
rect 28408 17660 28414 17672
rect 28721 17663 28779 17669
rect 28721 17660 28733 17663
rect 28408 17632 28733 17660
rect 28408 17620 28414 17632
rect 28721 17629 28733 17632
rect 28767 17629 28779 17663
rect 29546 17660 29552 17672
rect 29507 17632 29552 17660
rect 28721 17623 28779 17629
rect 29546 17620 29552 17632
rect 29604 17620 29610 17672
rect 29656 17660 29684 17700
rect 31389 17697 31401 17731
rect 31435 17728 31447 17731
rect 32030 17728 32036 17740
rect 31435 17700 32036 17728
rect 31435 17697 31447 17700
rect 31389 17691 31447 17697
rect 32030 17688 32036 17700
rect 32088 17688 32094 17740
rect 38286 17728 38292 17740
rect 38120 17700 38292 17728
rect 31665 17663 31723 17669
rect 29656 17632 31064 17660
rect 26418 17592 26424 17604
rect 25792 17564 26424 17592
rect 26418 17552 26424 17564
rect 26476 17552 26482 17604
rect 26513 17595 26571 17601
rect 26513 17561 26525 17595
rect 26559 17592 26571 17595
rect 28368 17592 28396 17620
rect 29822 17601 29828 17604
rect 26559 17564 28396 17592
rect 26559 17561 26571 17564
rect 26513 17555 26571 17561
rect 29816 17555 29828 17601
rect 29880 17592 29886 17604
rect 29880 17564 29916 17592
rect 20487 17496 22094 17524
rect 20487 17493 20499 17496
rect 20441 17487 20499 17493
rect 22922 17484 22928 17536
rect 22980 17524 22986 17536
rect 23290 17524 23296 17536
rect 22980 17496 23296 17524
rect 22980 17484 22986 17496
rect 23290 17484 23296 17496
rect 23348 17484 23354 17536
rect 25774 17484 25780 17536
rect 25832 17524 25838 17536
rect 26528 17524 26556 17555
rect 29822 17552 29828 17555
rect 29880 17552 29886 17564
rect 25832 17496 26556 17524
rect 25832 17484 25838 17496
rect 29362 17484 29368 17536
rect 29420 17524 29426 17536
rect 30929 17527 30987 17533
rect 30929 17524 30941 17527
rect 29420 17496 30941 17524
rect 29420 17484 29426 17496
rect 30929 17493 30941 17496
rect 30975 17493 30987 17527
rect 31036 17524 31064 17632
rect 31665 17629 31677 17663
rect 31711 17660 31723 17663
rect 32769 17663 32827 17669
rect 31711 17632 31745 17660
rect 31711 17629 31723 17632
rect 31665 17623 31723 17629
rect 32769 17629 32781 17663
rect 32815 17660 32827 17663
rect 34146 17660 34152 17672
rect 32815 17632 34152 17660
rect 32815 17629 32827 17632
rect 32769 17623 32827 17629
rect 31478 17552 31484 17604
rect 31536 17592 31542 17604
rect 31680 17592 31708 17623
rect 34146 17620 34152 17632
rect 34204 17620 34210 17672
rect 37918 17660 37924 17672
rect 37879 17632 37924 17660
rect 37918 17620 37924 17632
rect 37976 17620 37982 17672
rect 38120 17669 38148 17700
rect 38286 17688 38292 17700
rect 38344 17728 38350 17740
rect 39945 17731 40003 17737
rect 39945 17728 39957 17731
rect 38344 17700 39957 17728
rect 38344 17688 38350 17700
rect 39945 17697 39957 17700
rect 39991 17728 40003 17731
rect 40770 17728 40776 17740
rect 39991 17700 40776 17728
rect 39991 17697 40003 17700
rect 39945 17691 40003 17697
rect 40770 17688 40776 17700
rect 40828 17688 40834 17740
rect 40880 17700 41460 17728
rect 38105 17663 38163 17669
rect 38105 17629 38117 17663
rect 38151 17629 38163 17663
rect 38105 17623 38163 17629
rect 40034 17620 40040 17672
rect 40092 17660 40098 17672
rect 40221 17663 40279 17669
rect 40221 17660 40233 17663
rect 40092 17632 40233 17660
rect 40092 17620 40098 17632
rect 40221 17629 40233 17632
rect 40267 17660 40279 17663
rect 40402 17660 40408 17672
rect 40267 17632 40408 17660
rect 40267 17629 40279 17632
rect 40221 17623 40279 17629
rect 40402 17620 40408 17632
rect 40460 17660 40466 17672
rect 40880 17660 40908 17700
rect 40460 17632 40908 17660
rect 40460 17620 40466 17632
rect 41046 17620 41052 17672
rect 41104 17660 41110 17672
rect 41432 17669 41460 17700
rect 44450 17688 44456 17740
rect 44508 17728 44514 17740
rect 44508 17700 45508 17728
rect 44508 17688 44514 17700
rect 41233 17663 41291 17669
rect 41233 17660 41245 17663
rect 41104 17632 41245 17660
rect 41104 17620 41110 17632
rect 41233 17629 41245 17632
rect 41279 17629 41291 17663
rect 41233 17623 41291 17629
rect 41417 17663 41475 17669
rect 41417 17629 41429 17663
rect 41463 17629 41475 17663
rect 42150 17660 42156 17672
rect 42111 17632 42156 17660
rect 41417 17623 41475 17629
rect 42150 17620 42156 17632
rect 42208 17620 42214 17672
rect 43254 17660 43260 17672
rect 43215 17632 43260 17660
rect 43254 17620 43260 17632
rect 43312 17620 43318 17672
rect 45480 17669 45508 17700
rect 45664 17669 45692 17756
rect 46290 17728 46296 17740
rect 46251 17700 46296 17728
rect 46290 17688 46296 17700
rect 46348 17688 46354 17740
rect 46477 17731 46535 17737
rect 46477 17697 46489 17731
rect 46523 17728 46535 17731
rect 47670 17728 47676 17740
rect 46523 17700 47676 17728
rect 46523 17697 46535 17700
rect 46477 17691 46535 17697
rect 47670 17688 47676 17700
rect 47728 17688 47734 17740
rect 48130 17728 48136 17740
rect 48091 17700 48136 17728
rect 48130 17688 48136 17700
rect 48188 17688 48194 17740
rect 45235 17663 45293 17669
rect 45235 17629 45247 17663
rect 45281 17629 45293 17663
rect 45235 17623 45293 17629
rect 45373 17663 45431 17669
rect 45373 17629 45385 17663
rect 45419 17629 45431 17663
rect 45373 17623 45431 17629
rect 45470 17663 45528 17669
rect 45470 17629 45482 17663
rect 45516 17629 45528 17663
rect 45470 17623 45528 17629
rect 45649 17663 45707 17669
rect 45649 17629 45661 17663
rect 45695 17629 45707 17663
rect 45649 17623 45707 17629
rect 32122 17592 32128 17604
rect 31536 17564 32128 17592
rect 31536 17552 31542 17564
rect 32122 17552 32128 17564
rect 32180 17592 32186 17604
rect 33781 17595 33839 17601
rect 33781 17592 33793 17595
rect 32180 17564 33793 17592
rect 32180 17552 32186 17564
rect 33781 17561 33793 17564
rect 33827 17592 33839 17595
rect 33870 17592 33876 17604
rect 33827 17564 33876 17592
rect 33827 17561 33839 17564
rect 33781 17555 33839 17561
rect 33870 17552 33876 17564
rect 33928 17552 33934 17604
rect 33965 17595 34023 17601
rect 33965 17561 33977 17595
rect 34011 17592 34023 17595
rect 35342 17592 35348 17604
rect 34011 17564 35348 17592
rect 34011 17561 34023 17564
rect 33965 17555 34023 17561
rect 35342 17552 35348 17564
rect 35400 17552 35406 17604
rect 37642 17524 37648 17536
rect 31036 17496 37648 17524
rect 30929 17487 30987 17493
rect 37642 17484 37648 17496
rect 37700 17484 37706 17536
rect 41417 17527 41475 17533
rect 41417 17493 41429 17527
rect 41463 17524 41475 17527
rect 41598 17524 41604 17536
rect 41463 17496 41604 17524
rect 41463 17493 41475 17496
rect 41417 17487 41475 17493
rect 41598 17484 41604 17496
rect 41656 17484 41662 17536
rect 41874 17484 41880 17536
rect 41932 17524 41938 17536
rect 43073 17527 43131 17533
rect 43073 17524 43085 17527
rect 41932 17496 43085 17524
rect 41932 17484 41938 17496
rect 43073 17493 43085 17496
rect 43119 17524 43131 17527
rect 45250 17524 45278 17623
rect 45388 17536 45416 17623
rect 43119 17496 45278 17524
rect 43119 17493 43131 17496
rect 43073 17487 43131 17493
rect 45370 17484 45376 17536
rect 45428 17484 45434 17536
rect 1104 17434 48852 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 48852 17434
rect 1104 17360 48852 17382
rect 19058 17320 19064 17332
rect 6886 17292 19064 17320
rect 2041 17255 2099 17261
rect 2041 17221 2053 17255
rect 2087 17252 2099 17255
rect 6886 17252 6914 17292
rect 19058 17280 19064 17292
rect 19116 17280 19122 17332
rect 21726 17280 21732 17332
rect 21784 17320 21790 17332
rect 22278 17320 22284 17332
rect 21784 17292 22284 17320
rect 21784 17280 21790 17292
rect 22278 17280 22284 17292
rect 22336 17320 22342 17332
rect 23017 17323 23075 17329
rect 23017 17320 23029 17323
rect 22336 17292 23029 17320
rect 22336 17280 22342 17292
rect 23017 17289 23029 17292
rect 23063 17289 23075 17323
rect 23017 17283 23075 17289
rect 24486 17280 24492 17332
rect 24544 17320 24550 17332
rect 29362 17320 29368 17332
rect 24544 17292 29368 17320
rect 24544 17280 24550 17292
rect 29362 17280 29368 17292
rect 29420 17280 29426 17332
rect 29822 17320 29828 17332
rect 29783 17292 29828 17320
rect 29822 17280 29828 17292
rect 29880 17280 29886 17332
rect 35986 17320 35992 17332
rect 35947 17292 35992 17320
rect 35986 17280 35992 17292
rect 36044 17280 36050 17332
rect 40957 17323 41015 17329
rect 40957 17289 40969 17323
rect 41003 17320 41015 17323
rect 41617 17323 41675 17329
rect 41617 17320 41629 17323
rect 41003 17292 41629 17320
rect 41003 17289 41015 17292
rect 40957 17283 41015 17289
rect 41617 17289 41629 17292
rect 41663 17289 41675 17323
rect 45830 17320 45836 17332
rect 41617 17283 41675 17289
rect 43548 17292 45836 17320
rect 2087 17224 6914 17252
rect 16025 17255 16083 17261
rect 2087 17221 2099 17224
rect 2041 17215 2099 17221
rect 16025 17221 16037 17255
rect 16071 17252 16083 17255
rect 16853 17255 16911 17261
rect 16853 17252 16865 17255
rect 16071 17224 16865 17252
rect 16071 17221 16083 17224
rect 16025 17215 16083 17221
rect 16853 17221 16865 17224
rect 16899 17221 16911 17255
rect 16853 17215 16911 17221
rect 19978 17212 19984 17264
rect 20036 17252 20042 17264
rect 20254 17252 20260 17264
rect 20036 17224 20260 17252
rect 20036 17212 20042 17224
rect 20254 17212 20260 17224
rect 20312 17212 20318 17264
rect 22370 17212 22376 17264
rect 22428 17252 22434 17264
rect 23937 17255 23995 17261
rect 23937 17252 23949 17255
rect 22428 17224 23949 17252
rect 22428 17212 22434 17224
rect 23937 17221 23949 17224
rect 23983 17252 23995 17255
rect 24670 17252 24676 17264
rect 23983 17224 24676 17252
rect 23983 17221 23995 17224
rect 23937 17215 23995 17221
rect 24670 17212 24676 17224
rect 24728 17212 24734 17264
rect 26234 17252 26240 17264
rect 25240 17224 25912 17252
rect 26195 17224 26240 17252
rect 1854 17184 1860 17196
rect 1815 17156 1860 17184
rect 1854 17144 1860 17156
rect 1912 17144 1918 17196
rect 15930 17184 15936 17196
rect 15891 17156 15936 17184
rect 15930 17144 15936 17156
rect 15988 17144 15994 17196
rect 16666 17184 16672 17196
rect 16627 17156 16672 17184
rect 16666 17144 16672 17156
rect 16724 17144 16730 17196
rect 19236 17187 19294 17193
rect 19236 17153 19248 17187
rect 19282 17184 19294 17187
rect 20622 17184 20628 17196
rect 19282 17156 20628 17184
rect 19282 17153 19294 17156
rect 19236 17147 19294 17153
rect 20622 17144 20628 17156
rect 20680 17144 20686 17196
rect 22922 17184 22928 17196
rect 22883 17156 22928 17184
rect 22922 17144 22928 17156
rect 22980 17144 22986 17196
rect 23753 17187 23811 17193
rect 23753 17153 23765 17187
rect 23799 17184 23811 17187
rect 23842 17184 23848 17196
rect 23799 17156 23848 17184
rect 23799 17153 23811 17156
rect 23753 17147 23811 17153
rect 23842 17144 23848 17156
rect 23900 17184 23906 17196
rect 24302 17184 24308 17196
rect 23900 17156 24308 17184
rect 23900 17144 23906 17156
rect 24302 17144 24308 17156
rect 24360 17184 24366 17196
rect 25240 17184 25268 17224
rect 24360 17156 25268 17184
rect 24360 17144 24366 17156
rect 25406 17144 25412 17196
rect 25464 17184 25470 17196
rect 25501 17187 25559 17193
rect 25501 17184 25513 17187
rect 25464 17156 25513 17184
rect 25464 17144 25470 17156
rect 25501 17153 25513 17156
rect 25547 17153 25559 17187
rect 25501 17147 25559 17153
rect 25685 17187 25743 17193
rect 25685 17153 25697 17187
rect 25731 17184 25743 17187
rect 25774 17184 25780 17196
rect 25731 17156 25780 17184
rect 25731 17153 25743 17156
rect 25685 17147 25743 17153
rect 25774 17144 25780 17156
rect 25832 17144 25838 17196
rect 25884 17184 25912 17224
rect 26234 17212 26240 17224
rect 26292 17212 26298 17264
rect 26786 17212 26792 17264
rect 26844 17252 26850 17264
rect 29270 17252 29276 17264
rect 26844 17224 29276 17252
rect 26844 17212 26850 17224
rect 29270 17212 29276 17224
rect 29328 17212 29334 17264
rect 30834 17252 30840 17264
rect 30024 17224 30840 17252
rect 27709 17187 27767 17193
rect 25884 17156 27016 17184
rect 18322 17116 18328 17128
rect 18283 17088 18328 17116
rect 18322 17076 18328 17088
rect 18380 17076 18386 17128
rect 18969 17119 19027 17125
rect 18969 17085 18981 17119
rect 19015 17085 19027 17119
rect 26418 17116 26424 17128
rect 18969 17079 19027 17085
rect 21974 17088 26424 17116
rect 2130 16940 2136 16992
rect 2188 16980 2194 16992
rect 2685 16983 2743 16989
rect 2685 16980 2697 16983
rect 2188 16952 2697 16980
rect 2188 16940 2194 16952
rect 2685 16949 2697 16952
rect 2731 16949 2743 16983
rect 18984 16980 19012 17079
rect 21974 17048 22002 17088
rect 26418 17076 26424 17088
rect 26476 17076 26482 17128
rect 26878 17048 26884 17060
rect 20824 17020 22002 17048
rect 22066 17020 26884 17048
rect 19334 16980 19340 16992
rect 18984 16952 19340 16980
rect 2685 16943 2743 16949
rect 19334 16940 19340 16952
rect 19392 16980 19398 16992
rect 20254 16980 20260 16992
rect 19392 16952 20260 16980
rect 19392 16940 19398 16952
rect 20254 16940 20260 16952
rect 20312 16940 20318 16992
rect 20346 16940 20352 16992
rect 20404 16980 20410 16992
rect 20824 16980 20852 17020
rect 20404 16952 20852 16980
rect 20404 16940 20410 16952
rect 20898 16940 20904 16992
rect 20956 16980 20962 16992
rect 22066 16980 22094 17020
rect 26878 17008 26884 17020
rect 26936 17008 26942 17060
rect 26988 17048 27016 17156
rect 27709 17153 27721 17187
rect 27755 17184 27767 17187
rect 27890 17184 27896 17196
rect 27755 17156 27896 17184
rect 27755 17153 27767 17156
rect 27709 17147 27767 17153
rect 27890 17144 27896 17156
rect 27948 17144 27954 17196
rect 30024 17193 30052 17224
rect 30834 17212 30840 17224
rect 30892 17212 30898 17264
rect 31113 17255 31171 17261
rect 31113 17221 31125 17255
rect 31159 17252 31171 17255
rect 31846 17252 31852 17264
rect 31159 17224 31852 17252
rect 31159 17221 31171 17224
rect 31113 17215 31171 17221
rect 31846 17212 31852 17224
rect 31904 17252 31910 17264
rect 33042 17252 33048 17264
rect 31904 17224 33048 17252
rect 31904 17212 31910 17224
rect 33042 17212 33048 17224
rect 33100 17212 33106 17264
rect 33870 17252 33876 17264
rect 33831 17224 33876 17252
rect 33870 17212 33876 17224
rect 33928 17212 33934 17264
rect 34057 17255 34115 17261
rect 34057 17221 34069 17255
rect 34103 17252 34115 17255
rect 35526 17252 35532 17264
rect 34103 17224 35532 17252
rect 34103 17221 34115 17224
rect 34057 17215 34115 17221
rect 35526 17212 35532 17224
rect 35584 17212 35590 17264
rect 39853 17255 39911 17261
rect 39853 17221 39865 17255
rect 39899 17252 39911 17255
rect 40589 17255 40647 17261
rect 40589 17252 40601 17255
rect 39899 17224 40601 17252
rect 39899 17221 39911 17224
rect 39853 17215 39911 17221
rect 40589 17221 40601 17224
rect 40635 17252 40647 17255
rect 41046 17252 41052 17264
rect 40635 17224 41052 17252
rect 40635 17221 40647 17224
rect 40589 17215 40647 17221
rect 41046 17212 41052 17224
rect 41104 17212 41110 17264
rect 41417 17255 41475 17261
rect 41417 17221 41429 17255
rect 41463 17252 41475 17255
rect 41782 17252 41788 17264
rect 41463 17224 41788 17252
rect 41463 17221 41475 17224
rect 41417 17215 41475 17221
rect 41782 17212 41788 17224
rect 41840 17252 41846 17264
rect 41966 17252 41972 17264
rect 41840 17224 41972 17252
rect 41840 17212 41846 17224
rect 41966 17212 41972 17224
rect 42024 17212 42030 17264
rect 30009 17187 30067 17193
rect 30009 17153 30021 17187
rect 30055 17153 30067 17187
rect 30009 17147 30067 17153
rect 30101 17187 30159 17193
rect 30101 17153 30113 17187
rect 30147 17153 30159 17187
rect 30282 17184 30288 17196
rect 30243 17156 30288 17184
rect 30101 17147 30159 17153
rect 29914 17076 29920 17128
rect 29972 17116 29978 17128
rect 30116 17116 30144 17147
rect 30282 17144 30288 17156
rect 30340 17144 30346 17196
rect 30377 17187 30435 17193
rect 30377 17153 30389 17187
rect 30423 17153 30435 17187
rect 30929 17187 30987 17193
rect 30929 17184 30941 17187
rect 30377 17147 30435 17153
rect 30852 17156 30941 17184
rect 29972 17088 30144 17116
rect 29972 17076 29978 17088
rect 28534 17048 28540 17060
rect 26988 17020 28540 17048
rect 20956 16952 22094 16980
rect 20956 16940 20962 16952
rect 22554 16940 22560 16992
rect 22612 16980 22618 16992
rect 23658 16980 23664 16992
rect 22612 16952 23664 16980
rect 22612 16940 22618 16952
rect 23658 16940 23664 16952
rect 23716 16940 23722 16992
rect 25590 16980 25596 16992
rect 25551 16952 25596 16980
rect 25590 16940 25596 16952
rect 25648 16940 25654 16992
rect 26329 16983 26387 16989
rect 26329 16949 26341 16983
rect 26375 16980 26387 16983
rect 26988 16980 27016 17020
rect 28534 17008 28540 17020
rect 28592 17008 28598 17060
rect 28626 17008 28632 17060
rect 28684 17048 28690 17060
rect 30392 17048 30420 17147
rect 30852 17128 30880 17156
rect 30929 17153 30941 17156
rect 30975 17184 30987 17187
rect 31294 17184 31300 17196
rect 30975 17156 31300 17184
rect 30975 17153 30987 17156
rect 30929 17147 30987 17153
rect 31294 17144 31300 17156
rect 31352 17144 31358 17196
rect 34146 17144 34152 17196
rect 34204 17184 34210 17196
rect 35897 17187 35955 17193
rect 35897 17184 35909 17187
rect 34204 17156 35909 17184
rect 34204 17144 34210 17156
rect 35897 17153 35909 17156
rect 35943 17153 35955 17187
rect 35897 17147 35955 17153
rect 36170 17144 36176 17196
rect 36228 17184 36234 17196
rect 37737 17187 37795 17193
rect 37737 17184 37749 17187
rect 36228 17156 37749 17184
rect 36228 17144 36234 17156
rect 37737 17153 37749 17156
rect 37783 17153 37795 17187
rect 40034 17184 40040 17196
rect 39995 17156 40040 17184
rect 37737 17147 37795 17153
rect 40034 17144 40040 17156
rect 40092 17144 40098 17196
rect 40129 17187 40187 17193
rect 40129 17153 40141 17187
rect 40175 17184 40187 17187
rect 40494 17184 40500 17196
rect 40175 17156 40500 17184
rect 40175 17153 40187 17156
rect 40129 17147 40187 17153
rect 40494 17144 40500 17156
rect 40552 17144 40558 17196
rect 40770 17184 40776 17196
rect 40731 17156 40776 17184
rect 40770 17144 40776 17156
rect 40828 17144 40834 17196
rect 30834 17076 30840 17128
rect 30892 17076 30898 17128
rect 37642 17076 37648 17128
rect 37700 17116 37706 17128
rect 43548 17116 43576 17292
rect 45830 17280 45836 17292
rect 45888 17280 45894 17332
rect 45373 17255 45431 17261
rect 45373 17221 45385 17255
rect 45419 17252 45431 17255
rect 47673 17255 47731 17261
rect 47673 17252 47685 17255
rect 45419 17224 47685 17252
rect 45419 17221 45431 17224
rect 45373 17215 45431 17221
rect 47673 17221 47685 17224
rect 47719 17221 47731 17255
rect 47673 17215 47731 17221
rect 47578 17184 47584 17196
rect 47539 17156 47584 17184
rect 47578 17144 47584 17156
rect 47636 17144 47642 17196
rect 37700 17088 43576 17116
rect 45189 17119 45247 17125
rect 37700 17076 37706 17088
rect 45189 17085 45201 17119
rect 45235 17116 45247 17119
rect 45830 17116 45836 17128
rect 45235 17088 45836 17116
rect 45235 17085 45247 17088
rect 45189 17079 45247 17085
rect 45830 17076 45836 17088
rect 45888 17076 45894 17128
rect 46842 17116 46848 17128
rect 46803 17088 46848 17116
rect 46842 17076 46848 17088
rect 46900 17076 46906 17128
rect 28684 17020 30420 17048
rect 37921 17051 37979 17057
rect 28684 17008 28690 17020
rect 37921 17017 37933 17051
rect 37967 17048 37979 17051
rect 39390 17048 39396 17060
rect 37967 17020 39396 17048
rect 37967 17017 37979 17020
rect 37921 17011 37979 17017
rect 39390 17008 39396 17020
rect 39448 17008 39454 17060
rect 40129 17051 40187 17057
rect 40129 17017 40141 17051
rect 40175 17048 40187 17051
rect 40175 17020 41092 17048
rect 40175 17017 40187 17020
rect 40129 17011 40187 17017
rect 27982 16980 27988 16992
rect 26375 16952 27016 16980
rect 27895 16952 27988 16980
rect 26375 16949 26387 16952
rect 26329 16943 26387 16949
rect 27982 16940 27988 16952
rect 28040 16980 28046 16992
rect 29730 16980 29736 16992
rect 28040 16952 29736 16980
rect 28040 16940 28046 16952
rect 29730 16940 29736 16952
rect 29788 16940 29794 16992
rect 33870 16940 33876 16992
rect 33928 16980 33934 16992
rect 34241 16983 34299 16989
rect 34241 16980 34253 16983
rect 33928 16952 34253 16980
rect 33928 16940 33934 16952
rect 34241 16949 34253 16952
rect 34287 16949 34299 16983
rect 41064 16980 41092 17020
rect 41414 16980 41420 16992
rect 41064 16952 41420 16980
rect 34241 16943 34299 16949
rect 41414 16940 41420 16952
rect 41472 16940 41478 16992
rect 41598 16980 41604 16992
rect 41559 16952 41604 16980
rect 41598 16940 41604 16952
rect 41656 16940 41662 16992
rect 41782 16980 41788 16992
rect 41743 16952 41788 16980
rect 41782 16940 41788 16952
rect 41840 16940 41846 16992
rect 1104 16890 48852 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 48852 16890
rect 1104 16816 48852 16838
rect 16666 16776 16672 16788
rect 6886 16748 16672 16776
rect 1854 16668 1860 16720
rect 1912 16708 1918 16720
rect 1912 16680 2268 16708
rect 1912 16668 1918 16680
rect 1397 16643 1455 16649
rect 1397 16609 1409 16643
rect 1443 16640 1455 16643
rect 2130 16640 2136 16652
rect 1443 16612 2136 16640
rect 1443 16609 1455 16612
rect 1397 16603 1455 16609
rect 2130 16600 2136 16612
rect 2188 16600 2194 16652
rect 2240 16649 2268 16680
rect 2225 16643 2283 16649
rect 2225 16609 2237 16643
rect 2271 16609 2283 16643
rect 2225 16603 2283 16609
rect 3326 16600 3332 16652
rect 3384 16640 3390 16652
rect 6886 16640 6914 16748
rect 16666 16736 16672 16748
rect 16724 16776 16730 16788
rect 17865 16779 17923 16785
rect 17865 16776 17877 16779
rect 16724 16748 17877 16776
rect 16724 16736 16730 16748
rect 17865 16745 17877 16748
rect 17911 16776 17923 16779
rect 20898 16776 20904 16788
rect 17911 16748 20904 16776
rect 17911 16745 17923 16748
rect 17865 16739 17923 16745
rect 20898 16736 20904 16748
rect 20956 16736 20962 16788
rect 23109 16779 23167 16785
rect 23109 16745 23121 16779
rect 23155 16776 23167 16779
rect 23198 16776 23204 16788
rect 23155 16748 23204 16776
rect 23155 16745 23167 16748
rect 23109 16739 23167 16745
rect 23198 16736 23204 16748
rect 23256 16736 23262 16788
rect 23382 16736 23388 16788
rect 23440 16776 23446 16788
rect 25133 16779 25191 16785
rect 25133 16776 25145 16779
rect 23440 16748 25145 16776
rect 23440 16736 23446 16748
rect 25133 16745 25145 16748
rect 25179 16776 25191 16779
rect 26145 16779 26203 16785
rect 25179 16748 26096 16776
rect 25179 16745 25191 16748
rect 25133 16739 25191 16745
rect 23293 16711 23351 16717
rect 23293 16677 23305 16711
rect 23339 16708 23351 16711
rect 23566 16708 23572 16720
rect 23339 16680 23572 16708
rect 23339 16677 23351 16680
rect 23293 16671 23351 16677
rect 23566 16668 23572 16680
rect 23624 16668 23630 16720
rect 25958 16708 25964 16720
rect 25516 16680 25964 16708
rect 3384 16612 6914 16640
rect 3384 16600 3390 16612
rect 17954 16600 17960 16652
rect 18012 16640 18018 16652
rect 20254 16640 20260 16652
rect 18012 16612 19288 16640
rect 20215 16612 20260 16640
rect 18012 16600 18018 16612
rect 19260 16584 19288 16612
rect 20254 16600 20260 16612
rect 20312 16600 20318 16652
rect 23201 16643 23259 16649
rect 23201 16609 23213 16643
rect 23247 16640 23259 16643
rect 23382 16640 23388 16652
rect 23247 16612 23388 16640
rect 23247 16609 23259 16612
rect 23201 16603 23259 16609
rect 23382 16600 23388 16612
rect 23440 16600 23446 16652
rect 23750 16640 23756 16652
rect 23492 16612 23756 16640
rect 15194 16532 15200 16584
rect 15252 16572 15258 16584
rect 15378 16572 15384 16584
rect 15252 16544 15384 16572
rect 15252 16532 15258 16544
rect 15378 16532 15384 16544
rect 15436 16572 15442 16584
rect 15933 16575 15991 16581
rect 15933 16572 15945 16575
rect 15436 16544 15945 16572
rect 15436 16532 15442 16544
rect 15933 16541 15945 16544
rect 15979 16572 15991 16575
rect 19242 16572 19248 16584
rect 15979 16544 19104 16572
rect 19203 16544 19248 16572
rect 15979 16541 15991 16544
rect 15933 16535 15991 16541
rect 19076 16516 19104 16544
rect 19242 16532 19248 16544
rect 19300 16532 19306 16584
rect 22097 16575 22155 16581
rect 22097 16541 22109 16575
rect 22143 16572 22155 16575
rect 22186 16572 22192 16584
rect 22143 16544 22192 16572
rect 22143 16541 22155 16544
rect 22097 16535 22155 16541
rect 22186 16532 22192 16544
rect 22244 16532 22250 16584
rect 22281 16575 22339 16581
rect 22281 16541 22293 16575
rect 22327 16572 22339 16575
rect 23014 16572 23020 16584
rect 22327 16544 23020 16572
rect 22327 16541 22339 16544
rect 22281 16535 22339 16541
rect 23014 16532 23020 16544
rect 23072 16532 23078 16584
rect 23492 16581 23520 16612
rect 23750 16600 23756 16612
rect 23808 16600 23814 16652
rect 24946 16600 24952 16652
rect 25004 16640 25010 16652
rect 25004 16612 25084 16640
rect 25004 16600 25010 16612
rect 25056 16581 25084 16612
rect 23477 16575 23535 16581
rect 23477 16541 23489 16575
rect 23523 16541 23535 16575
rect 23477 16535 23535 16541
rect 25041 16575 25099 16581
rect 25041 16541 25053 16575
rect 25087 16572 25099 16575
rect 25516 16572 25544 16680
rect 25958 16668 25964 16680
rect 26016 16668 26022 16720
rect 25590 16600 25596 16652
rect 25648 16640 25654 16652
rect 26068 16640 26096 16748
rect 26145 16745 26157 16779
rect 26191 16776 26203 16779
rect 26234 16776 26240 16788
rect 26191 16748 26240 16776
rect 26191 16745 26203 16748
rect 26145 16739 26203 16745
rect 26234 16736 26240 16748
rect 26292 16736 26298 16788
rect 26878 16736 26884 16788
rect 26936 16776 26942 16788
rect 42150 16776 42156 16788
rect 26936 16748 41414 16776
rect 42111 16748 42156 16776
rect 26936 16736 26942 16748
rect 26973 16711 27031 16717
rect 26973 16677 26985 16711
rect 27019 16708 27031 16711
rect 27338 16708 27344 16720
rect 27019 16680 27344 16708
rect 27019 16677 27031 16680
rect 26973 16671 27031 16677
rect 27338 16668 27344 16680
rect 27396 16668 27402 16720
rect 27614 16668 27620 16720
rect 27672 16708 27678 16720
rect 27890 16708 27896 16720
rect 27672 16680 27896 16708
rect 27672 16668 27678 16680
rect 27890 16668 27896 16680
rect 27948 16668 27954 16720
rect 29178 16668 29184 16720
rect 29236 16708 29242 16720
rect 30926 16708 30932 16720
rect 29236 16680 30932 16708
rect 29236 16668 29242 16680
rect 30926 16668 30932 16680
rect 30984 16668 30990 16720
rect 33226 16668 33232 16720
rect 33284 16708 33290 16720
rect 34054 16708 34060 16720
rect 33284 16680 34060 16708
rect 33284 16668 33290 16680
rect 34054 16668 34060 16680
rect 34112 16668 34118 16720
rect 37642 16708 37648 16720
rect 37603 16680 37648 16708
rect 37642 16668 37648 16680
rect 37700 16668 37706 16720
rect 41386 16708 41414 16748
rect 42150 16736 42156 16748
rect 42208 16736 42214 16788
rect 45830 16776 45836 16788
rect 45791 16748 45836 16776
rect 45830 16736 45836 16748
rect 45888 16736 45894 16788
rect 47578 16708 47584 16720
rect 41386 16680 47584 16708
rect 47578 16668 47584 16680
rect 47636 16668 47642 16720
rect 27982 16640 27988 16652
rect 25648 16612 26004 16640
rect 26068 16612 27988 16640
rect 25648 16600 25654 16612
rect 25682 16572 25688 16584
rect 25087 16544 25544 16572
rect 25643 16544 25688 16572
rect 25087 16541 25099 16544
rect 25041 16535 25099 16541
rect 25682 16532 25688 16544
rect 25740 16532 25746 16584
rect 25866 16572 25872 16584
rect 25827 16544 25872 16572
rect 25866 16532 25872 16544
rect 25924 16532 25930 16584
rect 25976 16581 26004 16612
rect 25961 16575 26019 16581
rect 25961 16541 25973 16575
rect 26007 16541 26019 16575
rect 26234 16572 26240 16584
rect 26195 16544 26240 16572
rect 25961 16535 26019 16541
rect 26234 16532 26240 16544
rect 26292 16532 26298 16584
rect 27724 16581 27752 16612
rect 27982 16600 27988 16612
rect 28040 16600 28046 16652
rect 33042 16600 33048 16652
rect 33100 16640 33106 16652
rect 33100 16612 33824 16640
rect 33100 16600 33106 16612
rect 27709 16575 27767 16581
rect 27709 16541 27721 16575
rect 27755 16541 27767 16575
rect 27709 16535 27767 16541
rect 30745 16575 30803 16581
rect 30745 16541 30757 16575
rect 30791 16572 30803 16575
rect 31478 16572 31484 16584
rect 30791 16544 31484 16572
rect 30791 16541 30803 16544
rect 30745 16535 30803 16541
rect 31478 16532 31484 16544
rect 31536 16532 31542 16584
rect 31573 16575 31631 16581
rect 31573 16541 31585 16575
rect 31619 16572 31631 16575
rect 31662 16572 31668 16584
rect 31619 16544 31668 16572
rect 31619 16541 31631 16544
rect 31573 16535 31631 16541
rect 31662 16532 31668 16544
rect 31720 16532 31726 16584
rect 31772 16544 32996 16572
rect 1578 16504 1584 16516
rect 1539 16476 1584 16504
rect 1578 16464 1584 16476
rect 1636 16464 1642 16516
rect 2590 16464 2596 16516
rect 2648 16504 2654 16516
rect 15746 16504 15752 16516
rect 2648 16476 15752 16504
rect 2648 16464 2654 16476
rect 15746 16464 15752 16476
rect 15804 16464 15810 16516
rect 15838 16464 15844 16516
rect 15896 16504 15902 16516
rect 16577 16507 16635 16513
rect 16577 16504 16589 16507
rect 15896 16476 16589 16504
rect 15896 16464 15902 16476
rect 16577 16473 16589 16476
rect 16623 16473 16635 16507
rect 16577 16467 16635 16473
rect 19058 16464 19064 16516
rect 19116 16504 19122 16516
rect 19521 16507 19579 16513
rect 19521 16504 19533 16507
rect 19116 16476 19533 16504
rect 19116 16464 19122 16476
rect 19521 16473 19533 16476
rect 19567 16473 19579 16507
rect 19521 16467 19579 16473
rect 20524 16507 20582 16513
rect 20524 16473 20536 16507
rect 20570 16504 20582 16507
rect 22554 16504 22560 16516
rect 20570 16476 22560 16504
rect 20570 16473 20582 16476
rect 20524 16467 20582 16473
rect 22554 16464 22560 16476
rect 22612 16464 22618 16516
rect 22922 16464 22928 16516
rect 22980 16504 22986 16516
rect 26789 16507 26847 16513
rect 26789 16504 26801 16507
rect 22980 16476 26801 16504
rect 22980 16464 22986 16476
rect 26789 16473 26801 16476
rect 26835 16473 26847 16507
rect 26789 16467 26847 16473
rect 30374 16464 30380 16516
rect 30432 16504 30438 16516
rect 30929 16507 30987 16513
rect 30929 16504 30941 16507
rect 30432 16476 30941 16504
rect 30432 16464 30438 16476
rect 30929 16473 30941 16476
rect 30975 16504 30987 16507
rect 31772 16504 31800 16544
rect 30975 16476 31800 16504
rect 31840 16507 31898 16513
rect 30975 16473 30987 16476
rect 30929 16467 30987 16473
rect 31840 16473 31852 16507
rect 31886 16504 31898 16507
rect 32122 16504 32128 16516
rect 31886 16476 32128 16504
rect 31886 16473 31898 16476
rect 31840 16467 31898 16473
rect 32122 16464 32128 16476
rect 32180 16464 32186 16516
rect 13814 16396 13820 16448
rect 13872 16436 13878 16448
rect 15470 16436 15476 16448
rect 13872 16408 15476 16436
rect 13872 16396 13878 16408
rect 15470 16396 15476 16408
rect 15528 16396 15534 16448
rect 16025 16439 16083 16445
rect 16025 16405 16037 16439
rect 16071 16436 16083 16439
rect 17034 16436 17040 16448
rect 16071 16408 17040 16436
rect 16071 16405 16083 16408
rect 16025 16399 16083 16405
rect 17034 16396 17040 16408
rect 17092 16396 17098 16448
rect 21634 16436 21640 16448
rect 21595 16408 21640 16436
rect 21634 16396 21640 16408
rect 21692 16396 21698 16448
rect 21818 16396 21824 16448
rect 21876 16436 21882 16448
rect 22189 16439 22247 16445
rect 22189 16436 22201 16439
rect 21876 16408 22201 16436
rect 21876 16396 21882 16408
rect 22189 16405 22201 16408
rect 22235 16405 22247 16439
rect 22738 16436 22744 16448
rect 22699 16408 22744 16436
rect 22189 16399 22247 16405
rect 22738 16396 22744 16408
rect 22796 16396 22802 16448
rect 24394 16396 24400 16448
rect 24452 16436 24458 16448
rect 25130 16436 25136 16448
rect 24452 16408 25136 16436
rect 24452 16396 24458 16408
rect 25130 16396 25136 16408
rect 25188 16396 25194 16448
rect 31113 16439 31171 16445
rect 31113 16405 31125 16439
rect 31159 16436 31171 16439
rect 32582 16436 32588 16448
rect 31159 16408 32588 16436
rect 31159 16405 31171 16408
rect 31113 16399 31171 16405
rect 32582 16396 32588 16408
rect 32640 16396 32646 16448
rect 32968 16445 32996 16544
rect 33410 16532 33416 16584
rect 33468 16572 33474 16584
rect 33796 16581 33824 16612
rect 33689 16575 33747 16581
rect 33689 16572 33701 16575
rect 33468 16544 33701 16572
rect 33468 16532 33474 16544
rect 33689 16541 33701 16544
rect 33735 16541 33747 16575
rect 33689 16535 33747 16541
rect 33781 16575 33839 16581
rect 33781 16541 33793 16575
rect 33827 16541 33839 16575
rect 33781 16535 33839 16541
rect 33870 16532 33876 16584
rect 33928 16572 33934 16584
rect 34072 16581 34100 16668
rect 35986 16600 35992 16652
rect 36044 16640 36050 16652
rect 40126 16640 40132 16652
rect 36044 16612 40132 16640
rect 36044 16600 36050 16612
rect 40126 16600 40132 16612
rect 40184 16600 40190 16652
rect 45922 16600 45928 16652
rect 45980 16640 45986 16652
rect 46293 16643 46351 16649
rect 46293 16640 46305 16643
rect 45980 16612 46305 16640
rect 45980 16600 45986 16612
rect 46293 16609 46305 16612
rect 46339 16609 46351 16643
rect 46293 16603 46351 16609
rect 34057 16575 34115 16581
rect 33928 16544 33973 16572
rect 33928 16532 33934 16544
rect 34057 16541 34069 16575
rect 34103 16541 34115 16575
rect 34057 16535 34115 16541
rect 38657 16575 38715 16581
rect 38657 16541 38669 16575
rect 38703 16541 38715 16575
rect 38657 16535 38715 16541
rect 39209 16575 39267 16581
rect 39209 16541 39221 16575
rect 39255 16572 39267 16575
rect 45830 16572 45836 16584
rect 39255 16544 45836 16572
rect 39255 16541 39267 16544
rect 39209 16535 39267 16541
rect 33594 16464 33600 16516
rect 33652 16504 33658 16516
rect 36357 16507 36415 16513
rect 36357 16504 36369 16507
rect 33652 16476 36369 16504
rect 33652 16464 33658 16476
rect 36357 16473 36369 16476
rect 36403 16504 36415 16507
rect 37458 16504 37464 16516
rect 36403 16476 37464 16504
rect 36403 16473 36415 16476
rect 36357 16467 36415 16473
rect 37458 16464 37464 16476
rect 37516 16504 37522 16516
rect 38672 16504 38700 16535
rect 45830 16532 45836 16544
rect 45888 16532 45894 16584
rect 37516 16476 38700 16504
rect 40396 16507 40454 16513
rect 37516 16464 37522 16476
rect 40396 16473 40408 16507
rect 40442 16504 40454 16507
rect 41230 16504 41236 16516
rect 40442 16476 41236 16504
rect 40442 16473 40454 16476
rect 40396 16467 40454 16473
rect 41230 16464 41236 16476
rect 41288 16464 41294 16516
rect 41414 16464 41420 16516
rect 41472 16504 41478 16516
rect 41966 16504 41972 16516
rect 41472 16476 41644 16504
rect 41927 16476 41972 16504
rect 41472 16464 41478 16476
rect 32953 16439 33011 16445
rect 32953 16405 32965 16439
rect 32999 16405 33011 16439
rect 32953 16399 33011 16405
rect 33413 16439 33471 16445
rect 33413 16405 33425 16439
rect 33459 16436 33471 16439
rect 34238 16436 34244 16448
rect 33459 16408 34244 16436
rect 33459 16405 33471 16408
rect 33413 16399 33471 16405
rect 34238 16396 34244 16408
rect 34296 16396 34302 16448
rect 40770 16396 40776 16448
rect 40828 16436 40834 16448
rect 41509 16439 41567 16445
rect 41509 16436 41521 16439
rect 40828 16408 41521 16436
rect 40828 16396 40834 16408
rect 41509 16405 41521 16408
rect 41555 16405 41567 16439
rect 41616 16436 41644 16476
rect 41966 16464 41972 16476
rect 42024 16464 42030 16516
rect 46474 16504 46480 16516
rect 46435 16476 46480 16504
rect 46474 16464 46480 16476
rect 46532 16464 46538 16516
rect 48133 16507 48191 16513
rect 48133 16473 48145 16507
rect 48179 16473 48191 16507
rect 48133 16467 48191 16473
rect 42169 16439 42227 16445
rect 42169 16436 42181 16439
rect 41616 16408 42181 16436
rect 41509 16399 41567 16405
rect 42169 16405 42181 16408
rect 42215 16405 42227 16439
rect 42169 16399 42227 16405
rect 42337 16439 42395 16445
rect 42337 16405 42349 16439
rect 42383 16436 42395 16439
rect 42610 16436 42616 16448
rect 42383 16408 42616 16436
rect 42383 16405 42395 16408
rect 42337 16399 42395 16405
rect 42610 16396 42616 16408
rect 42668 16396 42674 16448
rect 46014 16396 46020 16448
rect 46072 16436 46078 16448
rect 48148 16436 48176 16467
rect 46072 16408 48176 16436
rect 46072 16396 46078 16408
rect 1104 16346 48852 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 48852 16346
rect 1104 16272 48852 16294
rect 1578 16192 1584 16244
rect 1636 16232 1642 16244
rect 2225 16235 2283 16241
rect 2225 16232 2237 16235
rect 1636 16204 2237 16232
rect 1636 16192 1642 16204
rect 2225 16201 2237 16204
rect 2271 16201 2283 16235
rect 20622 16232 20628 16244
rect 2225 16195 2283 16201
rect 13924 16204 20484 16232
rect 20583 16204 20628 16232
rect 13814 16164 13820 16176
rect 6886 16136 13820 16164
rect 1486 16056 1492 16108
rect 1544 16096 1550 16108
rect 2133 16099 2191 16105
rect 2133 16096 2145 16099
rect 1544 16068 2145 16096
rect 1544 16056 1550 16068
rect 2133 16065 2145 16068
rect 2179 16096 2191 16099
rect 6886 16096 6914 16136
rect 13814 16124 13820 16136
rect 13872 16124 13878 16176
rect 2179 16068 6914 16096
rect 13924 16096 13952 16204
rect 15470 16124 15476 16176
rect 15528 16164 15534 16176
rect 16206 16164 16212 16176
rect 15528 16136 16212 16164
rect 15528 16124 15534 16136
rect 16206 16124 16212 16136
rect 16264 16124 16270 16176
rect 17034 16164 17040 16176
rect 16995 16136 17040 16164
rect 17034 16124 17040 16136
rect 17092 16124 17098 16176
rect 20456 16164 20484 16204
rect 20622 16192 20628 16204
rect 20680 16192 20686 16244
rect 20732 16204 22968 16232
rect 20732 16164 20760 16204
rect 20456 16136 20760 16164
rect 21634 16124 21640 16176
rect 21692 16164 21698 16176
rect 22940 16164 22968 16204
rect 23014 16192 23020 16244
rect 23072 16232 23078 16244
rect 23661 16235 23719 16241
rect 23661 16232 23673 16235
rect 23072 16204 23673 16232
rect 23072 16192 23078 16204
rect 23661 16201 23673 16204
rect 23707 16201 23719 16235
rect 23661 16195 23719 16201
rect 24118 16192 24124 16244
rect 24176 16232 24182 16244
rect 24578 16232 24584 16244
rect 24176 16204 24584 16232
rect 24176 16192 24182 16204
rect 24578 16192 24584 16204
rect 24636 16192 24642 16244
rect 32122 16232 32128 16244
rect 32083 16204 32128 16232
rect 32122 16192 32128 16204
rect 32180 16192 32186 16244
rect 35526 16232 35532 16244
rect 35487 16204 35532 16232
rect 35526 16192 35532 16204
rect 35584 16192 35590 16244
rect 40034 16192 40040 16244
rect 40092 16232 40098 16244
rect 40681 16235 40739 16241
rect 40681 16232 40693 16235
rect 40092 16204 40693 16232
rect 40092 16192 40098 16204
rect 40681 16201 40693 16204
rect 40727 16201 40739 16235
rect 41230 16232 41236 16244
rect 41191 16204 41236 16232
rect 40681 16195 40739 16201
rect 41230 16192 41236 16204
rect 41288 16192 41294 16244
rect 46474 16232 46480 16244
rect 46435 16204 46480 16232
rect 46474 16192 46480 16204
rect 46532 16192 46538 16244
rect 30374 16164 30380 16176
rect 21692 16136 22232 16164
rect 22940 16136 30380 16164
rect 21692 16124 21698 16136
rect 14001 16099 14059 16105
rect 14001 16096 14013 16099
rect 13924 16068 14013 16096
rect 2179 16065 2191 16068
rect 2133 16059 2191 16065
rect 14001 16065 14013 16068
rect 14047 16065 14059 16099
rect 19242 16096 19248 16108
rect 19203 16068 19248 16096
rect 14001 16059 14059 16065
rect 19242 16056 19248 16068
rect 19300 16056 19306 16108
rect 20806 16096 20812 16108
rect 20767 16068 20812 16096
rect 20806 16056 20812 16068
rect 20864 16056 20870 16108
rect 21818 16096 21824 16108
rect 21779 16068 21824 16096
rect 21818 16056 21824 16068
rect 21876 16056 21882 16108
rect 21993 16099 22051 16105
rect 21993 16096 22005 16099
rect 21974 16065 22005 16096
rect 22039 16065 22051 16099
rect 21974 16059 22051 16065
rect 22106 16099 22164 16105
rect 22106 16065 22118 16099
rect 22152 16096 22164 16099
rect 22204 16096 22232 16136
rect 30374 16124 30380 16136
rect 30432 16124 30438 16176
rect 31018 16164 31024 16176
rect 30668 16136 31024 16164
rect 22388 16106 22600 16120
rect 22152 16068 22232 16096
rect 22296 16099 22600 16106
rect 22296 16068 22339 16099
rect 22152 16065 22164 16068
rect 22106 16059 22164 16065
rect 22327 16065 22339 16068
rect 22373 16096 22600 16099
rect 23106 16096 23112 16108
rect 22373 16092 23112 16096
rect 22373 16078 22416 16092
rect 22373 16065 22385 16078
rect 22572 16068 23112 16092
rect 22327 16059 22385 16065
rect 290 15988 296 16040
rect 348 16028 354 16040
rect 14182 16028 14188 16040
rect 348 16000 6914 16028
rect 14143 16000 14188 16028
rect 348 15988 354 16000
rect 6886 15960 6914 16000
rect 14182 15988 14188 16000
rect 14240 15988 14246 16040
rect 14461 16031 14519 16037
rect 14461 15997 14473 16031
rect 14507 15997 14519 16031
rect 14461 15991 14519 15997
rect 16853 16031 16911 16037
rect 16853 15997 16865 16031
rect 16899 15997 16911 16031
rect 16853 15991 16911 15997
rect 18233 16031 18291 16037
rect 18233 15997 18245 16031
rect 18279 15997 18291 16031
rect 19886 16028 19892 16040
rect 19847 16000 19892 16028
rect 18233 15991 18291 15997
rect 14476 15960 14504 15991
rect 6886 15932 14504 15960
rect 16868 15960 16896 15991
rect 18138 15960 18144 15972
rect 16868 15932 18144 15960
rect 18138 15920 18144 15932
rect 18196 15920 18202 15972
rect 12986 15852 12992 15904
rect 13044 15892 13050 15904
rect 18248 15892 18276 15991
rect 19886 15988 19892 16000
rect 19944 15988 19950 16040
rect 21726 15988 21732 16040
rect 21784 16028 21790 16040
rect 21974 16028 22002 16059
rect 23106 16056 23112 16068
rect 23164 16056 23170 16108
rect 23477 16099 23535 16105
rect 23477 16065 23489 16099
rect 23523 16096 23535 16099
rect 24118 16096 24124 16108
rect 23523 16068 24124 16096
rect 23523 16065 23535 16068
rect 23477 16059 23535 16065
rect 24118 16056 24124 16068
rect 24176 16056 24182 16108
rect 24305 16099 24363 16105
rect 24305 16065 24317 16099
rect 24351 16096 24363 16099
rect 24394 16096 24400 16108
rect 24351 16068 24400 16096
rect 24351 16065 24363 16068
rect 24305 16059 24363 16065
rect 24394 16056 24400 16068
rect 24452 16056 24458 16108
rect 24946 16096 24952 16108
rect 24907 16068 24952 16096
rect 24946 16056 24952 16068
rect 25004 16056 25010 16108
rect 29454 16096 29460 16108
rect 29415 16068 29460 16096
rect 29454 16056 29460 16068
rect 29512 16056 29518 16108
rect 30558 16096 30564 16108
rect 30519 16068 30564 16096
rect 30558 16056 30564 16068
rect 30616 16056 30622 16108
rect 30668 16105 30696 16136
rect 31018 16124 31024 16136
rect 31076 16124 31082 16176
rect 33042 16164 33048 16176
rect 32508 16136 33048 16164
rect 30653 16099 30711 16105
rect 30653 16065 30665 16099
rect 30699 16065 30711 16099
rect 30653 16059 30711 16065
rect 30742 16056 30748 16108
rect 30800 16096 30806 16108
rect 30929 16099 30987 16105
rect 30800 16068 30845 16096
rect 30800 16056 30806 16068
rect 30929 16065 30941 16099
rect 30975 16065 30987 16099
rect 30929 16059 30987 16065
rect 21784 16000 22002 16028
rect 22189 16031 22247 16037
rect 21784 15988 21790 16000
rect 22189 15997 22201 16031
rect 22235 16028 22247 16031
rect 22235 16000 22324 16028
rect 22235 15997 22247 16000
rect 22189 15991 22247 15997
rect 22296 15960 22324 16000
rect 22554 15988 22560 16040
rect 22612 16028 22618 16040
rect 23293 16031 23351 16037
rect 22612 16000 22657 16028
rect 22612 15988 22618 16000
rect 23293 15997 23305 16031
rect 23339 15997 23351 16031
rect 24412 16028 24440 16056
rect 25041 16031 25099 16037
rect 25041 16028 25053 16031
rect 24412 16000 25053 16028
rect 23293 15991 23351 15997
rect 25041 15997 25053 16000
rect 25087 15997 25099 16031
rect 25041 15991 25099 15997
rect 29641 16031 29699 16037
rect 29641 15997 29653 16031
rect 29687 16028 29699 16031
rect 30944 16028 30972 16059
rect 31938 16056 31944 16108
rect 31996 16096 32002 16108
rect 32508 16105 32536 16136
rect 33042 16124 33048 16136
rect 33100 16124 33106 16176
rect 33689 16167 33747 16173
rect 33689 16133 33701 16167
rect 33735 16164 33747 16167
rect 34146 16164 34152 16176
rect 33735 16136 34152 16164
rect 33735 16133 33747 16136
rect 33689 16127 33747 16133
rect 34146 16124 34152 16136
rect 34204 16124 34210 16176
rect 40052 16164 40080 16192
rect 39040 16136 40080 16164
rect 32401 16099 32459 16105
rect 32401 16096 32413 16099
rect 31996 16068 32413 16096
rect 31996 16056 32002 16068
rect 32401 16065 32413 16068
rect 32447 16065 32459 16099
rect 32401 16059 32459 16065
rect 32493 16099 32551 16105
rect 32493 16065 32505 16099
rect 32539 16065 32551 16099
rect 32493 16059 32551 16065
rect 32582 16056 32588 16108
rect 32640 16096 32646 16108
rect 32769 16099 32827 16105
rect 32640 16068 32685 16096
rect 32640 16056 32646 16068
rect 32769 16065 32781 16099
rect 32815 16096 32827 16099
rect 33226 16096 33232 16108
rect 32815 16068 33232 16096
rect 32815 16065 32827 16068
rect 32769 16059 32827 16065
rect 33226 16056 33232 16068
rect 33284 16056 33290 16108
rect 33502 16096 33508 16108
rect 33463 16068 33508 16096
rect 33502 16056 33508 16068
rect 33560 16056 33566 16108
rect 34238 16056 34244 16108
rect 34296 16096 34302 16108
rect 34405 16099 34463 16105
rect 34405 16096 34417 16099
rect 34296 16068 34417 16096
rect 34296 16056 34302 16068
rect 34405 16065 34417 16068
rect 34451 16065 34463 16099
rect 37458 16096 37464 16108
rect 37419 16068 37464 16096
rect 34405 16059 34463 16065
rect 37458 16056 37464 16068
rect 37516 16056 37522 16108
rect 39040 16105 39068 16136
rect 45830 16124 45836 16176
rect 45888 16164 45894 16176
rect 46566 16164 46572 16176
rect 45888 16136 46572 16164
rect 45888 16124 45894 16136
rect 46566 16124 46572 16136
rect 46624 16124 46630 16176
rect 39025 16099 39083 16105
rect 39025 16065 39037 16099
rect 39071 16065 39083 16099
rect 39025 16059 39083 16065
rect 39114 16102 39172 16108
rect 39114 16068 39126 16102
rect 39160 16068 39172 16102
rect 39114 16062 39172 16068
rect 31478 16028 31484 16040
rect 29687 16000 31484 16028
rect 29687 15997 29699 16000
rect 29641 15991 29699 15997
rect 22370 15960 22376 15972
rect 22296 15932 22376 15960
rect 22370 15920 22376 15932
rect 22428 15920 22434 15972
rect 13044 15864 18276 15892
rect 23308 15892 23336 15991
rect 31478 15988 31484 16000
rect 31536 15988 31542 16040
rect 33594 16028 33600 16040
rect 31726 16000 33600 16028
rect 23658 15920 23664 15972
rect 23716 15960 23722 15972
rect 24489 15963 24547 15969
rect 24489 15960 24501 15963
rect 23716 15932 24501 15960
rect 23716 15920 23722 15932
rect 24489 15929 24501 15932
rect 24535 15929 24547 15963
rect 24489 15923 24547 15929
rect 26878 15920 26884 15972
rect 26936 15960 26942 15972
rect 31726 15960 31754 16000
rect 33594 15988 33600 16000
rect 33652 15988 33658 16040
rect 34149 16031 34207 16037
rect 34149 15997 34161 16031
rect 34195 15997 34207 16031
rect 34149 15991 34207 15997
rect 26936 15932 31754 15960
rect 26936 15920 26942 15932
rect 34164 15904 34192 15991
rect 38930 15988 38936 16040
rect 38988 16028 38994 16040
rect 39132 16028 39160 16062
rect 39206 16056 39212 16108
rect 39264 16096 39270 16108
rect 39264 16068 39309 16096
rect 39264 16056 39270 16068
rect 39390 16056 39396 16108
rect 39448 16096 39454 16108
rect 40494 16096 40500 16108
rect 39448 16068 39493 16096
rect 40455 16068 40500 16096
rect 39448 16056 39454 16068
rect 40494 16056 40500 16068
rect 40552 16056 40558 16108
rect 40773 16099 40831 16105
rect 40773 16065 40785 16099
rect 40819 16096 40831 16099
rect 41046 16096 41052 16108
rect 40819 16068 41052 16096
rect 40819 16065 40831 16068
rect 40773 16059 40831 16065
rect 41046 16056 41052 16068
rect 41104 16056 41110 16108
rect 41417 16099 41475 16105
rect 41417 16065 41429 16099
rect 41463 16096 41475 16099
rect 41782 16096 41788 16108
rect 41463 16068 41788 16096
rect 41463 16065 41475 16068
rect 41417 16059 41475 16065
rect 41782 16056 41788 16068
rect 41840 16056 41846 16108
rect 42610 16096 42616 16108
rect 42571 16068 42616 16096
rect 42610 16056 42616 16068
rect 42668 16056 42674 16108
rect 46385 16099 46443 16105
rect 46385 16096 46397 16099
rect 45756 16068 46397 16096
rect 38988 16000 39160 16028
rect 40313 16031 40371 16037
rect 38988 15988 38994 16000
rect 40313 15997 40325 16031
rect 40359 16028 40371 16031
rect 42150 16028 42156 16040
rect 40359 16000 42156 16028
rect 40359 15997 40371 16000
rect 40313 15991 40371 15997
rect 42150 15988 42156 16000
rect 42208 15988 42214 16040
rect 37645 15963 37703 15969
rect 37645 15929 37657 15963
rect 37691 15960 37703 15963
rect 38378 15960 38384 15972
rect 37691 15932 38384 15960
rect 37691 15929 37703 15932
rect 37645 15923 37703 15929
rect 38378 15920 38384 15932
rect 38436 15960 38442 15972
rect 45756 15960 45784 16068
rect 46385 16065 46397 16068
rect 46431 16096 46443 16099
rect 47302 16096 47308 16108
rect 46431 16068 47308 16096
rect 46431 16065 46443 16068
rect 46385 16059 46443 16065
rect 47302 16056 47308 16068
rect 47360 16056 47366 16108
rect 47394 16056 47400 16108
rect 47452 16096 47458 16108
rect 47581 16099 47639 16105
rect 47581 16096 47593 16099
rect 47452 16068 47593 16096
rect 47452 16056 47458 16068
rect 47581 16065 47593 16068
rect 47627 16065 47639 16099
rect 47581 16059 47639 16065
rect 38436 15932 45784 15960
rect 38436 15920 38442 15932
rect 23750 15892 23756 15904
rect 23308 15864 23756 15892
rect 13044 15852 13050 15864
rect 23750 15852 23756 15864
rect 23808 15892 23814 15904
rect 26786 15892 26792 15904
rect 23808 15864 26792 15892
rect 23808 15852 23814 15864
rect 26786 15852 26792 15864
rect 26844 15852 26850 15904
rect 30285 15895 30343 15901
rect 30285 15861 30297 15895
rect 30331 15892 30343 15895
rect 30650 15892 30656 15904
rect 30331 15864 30656 15892
rect 30331 15861 30343 15864
rect 30285 15855 30343 15861
rect 30650 15852 30656 15864
rect 30708 15852 30714 15904
rect 31662 15852 31668 15904
rect 31720 15892 31726 15904
rect 34146 15892 34152 15904
rect 31720 15864 34152 15892
rect 31720 15852 31726 15864
rect 34146 15852 34152 15864
rect 34204 15852 34210 15904
rect 38749 15895 38807 15901
rect 38749 15861 38761 15895
rect 38795 15892 38807 15895
rect 39666 15892 39672 15904
rect 38795 15864 39672 15892
rect 38795 15861 38807 15864
rect 38749 15855 38807 15861
rect 39666 15852 39672 15864
rect 39724 15852 39730 15904
rect 42426 15892 42432 15904
rect 42387 15864 42432 15892
rect 42426 15852 42432 15864
rect 42484 15852 42490 15904
rect 45925 15895 45983 15901
rect 45925 15861 45937 15895
rect 45971 15892 45983 15895
rect 46290 15892 46296 15904
rect 45971 15864 46296 15892
rect 45971 15861 45983 15864
rect 45925 15855 45983 15861
rect 46290 15852 46296 15864
rect 46348 15852 46354 15904
rect 46474 15852 46480 15904
rect 46532 15892 46538 15904
rect 47673 15895 47731 15901
rect 47673 15892 47685 15895
rect 46532 15864 47685 15892
rect 46532 15852 46538 15864
rect 47673 15861 47685 15864
rect 47719 15861 47731 15895
rect 47673 15855 47731 15861
rect 1104 15802 48852 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 48852 15802
rect 1104 15728 48852 15750
rect 4614 15648 4620 15700
rect 4672 15688 4678 15700
rect 14182 15688 14188 15700
rect 4672 15660 6914 15688
rect 14143 15660 14188 15688
rect 4672 15648 4678 15660
rect 6886 15620 6914 15660
rect 14182 15648 14188 15660
rect 14240 15648 14246 15700
rect 15746 15648 15752 15700
rect 15804 15688 15810 15700
rect 17678 15688 17684 15700
rect 15804 15660 17684 15688
rect 15804 15648 15810 15660
rect 17678 15648 17684 15660
rect 17736 15688 17742 15700
rect 19886 15688 19892 15700
rect 17736 15660 19892 15688
rect 17736 15648 17742 15660
rect 19886 15648 19892 15660
rect 19944 15648 19950 15700
rect 20254 15648 20260 15700
rect 20312 15688 20318 15700
rect 21913 15691 21971 15697
rect 21913 15688 21925 15691
rect 20312 15660 21925 15688
rect 20312 15648 20318 15660
rect 21913 15657 21925 15660
rect 21959 15657 21971 15691
rect 30558 15688 30564 15700
rect 21913 15651 21971 15657
rect 22066 15660 30564 15688
rect 22066 15620 22094 15660
rect 30558 15648 30564 15660
rect 30616 15648 30622 15700
rect 31938 15688 31944 15700
rect 31726 15660 31944 15688
rect 6886 15592 22094 15620
rect 23658 15580 23664 15632
rect 23716 15620 23722 15632
rect 24210 15620 24216 15632
rect 23716 15592 24216 15620
rect 23716 15580 23722 15592
rect 24210 15580 24216 15592
rect 24268 15620 24274 15632
rect 24673 15623 24731 15629
rect 24673 15620 24685 15623
rect 24268 15592 24685 15620
rect 24268 15580 24274 15592
rect 24673 15589 24685 15592
rect 24719 15589 24731 15623
rect 24673 15583 24731 15589
rect 25317 15623 25375 15629
rect 25317 15589 25329 15623
rect 25363 15620 25375 15623
rect 26694 15620 26700 15632
rect 25363 15592 26700 15620
rect 25363 15589 25375 15592
rect 25317 15583 25375 15589
rect 26694 15580 26700 15592
rect 26752 15580 26758 15632
rect 16761 15555 16819 15561
rect 16761 15521 16773 15555
rect 16807 15552 16819 15555
rect 17862 15552 17868 15564
rect 16807 15524 17868 15552
rect 16807 15521 16819 15524
rect 16761 15515 16819 15521
rect 17862 15512 17868 15524
rect 17920 15512 17926 15564
rect 18138 15552 18144 15564
rect 18099 15524 18144 15552
rect 18138 15512 18144 15524
rect 18196 15512 18202 15564
rect 20625 15555 20683 15561
rect 20625 15521 20637 15555
rect 20671 15552 20683 15555
rect 20990 15552 20996 15564
rect 20671 15524 20996 15552
rect 20671 15521 20683 15524
rect 20625 15515 20683 15521
rect 20990 15512 20996 15524
rect 21048 15512 21054 15564
rect 21634 15512 21640 15564
rect 21692 15552 21698 15564
rect 22278 15552 22284 15564
rect 21692 15524 22284 15552
rect 21692 15512 21698 15524
rect 22278 15512 22284 15524
rect 22336 15512 22342 15564
rect 24946 15512 24952 15564
rect 25004 15552 25010 15564
rect 25004 15524 25452 15552
rect 25004 15512 25010 15524
rect 13262 15444 13268 15496
rect 13320 15484 13326 15496
rect 14090 15484 14096 15496
rect 13320 15456 14096 15484
rect 13320 15444 13326 15456
rect 14090 15444 14096 15456
rect 14148 15444 14154 15496
rect 15378 15484 15384 15496
rect 15339 15456 15384 15484
rect 15378 15444 15384 15456
rect 15436 15444 15442 15496
rect 16025 15487 16083 15493
rect 16025 15453 16037 15487
rect 16071 15484 16083 15487
rect 16574 15484 16580 15496
rect 16071 15456 16580 15484
rect 16071 15453 16083 15456
rect 16025 15447 16083 15453
rect 16574 15444 16580 15456
rect 16632 15444 16638 15496
rect 19242 15444 19248 15496
rect 19300 15484 19306 15496
rect 22465 15487 22523 15493
rect 19300 15456 21956 15484
rect 19300 15444 19306 15456
rect 15473 15419 15531 15425
rect 15473 15385 15485 15419
rect 15519 15416 15531 15419
rect 16945 15419 17003 15425
rect 15519 15388 16712 15416
rect 15519 15385 15531 15388
rect 15473 15379 15531 15385
rect 16209 15351 16267 15357
rect 16209 15317 16221 15351
rect 16255 15348 16267 15351
rect 16574 15348 16580 15360
rect 16255 15320 16580 15348
rect 16255 15317 16267 15320
rect 16209 15311 16267 15317
rect 16574 15308 16580 15320
rect 16632 15308 16638 15360
rect 16684 15348 16712 15388
rect 16945 15385 16957 15419
rect 16991 15385 17003 15419
rect 16945 15379 17003 15385
rect 20441 15419 20499 15425
rect 20441 15385 20453 15419
rect 20487 15416 20499 15419
rect 21450 15416 21456 15428
rect 20487 15388 21456 15416
rect 20487 15385 20499 15388
rect 20441 15379 20499 15385
rect 16960 15348 16988 15379
rect 21450 15376 21456 15388
rect 21508 15376 21514 15428
rect 21818 15416 21824 15428
rect 21779 15388 21824 15416
rect 21818 15376 21824 15388
rect 21876 15376 21882 15428
rect 21928 15416 21956 15456
rect 22465 15453 22477 15487
rect 22511 15484 22523 15487
rect 22554 15484 22560 15496
rect 22511 15456 22560 15484
rect 22511 15453 22523 15456
rect 22465 15447 22523 15453
rect 22554 15444 22560 15456
rect 22612 15444 22618 15496
rect 22738 15493 22744 15496
rect 22732 15484 22744 15493
rect 22699 15456 22744 15484
rect 22732 15447 22744 15456
rect 22738 15444 22744 15447
rect 22796 15444 22802 15496
rect 24394 15484 24400 15496
rect 24355 15456 24400 15484
rect 24394 15444 24400 15456
rect 24452 15444 24458 15496
rect 24578 15484 24584 15496
rect 24539 15456 24584 15484
rect 24578 15444 24584 15456
rect 24636 15484 24642 15496
rect 25424 15493 25452 15524
rect 25774 15512 25780 15564
rect 25832 15552 25838 15564
rect 26142 15552 26148 15564
rect 25832 15524 26148 15552
rect 25832 15512 25838 15524
rect 26142 15512 26148 15524
rect 26200 15552 26206 15564
rect 26513 15555 26571 15561
rect 26513 15552 26525 15555
rect 26200 15524 26525 15552
rect 26200 15512 26206 15524
rect 26513 15521 26525 15524
rect 26559 15521 26571 15555
rect 26513 15515 26571 15521
rect 25225 15487 25283 15493
rect 25225 15484 25237 15487
rect 24636 15456 25237 15484
rect 24636 15444 24642 15456
rect 25225 15453 25237 15456
rect 25271 15453 25283 15487
rect 25225 15447 25283 15453
rect 25409 15487 25467 15493
rect 25409 15453 25421 15487
rect 25455 15453 25467 15487
rect 25409 15447 25467 15453
rect 26234 15444 26240 15496
rect 26292 15484 26298 15496
rect 26329 15487 26387 15493
rect 26329 15484 26341 15487
rect 26292 15456 26341 15484
rect 26292 15444 26298 15456
rect 26329 15453 26341 15456
rect 26375 15484 26387 15487
rect 27617 15487 27675 15493
rect 26375 15456 27568 15484
rect 26375 15453 26387 15456
rect 26329 15447 26387 15453
rect 26878 15416 26884 15428
rect 21928 15388 26884 15416
rect 26878 15376 26884 15388
rect 26936 15376 26942 15428
rect 16684 15320 16988 15348
rect 19981 15351 20039 15357
rect 19981 15317 19993 15351
rect 20027 15348 20039 15351
rect 20254 15348 20260 15360
rect 20027 15320 20260 15348
rect 20027 15317 20039 15320
rect 19981 15311 20039 15317
rect 20254 15308 20260 15320
rect 20312 15308 20318 15360
rect 20346 15308 20352 15360
rect 20404 15348 20410 15360
rect 20404 15320 20449 15348
rect 20404 15308 20410 15320
rect 22186 15308 22192 15360
rect 22244 15348 22250 15360
rect 23198 15348 23204 15360
rect 22244 15320 23204 15348
rect 22244 15308 22250 15320
rect 23198 15308 23204 15320
rect 23256 15308 23262 15360
rect 23842 15348 23848 15360
rect 23803 15320 23848 15348
rect 23842 15308 23848 15320
rect 23900 15308 23906 15360
rect 24578 15308 24584 15360
rect 24636 15348 24642 15360
rect 25774 15348 25780 15360
rect 24636 15320 25780 15348
rect 24636 15308 24642 15320
rect 25774 15308 25780 15320
rect 25832 15308 25838 15360
rect 25958 15348 25964 15360
rect 25919 15320 25964 15348
rect 25958 15308 25964 15320
rect 26016 15308 26022 15360
rect 26418 15348 26424 15360
rect 26379 15320 26424 15348
rect 26418 15308 26424 15320
rect 26476 15308 26482 15360
rect 27540 15348 27568 15456
rect 27617 15453 27629 15487
rect 27663 15484 27675 15487
rect 29546 15484 29552 15496
rect 27663 15456 29552 15484
rect 27663 15453 27675 15456
rect 27617 15447 27675 15453
rect 29546 15444 29552 15456
rect 29604 15444 29610 15496
rect 30558 15484 30564 15496
rect 30519 15456 30564 15484
rect 30558 15444 30564 15456
rect 30616 15444 30622 15496
rect 30650 15444 30656 15496
rect 30708 15484 30714 15496
rect 30817 15487 30875 15493
rect 30817 15484 30829 15487
rect 30708 15456 30829 15484
rect 30708 15444 30714 15456
rect 30817 15453 30829 15456
rect 30863 15453 30875 15487
rect 30817 15447 30875 15453
rect 27884 15419 27942 15425
rect 27884 15385 27896 15419
rect 27930 15416 27942 15419
rect 28258 15416 28264 15428
rect 27930 15388 28264 15416
rect 27930 15385 27942 15388
rect 27884 15379 27942 15385
rect 28258 15376 28264 15388
rect 28316 15376 28322 15428
rect 30098 15416 30104 15428
rect 28828 15388 30104 15416
rect 28828 15348 28856 15388
rect 30098 15376 30104 15388
rect 30156 15416 30162 15428
rect 31726 15416 31754 15660
rect 31938 15648 31944 15660
rect 31996 15648 32002 15700
rect 39025 15691 39083 15697
rect 39025 15657 39037 15691
rect 39071 15688 39083 15691
rect 39206 15688 39212 15700
rect 39071 15660 39212 15688
rect 39071 15657 39083 15660
rect 39025 15651 39083 15657
rect 39206 15648 39212 15660
rect 39264 15648 39270 15700
rect 38930 15620 38936 15632
rect 37016 15592 38936 15620
rect 37016 15493 37044 15592
rect 38930 15580 38936 15592
rect 38988 15580 38994 15632
rect 38105 15555 38163 15561
rect 38105 15552 38117 15555
rect 37108 15524 38117 15552
rect 37108 15493 37136 15524
rect 38105 15521 38117 15524
rect 38151 15521 38163 15555
rect 38105 15515 38163 15521
rect 40126 15512 40132 15564
rect 40184 15552 40190 15564
rect 40313 15555 40371 15561
rect 40313 15552 40325 15555
rect 40184 15524 40325 15552
rect 40184 15512 40190 15524
rect 40313 15521 40325 15524
rect 40359 15521 40371 15555
rect 46290 15552 46296 15564
rect 46251 15524 46296 15552
rect 40313 15515 40371 15521
rect 46290 15512 46296 15524
rect 46348 15512 46354 15564
rect 46474 15552 46480 15564
rect 46435 15524 46480 15552
rect 46474 15512 46480 15524
rect 46532 15512 46538 15564
rect 48130 15552 48136 15564
rect 48091 15524 48136 15552
rect 48130 15512 48136 15524
rect 48188 15512 48194 15564
rect 36909 15487 36967 15493
rect 36909 15453 36921 15487
rect 36955 15453 36967 15487
rect 36909 15447 36967 15453
rect 37001 15487 37059 15493
rect 37001 15453 37013 15487
rect 37047 15453 37059 15487
rect 37001 15447 37059 15453
rect 37093 15487 37151 15493
rect 37093 15453 37105 15487
rect 37139 15453 37151 15487
rect 37093 15447 37151 15453
rect 34698 15416 34704 15428
rect 30156 15388 31754 15416
rect 34659 15388 34704 15416
rect 30156 15376 30162 15388
rect 34698 15376 34704 15388
rect 34756 15376 34762 15428
rect 34885 15419 34943 15425
rect 34885 15385 34897 15419
rect 34931 15416 34943 15419
rect 35710 15416 35716 15428
rect 34931 15388 35716 15416
rect 34931 15385 34943 15388
rect 34885 15379 34943 15385
rect 28994 15348 29000 15360
rect 27540 15320 28856 15348
rect 28955 15320 29000 15348
rect 28994 15308 29000 15320
rect 29052 15308 29058 15360
rect 30650 15308 30656 15360
rect 30708 15348 30714 15360
rect 34900 15348 34928 15379
rect 35710 15376 35716 15388
rect 35768 15376 35774 15428
rect 30708 15320 34928 15348
rect 35069 15351 35127 15357
rect 30708 15308 30714 15320
rect 35069 15317 35081 15351
rect 35115 15348 35127 15351
rect 35342 15348 35348 15360
rect 35115 15320 35348 15348
rect 35115 15317 35127 15320
rect 35069 15311 35127 15317
rect 35342 15308 35348 15320
rect 35400 15308 35406 15360
rect 36633 15351 36691 15357
rect 36633 15317 36645 15351
rect 36679 15348 36691 15351
rect 36722 15348 36728 15360
rect 36679 15320 36728 15348
rect 36679 15317 36691 15320
rect 36633 15311 36691 15317
rect 36722 15308 36728 15320
rect 36780 15308 36786 15360
rect 36924 15348 36952 15447
rect 37182 15444 37188 15496
rect 37240 15484 37246 15496
rect 37277 15487 37335 15493
rect 37277 15484 37289 15487
rect 37240 15456 37289 15484
rect 37240 15444 37246 15456
rect 37277 15453 37289 15456
rect 37323 15453 37335 15487
rect 37277 15447 37335 15453
rect 37737 15487 37795 15493
rect 37737 15453 37749 15487
rect 37783 15484 37795 15487
rect 38657 15487 38715 15493
rect 38657 15484 38669 15487
rect 37783 15456 38669 15484
rect 37783 15453 37795 15456
rect 37737 15447 37795 15453
rect 38657 15453 38669 15456
rect 38703 15484 38715 15487
rect 40580 15487 40638 15493
rect 38703 15456 39252 15484
rect 38703 15453 38715 15456
rect 38657 15447 38715 15453
rect 37918 15416 37924 15428
rect 37879 15388 37924 15416
rect 37918 15376 37924 15388
rect 37976 15376 37982 15428
rect 38838 15416 38844 15428
rect 38799 15388 38844 15416
rect 38838 15376 38844 15388
rect 38896 15376 38902 15428
rect 39224 15416 39252 15456
rect 40580 15453 40592 15487
rect 40626 15484 40638 15487
rect 42426 15484 42432 15496
rect 40626 15456 42432 15484
rect 40626 15453 40638 15456
rect 40580 15447 40638 15453
rect 42426 15444 42432 15456
rect 42484 15444 42490 15496
rect 42702 15416 42708 15428
rect 39224 15388 42708 15416
rect 42702 15376 42708 15388
rect 42760 15376 42766 15428
rect 40494 15348 40500 15360
rect 36924 15320 40500 15348
rect 40494 15308 40500 15320
rect 40552 15348 40558 15360
rect 41693 15351 41751 15357
rect 41693 15348 41705 15351
rect 40552 15320 41705 15348
rect 40552 15308 40558 15320
rect 41693 15317 41705 15320
rect 41739 15317 41751 15351
rect 41693 15311 41751 15317
rect 1104 15258 48852 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 48852 15258
rect 1104 15184 48852 15206
rect 1670 15104 1676 15156
rect 1728 15144 1734 15156
rect 1728 15116 24992 15144
rect 1728 15104 1734 15116
rect 16025 15079 16083 15085
rect 16025 15045 16037 15079
rect 16071 15076 16083 15079
rect 16853 15079 16911 15085
rect 16853 15076 16865 15079
rect 16071 15048 16865 15076
rect 16071 15045 16083 15048
rect 16025 15039 16083 15045
rect 16853 15045 16865 15048
rect 16899 15045 16911 15079
rect 16853 15039 16911 15045
rect 17678 15036 17684 15088
rect 17736 15076 17742 15088
rect 18969 15079 19027 15085
rect 18969 15076 18981 15079
rect 17736 15048 18981 15076
rect 17736 15036 17742 15048
rect 18969 15045 18981 15048
rect 19015 15045 19027 15079
rect 18969 15039 19027 15045
rect 20070 15036 20076 15088
rect 20128 15076 20134 15088
rect 20622 15076 20628 15088
rect 20128 15048 20628 15076
rect 20128 15036 20134 15048
rect 20622 15036 20628 15048
rect 20680 15036 20686 15088
rect 21450 15036 21456 15088
rect 21508 15076 21514 15088
rect 21821 15079 21879 15085
rect 21821 15076 21833 15079
rect 21508 15048 21833 15076
rect 21508 15036 21514 15048
rect 21821 15045 21833 15048
rect 21867 15045 21879 15079
rect 22833 15079 22891 15085
rect 22833 15076 22845 15079
rect 21821 15039 21879 15045
rect 22112 15048 22845 15076
rect 15838 14968 15844 15020
rect 15896 15008 15902 15020
rect 15933 15011 15991 15017
rect 15933 15008 15945 15011
rect 15896 14980 15945 15008
rect 15896 14968 15902 14980
rect 15933 14977 15945 14980
rect 15979 14977 15991 15011
rect 15933 14971 15991 14977
rect 21174 14968 21180 15020
rect 21232 15008 21238 15020
rect 22112 15017 22140 15048
rect 22833 15045 22845 15048
rect 22879 15045 22891 15079
rect 22833 15039 22891 15045
rect 23032 15048 23796 15076
rect 23032 15017 23060 15048
rect 22005 15011 22063 15017
rect 22005 15008 22017 15011
rect 21232 14980 22017 15008
rect 21232 14968 21238 14980
rect 22005 14977 22017 14980
rect 22051 14977 22063 15011
rect 22005 14971 22063 14977
rect 22097 15011 22155 15017
rect 22097 14977 22109 15011
rect 22143 14977 22155 15011
rect 22097 14971 22155 14977
rect 22373 15011 22431 15017
rect 22373 14977 22385 15011
rect 22419 14977 22431 15011
rect 22373 14971 22431 14977
rect 23017 15011 23075 15017
rect 23017 14977 23029 15011
rect 23063 14977 23075 15011
rect 23198 15008 23204 15020
rect 23159 14980 23204 15008
rect 23017 14971 23075 14977
rect 16669 14943 16727 14949
rect 16669 14909 16681 14943
rect 16715 14940 16727 14943
rect 16942 14940 16948 14952
rect 16715 14912 16948 14940
rect 16715 14909 16727 14912
rect 16669 14903 16727 14909
rect 16942 14900 16948 14912
rect 17000 14900 17006 14952
rect 18230 14940 18236 14952
rect 18191 14912 18236 14940
rect 18230 14900 18236 14912
rect 18288 14900 18294 14952
rect 21910 14900 21916 14952
rect 21968 14940 21974 14952
rect 22388 14940 22416 14971
rect 23198 14968 23204 14980
rect 23256 14968 23262 15020
rect 23293 15011 23351 15017
rect 23293 14977 23305 15011
rect 23339 14977 23351 15011
rect 23768 15008 23796 15048
rect 23842 15036 23848 15088
rect 23900 15076 23906 15088
rect 24857 15079 24915 15085
rect 24857 15076 24869 15079
rect 23900 15048 24869 15076
rect 23900 15036 23906 15048
rect 24857 15045 24869 15048
rect 24903 15045 24915 15079
rect 24857 15039 24915 15045
rect 24029 15011 24087 15017
rect 24029 15008 24041 15011
rect 23768 14980 24041 15008
rect 23293 14971 23351 14977
rect 24029 14977 24041 14980
rect 24075 15008 24087 15011
rect 24394 15008 24400 15020
rect 24075 14980 24400 15008
rect 24075 14977 24087 14980
rect 24029 14971 24087 14977
rect 21968 14912 22416 14940
rect 21968 14900 21974 14912
rect 4062 14832 4068 14884
rect 4120 14872 4126 14884
rect 4120 14844 6914 14872
rect 4120 14832 4126 14844
rect 6886 14804 6914 14844
rect 18046 14832 18052 14884
rect 18104 14872 18110 14884
rect 21450 14872 21456 14884
rect 18104 14844 21456 14872
rect 18104 14832 18110 14844
rect 21450 14832 21456 14844
rect 21508 14832 21514 14884
rect 22002 14832 22008 14884
rect 22060 14872 22066 14884
rect 23308 14872 23336 14971
rect 24394 14968 24400 14980
rect 24452 14968 24458 15020
rect 24964 15008 24992 15116
rect 25130 15104 25136 15156
rect 25188 15144 25194 15156
rect 27062 15144 27068 15156
rect 25188 15116 27068 15144
rect 25188 15104 25194 15116
rect 27062 15104 27068 15116
rect 27120 15104 27126 15156
rect 27433 15147 27491 15153
rect 27433 15113 27445 15147
rect 27479 15113 27491 15147
rect 27433 15107 27491 15113
rect 25041 15079 25099 15085
rect 25041 15045 25053 15079
rect 25087 15076 25099 15079
rect 27246 15076 27252 15088
rect 25087 15048 27252 15076
rect 25087 15045 25099 15048
rect 25041 15039 25099 15045
rect 27246 15036 27252 15048
rect 27304 15036 27310 15088
rect 24964 14980 25360 15008
rect 23382 14900 23388 14952
rect 23440 14940 23446 14952
rect 25222 14940 25228 14952
rect 23440 14912 25228 14940
rect 23440 14900 23446 14912
rect 25222 14900 25228 14912
rect 25280 14900 25286 14952
rect 22060 14844 23336 14872
rect 25332 14872 25360 14980
rect 25774 14968 25780 15020
rect 25832 15008 25838 15020
rect 26053 15011 26111 15017
rect 26053 15008 26065 15011
rect 25832 14980 26065 15008
rect 25832 14968 25838 14980
rect 26053 14977 26065 14980
rect 26099 15008 26111 15011
rect 27448 15008 27476 15107
rect 27522 15104 27528 15156
rect 27580 15144 27586 15156
rect 30285 15147 30343 15153
rect 27580 15116 30236 15144
rect 27580 15104 27586 15116
rect 27893 15079 27951 15085
rect 27893 15045 27905 15079
rect 27939 15076 27951 15079
rect 28629 15079 28687 15085
rect 28629 15076 28641 15079
rect 27939 15048 28641 15076
rect 27939 15045 27951 15048
rect 27893 15039 27951 15045
rect 28629 15045 28641 15048
rect 28675 15076 28687 15079
rect 28994 15076 29000 15088
rect 28675 15048 29000 15076
rect 28675 15045 28687 15048
rect 28629 15039 28687 15045
rect 28994 15036 29000 15048
rect 29052 15036 29058 15088
rect 30098 15076 30104 15088
rect 30059 15048 30104 15076
rect 30098 15036 30104 15048
rect 30156 15036 30162 15088
rect 30208 15076 30236 15116
rect 30285 15113 30297 15147
rect 30331 15144 30343 15147
rect 30742 15144 30748 15156
rect 30331 15116 30748 15144
rect 30331 15113 30343 15116
rect 30285 15107 30343 15113
rect 30742 15104 30748 15116
rect 30800 15104 30806 15156
rect 46198 15144 46204 15156
rect 30852 15116 46204 15144
rect 30852 15076 30880 15116
rect 46198 15104 46204 15116
rect 46256 15104 46262 15156
rect 46382 15104 46388 15156
rect 46440 15144 46446 15156
rect 46845 15147 46903 15153
rect 46845 15144 46857 15147
rect 46440 15116 46857 15144
rect 46440 15104 46446 15116
rect 46845 15113 46857 15116
rect 46891 15113 46903 15147
rect 46845 15107 46903 15113
rect 30208 15048 30880 15076
rect 31018 15036 31024 15088
rect 31076 15076 31082 15088
rect 31076 15048 31337 15076
rect 31076 15036 31082 15048
rect 31309 15020 31337 15048
rect 31478 15036 31484 15088
rect 31536 15076 31542 15088
rect 35434 15076 35440 15088
rect 31536 15048 35440 15076
rect 31536 15036 31542 15048
rect 26099 14980 27476 15008
rect 27801 15011 27859 15017
rect 26099 14977 26111 14980
rect 26053 14971 26111 14977
rect 27801 14977 27813 15011
rect 27847 15008 27859 15011
rect 28166 15008 28172 15020
rect 27847 14980 28172 15008
rect 27847 14977 27859 14980
rect 27801 14971 27859 14977
rect 28166 14968 28172 14980
rect 28224 14968 28230 15020
rect 28810 14968 28816 15020
rect 28868 15008 28874 15020
rect 28905 15011 28963 15017
rect 28905 15008 28917 15011
rect 28868 14980 28917 15008
rect 28868 14968 28874 14980
rect 28905 14977 28917 14980
rect 28951 14977 28963 15011
rect 28905 14971 28963 14977
rect 29917 15011 29975 15017
rect 29917 14977 29929 15011
rect 29963 14977 29975 15011
rect 31185 15011 31243 15017
rect 31185 15008 31197 15011
rect 29917 14971 29975 14977
rect 30576 14980 31197 15008
rect 26145 14943 26203 14949
rect 26145 14909 26157 14943
rect 26191 14940 26203 14943
rect 26234 14940 26240 14952
rect 26191 14912 26240 14940
rect 26191 14909 26203 14912
rect 26145 14903 26203 14909
rect 26234 14900 26240 14912
rect 26292 14900 26298 14952
rect 27246 14900 27252 14952
rect 27304 14940 27310 14952
rect 27985 14943 28043 14949
rect 27985 14940 27997 14943
rect 27304 14912 27997 14940
rect 27304 14900 27310 14912
rect 27985 14909 27997 14912
rect 28031 14940 28043 14943
rect 28350 14940 28356 14952
rect 28031 14912 28356 14940
rect 28031 14909 28043 14912
rect 27985 14903 28043 14909
rect 28350 14900 28356 14912
rect 28408 14900 28414 14952
rect 28718 14940 28724 14952
rect 28679 14912 28724 14940
rect 28718 14900 28724 14912
rect 28776 14900 28782 14952
rect 29932 14940 29960 14971
rect 30374 14940 30380 14952
rect 29932 14912 30380 14940
rect 30374 14900 30380 14912
rect 30432 14900 30438 14952
rect 30576 14881 30604 14980
rect 31185 14977 31197 14980
rect 31231 14977 31243 15011
rect 31185 14971 31243 14977
rect 31294 15014 31352 15020
rect 31294 14980 31306 15014
rect 31340 14980 31352 15014
rect 31294 14974 31352 14980
rect 31386 14968 31392 15020
rect 31444 15017 31450 15020
rect 31588 15017 31616 15048
rect 35434 15036 35440 15048
rect 35492 15036 35498 15088
rect 36633 15079 36691 15085
rect 36633 15045 36645 15079
rect 36679 15076 36691 15079
rect 37461 15079 37519 15085
rect 37461 15076 37473 15079
rect 36679 15048 37473 15076
rect 36679 15045 36691 15048
rect 36633 15039 36691 15045
rect 37461 15045 37473 15048
rect 37507 15045 37519 15079
rect 40126 15076 40132 15088
rect 37461 15039 37519 15045
rect 39592 15048 40132 15076
rect 31444 15008 31452 15017
rect 31573 15011 31631 15017
rect 31444 14980 31489 15008
rect 31444 14971 31452 14980
rect 31573 14977 31585 15011
rect 31619 14977 31631 15011
rect 31573 14971 31631 14977
rect 31444 14968 31450 14971
rect 31662 14968 31668 15020
rect 31720 15008 31726 15020
rect 32125 15011 32183 15017
rect 32125 15008 32137 15011
rect 31720 14980 32137 15008
rect 31720 14968 31726 14980
rect 32125 14977 32137 14980
rect 32171 14977 32183 15011
rect 32381 15011 32439 15017
rect 32381 15008 32393 15011
rect 32125 14971 32183 14977
rect 32232 14980 32393 15008
rect 32232 14940 32260 14980
rect 32381 14977 32393 14980
rect 32427 14977 32439 15011
rect 32381 14971 32439 14977
rect 34146 14968 34152 15020
rect 34204 15008 34210 15020
rect 34606 15017 34612 15020
rect 34333 15011 34391 15017
rect 34333 15008 34345 15011
rect 34204 14980 34345 15008
rect 34204 14968 34210 14980
rect 34333 14977 34345 14980
rect 34379 14977 34391 15011
rect 34333 14971 34391 14977
rect 34600 14971 34612 15017
rect 34664 15008 34670 15020
rect 39592 15017 39620 15048
rect 40126 15036 40132 15048
rect 40184 15036 40190 15088
rect 36541 15011 36599 15017
rect 34664 14980 34700 15008
rect 34606 14968 34612 14971
rect 34664 14968 34670 14980
rect 36541 14977 36553 15011
rect 36587 15008 36599 15011
rect 39577 15011 39635 15017
rect 36587 14980 37228 15008
rect 36587 14977 36599 14980
rect 36541 14971 36599 14977
rect 32140 14912 32260 14940
rect 30561 14875 30619 14881
rect 30561 14872 30573 14875
rect 25332 14844 30573 14872
rect 22060 14832 22066 14844
rect 30561 14841 30573 14844
rect 30607 14841 30619 14875
rect 30561 14835 30619 14841
rect 30929 14875 30987 14881
rect 30929 14841 30941 14875
rect 30975 14872 30987 14875
rect 32140 14872 32168 14912
rect 35710 14872 35716 14884
rect 30975 14844 32168 14872
rect 35671 14844 35716 14872
rect 30975 14841 30987 14844
rect 30929 14835 30987 14841
rect 35710 14832 35716 14844
rect 35768 14832 35774 14884
rect 37200 14872 37228 14980
rect 39577 14977 39589 15011
rect 39623 14977 39635 15011
rect 39577 14971 39635 14977
rect 39666 14968 39672 15020
rect 39724 15008 39730 15020
rect 39833 15011 39891 15017
rect 39833 15008 39845 15011
rect 39724 14980 39845 15008
rect 39724 14968 39730 14980
rect 39833 14977 39845 14980
rect 39879 14977 39891 15011
rect 39833 14971 39891 14977
rect 46842 14968 46848 15020
rect 46900 15008 46906 15020
rect 47029 15011 47087 15017
rect 47029 15008 47041 15011
rect 46900 14980 47041 15008
rect 46900 14968 46906 14980
rect 47029 14977 47041 14980
rect 47075 14977 47087 15011
rect 47029 14971 47087 14977
rect 37277 14943 37335 14949
rect 37277 14909 37289 14943
rect 37323 14940 37335 14943
rect 37918 14940 37924 14952
rect 37323 14912 37924 14940
rect 37323 14909 37335 14912
rect 37277 14903 37335 14909
rect 37918 14900 37924 14912
rect 37976 14900 37982 14952
rect 39022 14940 39028 14952
rect 38983 14912 39028 14940
rect 39022 14900 39028 14912
rect 39080 14900 39086 14952
rect 38378 14872 38384 14884
rect 37200 14844 38384 14872
rect 38378 14832 38384 14844
rect 38436 14832 38442 14884
rect 20070 14804 20076 14816
rect 6886 14776 20076 14804
rect 20070 14764 20076 14776
rect 20128 14804 20134 14816
rect 20257 14807 20315 14813
rect 20257 14804 20269 14807
rect 20128 14776 20269 14804
rect 20128 14764 20134 14776
rect 20257 14773 20269 14776
rect 20303 14773 20315 14807
rect 20257 14767 20315 14773
rect 21634 14764 21640 14816
rect 21692 14804 21698 14816
rect 22186 14804 22192 14816
rect 21692 14776 22192 14804
rect 21692 14764 21698 14776
rect 22186 14764 22192 14776
rect 22244 14764 22250 14816
rect 22281 14807 22339 14813
rect 22281 14773 22293 14807
rect 22327 14804 22339 14807
rect 23290 14804 23296 14816
rect 22327 14776 23296 14804
rect 22327 14773 22339 14776
rect 22281 14767 22339 14773
rect 23290 14764 23296 14776
rect 23348 14764 23354 14816
rect 24026 14764 24032 14816
rect 24084 14804 24090 14816
rect 24213 14807 24271 14813
rect 24213 14804 24225 14807
rect 24084 14776 24225 14804
rect 24084 14764 24090 14776
rect 24213 14773 24225 14776
rect 24259 14773 24271 14807
rect 26142 14804 26148 14816
rect 26103 14776 26148 14804
rect 24213 14767 24271 14773
rect 26142 14764 26148 14776
rect 26200 14764 26206 14816
rect 26418 14804 26424 14816
rect 26379 14776 26424 14804
rect 26418 14764 26424 14776
rect 26476 14764 26482 14816
rect 28718 14804 28724 14816
rect 28679 14776 28724 14804
rect 28718 14764 28724 14776
rect 28776 14764 28782 14816
rect 29086 14804 29092 14816
rect 29047 14776 29092 14804
rect 29086 14764 29092 14776
rect 29144 14764 29150 14816
rect 31202 14764 31208 14816
rect 31260 14804 31266 14816
rect 33410 14804 33416 14816
rect 31260 14776 33416 14804
rect 31260 14764 31266 14776
rect 33410 14764 33416 14776
rect 33468 14804 33474 14816
rect 33505 14807 33563 14813
rect 33505 14804 33517 14807
rect 33468 14776 33517 14804
rect 33468 14764 33474 14776
rect 33505 14773 33517 14776
rect 33551 14773 33563 14807
rect 33505 14767 33563 14773
rect 38838 14764 38844 14816
rect 38896 14804 38902 14816
rect 40957 14807 41015 14813
rect 40957 14804 40969 14807
rect 38896 14776 40969 14804
rect 38896 14764 38902 14776
rect 40957 14773 40969 14776
rect 41003 14773 41015 14807
rect 47762 14804 47768 14816
rect 47723 14776 47768 14804
rect 40957 14767 41015 14773
rect 47762 14764 47768 14776
rect 47820 14764 47826 14816
rect 1104 14714 48852 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 48852 14714
rect 1104 14640 48852 14662
rect 16758 14560 16764 14612
rect 16816 14600 16822 14612
rect 16945 14603 17003 14609
rect 16945 14600 16957 14603
rect 16816 14572 16957 14600
rect 16816 14560 16822 14572
rect 16945 14569 16957 14572
rect 16991 14569 17003 14603
rect 21358 14600 21364 14612
rect 16945 14563 17003 14569
rect 19260 14572 21364 14600
rect 17954 14424 17960 14476
rect 18012 14464 18018 14476
rect 18874 14464 18880 14476
rect 18012 14436 18880 14464
rect 18012 14424 18018 14436
rect 18874 14424 18880 14436
rect 18932 14464 18938 14476
rect 19260 14473 19288 14572
rect 21358 14560 21364 14572
rect 21416 14560 21422 14612
rect 25409 14603 25467 14609
rect 25409 14569 25421 14603
rect 25455 14600 25467 14603
rect 25866 14600 25872 14612
rect 25455 14572 25872 14600
rect 25455 14569 25467 14572
rect 25409 14563 25467 14569
rect 25866 14560 25872 14572
rect 25924 14560 25930 14612
rect 26694 14600 26700 14612
rect 26655 14572 26700 14600
rect 26694 14560 26700 14572
rect 26752 14560 26758 14612
rect 29086 14600 29092 14612
rect 26804 14572 29092 14600
rect 20346 14492 20352 14544
rect 20404 14532 20410 14544
rect 20625 14535 20683 14541
rect 20625 14532 20637 14535
rect 20404 14504 20637 14532
rect 20404 14492 20410 14504
rect 20625 14501 20637 14504
rect 20671 14532 20683 14535
rect 21450 14532 21456 14544
rect 20671 14504 21456 14532
rect 20671 14501 20683 14504
rect 20625 14495 20683 14501
rect 21450 14492 21456 14504
rect 21508 14492 21514 14544
rect 21634 14492 21640 14544
rect 21692 14532 21698 14544
rect 22005 14535 22063 14541
rect 22005 14532 22017 14535
rect 21692 14504 22017 14532
rect 21692 14492 21698 14504
rect 22005 14501 22017 14504
rect 22051 14501 22063 14535
rect 22005 14495 22063 14501
rect 23474 14492 23480 14544
rect 23532 14532 23538 14544
rect 26804 14532 26832 14572
rect 29086 14560 29092 14572
rect 29144 14560 29150 14612
rect 31386 14560 31392 14612
rect 31444 14600 31450 14612
rect 31481 14603 31539 14609
rect 31481 14600 31493 14603
rect 31444 14572 31493 14600
rect 31444 14560 31450 14572
rect 31481 14569 31493 14572
rect 31527 14569 31539 14603
rect 31481 14563 31539 14569
rect 34606 14560 34612 14612
rect 34664 14600 34670 14612
rect 34701 14603 34759 14609
rect 34701 14600 34713 14603
rect 34664 14572 34713 14600
rect 34664 14560 34670 14572
rect 34701 14569 34713 14572
rect 34747 14569 34759 14603
rect 37829 14603 37887 14609
rect 34701 14563 34759 14569
rect 34992 14572 36492 14600
rect 23532 14504 26832 14532
rect 26973 14535 27031 14541
rect 23532 14492 23538 14504
rect 26973 14501 26985 14535
rect 27019 14501 27031 14535
rect 26973 14495 27031 14501
rect 19245 14467 19303 14473
rect 19245 14464 19257 14467
rect 18932 14436 19257 14464
rect 18932 14424 18938 14436
rect 19245 14433 19257 14436
rect 19291 14433 19303 14467
rect 19245 14427 19303 14433
rect 22278 14424 22284 14476
rect 22336 14464 22342 14476
rect 22465 14467 22523 14473
rect 22465 14464 22477 14467
rect 22336 14436 22477 14464
rect 22336 14424 22342 14436
rect 22465 14433 22477 14436
rect 22511 14433 22523 14467
rect 22465 14427 22523 14433
rect 22649 14467 22707 14473
rect 22649 14433 22661 14467
rect 22695 14464 22707 14467
rect 23842 14464 23848 14476
rect 22695 14436 23848 14464
rect 22695 14433 22707 14436
rect 22649 14427 22707 14433
rect 23842 14424 23848 14436
rect 23900 14424 23906 14476
rect 25685 14467 25743 14473
rect 25685 14433 25697 14467
rect 25731 14464 25743 14467
rect 26142 14464 26148 14476
rect 25731 14436 26148 14464
rect 25731 14433 25743 14436
rect 25685 14427 25743 14433
rect 26142 14424 26148 14436
rect 26200 14424 26206 14476
rect 1762 14356 1768 14408
rect 1820 14396 1826 14408
rect 2041 14399 2099 14405
rect 2041 14396 2053 14399
rect 1820 14368 2053 14396
rect 1820 14356 1826 14368
rect 2041 14365 2053 14368
rect 2087 14365 2099 14399
rect 2041 14359 2099 14365
rect 16574 14356 16580 14408
rect 16632 14396 16638 14408
rect 16853 14399 16911 14405
rect 16853 14396 16865 14399
rect 16632 14368 16865 14396
rect 16632 14356 16638 14368
rect 16853 14365 16865 14368
rect 16899 14396 16911 14399
rect 17678 14396 17684 14408
rect 16899 14368 17684 14396
rect 16899 14365 16911 14368
rect 16853 14359 16911 14365
rect 17678 14356 17684 14368
rect 17736 14356 17742 14408
rect 21269 14399 21327 14405
rect 21269 14365 21281 14399
rect 21315 14396 21327 14399
rect 21818 14396 21824 14408
rect 21315 14368 21824 14396
rect 21315 14365 21327 14368
rect 21269 14359 21327 14365
rect 21818 14356 21824 14368
rect 21876 14356 21882 14408
rect 22186 14356 22192 14408
rect 22244 14396 22250 14408
rect 22373 14399 22431 14405
rect 22373 14396 22385 14399
rect 22244 14368 22385 14396
rect 22244 14356 22250 14368
rect 22373 14365 22385 14368
rect 22419 14396 22431 14399
rect 23106 14396 23112 14408
rect 22419 14368 23112 14396
rect 22419 14365 22431 14368
rect 22373 14359 22431 14365
rect 23106 14356 23112 14368
rect 23164 14356 23170 14408
rect 23860 14396 23888 14424
rect 24765 14399 24823 14405
rect 24765 14396 24777 14399
rect 23860 14368 24777 14396
rect 24765 14365 24777 14368
rect 24811 14365 24823 14399
rect 24765 14359 24823 14365
rect 25593 14399 25651 14405
rect 25593 14365 25605 14399
rect 25639 14365 25651 14399
rect 25774 14396 25780 14408
rect 25735 14368 25780 14396
rect 25593 14359 25651 14365
rect 18509 14331 18567 14337
rect 18509 14297 18521 14331
rect 18555 14328 18567 14331
rect 18598 14328 18604 14340
rect 18555 14300 18604 14328
rect 18555 14297 18567 14300
rect 18509 14291 18567 14297
rect 18598 14288 18604 14300
rect 18656 14288 18662 14340
rect 19512 14331 19570 14337
rect 19512 14297 19524 14331
rect 19558 14328 19570 14331
rect 20070 14328 20076 14340
rect 19558 14300 20076 14328
rect 19558 14297 19570 14300
rect 19512 14291 19570 14297
rect 20070 14288 20076 14300
rect 20128 14288 20134 14340
rect 21358 14288 21364 14340
rect 21416 14328 21422 14340
rect 21453 14331 21511 14337
rect 21453 14328 21465 14331
rect 21416 14300 21465 14328
rect 21416 14288 21422 14300
rect 21453 14297 21465 14300
rect 21499 14297 21511 14331
rect 25608 14328 25636 14359
rect 25774 14356 25780 14368
rect 25832 14356 25838 14408
rect 25869 14399 25927 14405
rect 25869 14365 25881 14399
rect 25915 14396 25927 14399
rect 25958 14396 25964 14408
rect 25915 14368 25964 14396
rect 25915 14365 25927 14368
rect 25869 14359 25927 14365
rect 25958 14356 25964 14368
rect 26016 14356 26022 14408
rect 26418 14396 26424 14408
rect 26379 14368 26424 14396
rect 26418 14356 26424 14368
rect 26476 14356 26482 14408
rect 26694 14396 26700 14408
rect 26655 14368 26700 14396
rect 26694 14356 26700 14368
rect 26752 14356 26758 14408
rect 26988 14396 27016 14495
rect 27062 14492 27068 14544
rect 27120 14532 27126 14544
rect 27982 14532 27988 14544
rect 27120 14504 27988 14532
rect 27120 14492 27126 14504
rect 27982 14492 27988 14504
rect 28040 14492 28046 14544
rect 28166 14492 28172 14544
rect 28224 14532 28230 14544
rect 31202 14532 31208 14544
rect 28224 14504 31208 14532
rect 28224 14492 28230 14504
rect 31202 14492 31208 14504
rect 31260 14492 31266 14544
rect 32677 14535 32735 14541
rect 32677 14501 32689 14535
rect 32723 14532 32735 14535
rect 33134 14532 33140 14544
rect 32723 14504 33140 14532
rect 32723 14501 32735 14504
rect 32677 14495 32735 14501
rect 33134 14492 33140 14504
rect 33192 14532 33198 14544
rect 33502 14532 33508 14544
rect 33192 14504 33508 14532
rect 33192 14492 33198 14504
rect 33502 14492 33508 14504
rect 33560 14492 33566 14544
rect 34146 14532 34152 14544
rect 34107 14504 34152 14532
rect 34146 14492 34152 14504
rect 34204 14532 34210 14544
rect 34992 14532 35020 14572
rect 34204 14504 35020 14532
rect 34204 14492 34210 14504
rect 27338 14424 27344 14476
rect 27396 14464 27402 14476
rect 27801 14467 27859 14473
rect 27396 14436 27752 14464
rect 27396 14424 27402 14436
rect 27724 14405 27752 14436
rect 27801 14433 27813 14467
rect 27847 14464 27859 14467
rect 28994 14464 29000 14476
rect 27847 14436 29000 14464
rect 27847 14433 27859 14436
rect 27801 14427 27859 14433
rect 28994 14424 29000 14436
rect 29052 14424 29058 14476
rect 31110 14424 31116 14476
rect 31168 14464 31174 14476
rect 34422 14464 34428 14476
rect 31168 14436 34428 14464
rect 31168 14424 31174 14436
rect 34422 14424 34428 14436
rect 34480 14464 34486 14476
rect 36464 14473 36492 14572
rect 37829 14569 37841 14603
rect 37875 14600 37887 14603
rect 37918 14600 37924 14612
rect 37875 14572 37924 14600
rect 37875 14569 37887 14572
rect 37829 14563 37887 14569
rect 37918 14560 37924 14572
rect 37976 14560 37982 14612
rect 36449 14467 36507 14473
rect 34480 14436 35112 14464
rect 34480 14424 34486 14436
rect 27525 14399 27583 14405
rect 27525 14396 27537 14399
rect 26988 14368 27537 14396
rect 27525 14365 27537 14368
rect 27571 14365 27583 14399
rect 27525 14359 27583 14365
rect 27709 14399 27767 14405
rect 27709 14365 27721 14399
rect 27755 14365 27767 14399
rect 27890 14396 27896 14408
rect 27851 14368 27896 14396
rect 27709 14359 27767 14365
rect 26234 14328 26240 14340
rect 25608 14300 26240 14328
rect 21453 14291 21511 14297
rect 26234 14288 26240 14300
rect 26292 14288 26298 14340
rect 18616 14260 18644 14288
rect 27724 14272 27752 14359
rect 27890 14356 27896 14368
rect 27948 14356 27954 14408
rect 28077 14399 28135 14405
rect 28077 14365 28089 14399
rect 28123 14396 28135 14399
rect 28166 14396 28172 14408
rect 28123 14368 28172 14396
rect 28123 14365 28135 14368
rect 28077 14359 28135 14365
rect 28166 14356 28172 14368
rect 28224 14356 28230 14408
rect 28258 14356 28264 14408
rect 28316 14396 28322 14408
rect 28316 14368 28361 14396
rect 28316 14356 28322 14368
rect 29086 14356 29092 14408
rect 29144 14396 29150 14408
rect 32493 14399 32551 14405
rect 31220 14396 31340 14398
rect 32493 14396 32505 14399
rect 29144 14370 32505 14396
rect 29144 14368 31248 14370
rect 31312 14368 32505 14370
rect 29144 14356 29150 14368
rect 32493 14365 32505 14368
rect 32539 14365 32551 14399
rect 32493 14359 32551 14365
rect 34882 14356 34888 14408
rect 34940 14405 34946 14408
rect 35084 14405 35112 14436
rect 36449 14433 36461 14467
rect 36495 14433 36507 14467
rect 36449 14427 36507 14433
rect 37458 14424 37464 14476
rect 37516 14464 37522 14476
rect 44266 14464 44272 14476
rect 37516 14436 44272 14464
rect 37516 14424 37522 14436
rect 44266 14424 44272 14436
rect 44324 14424 44330 14476
rect 46293 14467 46351 14473
rect 46293 14433 46305 14467
rect 46339 14464 46351 14467
rect 47762 14464 47768 14476
rect 46339 14436 47768 14464
rect 46339 14433 46351 14436
rect 46293 14427 46351 14433
rect 47762 14424 47768 14436
rect 47820 14424 47826 14476
rect 34940 14399 34989 14405
rect 34940 14365 34943 14399
rect 34977 14365 34989 14399
rect 34940 14359 34989 14365
rect 35069 14399 35127 14405
rect 35069 14365 35081 14399
rect 35115 14365 35127 14399
rect 35069 14359 35127 14365
rect 34940 14356 34946 14359
rect 35158 14356 35164 14408
rect 35216 14402 35222 14408
rect 35216 14393 35224 14402
rect 35345 14399 35403 14405
rect 35216 14365 35258 14393
rect 35345 14365 35357 14399
rect 35391 14396 35403 14399
rect 35434 14396 35440 14408
rect 35391 14368 35440 14396
rect 35391 14365 35403 14368
rect 35216 14356 35224 14365
rect 35345 14359 35403 14365
rect 35434 14356 35440 14368
rect 35492 14356 35498 14408
rect 36722 14405 36728 14408
rect 36716 14396 36728 14405
rect 36683 14368 36728 14396
rect 36716 14359 36728 14368
rect 36722 14356 36728 14359
rect 36780 14356 36786 14408
rect 38378 14396 38384 14408
rect 38339 14368 38384 14396
rect 38378 14356 38384 14368
rect 38436 14356 38442 14408
rect 30374 14288 30380 14340
rect 30432 14328 30438 14340
rect 31113 14331 31171 14337
rect 31113 14328 31125 14331
rect 30432 14300 31125 14328
rect 30432 14288 30438 14300
rect 31113 14297 31125 14300
rect 31159 14297 31171 14331
rect 31113 14291 31171 14297
rect 22646 14260 22652 14272
rect 18616 14232 22652 14260
rect 22646 14220 22652 14232
rect 22704 14220 22710 14272
rect 22738 14220 22744 14272
rect 22796 14260 22802 14272
rect 23382 14260 23388 14272
rect 22796 14232 23388 14260
rect 22796 14220 22802 14232
rect 23382 14220 23388 14232
rect 23440 14220 23446 14272
rect 24394 14220 24400 14272
rect 24452 14260 24458 14272
rect 24857 14263 24915 14269
rect 24857 14260 24869 14263
rect 24452 14232 24869 14260
rect 24452 14220 24458 14232
rect 24857 14229 24869 14232
rect 24903 14229 24915 14263
rect 27706 14260 27712 14272
rect 27619 14232 27712 14260
rect 24857 14223 24915 14229
rect 27706 14220 27712 14232
rect 27764 14260 27770 14272
rect 28166 14260 28172 14272
rect 27764 14232 28172 14260
rect 27764 14220 27770 14232
rect 28166 14220 28172 14232
rect 28224 14220 28230 14272
rect 31128 14260 31156 14291
rect 31202 14288 31208 14340
rect 31260 14328 31266 14340
rect 31297 14331 31355 14337
rect 31297 14328 31309 14331
rect 31260 14300 31309 14328
rect 31260 14288 31266 14300
rect 31297 14297 31309 14300
rect 31343 14297 31355 14331
rect 31297 14291 31355 14297
rect 33042 14288 33048 14340
rect 33100 14328 33106 14340
rect 33965 14331 34023 14337
rect 33965 14328 33977 14331
rect 33100 14300 33977 14328
rect 33100 14288 33106 14300
rect 33965 14297 33977 14300
rect 34011 14297 34023 14331
rect 33965 14291 34023 14297
rect 38286 14288 38292 14340
rect 38344 14328 38350 14340
rect 46477 14331 46535 14337
rect 38344 14300 41414 14328
rect 38344 14288 38350 14300
rect 33502 14260 33508 14272
rect 31128 14232 33508 14260
rect 33502 14220 33508 14232
rect 33560 14260 33566 14272
rect 34698 14260 34704 14272
rect 33560 14232 34704 14260
rect 33560 14220 33566 14232
rect 34698 14220 34704 14232
rect 34756 14260 34762 14272
rect 35434 14260 35440 14272
rect 34756 14232 35440 14260
rect 34756 14220 34762 14232
rect 35434 14220 35440 14232
rect 35492 14220 35498 14272
rect 38470 14260 38476 14272
rect 38431 14232 38476 14260
rect 38470 14220 38476 14232
rect 38528 14220 38534 14272
rect 41386 14260 41414 14300
rect 46477 14297 46489 14331
rect 46523 14328 46535 14331
rect 46750 14328 46756 14340
rect 46523 14300 46756 14328
rect 46523 14297 46535 14300
rect 46477 14291 46535 14297
rect 46750 14288 46756 14300
rect 46808 14288 46814 14340
rect 48130 14328 48136 14340
rect 48091 14300 48136 14328
rect 48130 14288 48136 14300
rect 48188 14288 48194 14340
rect 47210 14260 47216 14272
rect 41386 14232 47216 14260
rect 47210 14220 47216 14232
rect 47268 14220 47274 14272
rect 1104 14170 48852 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 48852 14170
rect 1104 14096 48852 14118
rect 20070 14056 20076 14068
rect 20031 14028 20076 14056
rect 20070 14016 20076 14028
rect 20128 14016 20134 14068
rect 21174 14056 21180 14068
rect 21135 14028 21180 14056
rect 21174 14016 21180 14028
rect 21232 14016 21238 14068
rect 21818 14016 21824 14068
rect 21876 14056 21882 14068
rect 23201 14059 23259 14065
rect 23201 14056 23213 14059
rect 21876 14028 23213 14056
rect 21876 14016 21882 14028
rect 23201 14025 23213 14028
rect 23247 14025 23259 14059
rect 23201 14019 23259 14025
rect 24964 14028 27844 14056
rect 19613 13991 19671 13997
rect 19613 13957 19625 13991
rect 19659 13988 19671 13991
rect 24964 13988 24992 14028
rect 19659 13960 24992 13988
rect 25041 13991 25099 13997
rect 19659 13957 19671 13960
rect 19613 13951 19671 13957
rect 25041 13957 25053 13991
rect 25087 13988 25099 13991
rect 25958 13988 25964 14000
rect 25087 13960 25964 13988
rect 25087 13957 25099 13960
rect 25041 13951 25099 13957
rect 25958 13948 25964 13960
rect 26016 13948 26022 14000
rect 1762 13920 1768 13932
rect 1723 13892 1768 13920
rect 1762 13880 1768 13892
rect 1820 13880 1826 13932
rect 15838 13880 15844 13932
rect 15896 13920 15902 13932
rect 16669 13923 16727 13929
rect 16669 13920 16681 13923
rect 15896 13892 16681 13920
rect 15896 13880 15902 13892
rect 16669 13889 16681 13892
rect 16715 13889 16727 13923
rect 17678 13920 17684 13932
rect 17639 13892 17684 13920
rect 16669 13883 16727 13889
rect 17678 13880 17684 13892
rect 17736 13920 17742 13932
rect 19245 13923 19303 13929
rect 19245 13920 19257 13923
rect 17736 13892 19257 13920
rect 17736 13880 17742 13892
rect 19245 13889 19257 13892
rect 19291 13889 19303 13923
rect 20254 13920 20260 13932
rect 20215 13892 20260 13920
rect 19245 13883 19303 13889
rect 20254 13880 20260 13892
rect 20312 13880 20318 13932
rect 21085 13923 21143 13929
rect 21085 13889 21097 13923
rect 21131 13889 21143 13923
rect 21085 13883 21143 13889
rect 21269 13923 21327 13929
rect 21269 13889 21281 13923
rect 21315 13920 21327 13923
rect 21634 13920 21640 13932
rect 21315 13892 21640 13920
rect 21315 13889 21327 13892
rect 21269 13883 21327 13889
rect 1946 13852 1952 13864
rect 1907 13824 1952 13852
rect 1946 13812 1952 13824
rect 2004 13812 2010 13864
rect 2774 13852 2780 13864
rect 2735 13824 2780 13852
rect 2774 13812 2780 13824
rect 2832 13812 2838 13864
rect 14090 13812 14096 13864
rect 14148 13852 14154 13864
rect 18046 13852 18052 13864
rect 14148 13824 18052 13852
rect 14148 13812 14154 13824
rect 18046 13812 18052 13824
rect 18104 13852 18110 13864
rect 18414 13852 18420 13864
rect 18104 13824 18420 13852
rect 18104 13812 18110 13824
rect 18414 13812 18420 13824
rect 18472 13812 18478 13864
rect 3050 13744 3056 13796
rect 3108 13784 3114 13796
rect 18138 13784 18144 13796
rect 3108 13756 18144 13784
rect 3108 13744 3114 13756
rect 18138 13744 18144 13756
rect 18196 13744 18202 13796
rect 21100 13784 21128 13883
rect 21634 13880 21640 13892
rect 21692 13880 21698 13932
rect 21910 13880 21916 13932
rect 21968 13920 21974 13932
rect 22189 13923 22247 13929
rect 22189 13920 22201 13923
rect 21968 13892 22201 13920
rect 21968 13880 21974 13892
rect 22189 13889 22201 13892
rect 22235 13889 22247 13923
rect 22189 13883 22247 13889
rect 23109 13923 23167 13929
rect 23109 13889 23121 13923
rect 23155 13920 23167 13923
rect 24302 13920 24308 13932
rect 23155 13892 24308 13920
rect 23155 13889 23167 13892
rect 23109 13883 23167 13889
rect 24302 13880 24308 13892
rect 24360 13880 24366 13932
rect 24394 13880 24400 13932
rect 24452 13920 24458 13932
rect 25314 13920 25320 13932
rect 24452 13892 24497 13920
rect 25275 13892 25320 13920
rect 24452 13880 24458 13892
rect 25314 13880 25320 13892
rect 25372 13880 25378 13932
rect 25774 13880 25780 13932
rect 25832 13920 25838 13932
rect 26145 13923 26203 13929
rect 26145 13920 26157 13923
rect 25832 13892 26157 13920
rect 25832 13880 25838 13892
rect 26145 13889 26157 13892
rect 26191 13889 26203 13923
rect 26145 13883 26203 13889
rect 27709 13923 27767 13929
rect 27709 13889 27721 13923
rect 27755 13889 27767 13923
rect 27816 13920 27844 14028
rect 27982 14016 27988 14068
rect 28040 14056 28046 14068
rect 46750 14056 46756 14068
rect 28040 14028 41414 14056
rect 46711 14028 46756 14056
rect 28040 14016 28046 14028
rect 28905 13991 28963 13997
rect 28905 13957 28917 13991
rect 28951 13988 28963 13991
rect 31570 13988 31576 14000
rect 28951 13960 31576 13988
rect 28951 13957 28963 13960
rect 28905 13951 28963 13957
rect 31570 13948 31576 13960
rect 31628 13948 31634 14000
rect 32861 13991 32919 13997
rect 32861 13957 32873 13991
rect 32907 13988 32919 13991
rect 33134 13988 33140 14000
rect 32907 13960 33140 13988
rect 32907 13957 32919 13960
rect 32861 13951 32919 13957
rect 33134 13948 33140 13960
rect 33192 13948 33198 14000
rect 33502 13988 33508 14000
rect 33463 13960 33508 13988
rect 33502 13948 33508 13960
rect 33560 13948 33566 14000
rect 33873 13991 33931 13997
rect 33873 13957 33885 13991
rect 33919 13988 33931 13991
rect 33919 13960 34836 13988
rect 33919 13957 33931 13960
rect 33873 13951 33931 13957
rect 34808 13932 34836 13960
rect 35342 13948 35348 14000
rect 35400 13988 35406 14000
rect 35621 13991 35679 13997
rect 35621 13988 35633 13991
rect 35400 13960 35633 13988
rect 35400 13948 35406 13960
rect 35621 13957 35633 13960
rect 35667 13957 35679 13991
rect 38470 13988 38476 14000
rect 38431 13960 38476 13988
rect 35621 13951 35679 13957
rect 38470 13948 38476 13960
rect 38528 13948 38534 14000
rect 41386 13988 41414 14028
rect 46750 14016 46756 14028
rect 46808 14016 46814 14068
rect 48041 14059 48099 14065
rect 48041 14025 48053 14059
rect 48087 14025 48099 14059
rect 48041 14019 48099 14025
rect 48056 13988 48084 14019
rect 41386 13960 48084 13988
rect 32125 13923 32183 13929
rect 27816 13892 31754 13920
rect 27709 13883 27767 13889
rect 21450 13812 21456 13864
rect 21508 13852 21514 13864
rect 22278 13852 22284 13864
rect 21508 13824 22284 13852
rect 21508 13812 21514 13824
rect 22278 13812 22284 13824
rect 22336 13812 22342 13864
rect 22465 13855 22523 13861
rect 22465 13821 22477 13855
rect 22511 13821 22523 13855
rect 22465 13815 22523 13821
rect 21821 13787 21879 13793
rect 21821 13784 21833 13787
rect 21100 13756 21833 13784
rect 21821 13753 21833 13756
rect 21867 13784 21879 13787
rect 22002 13784 22008 13796
rect 21867 13756 22008 13784
rect 21867 13753 21879 13756
rect 21821 13747 21879 13753
rect 22002 13744 22008 13756
rect 22060 13744 22066 13796
rect 22480 13784 22508 13815
rect 23474 13784 23480 13796
rect 22480 13756 23480 13784
rect 23474 13744 23480 13756
rect 23532 13784 23538 13796
rect 24412 13784 24440 13880
rect 25225 13855 25283 13861
rect 25225 13821 25237 13855
rect 25271 13852 25283 13855
rect 25792 13852 25820 13880
rect 25271 13824 25820 13852
rect 25271 13821 25283 13824
rect 25225 13815 25283 13821
rect 26234 13812 26240 13864
rect 26292 13852 26298 13864
rect 26421 13855 26479 13861
rect 26421 13852 26433 13855
rect 26292 13824 26433 13852
rect 26292 13812 26298 13824
rect 26421 13821 26433 13824
rect 26467 13821 26479 13855
rect 26421 13815 26479 13821
rect 24578 13784 24584 13796
rect 23532 13756 24440 13784
rect 24539 13756 24584 13784
rect 23532 13744 23538 13756
rect 24578 13744 24584 13756
rect 24636 13744 24642 13796
rect 25961 13787 26019 13793
rect 25332 13756 25636 13784
rect 16761 13719 16819 13725
rect 16761 13685 16773 13719
rect 16807 13716 16819 13719
rect 16850 13716 16856 13728
rect 16807 13688 16856 13716
rect 16807 13685 16819 13688
rect 16761 13679 16819 13685
rect 16850 13676 16856 13688
rect 16908 13676 16914 13728
rect 20530 13676 20536 13728
rect 20588 13716 20594 13728
rect 21174 13716 21180 13728
rect 20588 13688 21180 13716
rect 20588 13676 20594 13688
rect 21174 13676 21180 13688
rect 21232 13676 21238 13728
rect 21358 13676 21364 13728
rect 21416 13716 21422 13728
rect 22554 13716 22560 13728
rect 21416 13688 22560 13716
rect 21416 13676 21422 13688
rect 22554 13676 22560 13688
rect 22612 13716 22618 13728
rect 24946 13716 24952 13728
rect 22612 13688 24952 13716
rect 22612 13676 22618 13688
rect 24946 13676 24952 13688
rect 25004 13676 25010 13728
rect 25332 13725 25360 13756
rect 25317 13719 25375 13725
rect 25317 13685 25329 13719
rect 25363 13685 25375 13719
rect 25498 13716 25504 13728
rect 25459 13688 25504 13716
rect 25317 13679 25375 13685
rect 25498 13676 25504 13688
rect 25556 13676 25562 13728
rect 25608 13716 25636 13756
rect 25961 13753 25973 13787
rect 26007 13784 26019 13787
rect 26694 13784 26700 13796
rect 26007 13756 26700 13784
rect 26007 13753 26019 13756
rect 25961 13747 26019 13753
rect 26694 13744 26700 13756
rect 26752 13744 26758 13796
rect 26142 13716 26148 13728
rect 25608 13688 26148 13716
rect 26142 13676 26148 13688
rect 26200 13716 26206 13728
rect 26329 13719 26387 13725
rect 26329 13716 26341 13719
rect 26200 13688 26341 13716
rect 26200 13676 26206 13688
rect 26329 13685 26341 13688
rect 26375 13716 26387 13719
rect 27341 13719 27399 13725
rect 27341 13716 27353 13719
rect 26375 13688 27353 13716
rect 26375 13685 26387 13688
rect 26329 13679 26387 13685
rect 27341 13685 27353 13688
rect 27387 13685 27399 13719
rect 27724 13716 27752 13883
rect 27801 13855 27859 13861
rect 27801 13821 27813 13855
rect 27847 13821 27859 13855
rect 27801 13815 27859 13821
rect 27893 13855 27951 13861
rect 27893 13821 27905 13855
rect 27939 13852 27951 13855
rect 28350 13852 28356 13864
rect 27939 13824 28356 13852
rect 27939 13821 27951 13824
rect 27893 13815 27951 13821
rect 27816 13784 27844 13815
rect 28350 13812 28356 13824
rect 28408 13812 28414 13864
rect 29086 13852 29092 13864
rect 29047 13824 29092 13852
rect 29086 13812 29092 13824
rect 29144 13812 29150 13864
rect 29822 13812 29828 13864
rect 29880 13852 29886 13864
rect 30101 13855 30159 13861
rect 30101 13852 30113 13855
rect 29880 13824 30113 13852
rect 29880 13812 29886 13824
rect 30101 13821 30113 13824
rect 30147 13821 30159 13855
rect 30374 13852 30380 13864
rect 30335 13824 30380 13852
rect 30101 13815 30159 13821
rect 30374 13812 30380 13824
rect 30432 13812 30438 13864
rect 31726 13852 31754 13892
rect 32125 13889 32137 13923
rect 32171 13920 32183 13923
rect 33318 13920 33324 13932
rect 32171 13892 33324 13920
rect 32171 13889 32183 13892
rect 32125 13883 32183 13889
rect 32140 13852 32168 13883
rect 33318 13880 33324 13892
rect 33376 13880 33382 13932
rect 33689 13923 33747 13929
rect 33689 13889 33701 13923
rect 33735 13889 33747 13923
rect 33689 13883 33747 13889
rect 31726 13824 32168 13852
rect 32214 13812 32220 13864
rect 32272 13852 32278 13864
rect 33042 13852 33048 13864
rect 32272 13824 33048 13852
rect 32272 13812 32278 13824
rect 33042 13812 33048 13824
rect 33100 13812 33106 13864
rect 27982 13784 27988 13796
rect 27816 13756 27988 13784
rect 27982 13744 27988 13756
rect 28040 13744 28046 13796
rect 31018 13744 31024 13796
rect 31076 13784 31082 13796
rect 33704 13784 33732 13883
rect 34514 13880 34520 13932
rect 34572 13929 34578 13932
rect 34572 13923 34621 13929
rect 34572 13889 34575 13923
rect 34609 13889 34621 13923
rect 34572 13883 34621 13889
rect 34682 13923 34740 13929
rect 34682 13889 34694 13923
rect 34728 13889 34740 13923
rect 34682 13883 34740 13889
rect 34793 13926 34851 13932
rect 34793 13892 34805 13926
rect 34839 13892 34851 13926
rect 34793 13886 34851 13892
rect 34977 13923 35035 13929
rect 34977 13889 34989 13923
rect 35023 13920 35035 13923
rect 35250 13920 35256 13932
rect 35023 13892 35256 13920
rect 35023 13889 35035 13892
rect 34977 13883 35035 13889
rect 34572 13880 34578 13883
rect 34422 13812 34428 13864
rect 34480 13852 34486 13864
rect 34697 13852 34725 13883
rect 35250 13880 35256 13892
rect 35308 13880 35314 13932
rect 35434 13920 35440 13932
rect 35395 13892 35440 13920
rect 35434 13880 35440 13892
rect 35492 13880 35498 13932
rect 46198 13880 46204 13932
rect 46256 13920 46262 13932
rect 46661 13923 46719 13929
rect 46661 13920 46673 13923
rect 46256 13892 46673 13920
rect 46256 13880 46262 13892
rect 46661 13889 46673 13892
rect 46707 13889 46719 13923
rect 47854 13920 47860 13932
rect 47815 13892 47860 13920
rect 46661 13883 46719 13889
rect 47854 13880 47860 13892
rect 47912 13880 47918 13932
rect 35802 13852 35808 13864
rect 34480 13824 34725 13852
rect 35763 13824 35808 13852
rect 34480 13812 34486 13824
rect 35802 13812 35808 13824
rect 35860 13812 35866 13864
rect 38289 13855 38347 13861
rect 38289 13821 38301 13855
rect 38335 13852 38347 13855
rect 38838 13852 38844 13864
rect 38335 13824 38844 13852
rect 38335 13821 38347 13824
rect 38289 13815 38347 13821
rect 38838 13812 38844 13824
rect 38896 13812 38902 13864
rect 39942 13852 39948 13864
rect 39903 13824 39948 13852
rect 39942 13812 39948 13824
rect 40000 13812 40006 13864
rect 35618 13784 35624 13796
rect 31076 13756 35624 13784
rect 31076 13744 31082 13756
rect 35618 13744 35624 13756
rect 35676 13744 35682 13796
rect 28718 13716 28724 13728
rect 27724 13688 28724 13716
rect 27341 13679 27399 13685
rect 28718 13676 28724 13688
rect 28776 13676 28782 13728
rect 32217 13719 32275 13725
rect 32217 13685 32229 13719
rect 32263 13716 32275 13719
rect 32490 13716 32496 13728
rect 32263 13688 32496 13716
rect 32263 13685 32275 13688
rect 32217 13679 32275 13685
rect 32490 13676 32496 13688
rect 32548 13676 32554 13728
rect 34333 13719 34391 13725
rect 34333 13685 34345 13719
rect 34379 13716 34391 13719
rect 34514 13716 34520 13728
rect 34379 13688 34520 13716
rect 34379 13685 34391 13688
rect 34333 13679 34391 13685
rect 34514 13676 34520 13688
rect 34572 13676 34578 13728
rect 1104 13626 48852 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 48852 13626
rect 1104 13552 48852 13574
rect 1946 13472 1952 13524
rect 2004 13512 2010 13524
rect 2133 13515 2191 13521
rect 2133 13512 2145 13515
rect 2004 13484 2145 13512
rect 2004 13472 2010 13484
rect 2133 13481 2145 13484
rect 2179 13481 2191 13515
rect 2133 13475 2191 13481
rect 16758 13472 16764 13524
rect 16816 13512 16822 13524
rect 18138 13512 18144 13524
rect 16816 13484 18144 13512
rect 16816 13472 16822 13484
rect 18138 13472 18144 13484
rect 18196 13472 18202 13524
rect 21453 13515 21511 13521
rect 21453 13481 21465 13515
rect 21499 13512 21511 13515
rect 21818 13512 21824 13524
rect 21499 13484 21824 13512
rect 21499 13481 21511 13484
rect 21453 13475 21511 13481
rect 21818 13472 21824 13484
rect 21876 13512 21882 13524
rect 22002 13512 22008 13524
rect 21876 13484 22008 13512
rect 21876 13472 21882 13484
rect 22002 13472 22008 13484
rect 22060 13472 22066 13524
rect 22557 13515 22615 13521
rect 22557 13481 22569 13515
rect 22603 13512 22615 13515
rect 23290 13512 23296 13524
rect 22603 13484 23296 13512
rect 22603 13481 22615 13484
rect 22557 13475 22615 13481
rect 23290 13472 23296 13484
rect 23348 13472 23354 13524
rect 23566 13512 23572 13524
rect 23527 13484 23572 13512
rect 23566 13472 23572 13484
rect 23624 13472 23630 13524
rect 24210 13472 24216 13524
rect 24268 13512 24274 13524
rect 24268 13484 27108 13512
rect 24268 13472 24274 13484
rect 26973 13447 27031 13453
rect 6886 13416 23244 13444
rect 1578 13336 1584 13388
rect 1636 13376 1642 13388
rect 6886 13376 6914 13416
rect 19150 13376 19156 13388
rect 1636 13348 6914 13376
rect 18432 13348 19156 13376
rect 1636 13336 1642 13348
rect 2038 13308 2044 13320
rect 1999 13280 2044 13308
rect 2038 13268 2044 13280
rect 2096 13268 2102 13320
rect 18432 13317 18460 13348
rect 19150 13336 19156 13348
rect 19208 13336 19214 13388
rect 19245 13379 19303 13385
rect 19245 13345 19257 13379
rect 19291 13376 19303 13379
rect 19334 13376 19340 13388
rect 19291 13348 19340 13376
rect 19291 13345 19303 13348
rect 19245 13339 19303 13345
rect 19334 13336 19340 13348
rect 19392 13336 19398 13388
rect 21361 13379 21419 13385
rect 21361 13345 21373 13379
rect 21407 13376 21419 13379
rect 21634 13376 21640 13388
rect 21407 13348 21640 13376
rect 21407 13345 21419 13348
rect 21361 13339 21419 13345
rect 21634 13336 21640 13348
rect 21692 13336 21698 13388
rect 22278 13336 22284 13388
rect 22336 13376 22342 13388
rect 22336 13348 22600 13376
rect 22336 13336 22342 13348
rect 18325 13311 18383 13317
rect 18325 13277 18337 13311
rect 18371 13277 18383 13311
rect 18325 13271 18383 13277
rect 18417 13311 18475 13317
rect 18417 13277 18429 13311
rect 18463 13277 18475 13311
rect 18417 13271 18475 13277
rect 18046 13172 18052 13184
rect 18007 13144 18052 13172
rect 18046 13132 18052 13144
rect 18104 13132 18110 13184
rect 18340 13172 18368 13271
rect 18506 13268 18512 13320
rect 18564 13308 18570 13320
rect 18693 13311 18751 13317
rect 18564 13280 18609 13308
rect 18564 13268 18570 13280
rect 18693 13277 18705 13311
rect 18739 13277 18751 13311
rect 18693 13271 18751 13277
rect 18708 13240 18736 13271
rect 19426 13268 19432 13320
rect 19484 13308 19490 13320
rect 19521 13311 19579 13317
rect 19521 13308 19533 13311
rect 19484 13280 19533 13308
rect 19484 13268 19490 13280
rect 19521 13277 19533 13280
rect 19567 13277 19579 13311
rect 19521 13271 19579 13277
rect 21269 13311 21327 13317
rect 21269 13277 21281 13311
rect 21315 13308 21327 13311
rect 22002 13308 22008 13320
rect 21315 13280 22008 13308
rect 21315 13277 21327 13280
rect 21269 13271 21327 13277
rect 22002 13268 22008 13280
rect 22060 13268 22066 13320
rect 22094 13268 22100 13320
rect 22152 13308 22158 13320
rect 22370 13308 22376 13320
rect 22152 13280 22197 13308
rect 22331 13280 22376 13308
rect 22152 13268 22158 13280
rect 22370 13268 22376 13280
rect 22428 13268 22434 13320
rect 22572 13317 22600 13348
rect 22557 13311 22615 13317
rect 22557 13277 22569 13311
rect 22603 13277 22615 13311
rect 23216 13308 23244 13416
rect 26973 13413 26985 13447
rect 27019 13413 27031 13447
rect 27080 13444 27108 13484
rect 27430 13472 27436 13524
rect 27488 13512 27494 13524
rect 28997 13515 29055 13521
rect 28997 13512 29009 13515
rect 27488 13484 29009 13512
rect 27488 13472 27494 13484
rect 28997 13481 29009 13484
rect 29043 13481 29055 13515
rect 28997 13475 29055 13481
rect 30558 13472 30564 13524
rect 30616 13512 30622 13524
rect 31662 13512 31668 13524
rect 30616 13484 31668 13512
rect 30616 13472 30622 13484
rect 31662 13472 31668 13484
rect 31720 13512 31726 13524
rect 31757 13515 31815 13521
rect 31757 13512 31769 13515
rect 31720 13484 31769 13512
rect 31720 13472 31726 13484
rect 31757 13481 31769 13484
rect 31803 13481 31815 13515
rect 31757 13475 31815 13481
rect 27080 13416 31754 13444
rect 26973 13407 27031 13413
rect 23290 13336 23296 13388
rect 23348 13376 23354 13388
rect 23842 13376 23848 13388
rect 23348 13348 23848 13376
rect 23348 13336 23354 13348
rect 23842 13336 23848 13348
rect 23900 13376 23906 13388
rect 24857 13379 24915 13385
rect 24857 13376 24869 13379
rect 23900 13348 24869 13376
rect 23900 13336 23906 13348
rect 24857 13345 24869 13348
rect 24903 13345 24915 13379
rect 24857 13339 24915 13345
rect 24949 13379 25007 13385
rect 24949 13345 24961 13379
rect 24995 13345 25007 13379
rect 24949 13339 25007 13345
rect 23385 13311 23443 13317
rect 23216 13280 23336 13308
rect 22557 13271 22615 13277
rect 19334 13240 19340 13252
rect 18708 13212 19340 13240
rect 19334 13200 19340 13212
rect 19392 13200 19398 13252
rect 22186 13240 22192 13252
rect 19444 13212 22192 13240
rect 19444 13172 19472 13212
rect 22186 13200 22192 13212
rect 22244 13200 22250 13252
rect 23201 13243 23259 13249
rect 23201 13209 23213 13243
rect 23247 13209 23259 13243
rect 23308 13240 23336 13280
rect 23385 13277 23397 13311
rect 23431 13308 23443 13311
rect 24762 13308 24768 13320
rect 23431 13280 24768 13308
rect 23431 13277 23443 13280
rect 23385 13271 23443 13277
rect 24762 13268 24768 13280
rect 24820 13268 24826 13320
rect 24210 13240 24216 13252
rect 23308 13212 24216 13240
rect 23201 13203 23259 13209
rect 18340 13144 19472 13172
rect 21637 13175 21695 13181
rect 21637 13141 21649 13175
rect 21683 13172 21695 13175
rect 22646 13172 22652 13184
rect 21683 13144 22652 13172
rect 21683 13141 21695 13144
rect 21637 13135 21695 13141
rect 22646 13132 22652 13144
rect 22704 13132 22710 13184
rect 22741 13175 22799 13181
rect 22741 13141 22753 13175
rect 22787 13172 22799 13175
rect 23216 13172 23244 13203
rect 24210 13200 24216 13212
rect 24268 13200 24274 13252
rect 24578 13200 24584 13252
rect 24636 13240 24642 13252
rect 24964 13240 24992 13339
rect 26142 13336 26148 13388
rect 26200 13376 26206 13388
rect 26513 13379 26571 13385
rect 26513 13376 26525 13379
rect 26200 13348 26525 13376
rect 26200 13336 26206 13348
rect 26513 13345 26525 13348
rect 26559 13345 26571 13379
rect 26988 13376 27016 13407
rect 27709 13379 27767 13385
rect 26988 13348 27660 13376
rect 26513 13339 26571 13345
rect 26234 13268 26240 13320
rect 26292 13308 26298 13320
rect 26605 13311 26663 13317
rect 26605 13308 26617 13311
rect 26292 13280 26617 13308
rect 26292 13268 26298 13280
rect 26605 13277 26617 13280
rect 26651 13277 26663 13311
rect 27430 13308 27436 13320
rect 27391 13280 27436 13308
rect 26605 13271 26663 13277
rect 27430 13268 27436 13280
rect 27488 13268 27494 13320
rect 27632 13317 27660 13348
rect 27709 13345 27721 13379
rect 27755 13345 27767 13379
rect 27709 13339 27767 13345
rect 27801 13379 27859 13385
rect 27801 13345 27813 13379
rect 27847 13376 27859 13379
rect 28166 13376 28172 13388
rect 27847 13348 28172 13376
rect 27847 13345 27859 13348
rect 27801 13339 27859 13345
rect 27617 13311 27675 13317
rect 27617 13277 27629 13311
rect 27663 13277 27675 13311
rect 27617 13271 27675 13277
rect 24636 13212 24992 13240
rect 24636 13200 24642 13212
rect 24394 13172 24400 13184
rect 22787 13144 23244 13172
rect 24355 13144 24400 13172
rect 22787 13141 22799 13144
rect 22741 13135 22799 13141
rect 24394 13132 24400 13144
rect 24452 13132 24458 13184
rect 24486 13132 24492 13184
rect 24544 13172 24550 13184
rect 24765 13175 24823 13181
rect 24765 13172 24777 13175
rect 24544 13144 24777 13172
rect 24544 13132 24550 13144
rect 24765 13141 24777 13144
rect 24811 13141 24823 13175
rect 24765 13135 24823 13141
rect 27614 13132 27620 13184
rect 27672 13172 27678 13184
rect 27724 13172 27752 13339
rect 28166 13336 28172 13348
rect 28224 13336 28230 13388
rect 30653 13379 30711 13385
rect 30653 13345 30665 13379
rect 30699 13376 30711 13379
rect 31110 13376 31116 13388
rect 30699 13348 31116 13376
rect 30699 13345 30711 13348
rect 30653 13339 30711 13345
rect 31110 13336 31116 13348
rect 31168 13336 31174 13388
rect 31726 13376 31754 13416
rect 31846 13376 31852 13388
rect 31726 13348 31852 13376
rect 31846 13336 31852 13348
rect 31904 13336 31910 13388
rect 32306 13376 32312 13388
rect 32267 13348 32312 13376
rect 32306 13336 32312 13348
rect 32364 13336 32370 13388
rect 32490 13376 32496 13388
rect 32451 13348 32496 13376
rect 32490 13336 32496 13348
rect 32548 13336 32554 13388
rect 33686 13376 33692 13388
rect 33647 13348 33692 13376
rect 33686 13336 33692 13348
rect 33744 13336 33750 13388
rect 34146 13336 34152 13388
rect 34204 13376 34210 13388
rect 34701 13379 34759 13385
rect 34701 13376 34713 13379
rect 34204 13348 34713 13376
rect 34204 13336 34210 13348
rect 34701 13345 34713 13348
rect 34747 13345 34759 13379
rect 34701 13339 34759 13345
rect 27982 13308 27988 13320
rect 27943 13280 27988 13308
rect 27982 13268 27988 13280
rect 28040 13268 28046 13320
rect 30006 13268 30012 13320
rect 30064 13308 30070 13320
rect 30469 13311 30527 13317
rect 30469 13308 30481 13311
rect 30064 13280 30481 13308
rect 30064 13268 30070 13280
rect 30469 13277 30481 13280
rect 30515 13277 30527 13311
rect 30469 13271 30527 13277
rect 31665 13311 31723 13317
rect 31665 13277 31677 13311
rect 31711 13308 31723 13311
rect 32214 13308 32220 13320
rect 31711 13280 32220 13308
rect 31711 13277 31723 13280
rect 31665 13271 31723 13277
rect 32214 13268 32220 13280
rect 32272 13268 32278 13320
rect 28534 13200 28540 13252
rect 28592 13240 28598 13252
rect 28629 13243 28687 13249
rect 28629 13240 28641 13243
rect 28592 13212 28641 13240
rect 28592 13200 28598 13212
rect 28629 13209 28641 13212
rect 28675 13209 28687 13243
rect 28629 13203 28687 13209
rect 28718 13200 28724 13252
rect 28776 13240 28782 13252
rect 28813 13243 28871 13249
rect 28813 13240 28825 13243
rect 28776 13212 28825 13240
rect 28776 13200 28782 13212
rect 28813 13209 28825 13212
rect 28859 13240 28871 13243
rect 31570 13240 31576 13252
rect 28859 13212 31576 13240
rect 28859 13209 28871 13212
rect 28813 13203 28871 13209
rect 31570 13200 31576 13212
rect 31628 13240 31634 13252
rect 31628 13212 31754 13240
rect 31628 13200 31634 13212
rect 28166 13172 28172 13184
rect 27672 13144 27752 13172
rect 28127 13144 28172 13172
rect 27672 13132 27678 13144
rect 28166 13132 28172 13144
rect 28224 13132 28230 13184
rect 31726 13172 31754 13212
rect 34698 13200 34704 13252
rect 34756 13240 34762 13252
rect 34946 13243 35004 13249
rect 34946 13240 34958 13243
rect 34756 13212 34958 13240
rect 34756 13200 34762 13212
rect 34946 13209 34958 13212
rect 34992 13209 35004 13243
rect 34946 13203 35004 13209
rect 35342 13172 35348 13184
rect 31726 13144 35348 13172
rect 35342 13132 35348 13144
rect 35400 13172 35406 13184
rect 36081 13175 36139 13181
rect 36081 13172 36093 13175
rect 35400 13144 36093 13172
rect 35400 13132 35406 13144
rect 36081 13141 36093 13144
rect 36127 13141 36139 13175
rect 36081 13135 36139 13141
rect 1104 13082 48852 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 48852 13082
rect 1104 13008 48852 13030
rect 1578 12968 1584 12980
rect 1539 12940 1584 12968
rect 1578 12928 1584 12940
rect 1636 12928 1642 12980
rect 2038 12928 2044 12980
rect 2096 12968 2102 12980
rect 18598 12968 18604 12980
rect 2096 12940 18604 12968
rect 2096 12928 2102 12940
rect 18598 12928 18604 12940
rect 18656 12928 18662 12980
rect 21634 12928 21640 12980
rect 21692 12928 21698 12980
rect 24302 12928 24308 12980
rect 24360 12968 24366 12980
rect 26237 12971 26295 12977
rect 26237 12968 26249 12971
rect 24360 12940 26249 12968
rect 24360 12928 24366 12940
rect 26237 12937 26249 12940
rect 26283 12937 26295 12971
rect 26237 12931 26295 12937
rect 27982 12928 27988 12980
rect 28040 12968 28046 12980
rect 28810 12968 28816 12980
rect 28040 12940 28816 12968
rect 28040 12928 28046 12940
rect 28810 12928 28816 12940
rect 28868 12968 28874 12980
rect 29641 12971 29699 12977
rect 29641 12968 29653 12971
rect 28868 12940 29653 12968
rect 28868 12928 28874 12940
rect 29641 12937 29653 12940
rect 29687 12937 29699 12971
rect 29641 12931 29699 12937
rect 16850 12900 16856 12912
rect 16811 12872 16856 12900
rect 16850 12860 16856 12872
rect 16908 12860 16914 12912
rect 18138 12860 18144 12912
rect 18196 12900 18202 12912
rect 21652 12900 21680 12928
rect 25041 12903 25099 12909
rect 18196 12872 20668 12900
rect 21652 12872 22324 12900
rect 18196 12860 18202 12872
rect 1394 12832 1400 12844
rect 1355 12804 1400 12832
rect 1394 12792 1400 12804
rect 1452 12792 1458 12844
rect 19150 12792 19156 12844
rect 19208 12832 19214 12844
rect 20640 12841 20668 12872
rect 20625 12835 20683 12841
rect 19208 12804 19656 12832
rect 19208 12792 19214 12804
rect 3510 12724 3516 12776
rect 3568 12764 3574 12776
rect 16666 12764 16672 12776
rect 3568 12736 6914 12764
rect 16627 12736 16672 12764
rect 3568 12724 3574 12736
rect 6886 12696 6914 12736
rect 16666 12724 16672 12736
rect 16724 12724 16730 12776
rect 17129 12767 17187 12773
rect 17129 12733 17141 12767
rect 17175 12733 17187 12767
rect 17129 12727 17187 12733
rect 17144 12696 17172 12727
rect 18966 12724 18972 12776
rect 19024 12764 19030 12776
rect 19628 12773 19656 12804
rect 20625 12801 20637 12835
rect 20671 12801 20683 12835
rect 20625 12795 20683 12801
rect 21634 12792 21640 12844
rect 21692 12832 21698 12844
rect 22002 12832 22008 12844
rect 21692 12804 22008 12832
rect 21692 12792 21698 12804
rect 22002 12792 22008 12804
rect 22060 12792 22066 12844
rect 22296 12841 22324 12872
rect 25041 12869 25053 12903
rect 25087 12900 25099 12903
rect 25498 12900 25504 12912
rect 25087 12872 25504 12900
rect 25087 12869 25099 12872
rect 25041 12863 25099 12869
rect 25498 12860 25504 12872
rect 25556 12860 25562 12912
rect 26145 12903 26203 12909
rect 26145 12869 26157 12903
rect 26191 12900 26203 12903
rect 29086 12900 29092 12912
rect 26191 12872 29092 12900
rect 26191 12869 26203 12872
rect 26145 12863 26203 12869
rect 29086 12860 29092 12872
rect 29144 12860 29150 12912
rect 32030 12900 32036 12912
rect 30392 12872 32036 12900
rect 22281 12835 22339 12841
rect 22281 12801 22293 12835
rect 22327 12801 22339 12835
rect 22281 12795 22339 12801
rect 22646 12792 22652 12844
rect 22704 12832 22710 12844
rect 23109 12835 23167 12841
rect 23109 12832 23121 12835
rect 22704 12804 23121 12832
rect 22704 12792 22710 12804
rect 23109 12801 23121 12804
rect 23155 12832 23167 12835
rect 25317 12835 25375 12841
rect 25317 12832 25329 12835
rect 23155 12804 25329 12832
rect 23155 12801 23167 12804
rect 23109 12795 23167 12801
rect 25317 12801 25329 12804
rect 25363 12801 25375 12835
rect 25317 12795 25375 12801
rect 26234 12792 26240 12844
rect 26292 12832 26298 12844
rect 26973 12835 27031 12841
rect 26973 12832 26985 12835
rect 26292 12804 26985 12832
rect 26292 12792 26298 12804
rect 26973 12801 26985 12804
rect 27019 12801 27031 12835
rect 26973 12795 27031 12801
rect 28166 12792 28172 12844
rect 28224 12832 28230 12844
rect 30392 12841 30420 12872
rect 32030 12860 32036 12872
rect 32088 12860 32094 12912
rect 34514 12860 34520 12912
rect 34572 12900 34578 12912
rect 34670 12903 34728 12909
rect 34670 12900 34682 12903
rect 34572 12872 34682 12900
rect 34572 12860 34578 12872
rect 34670 12869 34682 12872
rect 34716 12869 34728 12903
rect 34670 12863 34728 12869
rect 28517 12835 28575 12841
rect 28517 12832 28529 12835
rect 28224 12804 28529 12832
rect 28224 12792 28230 12804
rect 28517 12801 28529 12804
rect 28563 12801 28575 12835
rect 28517 12795 28575 12801
rect 30377 12835 30435 12841
rect 30377 12801 30389 12835
rect 30423 12801 30435 12835
rect 30377 12795 30435 12801
rect 31662 12792 31668 12844
rect 31720 12832 31726 12844
rect 32125 12835 32183 12841
rect 32125 12832 32137 12835
rect 31720 12804 32137 12832
rect 31720 12792 31726 12804
rect 32125 12801 32137 12804
rect 32171 12801 32183 12835
rect 32125 12795 32183 12801
rect 32214 12792 32220 12844
rect 32272 12832 32278 12844
rect 32381 12835 32439 12841
rect 32381 12832 32393 12835
rect 32272 12804 32393 12832
rect 32272 12792 32278 12804
rect 32381 12801 32393 12804
rect 32427 12801 32439 12835
rect 32381 12795 32439 12801
rect 34146 12792 34152 12844
rect 34204 12832 34210 12844
rect 34425 12835 34483 12841
rect 34425 12832 34437 12835
rect 34204 12804 34437 12832
rect 34204 12792 34210 12804
rect 34425 12801 34437 12804
rect 34471 12801 34483 12835
rect 34425 12795 34483 12801
rect 19337 12767 19395 12773
rect 19337 12764 19349 12767
rect 19024 12736 19349 12764
rect 19024 12724 19030 12736
rect 19337 12733 19349 12736
rect 19383 12733 19395 12767
rect 19337 12727 19395 12733
rect 19613 12767 19671 12773
rect 19613 12733 19625 12767
rect 19659 12764 19671 12767
rect 20254 12764 20260 12776
rect 19659 12736 20260 12764
rect 19659 12733 19671 12736
rect 19613 12727 19671 12733
rect 20254 12724 20260 12736
rect 20312 12724 20318 12776
rect 21818 12724 21824 12776
rect 21876 12764 21882 12776
rect 22189 12767 22247 12773
rect 22189 12764 22201 12767
rect 21876 12736 22201 12764
rect 21876 12724 21882 12736
rect 22189 12733 22201 12736
rect 22235 12733 22247 12767
rect 22189 12727 22247 12733
rect 22830 12724 22836 12776
rect 22888 12764 22894 12776
rect 23385 12767 23443 12773
rect 23385 12764 23397 12767
rect 22888 12736 23397 12764
rect 22888 12724 22894 12736
rect 23385 12733 23397 12736
rect 23431 12764 23443 12767
rect 24854 12764 24860 12776
rect 23431 12736 24860 12764
rect 23431 12733 23443 12736
rect 23385 12727 23443 12733
rect 24854 12724 24860 12736
rect 24912 12724 24918 12776
rect 25225 12767 25283 12773
rect 25225 12733 25237 12767
rect 25271 12764 25283 12767
rect 25682 12764 25688 12776
rect 25271 12736 25688 12764
rect 25271 12733 25283 12736
rect 25225 12727 25283 12733
rect 25682 12724 25688 12736
rect 25740 12724 25746 12776
rect 26694 12724 26700 12776
rect 26752 12764 26758 12776
rect 27249 12767 27307 12773
rect 27249 12764 27261 12767
rect 26752 12736 27261 12764
rect 26752 12724 26758 12736
rect 27249 12733 27261 12736
rect 27295 12733 27307 12767
rect 27249 12727 27307 12733
rect 28261 12767 28319 12773
rect 28261 12733 28273 12767
rect 28307 12733 28319 12767
rect 28261 12727 28319 12733
rect 30653 12767 30711 12773
rect 30653 12733 30665 12767
rect 30699 12764 30711 12767
rect 30699 12736 31754 12764
rect 30699 12733 30711 12736
rect 30653 12727 30711 12733
rect 6886 12668 17172 12696
rect 20622 12656 20628 12708
rect 20680 12696 20686 12708
rect 20898 12696 20904 12708
rect 20680 12668 20904 12696
rect 20680 12656 20686 12668
rect 20898 12656 20904 12668
rect 20956 12656 20962 12708
rect 23198 12696 23204 12708
rect 22066 12668 23204 12696
rect 19426 12588 19432 12640
rect 19484 12628 19490 12640
rect 19702 12628 19708 12640
rect 19484 12600 19708 12628
rect 19484 12588 19490 12600
rect 19702 12588 19708 12600
rect 19760 12588 19766 12640
rect 20714 12628 20720 12640
rect 20675 12600 20720 12628
rect 20714 12588 20720 12600
rect 20772 12588 20778 12640
rect 21821 12631 21879 12637
rect 21821 12597 21833 12631
rect 21867 12628 21879 12631
rect 22066 12628 22094 12668
rect 23198 12656 23204 12668
rect 23256 12656 23262 12708
rect 24946 12656 24952 12708
rect 25004 12696 25010 12708
rect 28276 12696 28304 12727
rect 25004 12668 28304 12696
rect 31726 12696 31754 12736
rect 32122 12696 32128 12708
rect 31726 12668 32128 12696
rect 25004 12656 25010 12668
rect 32122 12656 32128 12668
rect 32180 12656 32186 12708
rect 21867 12600 22094 12628
rect 21867 12597 21879 12600
rect 21821 12591 21879 12597
rect 24394 12588 24400 12640
rect 24452 12628 24458 12640
rect 24578 12628 24584 12640
rect 24452 12600 24584 12628
rect 24452 12588 24458 12600
rect 24578 12588 24584 12600
rect 24636 12628 24642 12640
rect 25041 12631 25099 12637
rect 25041 12628 25053 12631
rect 24636 12600 25053 12628
rect 24636 12588 24642 12600
rect 25041 12597 25053 12600
rect 25087 12597 25099 12631
rect 25041 12591 25099 12597
rect 25406 12588 25412 12640
rect 25464 12628 25470 12640
rect 25501 12631 25559 12637
rect 25501 12628 25513 12631
rect 25464 12600 25513 12628
rect 25464 12588 25470 12600
rect 25501 12597 25513 12600
rect 25547 12597 25559 12631
rect 25501 12591 25559 12597
rect 26786 12588 26792 12640
rect 26844 12628 26850 12640
rect 27065 12631 27123 12637
rect 27065 12628 27077 12631
rect 26844 12600 27077 12628
rect 26844 12588 26850 12600
rect 27065 12597 27077 12600
rect 27111 12597 27123 12631
rect 27065 12591 27123 12597
rect 27246 12588 27252 12640
rect 27304 12628 27310 12640
rect 27525 12631 27583 12637
rect 27525 12628 27537 12631
rect 27304 12600 27537 12628
rect 27304 12588 27310 12600
rect 27525 12597 27537 12600
rect 27571 12597 27583 12631
rect 27525 12591 27583 12597
rect 27614 12588 27620 12640
rect 27672 12628 27678 12640
rect 28258 12628 28264 12640
rect 27672 12600 28264 12628
rect 27672 12588 27678 12600
rect 28258 12588 28264 12600
rect 28316 12588 28322 12640
rect 32306 12588 32312 12640
rect 32364 12628 32370 12640
rect 33505 12631 33563 12637
rect 33505 12628 33517 12631
rect 32364 12600 33517 12628
rect 32364 12588 32370 12600
rect 33505 12597 33517 12600
rect 33551 12597 33563 12631
rect 33505 12591 33563 12597
rect 35618 12588 35624 12640
rect 35676 12628 35682 12640
rect 35805 12631 35863 12637
rect 35805 12628 35817 12631
rect 35676 12600 35817 12628
rect 35676 12588 35682 12600
rect 35805 12597 35817 12600
rect 35851 12597 35863 12631
rect 35805 12591 35863 12597
rect 1104 12538 48852 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 48852 12538
rect 1104 12464 48852 12486
rect 16666 12384 16672 12436
rect 16724 12424 16730 12436
rect 17865 12427 17923 12433
rect 17865 12424 17877 12427
rect 16724 12396 17877 12424
rect 16724 12384 16730 12396
rect 17865 12393 17877 12396
rect 17911 12393 17923 12427
rect 17865 12387 17923 12393
rect 17880 12288 17908 12387
rect 18506 12384 18512 12436
rect 18564 12424 18570 12436
rect 18693 12427 18751 12433
rect 18693 12424 18705 12427
rect 18564 12396 18705 12424
rect 18564 12384 18570 12396
rect 18693 12393 18705 12396
rect 18739 12393 18751 12427
rect 18693 12387 18751 12393
rect 20714 12384 20720 12436
rect 20772 12384 20778 12436
rect 21634 12424 21640 12436
rect 21595 12396 21640 12424
rect 21634 12384 21640 12396
rect 21692 12384 21698 12436
rect 22922 12424 22928 12436
rect 22883 12396 22928 12424
rect 22922 12384 22928 12396
rect 22980 12384 22986 12436
rect 24578 12384 24584 12436
rect 24636 12424 24642 12436
rect 25317 12427 25375 12433
rect 25317 12424 25329 12427
rect 24636 12396 25329 12424
rect 24636 12384 24642 12396
rect 25317 12393 25329 12396
rect 25363 12393 25375 12427
rect 25317 12387 25375 12393
rect 25777 12427 25835 12433
rect 25777 12393 25789 12427
rect 25823 12424 25835 12427
rect 26234 12424 26240 12436
rect 25823 12396 26240 12424
rect 25823 12393 25835 12396
rect 25777 12387 25835 12393
rect 26234 12384 26240 12396
rect 26292 12384 26298 12436
rect 31297 12427 31355 12433
rect 31297 12393 31309 12427
rect 31343 12424 31355 12427
rect 32214 12424 32220 12436
rect 31343 12396 32220 12424
rect 31343 12393 31355 12396
rect 31297 12387 31355 12393
rect 32214 12384 32220 12396
rect 32272 12384 32278 12436
rect 34698 12424 34704 12436
rect 34659 12396 34704 12424
rect 34698 12384 34704 12396
rect 34756 12384 34762 12436
rect 44726 12384 44732 12436
rect 44784 12424 44790 12436
rect 46842 12424 46848 12436
rect 44784 12396 46848 12424
rect 44784 12384 44790 12396
rect 46842 12384 46848 12396
rect 46900 12384 46906 12436
rect 19242 12316 19248 12368
rect 19300 12356 19306 12368
rect 20346 12356 20352 12368
rect 19300 12328 20352 12356
rect 19300 12316 19306 12328
rect 20346 12316 20352 12328
rect 20404 12316 20410 12368
rect 19429 12291 19487 12297
rect 17880 12260 18552 12288
rect 16485 12223 16543 12229
rect 16485 12189 16497 12223
rect 16531 12220 16543 12223
rect 17954 12220 17960 12232
rect 16531 12192 17960 12220
rect 16531 12189 16543 12192
rect 16485 12183 16543 12189
rect 17954 12180 17960 12192
rect 18012 12180 18018 12232
rect 18524 12229 18552 12260
rect 19429 12257 19441 12291
rect 19475 12288 19487 12291
rect 20732 12288 20760 12384
rect 29270 12356 29276 12368
rect 19475 12260 20760 12288
rect 20824 12328 29276 12356
rect 19475 12257 19487 12260
rect 19429 12251 19487 12257
rect 18509 12223 18567 12229
rect 18509 12189 18521 12223
rect 18555 12189 18567 12223
rect 18509 12183 18567 12189
rect 19150 12180 19156 12232
rect 19208 12220 19214 12232
rect 19245 12223 19303 12229
rect 19245 12220 19257 12223
rect 19208 12192 19257 12220
rect 19208 12180 19214 12192
rect 19245 12189 19257 12192
rect 19291 12189 19303 12223
rect 19245 12183 19303 12189
rect 16752 12155 16810 12161
rect 16752 12121 16764 12155
rect 16798 12152 16810 12155
rect 18046 12152 18052 12164
rect 16798 12124 18052 12152
rect 16798 12121 16810 12124
rect 16752 12115 16810 12121
rect 18046 12112 18052 12124
rect 18104 12112 18110 12164
rect 18325 12155 18383 12161
rect 18325 12121 18337 12155
rect 18371 12152 18383 12155
rect 19702 12152 19708 12164
rect 18371 12124 19708 12152
rect 18371 12121 18383 12124
rect 18325 12115 18383 12121
rect 19352 12096 19380 12124
rect 19702 12112 19708 12124
rect 19760 12112 19766 12164
rect 20346 12112 20352 12164
rect 20404 12152 20410 12164
rect 20824 12152 20852 12328
rect 29270 12316 29276 12328
rect 29328 12316 29334 12368
rect 22281 12291 22339 12297
rect 22281 12257 22293 12291
rect 22327 12288 22339 12291
rect 23566 12288 23572 12300
rect 22327 12260 23572 12288
rect 22327 12257 22339 12260
rect 22281 12251 22339 12257
rect 23566 12248 23572 12260
rect 23624 12248 23630 12300
rect 27338 12248 27344 12300
rect 27396 12288 27402 12300
rect 27801 12291 27859 12297
rect 27801 12288 27813 12291
rect 27396 12260 27813 12288
rect 27396 12248 27402 12260
rect 27801 12257 27813 12260
rect 27847 12257 27859 12291
rect 32769 12291 32827 12297
rect 32769 12288 32781 12291
rect 27801 12251 27859 12257
rect 31772 12260 32781 12288
rect 22094 12180 22100 12232
rect 22152 12220 22158 12232
rect 22370 12220 22376 12232
rect 22152 12192 22376 12220
rect 22152 12180 22158 12192
rect 22370 12180 22376 12192
rect 22428 12180 22434 12232
rect 22830 12220 22836 12232
rect 22791 12192 22836 12220
rect 22830 12180 22836 12192
rect 22888 12180 22894 12232
rect 23201 12223 23259 12229
rect 23201 12189 23213 12223
rect 23247 12220 23259 12223
rect 23290 12220 23296 12232
rect 23247 12192 23296 12220
rect 23247 12189 23259 12192
rect 23201 12183 23259 12189
rect 23290 12180 23296 12192
rect 23348 12180 23354 12232
rect 23750 12180 23756 12232
rect 23808 12220 23814 12232
rect 24673 12223 24731 12229
rect 24673 12220 24685 12223
rect 23808 12192 24685 12220
rect 23808 12180 23814 12192
rect 24673 12189 24685 12192
rect 24719 12189 24731 12223
rect 24673 12183 24731 12189
rect 24857 12223 24915 12229
rect 24857 12189 24869 12223
rect 24903 12220 24915 12223
rect 24946 12220 24952 12232
rect 24903 12192 24952 12220
rect 24903 12189 24915 12192
rect 24857 12183 24915 12189
rect 24946 12180 24952 12192
rect 25004 12180 25010 12232
rect 25148 12192 25452 12220
rect 20404 12124 20852 12152
rect 21085 12155 21143 12161
rect 20404 12112 20410 12124
rect 21085 12121 21097 12155
rect 21131 12152 21143 12155
rect 25148 12152 25176 12192
rect 25314 12152 25320 12164
rect 21131 12124 25176 12152
rect 25227 12124 25320 12152
rect 21131 12121 21143 12124
rect 21085 12115 21143 12121
rect 25314 12112 25320 12124
rect 25372 12112 25378 12164
rect 25424 12152 25452 12192
rect 25498 12180 25504 12232
rect 25556 12220 25562 12232
rect 25633 12223 25691 12229
rect 25556 12192 25601 12220
rect 25556 12180 25562 12192
rect 25633 12189 25645 12223
rect 25679 12220 25691 12223
rect 25774 12220 25780 12232
rect 25679 12192 25780 12220
rect 25679 12189 25691 12192
rect 25633 12183 25691 12189
rect 25774 12180 25780 12192
rect 25832 12180 25838 12232
rect 27614 12180 27620 12232
rect 27672 12220 27678 12232
rect 27709 12223 27767 12229
rect 27709 12220 27721 12223
rect 27672 12192 27721 12220
rect 27672 12180 27678 12192
rect 27709 12189 27721 12192
rect 27755 12220 27767 12223
rect 28626 12220 28632 12232
rect 27755 12192 28632 12220
rect 27755 12189 27767 12192
rect 27709 12183 27767 12189
rect 28626 12180 28632 12192
rect 28684 12180 28690 12232
rect 30469 12223 30527 12229
rect 30469 12189 30481 12223
rect 30515 12220 30527 12223
rect 30834 12220 30840 12232
rect 30515 12192 30840 12220
rect 30515 12189 30527 12192
rect 30469 12183 30527 12189
rect 30834 12180 30840 12192
rect 30892 12180 30898 12232
rect 31570 12220 31576 12232
rect 31531 12192 31576 12220
rect 31570 12180 31576 12192
rect 31628 12180 31634 12232
rect 31772 12229 31800 12260
rect 32769 12257 32781 12260
rect 32815 12257 32827 12291
rect 32769 12251 32827 12257
rect 34422 12248 34428 12300
rect 34480 12288 34486 12300
rect 35802 12288 35808 12300
rect 34480 12260 35112 12288
rect 34480 12248 34486 12260
rect 31665 12223 31723 12229
rect 31665 12189 31677 12223
rect 31711 12189 31723 12223
rect 31665 12183 31723 12189
rect 31757 12223 31815 12229
rect 31757 12189 31769 12223
rect 31803 12189 31815 12223
rect 31757 12183 31815 12189
rect 31941 12223 31999 12229
rect 31941 12189 31953 12223
rect 31987 12189 31999 12223
rect 31941 12183 31999 12189
rect 28258 12152 28264 12164
rect 25424 12124 28264 12152
rect 28258 12112 28264 12124
rect 28316 12112 28322 12164
rect 30653 12155 30711 12161
rect 30653 12121 30665 12155
rect 30699 12152 30711 12155
rect 31294 12152 31300 12164
rect 30699 12124 31300 12152
rect 30699 12121 30711 12124
rect 30653 12115 30711 12121
rect 31294 12112 31300 12124
rect 31352 12152 31358 12164
rect 31680 12152 31708 12183
rect 31352 12124 31708 12152
rect 31352 12112 31358 12124
rect 19334 12044 19340 12096
rect 19392 12044 19398 12096
rect 22005 12087 22063 12093
rect 22005 12053 22017 12087
rect 22051 12084 22063 12087
rect 22370 12084 22376 12096
rect 22051 12056 22376 12084
rect 22051 12053 22063 12056
rect 22005 12047 22063 12053
rect 22370 12044 22376 12056
rect 22428 12044 22434 12096
rect 23382 12084 23388 12096
rect 23343 12056 23388 12084
rect 23382 12044 23388 12056
rect 23440 12044 23446 12096
rect 25332 12084 25360 12112
rect 25682 12084 25688 12096
rect 25332 12056 25688 12084
rect 25682 12044 25688 12056
rect 25740 12084 25746 12096
rect 27249 12087 27307 12093
rect 27249 12084 27261 12087
rect 25740 12056 27261 12084
rect 25740 12044 25746 12056
rect 27249 12053 27261 12056
rect 27295 12053 27307 12087
rect 27249 12047 27307 12053
rect 27617 12087 27675 12093
rect 27617 12053 27629 12087
rect 27663 12084 27675 12087
rect 28166 12084 28172 12096
rect 27663 12056 28172 12084
rect 27663 12053 27675 12056
rect 27617 12047 27675 12053
rect 28166 12044 28172 12056
rect 28224 12044 28230 12096
rect 31956 12084 31984 12183
rect 32306 12180 32312 12232
rect 32364 12220 32370 12232
rect 32585 12223 32643 12229
rect 32585 12220 32597 12223
rect 32364 12192 32597 12220
rect 32364 12180 32370 12192
rect 32585 12189 32597 12192
rect 32631 12189 32643 12223
rect 32585 12183 32643 12189
rect 32674 12180 32680 12232
rect 32732 12220 32738 12232
rect 33229 12223 33287 12229
rect 33229 12220 33241 12223
rect 32732 12192 33241 12220
rect 32732 12180 32738 12192
rect 33229 12189 33241 12192
rect 33275 12220 33287 12223
rect 33318 12220 33324 12232
rect 33275 12192 33324 12220
rect 33275 12189 33287 12192
rect 33229 12183 33287 12189
rect 33318 12180 33324 12192
rect 33376 12180 33382 12232
rect 35084 12229 35112 12260
rect 35176 12260 35808 12288
rect 35176 12229 35204 12260
rect 35802 12248 35808 12260
rect 35860 12248 35866 12300
rect 34977 12223 35035 12229
rect 34977 12189 34989 12223
rect 35023 12189 35035 12223
rect 34977 12183 35035 12189
rect 35069 12223 35127 12229
rect 35069 12189 35081 12223
rect 35115 12189 35127 12223
rect 35069 12183 35127 12189
rect 35161 12223 35219 12229
rect 35161 12189 35173 12223
rect 35207 12189 35219 12223
rect 35161 12183 35219 12189
rect 35345 12223 35403 12229
rect 35345 12189 35357 12223
rect 35391 12220 35403 12223
rect 35526 12220 35532 12232
rect 35391 12192 35532 12220
rect 35391 12189 35403 12192
rect 35345 12183 35403 12189
rect 32122 12112 32128 12164
rect 32180 12152 32186 12164
rect 32401 12155 32459 12161
rect 32401 12152 32413 12155
rect 32180 12124 32413 12152
rect 32180 12112 32186 12124
rect 32401 12121 32413 12124
rect 32447 12121 32459 12155
rect 34992 12152 35020 12183
rect 35526 12180 35532 12192
rect 35584 12180 35590 12232
rect 35894 12220 35900 12232
rect 35855 12192 35900 12220
rect 35894 12180 35900 12192
rect 35952 12220 35958 12232
rect 36170 12220 36176 12232
rect 35952 12192 36176 12220
rect 35952 12180 35958 12192
rect 36170 12180 36176 12192
rect 36228 12180 36234 12232
rect 44818 12152 44824 12164
rect 34992 12124 44824 12152
rect 32401 12115 32459 12121
rect 44818 12112 44824 12124
rect 44876 12112 44882 12164
rect 33134 12084 33140 12096
rect 31956 12056 33140 12084
rect 33134 12044 33140 12056
rect 33192 12044 33198 12096
rect 33318 12084 33324 12096
rect 33279 12056 33324 12084
rect 33318 12044 33324 12056
rect 33376 12044 33382 12096
rect 36078 12084 36084 12096
rect 36039 12056 36084 12084
rect 36078 12044 36084 12056
rect 36136 12084 36142 12096
rect 37182 12084 37188 12096
rect 36136 12056 37188 12084
rect 36136 12044 36142 12056
rect 37182 12044 37188 12056
rect 37240 12044 37246 12096
rect 1104 11994 48852 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 48852 11994
rect 1104 11920 48852 11942
rect 19150 11880 19156 11892
rect 19111 11852 19156 11880
rect 19150 11840 19156 11852
rect 19208 11840 19214 11892
rect 22186 11840 22192 11892
rect 22244 11880 22250 11892
rect 24946 11880 24952 11892
rect 22244 11852 24952 11880
rect 22244 11840 22250 11852
rect 24946 11840 24952 11852
rect 25004 11840 25010 11892
rect 25501 11883 25559 11889
rect 25501 11849 25513 11883
rect 25547 11880 25559 11883
rect 26694 11880 26700 11892
rect 25547 11852 26700 11880
rect 25547 11849 25559 11852
rect 25501 11843 25559 11849
rect 26694 11840 26700 11852
rect 26752 11840 26758 11892
rect 28626 11840 28632 11892
rect 28684 11880 28690 11892
rect 29181 11883 29239 11889
rect 29181 11880 29193 11883
rect 28684 11852 29193 11880
rect 28684 11840 28690 11852
rect 29181 11849 29193 11852
rect 29227 11849 29239 11883
rect 29181 11843 29239 11849
rect 29270 11840 29276 11892
rect 29328 11880 29334 11892
rect 36078 11880 36084 11892
rect 29328 11852 36084 11880
rect 29328 11840 29334 11852
rect 36078 11840 36084 11852
rect 36136 11840 36142 11892
rect 18040 11815 18098 11821
rect 18040 11781 18052 11815
rect 18086 11812 18098 11815
rect 19613 11815 19671 11821
rect 19613 11812 19625 11815
rect 18086 11784 19625 11812
rect 18086 11781 18098 11784
rect 18040 11775 18098 11781
rect 19613 11781 19625 11784
rect 19659 11781 19671 11815
rect 20346 11812 20352 11824
rect 19613 11775 19671 11781
rect 19720 11784 20352 11812
rect 2041 11747 2099 11753
rect 2041 11713 2053 11747
rect 2087 11744 2099 11747
rect 15930 11744 15936 11756
rect 2087 11716 15936 11744
rect 2087 11713 2099 11716
rect 2041 11707 2099 11713
rect 15930 11704 15936 11716
rect 15988 11704 15994 11756
rect 19426 11704 19432 11756
rect 19484 11744 19490 11756
rect 19720 11744 19748 11784
rect 20346 11772 20352 11784
rect 20404 11772 20410 11824
rect 23382 11812 23388 11824
rect 21836 11784 23388 11812
rect 19484 11716 19748 11744
rect 19889 11747 19947 11753
rect 19484 11704 19490 11716
rect 19889 11713 19901 11747
rect 19935 11713 19947 11747
rect 19889 11707 19947 11713
rect 19981 11747 20039 11753
rect 19981 11713 19993 11747
rect 20027 11713 20039 11747
rect 19981 11707 20039 11713
rect 17586 11636 17592 11688
rect 17644 11676 17650 11688
rect 17773 11679 17831 11685
rect 17773 11676 17785 11679
rect 17644 11648 17785 11676
rect 17644 11636 17650 11648
rect 17773 11645 17785 11648
rect 17819 11645 17831 11679
rect 17773 11639 17831 11645
rect 19904 11608 19932 11707
rect 19996 11676 20024 11707
rect 20070 11704 20076 11756
rect 20128 11744 20134 11756
rect 20257 11747 20315 11753
rect 20128 11716 20173 11744
rect 20128 11704 20134 11716
rect 20257 11713 20269 11747
rect 20303 11744 20315 11747
rect 20364 11744 20392 11772
rect 21836 11753 21864 11784
rect 23382 11772 23388 11784
rect 23440 11772 23446 11824
rect 23750 11772 23756 11824
rect 23808 11812 23814 11824
rect 24118 11812 24124 11824
rect 23808 11784 24124 11812
rect 23808 11772 23814 11784
rect 24118 11772 24124 11784
rect 24176 11772 24182 11824
rect 28166 11772 28172 11824
rect 28224 11812 28230 11824
rect 31018 11812 31024 11824
rect 28224 11784 31024 11812
rect 28224 11772 28230 11784
rect 31018 11772 31024 11784
rect 31076 11772 31082 11824
rect 32493 11815 32551 11821
rect 32493 11812 32505 11815
rect 31496 11784 32505 11812
rect 20303 11716 20392 11744
rect 21821 11747 21879 11753
rect 20303 11713 20315 11716
rect 20257 11707 20315 11713
rect 21821 11713 21833 11747
rect 21867 11713 21879 11747
rect 21821 11707 21879 11713
rect 21910 11704 21916 11756
rect 21968 11744 21974 11756
rect 22005 11747 22063 11753
rect 22005 11744 22017 11747
rect 21968 11716 22017 11744
rect 21968 11704 21974 11716
rect 22005 11713 22017 11716
rect 22051 11713 22063 11747
rect 22005 11707 22063 11713
rect 22094 11704 22100 11756
rect 22152 11744 22158 11756
rect 22370 11744 22376 11756
rect 22152 11716 22197 11744
rect 22283 11716 22376 11744
rect 22152 11704 22158 11716
rect 22370 11704 22376 11716
rect 22428 11704 22434 11756
rect 23198 11744 23204 11756
rect 23159 11716 23204 11744
rect 23198 11704 23204 11716
rect 23256 11704 23262 11756
rect 23474 11744 23480 11756
rect 23387 11716 23480 11744
rect 23474 11704 23480 11716
rect 23532 11744 23538 11756
rect 24486 11744 24492 11756
rect 23532 11716 24492 11744
rect 23532 11704 23538 11716
rect 24486 11704 24492 11716
rect 24544 11704 24550 11756
rect 25682 11744 25688 11756
rect 25643 11716 25688 11744
rect 25682 11704 25688 11716
rect 25740 11704 25746 11756
rect 28074 11753 28080 11756
rect 28068 11707 28080 11753
rect 28132 11744 28138 11756
rect 28132 11716 28168 11744
rect 28074 11704 28080 11707
rect 28132 11704 28138 11716
rect 29730 11704 29736 11756
rect 29788 11744 29794 11756
rect 30282 11744 30288 11756
rect 29788 11716 30288 11744
rect 29788 11704 29794 11716
rect 30282 11704 30288 11716
rect 30340 11704 30346 11756
rect 31036 11744 31064 11772
rect 31159 11747 31217 11753
rect 31159 11744 31171 11747
rect 31036 11716 31171 11744
rect 31159 11713 31171 11716
rect 31205 11713 31217 11747
rect 31294 11744 31300 11756
rect 31255 11716 31300 11744
rect 31159 11707 31217 11713
rect 31294 11704 31300 11716
rect 31352 11704 31358 11756
rect 31410 11747 31468 11753
rect 31410 11713 31422 11747
rect 31456 11744 31468 11747
rect 31496 11744 31524 11784
rect 32493 11781 32505 11784
rect 32539 11781 32551 11815
rect 33318 11812 33324 11824
rect 33279 11784 33324 11812
rect 32493 11775 32551 11781
rect 33318 11772 33324 11784
rect 33376 11772 33382 11824
rect 31456 11716 31524 11744
rect 31573 11747 31631 11753
rect 31456 11713 31468 11716
rect 31410 11707 31468 11713
rect 31573 11713 31585 11747
rect 31619 11713 31631 11747
rect 32122 11744 32128 11756
rect 32083 11716 32128 11744
rect 31573 11707 31631 11713
rect 20346 11676 20352 11688
rect 19996 11648 20352 11676
rect 20346 11636 20352 11648
rect 20404 11636 20410 11688
rect 22186 11676 22192 11688
rect 22147 11648 22192 11676
rect 22186 11636 22192 11648
rect 22244 11636 22250 11688
rect 22388 11676 22416 11704
rect 24394 11676 24400 11688
rect 22388 11648 24400 11676
rect 22388 11608 22416 11648
rect 24394 11636 24400 11648
rect 24452 11636 24458 11688
rect 25958 11676 25964 11688
rect 25919 11648 25964 11676
rect 25958 11636 25964 11648
rect 26016 11636 26022 11688
rect 27430 11636 27436 11688
rect 27488 11676 27494 11688
rect 27801 11679 27859 11685
rect 27801 11676 27813 11679
rect 27488 11648 27813 11676
rect 27488 11636 27494 11648
rect 27801 11645 27813 11648
rect 27847 11645 27859 11679
rect 31588 11676 31616 11707
rect 32122 11704 32128 11716
rect 32180 11704 32186 11756
rect 32309 11747 32367 11753
rect 32309 11713 32321 11747
rect 32355 11744 32367 11747
rect 32858 11744 32864 11756
rect 32355 11716 32864 11744
rect 32355 11713 32367 11716
rect 32309 11707 32367 11713
rect 32858 11704 32864 11716
rect 32916 11744 32922 11756
rect 33137 11747 33195 11753
rect 33137 11744 33149 11747
rect 32916 11716 33149 11744
rect 32916 11704 32922 11716
rect 33137 11713 33149 11716
rect 33183 11713 33195 11747
rect 33137 11707 33195 11713
rect 34330 11676 34336 11688
rect 27801 11639 27859 11645
rect 31496 11648 31616 11676
rect 34291 11648 34336 11676
rect 31496 11620 31524 11648
rect 34330 11636 34336 11648
rect 34388 11636 34394 11688
rect 19904 11580 22416 11608
rect 30469 11611 30527 11617
rect 30469 11577 30481 11611
rect 30515 11608 30527 11611
rect 31478 11608 31484 11620
rect 30515 11580 31484 11608
rect 30515 11577 30527 11580
rect 30469 11571 30527 11577
rect 31478 11568 31484 11580
rect 31536 11568 31542 11620
rect 1578 11500 1584 11552
rect 1636 11540 1642 11552
rect 2133 11543 2191 11549
rect 2133 11540 2145 11543
rect 1636 11512 2145 11540
rect 1636 11500 1642 11512
rect 2133 11509 2145 11512
rect 2179 11509 2191 11543
rect 2133 11503 2191 11509
rect 21358 11500 21364 11552
rect 21416 11540 21422 11552
rect 22557 11543 22615 11549
rect 22557 11540 22569 11543
rect 21416 11512 22569 11540
rect 21416 11500 21422 11512
rect 22557 11509 22569 11512
rect 22603 11509 22615 11543
rect 22557 11503 22615 11509
rect 22830 11500 22836 11552
rect 22888 11540 22894 11552
rect 23017 11543 23075 11549
rect 23017 11540 23029 11543
rect 22888 11512 23029 11540
rect 22888 11500 22894 11512
rect 23017 11509 23029 11512
rect 23063 11509 23075 11543
rect 23017 11503 23075 11509
rect 23385 11543 23443 11549
rect 23385 11509 23397 11543
rect 23431 11540 23443 11543
rect 23750 11540 23756 11552
rect 23431 11512 23756 11540
rect 23431 11509 23443 11512
rect 23385 11503 23443 11509
rect 23750 11500 23756 11512
rect 23808 11540 23814 11552
rect 24026 11540 24032 11552
rect 23808 11512 24032 11540
rect 23808 11500 23814 11512
rect 24026 11500 24032 11512
rect 24084 11500 24090 11552
rect 25498 11500 25504 11552
rect 25556 11540 25562 11552
rect 25866 11540 25872 11552
rect 25556 11512 25872 11540
rect 25556 11500 25562 11512
rect 25866 11500 25872 11512
rect 25924 11500 25930 11552
rect 30929 11543 30987 11549
rect 30929 11509 30941 11543
rect 30975 11540 30987 11543
rect 31754 11540 31760 11552
rect 30975 11512 31760 11540
rect 30975 11509 30987 11512
rect 30929 11503 30987 11509
rect 31754 11500 31760 11512
rect 31812 11500 31818 11552
rect 46290 11500 46296 11552
rect 46348 11540 46354 11552
rect 47765 11543 47823 11549
rect 47765 11540 47777 11543
rect 46348 11512 47777 11540
rect 46348 11500 46354 11512
rect 47765 11509 47777 11512
rect 47811 11509 47823 11543
rect 47765 11503 47823 11509
rect 1104 11450 48852 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 48852 11450
rect 1104 11376 48852 11398
rect 19613 11339 19671 11345
rect 19613 11305 19625 11339
rect 19659 11336 19671 11339
rect 20070 11336 20076 11348
rect 19659 11308 20076 11336
rect 19659 11305 19671 11308
rect 19613 11299 19671 11305
rect 20070 11296 20076 11308
rect 20128 11296 20134 11348
rect 21821 11339 21879 11345
rect 21821 11305 21833 11339
rect 21867 11336 21879 11339
rect 22094 11336 22100 11348
rect 21867 11308 22100 11336
rect 21867 11305 21879 11308
rect 21821 11299 21879 11305
rect 22094 11296 22100 11308
rect 22152 11296 22158 11348
rect 23753 11339 23811 11345
rect 23753 11305 23765 11339
rect 23799 11336 23811 11339
rect 23842 11336 23848 11348
rect 23799 11308 23848 11336
rect 23799 11305 23811 11308
rect 23753 11299 23811 11305
rect 23842 11296 23848 11308
rect 23900 11296 23906 11348
rect 24026 11296 24032 11348
rect 24084 11336 24090 11348
rect 25777 11339 25835 11345
rect 25777 11336 25789 11339
rect 24084 11308 25789 11336
rect 24084 11296 24090 11308
rect 25777 11305 25789 11308
rect 25823 11305 25835 11339
rect 25777 11299 25835 11305
rect 27985 11339 28043 11345
rect 27985 11305 27997 11339
rect 28031 11336 28043 11339
rect 28074 11336 28080 11348
rect 28031 11308 28080 11336
rect 28031 11305 28043 11308
rect 27985 11299 28043 11305
rect 28074 11296 28080 11308
rect 28132 11296 28138 11348
rect 28258 11296 28264 11348
rect 28316 11336 28322 11348
rect 46566 11336 46572 11348
rect 28316 11308 46572 11336
rect 28316 11296 28322 11308
rect 46566 11296 46572 11308
rect 46624 11296 46630 11348
rect 27614 11268 27620 11280
rect 27540 11240 27620 11268
rect 1578 11200 1584 11212
rect 1539 11172 1584 11200
rect 1578 11160 1584 11172
rect 1636 11160 1642 11212
rect 2774 11200 2780 11212
rect 2735 11172 2780 11200
rect 2774 11160 2780 11172
rect 2832 11160 2838 11212
rect 23382 11160 23388 11212
rect 23440 11200 23446 11212
rect 27540 11209 27568 11240
rect 27614 11228 27620 11240
rect 27672 11228 27678 11280
rect 32858 11268 32864 11280
rect 32819 11240 32864 11268
rect 32858 11228 32864 11240
rect 32916 11228 32922 11280
rect 26605 11203 26663 11209
rect 26605 11200 26617 11203
rect 23440 11172 26617 11200
rect 23440 11160 23446 11172
rect 26605 11169 26617 11172
rect 26651 11169 26663 11203
rect 26605 11163 26663 11169
rect 27525 11203 27583 11209
rect 27525 11169 27537 11203
rect 27571 11169 27583 11203
rect 28166 11200 28172 11212
rect 27525 11163 27583 11169
rect 27816 11172 28172 11200
rect 1397 11135 1455 11141
rect 1397 11101 1409 11135
rect 1443 11101 1455 11135
rect 1397 11095 1455 11101
rect 1412 11064 1440 11095
rect 19150 11092 19156 11144
rect 19208 11132 19214 11144
rect 19429 11135 19487 11141
rect 19429 11132 19441 11135
rect 19208 11104 19441 11132
rect 19208 11092 19214 11104
rect 19429 11101 19441 11104
rect 19475 11101 19487 11135
rect 19429 11095 19487 11101
rect 20441 11135 20499 11141
rect 20441 11101 20453 11135
rect 20487 11132 20499 11135
rect 21818 11132 21824 11144
rect 20487 11104 21824 11132
rect 20487 11101 20499 11104
rect 20441 11095 20499 11101
rect 21818 11092 21824 11104
rect 21876 11132 21882 11144
rect 22373 11135 22431 11141
rect 22373 11132 22385 11135
rect 21876 11104 22385 11132
rect 21876 11092 21882 11104
rect 22373 11101 22385 11104
rect 22419 11101 22431 11135
rect 22373 11095 22431 11101
rect 23198 11092 23204 11144
rect 23256 11132 23262 11144
rect 25593 11135 25651 11141
rect 25593 11132 25605 11135
rect 23256 11104 25605 11132
rect 23256 11092 23262 11104
rect 25593 11101 25605 11104
rect 25639 11101 25651 11135
rect 25593 11095 25651 11101
rect 25869 11135 25927 11141
rect 25869 11101 25881 11135
rect 25915 11132 25927 11135
rect 26050 11132 26056 11144
rect 25915 11104 26056 11132
rect 25915 11101 25927 11104
rect 25869 11095 25927 11101
rect 26050 11092 26056 11104
rect 26108 11092 26114 11144
rect 27246 11132 27252 11144
rect 27207 11104 27252 11132
rect 27246 11092 27252 11104
rect 27304 11092 27310 11144
rect 27433 11135 27491 11141
rect 27433 11101 27445 11135
rect 27479 11101 27491 11135
rect 27614 11132 27620 11144
rect 27575 11104 27620 11132
rect 27433 11095 27491 11101
rect 2314 11064 2320 11076
rect 1412 11036 2320 11064
rect 2314 11024 2320 11036
rect 2372 11024 2378 11076
rect 19245 11067 19303 11073
rect 19245 11033 19257 11067
rect 19291 11064 19303 11067
rect 19334 11064 19340 11076
rect 19291 11036 19340 11064
rect 19291 11033 19303 11036
rect 19245 11027 19303 11033
rect 19334 11024 19340 11036
rect 19392 11024 19398 11076
rect 20708 11067 20766 11073
rect 20708 11033 20720 11067
rect 20754 11064 20766 11067
rect 21358 11064 21364 11076
rect 20754 11036 21364 11064
rect 20754 11033 20766 11036
rect 20708 11027 20766 11033
rect 21358 11024 21364 11036
rect 21416 11024 21422 11076
rect 22640 11067 22698 11073
rect 22640 11033 22652 11067
rect 22686 11064 22698 11067
rect 23382 11064 23388 11076
rect 22686 11036 23388 11064
rect 22686 11033 22698 11036
rect 22640 11027 22698 11033
rect 23382 11024 23388 11036
rect 23440 11024 23446 11076
rect 24578 11064 24584 11076
rect 24539 11036 24584 11064
rect 24578 11024 24584 11036
rect 24636 11024 24642 11076
rect 24765 11067 24823 11073
rect 24765 11033 24777 11067
rect 24811 11064 24823 11067
rect 24854 11064 24860 11076
rect 24811 11036 24860 11064
rect 24811 11033 24823 11036
rect 24765 11027 24823 11033
rect 24854 11024 24860 11036
rect 24912 11024 24918 11076
rect 24949 11067 25007 11073
rect 24949 11033 24961 11067
rect 24995 11064 25007 11067
rect 25958 11064 25964 11076
rect 24995 11036 25964 11064
rect 24995 11033 25007 11036
rect 24949 11027 25007 11033
rect 25958 11024 25964 11036
rect 26016 11064 26022 11076
rect 26421 11067 26479 11073
rect 26421 11064 26433 11067
rect 26016 11036 26433 11064
rect 26016 11024 26022 11036
rect 26421 11033 26433 11036
rect 26467 11033 26479 11067
rect 27448 11064 27476 11095
rect 27614 11092 27620 11104
rect 27672 11092 27678 11144
rect 27816 11141 27844 11172
rect 28166 11160 28172 11172
rect 28224 11160 28230 11212
rect 46290 11200 46296 11212
rect 46251 11172 46296 11200
rect 46290 11160 46296 11172
rect 46348 11160 46354 11212
rect 27801 11135 27859 11141
rect 27801 11101 27813 11135
rect 27847 11101 27859 11135
rect 27801 11095 27859 11101
rect 27890 11092 27896 11144
rect 27948 11132 27954 11144
rect 28537 11135 28595 11141
rect 28537 11132 28549 11135
rect 27948 11104 28549 11132
rect 27948 11092 27954 11104
rect 28537 11101 28549 11104
rect 28583 11101 28595 11135
rect 30006 11132 30012 11144
rect 29967 11104 30012 11132
rect 28537 11095 28595 11101
rect 30006 11092 30012 11104
rect 30064 11092 30070 11144
rect 31481 11135 31539 11141
rect 31481 11101 31493 11135
rect 31527 11132 31539 11135
rect 31570 11132 31576 11144
rect 31527 11104 31576 11132
rect 31527 11101 31539 11104
rect 31481 11095 31539 11101
rect 31570 11092 31576 11104
rect 31628 11092 31634 11144
rect 31754 11141 31760 11144
rect 31748 11095 31760 11141
rect 31812 11132 31818 11144
rect 31812 11104 31848 11132
rect 31754 11092 31760 11095
rect 31812 11092 31818 11104
rect 27706 11064 27712 11076
rect 27448 11036 27712 11064
rect 26421 11027 26479 11033
rect 27706 11024 27712 11036
rect 27764 11024 27770 11076
rect 28718 11064 28724 11076
rect 28679 11036 28724 11064
rect 28718 11024 28724 11036
rect 28776 11024 28782 11076
rect 30282 11024 30288 11076
rect 30340 11064 30346 11076
rect 35894 11064 35900 11076
rect 30340 11036 35900 11064
rect 30340 11024 30346 11036
rect 35894 11024 35900 11036
rect 35952 11024 35958 11076
rect 46477 11067 46535 11073
rect 46477 11033 46489 11067
rect 46523 11064 46535 11067
rect 46934 11064 46940 11076
rect 46523 11036 46940 11064
rect 46523 11033 46535 11036
rect 46477 11027 46535 11033
rect 46934 11024 46940 11036
rect 46992 11024 46998 11076
rect 48130 11064 48136 11076
rect 48091 11036 48136 11064
rect 48130 11024 48136 11036
rect 48188 11024 48194 11076
rect 18782 10956 18788 11008
rect 18840 10996 18846 11008
rect 23474 10996 23480 11008
rect 18840 10968 23480 10996
rect 18840 10956 18846 10968
rect 23474 10956 23480 10968
rect 23532 10956 23538 11008
rect 25038 10956 25044 11008
rect 25096 10996 25102 11008
rect 25409 10999 25467 11005
rect 25409 10996 25421 10999
rect 25096 10968 25421 10996
rect 25096 10956 25102 10968
rect 25409 10965 25421 10968
rect 25455 10965 25467 10999
rect 25409 10959 25467 10965
rect 28994 10956 29000 11008
rect 29052 10996 29058 11008
rect 30101 10999 30159 11005
rect 30101 10996 30113 10999
rect 29052 10968 30113 10996
rect 29052 10956 29058 10968
rect 30101 10965 30113 10968
rect 30147 10996 30159 10999
rect 30190 10996 30196 11008
rect 30147 10968 30196 10996
rect 30147 10965 30159 10968
rect 30101 10959 30159 10965
rect 30190 10956 30196 10968
rect 30248 10956 30254 11008
rect 1104 10906 48852 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 48852 10906
rect 1104 10832 48852 10854
rect 23382 10792 23388 10804
rect 23343 10764 23388 10792
rect 23382 10752 23388 10764
rect 23440 10752 23446 10804
rect 23842 10752 23848 10804
rect 23900 10752 23906 10804
rect 24029 10795 24087 10801
rect 24029 10761 24041 10795
rect 24075 10792 24087 10795
rect 24854 10792 24860 10804
rect 24075 10764 24860 10792
rect 24075 10761 24087 10764
rect 24029 10755 24087 10761
rect 24854 10752 24860 10764
rect 24912 10792 24918 10804
rect 25682 10792 25688 10804
rect 24912 10764 25688 10792
rect 24912 10752 24918 10764
rect 25682 10752 25688 10764
rect 25740 10752 25746 10804
rect 26510 10792 26516 10804
rect 26068 10764 26516 10792
rect 23109 10727 23167 10733
rect 23109 10693 23121 10727
rect 23155 10724 23167 10727
rect 23860 10724 23888 10752
rect 24210 10724 24216 10736
rect 23155 10696 23888 10724
rect 24044 10696 24216 10724
rect 23155 10693 23167 10696
rect 23109 10687 23167 10693
rect 1394 10656 1400 10668
rect 1355 10628 1400 10656
rect 1394 10616 1400 10628
rect 1452 10616 1458 10668
rect 2314 10656 2320 10668
rect 2275 10628 2320 10656
rect 2314 10616 2320 10628
rect 2372 10616 2378 10668
rect 18782 10656 18788 10668
rect 18743 10628 18788 10656
rect 18782 10616 18788 10628
rect 18840 10616 18846 10668
rect 18877 10659 18935 10665
rect 18877 10625 18889 10659
rect 18923 10625 18935 10659
rect 18877 10619 18935 10625
rect 18892 10588 18920 10619
rect 18966 10616 18972 10668
rect 19024 10656 19030 10668
rect 19153 10659 19211 10665
rect 19024 10628 19069 10656
rect 19024 10616 19030 10628
rect 19153 10625 19165 10659
rect 19199 10656 19211 10659
rect 19426 10656 19432 10668
rect 19199 10628 19432 10656
rect 19199 10625 19211 10628
rect 19153 10619 19211 10625
rect 19426 10616 19432 10628
rect 19484 10616 19490 10668
rect 22830 10656 22836 10668
rect 22791 10628 22836 10656
rect 22830 10616 22836 10628
rect 22888 10616 22894 10668
rect 23014 10656 23020 10668
rect 22975 10628 23020 10656
rect 23014 10616 23020 10628
rect 23072 10616 23078 10668
rect 23201 10659 23259 10665
rect 23201 10625 23213 10659
rect 23247 10625 23259 10659
rect 23201 10619 23259 10625
rect 23845 10659 23903 10665
rect 23845 10625 23857 10659
rect 23891 10656 23903 10659
rect 24044 10656 24072 10696
rect 24210 10684 24216 10696
rect 24268 10724 24274 10736
rect 24486 10724 24492 10736
rect 24268 10696 24492 10724
rect 24268 10684 24274 10696
rect 24486 10684 24492 10696
rect 24544 10684 24550 10736
rect 25225 10727 25283 10733
rect 25225 10693 25237 10727
rect 25271 10724 25283 10727
rect 25958 10724 25964 10736
rect 25271 10696 25964 10724
rect 25271 10693 25283 10696
rect 25225 10687 25283 10693
rect 25958 10684 25964 10696
rect 26016 10684 26022 10736
rect 26068 10733 26096 10764
rect 26510 10752 26516 10764
rect 26568 10752 26574 10804
rect 28718 10752 28724 10804
rect 28776 10792 28782 10804
rect 30558 10792 30564 10804
rect 28776 10764 30564 10792
rect 28776 10752 28782 10764
rect 30558 10752 30564 10764
rect 30616 10752 30622 10804
rect 46934 10792 46940 10804
rect 46895 10764 46940 10792
rect 46934 10752 46940 10764
rect 46992 10752 46998 10804
rect 26053 10727 26111 10733
rect 26053 10693 26065 10727
rect 26099 10693 26111 10727
rect 26053 10687 26111 10693
rect 26237 10727 26295 10733
rect 26237 10693 26249 10727
rect 26283 10724 26295 10727
rect 26694 10724 26700 10736
rect 26283 10696 26700 10724
rect 26283 10693 26295 10696
rect 26237 10687 26295 10693
rect 26694 10684 26700 10696
rect 26752 10684 26758 10736
rect 48038 10724 48044 10736
rect 30070 10696 48044 10724
rect 23891 10628 24072 10656
rect 24121 10659 24179 10665
rect 23891 10625 23903 10628
rect 23845 10619 23903 10625
rect 24121 10625 24133 10659
rect 24167 10656 24179 10659
rect 24578 10656 24584 10668
rect 24167 10628 24584 10656
rect 24167 10625 24179 10628
rect 24121 10619 24179 10625
rect 19518 10588 19524 10600
rect 18892 10560 19524 10588
rect 19518 10548 19524 10560
rect 19576 10588 19582 10600
rect 20254 10588 20260 10600
rect 19576 10560 20260 10588
rect 19576 10548 19582 10560
rect 20254 10548 20260 10560
rect 20312 10548 20318 10600
rect 23216 10588 23244 10619
rect 24578 10616 24584 10628
rect 24636 10616 24642 10668
rect 24949 10659 25007 10665
rect 24949 10625 24961 10659
rect 24995 10656 25007 10659
rect 25038 10656 25044 10668
rect 24995 10628 25044 10656
rect 24995 10625 25007 10628
rect 24949 10619 25007 10625
rect 25038 10616 25044 10628
rect 25096 10616 25102 10668
rect 25130 10616 25136 10668
rect 25188 10656 25194 10668
rect 25317 10659 25375 10665
rect 25188 10628 25233 10656
rect 25188 10616 25194 10628
rect 25317 10625 25329 10659
rect 25363 10625 25375 10659
rect 25317 10619 25375 10625
rect 23658 10588 23664 10600
rect 23216 10560 23664 10588
rect 23658 10548 23664 10560
rect 23716 10588 23722 10600
rect 25332 10588 25360 10619
rect 25406 10616 25412 10668
rect 25464 10656 25470 10668
rect 26326 10656 26332 10668
rect 25464 10628 26332 10656
rect 25464 10616 25470 10628
rect 26326 10616 26332 10628
rect 26384 10616 26390 10668
rect 26973 10659 27031 10665
rect 26973 10625 26985 10659
rect 27019 10625 27031 10659
rect 26973 10619 27031 10625
rect 26988 10588 27016 10619
rect 27062 10616 27068 10668
rect 27120 10656 27126 10668
rect 27157 10659 27215 10665
rect 27157 10656 27169 10659
rect 27120 10628 27169 10656
rect 27120 10616 27126 10628
rect 27157 10625 27169 10628
rect 27203 10625 27215 10659
rect 27157 10619 27215 10625
rect 28537 10659 28595 10665
rect 28537 10625 28549 10659
rect 28583 10656 28595 10659
rect 29822 10656 29828 10668
rect 28583 10628 29828 10656
rect 28583 10625 28595 10628
rect 28537 10619 28595 10625
rect 29822 10616 29828 10628
rect 29880 10616 29886 10668
rect 30070 10665 30098 10696
rect 48038 10684 48044 10696
rect 48096 10684 48102 10736
rect 30055 10659 30113 10665
rect 30055 10625 30067 10659
rect 30101 10625 30113 10659
rect 30190 10656 30196 10668
rect 30151 10628 30196 10656
rect 30055 10619 30113 10625
rect 30190 10616 30196 10628
rect 30248 10616 30254 10668
rect 30285 10659 30343 10665
rect 30285 10625 30297 10659
rect 30331 10654 30343 10659
rect 30374 10654 30380 10668
rect 30331 10626 30380 10654
rect 30331 10625 30343 10626
rect 30285 10619 30343 10625
rect 30374 10616 30380 10626
rect 30432 10616 30438 10668
rect 30469 10659 30527 10665
rect 30469 10625 30481 10659
rect 30515 10656 30527 10659
rect 30558 10656 30564 10668
rect 30515 10628 30564 10656
rect 30515 10625 30527 10628
rect 30469 10619 30527 10625
rect 30558 10616 30564 10628
rect 30616 10616 30622 10668
rect 32582 10656 32588 10668
rect 32543 10628 32588 10656
rect 32582 10616 32588 10628
rect 32640 10616 32646 10668
rect 46382 10616 46388 10668
rect 46440 10656 46446 10668
rect 46845 10659 46903 10665
rect 46845 10656 46857 10659
rect 46440 10628 46857 10656
rect 46440 10616 46446 10628
rect 46845 10625 46857 10628
rect 46891 10625 46903 10659
rect 47854 10656 47860 10668
rect 47815 10628 47860 10656
rect 46845 10619 46903 10625
rect 47854 10616 47860 10628
rect 47912 10616 47918 10668
rect 23716 10560 25360 10588
rect 26068 10560 27016 10588
rect 23716 10548 23722 10560
rect 1581 10523 1639 10529
rect 1581 10489 1593 10523
rect 1627 10520 1639 10523
rect 22738 10520 22744 10532
rect 1627 10492 22744 10520
rect 1627 10489 1639 10492
rect 1581 10483 1639 10489
rect 22738 10480 22744 10492
rect 22796 10480 22802 10532
rect 22922 10480 22928 10532
rect 22980 10520 22986 10532
rect 26068 10529 26096 10560
rect 28626 10548 28632 10600
rect 28684 10588 28690 10600
rect 28813 10591 28871 10597
rect 28813 10588 28825 10591
rect 28684 10560 28825 10588
rect 28684 10548 28690 10560
rect 28813 10557 28825 10560
rect 28859 10557 28871 10591
rect 28813 10551 28871 10557
rect 32950 10548 32956 10600
rect 33008 10588 33014 10600
rect 33229 10591 33287 10597
rect 33229 10588 33241 10591
rect 33008 10560 33241 10588
rect 33008 10548 33014 10560
rect 33229 10557 33241 10560
rect 33275 10557 33287 10591
rect 33229 10551 33287 10557
rect 33413 10591 33471 10597
rect 33413 10557 33425 10591
rect 33459 10557 33471 10591
rect 34606 10588 34612 10600
rect 34567 10560 34612 10588
rect 33413 10551 33471 10557
rect 26053 10523 26111 10529
rect 22980 10492 25636 10520
rect 22980 10480 22986 10492
rect 18506 10452 18512 10464
rect 18467 10424 18512 10452
rect 18506 10412 18512 10424
rect 18564 10412 18570 10464
rect 23474 10412 23480 10464
rect 23532 10452 23538 10464
rect 23845 10455 23903 10461
rect 23845 10452 23857 10455
rect 23532 10424 23857 10452
rect 23532 10412 23538 10424
rect 23845 10421 23857 10424
rect 23891 10421 23903 10455
rect 25498 10452 25504 10464
rect 25459 10424 25504 10452
rect 23845 10415 23903 10421
rect 25498 10412 25504 10424
rect 25556 10412 25562 10464
rect 25608 10452 25636 10492
rect 26053 10489 26065 10523
rect 26099 10489 26111 10523
rect 26053 10483 26111 10489
rect 32677 10523 32735 10529
rect 32677 10489 32689 10523
rect 32723 10520 32735 10523
rect 33428 10520 33456 10551
rect 34606 10548 34612 10560
rect 34664 10548 34670 10600
rect 48041 10523 48099 10529
rect 48041 10520 48053 10523
rect 32723 10492 33456 10520
rect 41386 10492 48053 10520
rect 32723 10489 32735 10492
rect 32677 10483 32735 10489
rect 26510 10452 26516 10464
rect 25608 10424 26516 10452
rect 26510 10412 26516 10424
rect 26568 10412 26574 10464
rect 27065 10455 27123 10461
rect 27065 10421 27077 10455
rect 27111 10452 27123 10455
rect 27154 10452 27160 10464
rect 27111 10424 27160 10452
rect 27111 10421 27123 10424
rect 27065 10415 27123 10421
rect 27154 10412 27160 10424
rect 27212 10412 27218 10464
rect 29822 10452 29828 10464
rect 29783 10424 29828 10452
rect 29822 10412 29828 10424
rect 29880 10412 29886 10464
rect 30926 10412 30932 10464
rect 30984 10452 30990 10464
rect 41386 10452 41414 10492
rect 48041 10489 48053 10492
rect 48087 10489 48099 10523
rect 48041 10483 48099 10489
rect 30984 10424 41414 10452
rect 30984 10412 30990 10424
rect 1104 10362 48852 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 48852 10362
rect 1104 10288 48852 10310
rect 23014 10248 23020 10260
rect 22975 10220 23020 10248
rect 23014 10208 23020 10220
rect 23072 10208 23078 10260
rect 24578 10208 24584 10260
rect 24636 10248 24642 10260
rect 24636 10220 24716 10248
rect 24636 10208 24642 10220
rect 24688 10180 24716 10220
rect 24946 10208 24952 10260
rect 25004 10248 25010 10260
rect 25409 10251 25467 10257
rect 25409 10248 25421 10251
rect 25004 10220 25421 10248
rect 25004 10208 25010 10220
rect 25409 10217 25421 10220
rect 25455 10248 25467 10251
rect 25590 10248 25596 10260
rect 25455 10220 25596 10248
rect 25455 10217 25467 10220
rect 25409 10211 25467 10217
rect 25590 10208 25596 10220
rect 25648 10208 25654 10260
rect 26237 10251 26295 10257
rect 26237 10217 26249 10251
rect 26283 10217 26295 10251
rect 26237 10211 26295 10217
rect 26252 10180 26280 10211
rect 26510 10208 26516 10260
rect 26568 10248 26574 10260
rect 27341 10251 27399 10257
rect 27341 10248 27353 10251
rect 26568 10220 27353 10248
rect 26568 10208 26574 10220
rect 27341 10217 27353 10220
rect 27387 10248 27399 10251
rect 28350 10248 28356 10260
rect 27387 10220 28356 10248
rect 27387 10217 27399 10220
rect 27341 10211 27399 10217
rect 28350 10208 28356 10220
rect 28408 10208 28414 10260
rect 28997 10251 29055 10257
rect 28997 10217 29009 10251
rect 29043 10248 29055 10251
rect 30282 10248 30288 10260
rect 29043 10220 30288 10248
rect 29043 10217 29055 10220
rect 28997 10211 29055 10217
rect 30282 10208 30288 10220
rect 30340 10208 30346 10260
rect 32950 10248 32956 10260
rect 32911 10220 32956 10248
rect 32950 10208 32956 10220
rect 33008 10208 33014 10260
rect 24688 10152 26280 10180
rect 19426 10072 19432 10124
rect 19484 10112 19490 10124
rect 20254 10112 20260 10124
rect 19484 10084 20260 10112
rect 19484 10072 19490 10084
rect 20254 10072 20260 10084
rect 20312 10072 20318 10124
rect 23474 10112 23480 10124
rect 22940 10084 23480 10112
rect 1762 10004 1768 10056
rect 1820 10044 1826 10056
rect 2041 10047 2099 10053
rect 2041 10044 2053 10047
rect 1820 10016 2053 10044
rect 1820 10004 1826 10016
rect 2041 10013 2053 10016
rect 2087 10013 2099 10047
rect 2041 10007 2099 10013
rect 16853 10047 16911 10053
rect 16853 10013 16865 10047
rect 16899 10044 16911 10047
rect 17586 10044 17592 10056
rect 16899 10016 17592 10044
rect 16899 10013 16911 10016
rect 16853 10007 16911 10013
rect 17586 10004 17592 10016
rect 17644 10004 17650 10056
rect 19334 10004 19340 10056
rect 19392 10044 19398 10056
rect 19702 10044 19708 10056
rect 19392 10016 19437 10044
rect 19663 10016 19708 10044
rect 19392 10004 19398 10016
rect 19702 10004 19708 10016
rect 19760 10004 19766 10056
rect 22940 10053 22968 10084
rect 23474 10072 23480 10084
rect 23532 10072 23538 10124
rect 25406 10112 25412 10124
rect 25367 10084 25412 10112
rect 25406 10072 25412 10084
rect 25464 10072 25470 10124
rect 26329 10115 26387 10121
rect 26329 10112 26341 10115
rect 25608 10084 26341 10112
rect 22925 10047 22983 10053
rect 22925 10013 22937 10047
rect 22971 10013 22983 10047
rect 22925 10007 22983 10013
rect 23109 10047 23167 10053
rect 23109 10013 23121 10047
rect 23155 10044 23167 10047
rect 23290 10044 23296 10056
rect 23155 10016 23296 10044
rect 23155 10013 23167 10016
rect 23109 10007 23167 10013
rect 23290 10004 23296 10016
rect 23348 10004 23354 10056
rect 24302 10004 24308 10056
rect 24360 10044 24366 10056
rect 24581 10047 24639 10053
rect 24581 10044 24593 10047
rect 24360 10016 24593 10044
rect 24360 10004 24366 10016
rect 24581 10013 24593 10016
rect 24627 10013 24639 10047
rect 25501 10047 25559 10053
rect 25501 10038 25513 10047
rect 24581 10007 24639 10013
rect 25424 10013 25513 10038
rect 25547 10046 25559 10047
rect 25608 10046 25636 10084
rect 26329 10081 26341 10084
rect 26375 10081 26387 10115
rect 31570 10112 31576 10124
rect 31531 10084 31576 10112
rect 26329 10075 26387 10081
rect 31570 10072 31576 10084
rect 31628 10072 31634 10124
rect 25547 10018 25636 10046
rect 25547 10013 25559 10018
rect 25424 10010 25559 10013
rect 17120 9979 17178 9985
rect 17120 9945 17132 9979
rect 17166 9976 17178 9979
rect 18506 9976 18512 9988
rect 17166 9948 18512 9976
rect 17166 9945 17178 9948
rect 17120 9939 17178 9945
rect 18506 9936 18512 9948
rect 18564 9936 18570 9988
rect 19426 9936 19432 9988
rect 19484 9976 19490 9988
rect 19521 9979 19579 9985
rect 19521 9976 19533 9979
rect 19484 9948 19533 9976
rect 19484 9936 19490 9948
rect 19521 9945 19533 9948
rect 19567 9945 19579 9979
rect 19521 9939 19579 9945
rect 22005 9979 22063 9985
rect 22005 9945 22017 9979
rect 22051 9976 22063 9979
rect 23661 9979 23719 9985
rect 23661 9976 23673 9979
rect 22051 9948 23673 9976
rect 22051 9945 22063 9948
rect 22005 9939 22063 9945
rect 23661 9945 23673 9948
rect 23707 9976 23719 9979
rect 24765 9979 24823 9985
rect 24765 9976 24777 9979
rect 23707 9948 24777 9976
rect 23707 9945 23719 9948
rect 23661 9939 23719 9945
rect 24765 9945 24777 9948
rect 24811 9945 24823 9979
rect 25222 9976 25228 9988
rect 25183 9948 25228 9976
rect 24765 9939 24823 9945
rect 25222 9936 25228 9948
rect 25280 9936 25286 9988
rect 18230 9908 18236 9920
rect 18191 9880 18236 9908
rect 18230 9868 18236 9880
rect 18288 9868 18294 9920
rect 21818 9868 21824 9920
rect 21876 9908 21882 9920
rect 22097 9911 22155 9917
rect 22097 9908 22109 9911
rect 21876 9880 22109 9908
rect 21876 9868 21882 9880
rect 22097 9877 22109 9880
rect 22143 9877 22155 9911
rect 22097 9871 22155 9877
rect 23474 9868 23480 9920
rect 23532 9908 23538 9920
rect 23753 9911 23811 9917
rect 23753 9908 23765 9911
rect 23532 9880 23765 9908
rect 23532 9868 23538 9880
rect 23753 9877 23765 9880
rect 23799 9877 23811 9911
rect 23753 9871 23811 9877
rect 24026 9868 24032 9920
rect 24084 9908 24090 9920
rect 25424 9908 25452 10010
rect 25501 10007 25559 10010
rect 25682 10004 25688 10056
rect 25740 10044 25746 10056
rect 26513 10047 26571 10053
rect 26513 10044 26525 10047
rect 25740 10016 26525 10044
rect 25740 10004 25746 10016
rect 26513 10013 26525 10016
rect 26559 10013 26571 10047
rect 26513 10007 26571 10013
rect 27614 10004 27620 10056
rect 27672 10044 27678 10056
rect 28813 10047 28871 10053
rect 28813 10044 28825 10047
rect 27672 10016 28825 10044
rect 27672 10004 27678 10016
rect 28813 10013 28825 10016
rect 28859 10013 28871 10047
rect 28813 10007 28871 10013
rect 29549 10047 29607 10053
rect 29549 10013 29561 10047
rect 29595 10044 29607 10047
rect 30190 10044 30196 10056
rect 29595 10016 30196 10044
rect 29595 10013 29607 10016
rect 29549 10007 29607 10013
rect 25590 9936 25596 9988
rect 25648 9976 25654 9988
rect 26237 9979 26295 9985
rect 26237 9976 26249 9979
rect 25648 9948 26249 9976
rect 25648 9936 25654 9948
rect 26237 9945 26249 9948
rect 26283 9945 26295 9979
rect 26237 9939 26295 9945
rect 26970 9936 26976 9988
rect 27028 9976 27034 9988
rect 27249 9979 27307 9985
rect 27249 9976 27261 9979
rect 27028 9948 27261 9976
rect 27028 9936 27034 9948
rect 27249 9945 27261 9948
rect 27295 9945 27307 9979
rect 28626 9976 28632 9988
rect 28587 9948 28632 9976
rect 27249 9939 27307 9945
rect 28626 9936 28632 9948
rect 28684 9936 28690 9988
rect 24084 9880 25452 9908
rect 25685 9911 25743 9917
rect 24084 9868 24090 9880
rect 25685 9877 25697 9911
rect 25731 9908 25743 9911
rect 25866 9908 25872 9920
rect 25731 9880 25872 9908
rect 25731 9877 25743 9880
rect 25685 9871 25743 9877
rect 25866 9868 25872 9880
rect 25924 9868 25930 9920
rect 26694 9908 26700 9920
rect 26655 9880 26700 9908
rect 26694 9868 26700 9880
rect 26752 9868 26758 9920
rect 28828 9908 28856 10007
rect 30190 10004 30196 10016
rect 30248 10044 30254 10056
rect 31588 10044 31616 10072
rect 30248 10016 31616 10044
rect 30248 10004 30254 10016
rect 29822 9985 29828 9988
rect 29816 9976 29828 9985
rect 29783 9948 29828 9976
rect 29816 9939 29828 9948
rect 29822 9936 29828 9939
rect 29880 9936 29886 9988
rect 31018 9936 31024 9988
rect 31076 9976 31082 9988
rect 31818 9979 31876 9985
rect 31818 9976 31830 9979
rect 31076 9948 31830 9976
rect 31076 9936 31082 9948
rect 31818 9945 31830 9948
rect 31864 9945 31876 9979
rect 31818 9939 31876 9945
rect 30926 9908 30932 9920
rect 28828 9880 30932 9908
rect 30926 9868 30932 9880
rect 30984 9868 30990 9920
rect 1104 9818 48852 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 48852 9818
rect 1104 9744 48852 9766
rect 18417 9707 18475 9713
rect 18417 9673 18429 9707
rect 18463 9704 18475 9707
rect 18966 9704 18972 9716
rect 18463 9676 18972 9704
rect 18463 9673 18475 9676
rect 18417 9667 18475 9673
rect 18966 9664 18972 9676
rect 19024 9664 19030 9716
rect 21174 9704 21180 9716
rect 19628 9686 21180 9704
rect 3142 9596 3148 9648
rect 3200 9636 3206 9648
rect 18138 9636 18144 9648
rect 3200 9608 18144 9636
rect 3200 9596 3206 9608
rect 18138 9596 18144 9608
rect 18196 9596 18202 9648
rect 19610 9634 19616 9686
rect 19668 9676 21180 9686
rect 19668 9634 19674 9676
rect 21174 9664 21180 9676
rect 21232 9664 21238 9716
rect 22462 9664 22468 9716
rect 22520 9704 22526 9716
rect 22557 9707 22615 9713
rect 22557 9704 22569 9707
rect 22520 9676 22569 9704
rect 22520 9664 22526 9676
rect 22557 9673 22569 9676
rect 22603 9704 22615 9707
rect 23290 9704 23296 9716
rect 22603 9676 23296 9704
rect 22603 9673 22615 9676
rect 22557 9667 22615 9673
rect 23290 9664 23296 9676
rect 23348 9704 23354 9716
rect 23348 9676 24164 9704
rect 23348 9664 23354 9676
rect 20990 9636 20996 9648
rect 19720 9608 20996 9636
rect 1762 9568 1768 9580
rect 1723 9540 1768 9568
rect 1762 9528 1768 9540
rect 1820 9528 1826 9580
rect 17405 9571 17463 9577
rect 17405 9537 17417 9571
rect 17451 9568 17463 9571
rect 17862 9568 17868 9580
rect 17451 9540 17868 9568
rect 17451 9537 17463 9540
rect 17405 9531 17463 9537
rect 17862 9528 17868 9540
rect 17920 9528 17926 9580
rect 18046 9568 18052 9580
rect 18007 9540 18052 9568
rect 18046 9528 18052 9540
rect 18104 9528 18110 9580
rect 18230 9568 18236 9580
rect 18191 9540 18236 9568
rect 18230 9528 18236 9540
rect 18288 9528 18294 9580
rect 19334 9528 19340 9580
rect 19392 9528 19398 9580
rect 19720 9577 19748 9608
rect 20990 9596 20996 9608
rect 21048 9636 21054 9648
rect 22002 9636 22008 9648
rect 21048 9608 22008 9636
rect 21048 9596 21054 9608
rect 22002 9596 22008 9608
rect 22060 9596 22066 9648
rect 24026 9636 24032 9648
rect 22664 9608 24032 9636
rect 22664 9580 22692 9608
rect 24026 9596 24032 9608
rect 24084 9596 24090 9648
rect 19705 9571 19763 9577
rect 19705 9537 19717 9571
rect 19751 9537 19763 9571
rect 19705 9531 19763 9537
rect 19797 9571 19855 9577
rect 19797 9537 19809 9571
rect 19843 9537 19855 9571
rect 19797 9531 19855 9537
rect 19889 9571 19947 9577
rect 19889 9537 19901 9571
rect 19935 9568 19947 9571
rect 19978 9568 19984 9580
rect 19935 9540 19984 9568
rect 19935 9537 19947 9540
rect 19889 9531 19947 9537
rect 1949 9503 2007 9509
rect 1949 9469 1961 9503
rect 1995 9500 2007 9503
rect 2222 9500 2228 9512
rect 1995 9472 2228 9500
rect 1995 9469 2007 9472
rect 1949 9463 2007 9469
rect 2222 9460 2228 9472
rect 2280 9460 2286 9512
rect 2774 9500 2780 9512
rect 2735 9472 2780 9500
rect 2774 9460 2780 9472
rect 2832 9460 2838 9512
rect 18064 9500 18092 9528
rect 19352 9500 19380 9528
rect 18064 9472 19380 9500
rect 19812 9500 19840 9531
rect 19978 9528 19984 9540
rect 20036 9528 20042 9580
rect 20073 9571 20131 9577
rect 20073 9537 20085 9571
rect 20119 9568 20131 9571
rect 20254 9568 20260 9580
rect 20119 9540 20260 9568
rect 20119 9537 20131 9540
rect 20073 9531 20131 9537
rect 20254 9528 20260 9540
rect 20312 9528 20318 9580
rect 22373 9571 22431 9577
rect 22373 9537 22385 9571
rect 22419 9537 22431 9571
rect 22646 9568 22652 9580
rect 22559 9540 22652 9568
rect 22373 9531 22431 9537
rect 22388 9500 22416 9531
rect 22646 9528 22652 9540
rect 22704 9528 22710 9580
rect 23753 9571 23811 9577
rect 23753 9537 23765 9571
rect 23799 9537 23811 9571
rect 23753 9531 23811 9537
rect 22922 9500 22928 9512
rect 19812 9472 20024 9500
rect 22388 9472 22928 9500
rect 19996 9444 20024 9472
rect 22922 9460 22928 9472
rect 22980 9460 22986 9512
rect 23768 9500 23796 9531
rect 23842 9528 23848 9580
rect 23900 9568 23906 9580
rect 23937 9571 23995 9577
rect 23937 9568 23949 9571
rect 23900 9540 23949 9568
rect 23900 9528 23906 9540
rect 23937 9537 23949 9540
rect 23983 9568 23995 9571
rect 24136 9568 24164 9676
rect 25222 9664 25228 9716
rect 25280 9704 25286 9716
rect 25685 9707 25743 9713
rect 25685 9704 25697 9707
rect 25280 9676 25697 9704
rect 25280 9664 25286 9676
rect 25685 9673 25697 9676
rect 25731 9704 25743 9707
rect 25774 9704 25780 9716
rect 25731 9676 25780 9704
rect 25731 9673 25743 9676
rect 25685 9667 25743 9673
rect 25774 9664 25780 9676
rect 25832 9664 25838 9716
rect 25958 9664 25964 9716
rect 26016 9704 26022 9716
rect 26145 9707 26203 9713
rect 26145 9704 26157 9707
rect 26016 9676 26157 9704
rect 26016 9664 26022 9676
rect 26145 9673 26157 9676
rect 26191 9673 26203 9707
rect 26145 9667 26203 9673
rect 26326 9664 26332 9716
rect 26384 9704 26390 9716
rect 27157 9707 27215 9713
rect 27157 9704 27169 9707
rect 26384 9676 27169 9704
rect 26384 9664 26390 9676
rect 27157 9673 27169 9676
rect 27203 9673 27215 9707
rect 27157 9667 27215 9673
rect 30929 9707 30987 9713
rect 30929 9673 30941 9707
rect 30975 9704 30987 9707
rect 31018 9704 31024 9716
rect 30975 9676 31024 9704
rect 30975 9673 30987 9676
rect 30929 9667 30987 9673
rect 31018 9664 31024 9676
rect 31076 9664 31082 9716
rect 31294 9664 31300 9716
rect 31352 9664 31358 9716
rect 31478 9664 31484 9716
rect 31536 9704 31542 9716
rect 31536 9676 31708 9704
rect 31536 9664 31542 9676
rect 26694 9636 26700 9648
rect 24412 9608 26700 9636
rect 24412 9577 24440 9608
rect 26694 9596 26700 9608
rect 26752 9596 26758 9648
rect 27525 9639 27583 9645
rect 27525 9605 27537 9639
rect 27571 9636 27583 9639
rect 27614 9636 27620 9648
rect 27571 9608 27620 9636
rect 27571 9605 27583 9608
rect 27525 9599 27583 9605
rect 27614 9596 27620 9608
rect 27672 9596 27678 9648
rect 31309 9583 31337 9664
rect 23983 9540 24164 9568
rect 24397 9571 24455 9577
rect 23983 9537 23995 9540
rect 23937 9531 23995 9537
rect 24397 9537 24409 9571
rect 24443 9537 24455 9571
rect 25866 9568 25872 9580
rect 24397 9531 24455 9537
rect 24596 9540 25872 9568
rect 24596 9500 24624 9540
rect 25866 9528 25872 9540
rect 25924 9528 25930 9580
rect 26050 9568 26056 9580
rect 26011 9540 26056 9568
rect 26050 9528 26056 9540
rect 26108 9528 26114 9580
rect 27338 9568 27344 9580
rect 26344 9540 27344 9568
rect 23768 9472 24624 9500
rect 24673 9503 24731 9509
rect 24673 9469 24685 9503
rect 24719 9500 24731 9503
rect 26234 9500 26240 9512
rect 24719 9472 26240 9500
rect 24719 9469 24731 9472
rect 24673 9463 24731 9469
rect 26234 9460 26240 9472
rect 26292 9460 26298 9512
rect 26344 9509 26372 9540
rect 27338 9528 27344 9540
rect 27396 9568 27402 9580
rect 27396 9540 27752 9568
rect 27396 9528 27402 9540
rect 26329 9503 26387 9509
rect 26329 9469 26341 9503
rect 26375 9469 26387 9503
rect 26329 9463 26387 9469
rect 27246 9460 27252 9512
rect 27304 9500 27310 9512
rect 27724 9509 27752 9540
rect 30926 9528 30932 9580
rect 30984 9568 30990 9580
rect 31294 9577 31352 9583
rect 31205 9571 31263 9577
rect 31205 9568 31217 9571
rect 30984 9540 31217 9568
rect 30984 9528 30990 9540
rect 31205 9537 31217 9540
rect 31251 9537 31263 9571
rect 31294 9543 31306 9577
rect 31340 9543 31352 9577
rect 31294 9537 31352 9543
rect 31394 9571 31452 9577
rect 31394 9537 31406 9571
rect 31440 9537 31452 9571
rect 31205 9531 31263 9537
rect 31394 9531 31452 9537
rect 31585 9571 31643 9577
rect 31585 9537 31597 9571
rect 31631 9568 31643 9571
rect 31680 9568 31708 9676
rect 32309 9639 32367 9645
rect 32309 9605 32321 9639
rect 32355 9636 32367 9639
rect 32950 9636 32956 9648
rect 32355 9608 32956 9636
rect 32355 9605 32367 9608
rect 32309 9599 32367 9605
rect 32950 9596 32956 9608
rect 33008 9596 33014 9648
rect 32122 9568 32128 9580
rect 31631 9540 31708 9568
rect 32083 9540 32128 9568
rect 31631 9537 31643 9540
rect 31585 9531 31643 9537
rect 27617 9503 27675 9509
rect 27617 9500 27629 9503
rect 27304 9472 27629 9500
rect 27304 9460 27310 9472
rect 27617 9469 27629 9472
rect 27663 9469 27675 9503
rect 27617 9463 27675 9469
rect 27709 9503 27767 9509
rect 27709 9469 27721 9503
rect 27755 9469 27767 9503
rect 27709 9463 27767 9469
rect 19978 9392 19984 9444
rect 20036 9392 20042 9444
rect 20622 9392 20628 9444
rect 20680 9432 20686 9444
rect 26878 9432 26884 9444
rect 20680 9404 26884 9432
rect 20680 9392 20686 9404
rect 26878 9392 26884 9404
rect 26936 9392 26942 9444
rect 31404 9432 31432 9531
rect 32122 9528 32128 9540
rect 32180 9528 32186 9580
rect 32493 9503 32551 9509
rect 32493 9469 32505 9503
rect 32539 9469 32551 9503
rect 32493 9463 32551 9469
rect 32508 9432 32536 9463
rect 31404 9404 32536 9432
rect 17034 9324 17040 9376
rect 17092 9364 17098 9376
rect 17497 9367 17555 9373
rect 17497 9364 17509 9367
rect 17092 9336 17509 9364
rect 17092 9324 17098 9336
rect 17497 9333 17509 9336
rect 17543 9333 17555 9367
rect 17497 9327 17555 9333
rect 19429 9367 19487 9373
rect 19429 9333 19441 9367
rect 19475 9364 19487 9367
rect 19518 9364 19524 9376
rect 19475 9336 19524 9364
rect 19475 9333 19487 9336
rect 19429 9327 19487 9333
rect 19518 9324 19524 9336
rect 19576 9324 19582 9376
rect 21542 9324 21548 9376
rect 21600 9364 21606 9376
rect 22373 9367 22431 9373
rect 22373 9364 22385 9367
rect 21600 9336 22385 9364
rect 21600 9324 21606 9336
rect 22373 9333 22385 9336
rect 22419 9333 22431 9367
rect 23750 9364 23756 9376
rect 23711 9336 23756 9364
rect 22373 9327 22431 9333
rect 23750 9324 23756 9336
rect 23808 9324 23814 9376
rect 24486 9364 24492 9376
rect 24447 9336 24492 9364
rect 24486 9324 24492 9336
rect 24544 9324 24550 9376
rect 24578 9324 24584 9376
rect 24636 9364 24642 9376
rect 24949 9367 25007 9373
rect 24949 9364 24961 9367
rect 24636 9336 24961 9364
rect 24636 9324 24642 9336
rect 24949 9333 24961 9336
rect 24995 9333 25007 9367
rect 24949 9327 25007 9333
rect 26234 9324 26240 9376
rect 26292 9364 26298 9376
rect 26970 9364 26976 9376
rect 26292 9336 26976 9364
rect 26292 9324 26298 9336
rect 26970 9324 26976 9336
rect 27028 9324 27034 9376
rect 1104 9274 48852 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 48852 9274
rect 1104 9200 48852 9222
rect 2222 9160 2228 9172
rect 2183 9132 2228 9160
rect 2222 9120 2228 9132
rect 2280 9120 2286 9172
rect 17402 9160 17408 9172
rect 6886 9132 17408 9160
rect 2133 8959 2191 8965
rect 2133 8925 2145 8959
rect 2179 8956 2191 8959
rect 6886 8956 6914 9132
rect 17402 9120 17408 9132
rect 17460 9120 17466 9172
rect 22462 9160 22468 9172
rect 19260 9132 20300 9160
rect 18230 9092 18236 9104
rect 16868 9064 18236 9092
rect 16868 9033 16896 9064
rect 18230 9052 18236 9064
rect 18288 9052 18294 9104
rect 16853 9027 16911 9033
rect 16853 8993 16865 9027
rect 16899 8993 16911 9027
rect 17034 9024 17040 9036
rect 16995 8996 17040 9024
rect 16853 8987 16911 8993
rect 17034 8984 17040 8996
rect 17092 8984 17098 9036
rect 17310 9024 17316 9036
rect 17271 8996 17316 9024
rect 17310 8984 17316 8996
rect 17368 8984 17374 9036
rect 17586 8984 17592 9036
rect 17644 9024 17650 9036
rect 19260 9024 19288 9132
rect 17644 8996 19288 9024
rect 17644 8984 17650 8996
rect 19260 8965 19288 8996
rect 19518 8965 19524 8968
rect 2179 8928 6914 8956
rect 19245 8959 19303 8965
rect 2179 8925 2191 8928
rect 2133 8919 2191 8925
rect 19245 8925 19257 8959
rect 19291 8925 19303 8959
rect 19512 8956 19524 8965
rect 19479 8928 19524 8956
rect 19245 8919 19303 8925
rect 19512 8919 19524 8928
rect 19518 8916 19524 8919
rect 19576 8916 19582 8968
rect 20272 8888 20300 9132
rect 21284 9132 22468 9160
rect 21284 8965 21312 9132
rect 22462 9120 22468 9132
rect 22520 9120 22526 9172
rect 23385 9163 23443 9169
rect 23385 9129 23397 9163
rect 23431 9160 23443 9163
rect 24486 9160 24492 9172
rect 23431 9132 24492 9160
rect 23431 9129 23443 9132
rect 23385 9123 23443 9129
rect 24486 9120 24492 9132
rect 24544 9120 24550 9172
rect 25130 9120 25136 9172
rect 25188 9160 25194 9172
rect 25593 9163 25651 9169
rect 25593 9160 25605 9163
rect 25188 9132 25605 9160
rect 25188 9120 25194 9132
rect 25593 9129 25605 9132
rect 25639 9129 25651 9163
rect 25593 9123 25651 9129
rect 25866 9120 25872 9172
rect 25924 9160 25930 9172
rect 25924 9132 26372 9160
rect 25924 9120 25930 9132
rect 21361 9095 21419 9101
rect 21361 9061 21373 9095
rect 21407 9092 21419 9095
rect 22094 9092 22100 9104
rect 21407 9064 22100 9092
rect 21407 9061 21419 9064
rect 21361 9055 21419 9061
rect 22094 9052 22100 9064
rect 22152 9092 22158 9104
rect 22646 9092 22652 9104
rect 22152 9064 22652 9092
rect 22152 9052 22158 9064
rect 22646 9052 22652 9064
rect 22704 9052 22710 9104
rect 22738 9052 22744 9104
rect 22796 9092 22802 9104
rect 22796 9064 22841 9092
rect 22796 9052 22802 9064
rect 25038 9052 25044 9104
rect 25096 9052 25102 9104
rect 25222 9052 25228 9104
rect 25280 9092 25286 9104
rect 26344 9092 26372 9132
rect 26878 9120 26884 9172
rect 26936 9160 26942 9172
rect 47857 9163 47915 9169
rect 47857 9160 47869 9163
rect 26936 9132 47869 9160
rect 26936 9120 26942 9132
rect 47857 9129 47869 9132
rect 47903 9129 47915 9163
rect 47857 9123 47915 9129
rect 26973 9095 27031 9101
rect 26973 9092 26985 9095
rect 25280 9064 26234 9092
rect 26344 9064 26985 9092
rect 25280 9052 25286 9064
rect 21542 9024 21548 9036
rect 21503 8996 21548 9024
rect 21542 8984 21548 8996
rect 21600 8984 21606 9036
rect 21910 8984 21916 9036
rect 21968 9024 21974 9036
rect 22281 9027 22339 9033
rect 21968 8996 22232 9024
rect 21968 8984 21974 8996
rect 22204 8968 22232 8996
rect 22281 8993 22293 9027
rect 22327 9024 22339 9027
rect 23198 9024 23204 9036
rect 22327 8996 23204 9024
rect 22327 8993 22339 8996
rect 22281 8987 22339 8993
rect 23198 8984 23204 8996
rect 23256 8984 23262 9036
rect 24026 9024 24032 9036
rect 23768 8996 24032 9024
rect 21269 8959 21327 8965
rect 21269 8925 21281 8959
rect 21315 8925 21327 8959
rect 21269 8919 21327 8925
rect 22005 8959 22063 8965
rect 22005 8925 22017 8959
rect 22051 8925 22063 8959
rect 22186 8956 22192 8968
rect 22147 8928 22192 8956
rect 22005 8919 22063 8925
rect 21818 8888 21824 8900
rect 20272 8860 21824 8888
rect 21818 8848 21824 8860
rect 21876 8848 21882 8900
rect 19334 8780 19340 8832
rect 19392 8820 19398 8832
rect 20625 8823 20683 8829
rect 20625 8820 20637 8823
rect 19392 8792 20637 8820
rect 19392 8780 19398 8792
rect 20625 8789 20637 8792
rect 20671 8789 20683 8823
rect 20625 8783 20683 8789
rect 21545 8823 21603 8829
rect 21545 8789 21557 8823
rect 21591 8820 21603 8823
rect 22020 8820 22048 8919
rect 22186 8916 22192 8928
rect 22244 8916 22250 8968
rect 22370 8956 22376 8968
rect 22331 8928 22376 8956
rect 22370 8916 22376 8928
rect 22428 8916 22434 8968
rect 22462 8916 22468 8968
rect 22520 8956 22526 8968
rect 22557 8959 22615 8965
rect 22557 8956 22569 8959
rect 22520 8928 22569 8956
rect 22520 8916 22526 8928
rect 22557 8925 22569 8928
rect 22603 8925 22615 8959
rect 23566 8956 23572 8968
rect 23527 8928 23572 8956
rect 22557 8919 22615 8925
rect 23566 8916 23572 8928
rect 23624 8916 23630 8968
rect 23768 8965 23796 8996
rect 24026 8984 24032 8996
rect 24084 8984 24090 9036
rect 24302 8984 24308 9036
rect 24360 9024 24366 9036
rect 25056 9024 25084 9052
rect 24360 8996 25084 9024
rect 24360 8984 24366 8996
rect 23753 8959 23811 8965
rect 23753 8925 23765 8959
rect 23799 8925 23811 8959
rect 23753 8919 23811 8925
rect 23842 8916 23848 8968
rect 23900 8956 23906 8968
rect 24394 8956 24400 8968
rect 23900 8928 23945 8956
rect 24355 8928 24400 8956
rect 23900 8916 23906 8928
rect 24394 8916 24400 8928
rect 24452 8916 24458 8968
rect 24780 8965 24808 8996
rect 24581 8959 24639 8965
rect 24581 8925 24593 8959
rect 24627 8925 24639 8959
rect 24581 8919 24639 8925
rect 24673 8959 24731 8965
rect 24673 8925 24685 8959
rect 24719 8925 24731 8959
rect 24673 8919 24731 8925
rect 24765 8959 24823 8965
rect 24765 8925 24777 8959
rect 24811 8925 24823 8959
rect 24765 8919 24823 8925
rect 24960 8959 25018 8965
rect 24960 8925 24972 8959
rect 25006 8956 25018 8959
rect 25774 8956 25780 8968
rect 25006 8928 25084 8956
rect 25735 8928 25780 8956
rect 25006 8925 25018 8928
rect 24960 8919 25018 8925
rect 22646 8848 22652 8900
rect 22704 8888 22710 8900
rect 24596 8888 24624 8919
rect 22704 8860 24624 8888
rect 24688 8888 24716 8919
rect 24854 8888 24860 8900
rect 24688 8860 24860 8888
rect 22704 8848 22710 8860
rect 24854 8848 24860 8860
rect 24912 8848 24918 8900
rect 25056 8832 25084 8928
rect 25774 8916 25780 8928
rect 25832 8916 25838 8968
rect 25866 8916 25872 8968
rect 25924 8956 25930 8968
rect 26206 8965 26234 9064
rect 26973 9061 26985 9064
rect 27019 9092 27031 9095
rect 27062 9092 27068 9104
rect 27019 9064 27068 9092
rect 27019 9061 27031 9064
rect 26973 9055 27031 9061
rect 27062 9052 27068 9064
rect 27120 9052 27126 9104
rect 29454 9052 29460 9104
rect 29512 9092 29518 9104
rect 31294 9092 31300 9104
rect 29512 9064 31300 9092
rect 29512 9052 29518 9064
rect 27430 9024 27436 9036
rect 27391 8996 27436 9024
rect 27430 8984 27436 8996
rect 27488 8984 27494 9036
rect 31128 9024 31156 9064
rect 31294 9052 31300 9064
rect 31352 9052 31358 9104
rect 41690 9052 41696 9104
rect 41748 9092 41754 9104
rect 46842 9092 46848 9104
rect 41748 9064 46848 9092
rect 41748 9052 41754 9064
rect 46842 9052 46848 9064
rect 46900 9052 46906 9104
rect 32490 9024 32496 9036
rect 31036 8996 31156 9024
rect 31220 8996 32496 9024
rect 26053 8959 26111 8965
rect 25924 8928 25969 8956
rect 25924 8916 25930 8928
rect 26053 8925 26065 8959
rect 26099 8925 26111 8959
rect 26053 8919 26111 8925
rect 26155 8959 26234 8965
rect 26155 8925 26167 8959
rect 26201 8928 26234 8959
rect 30650 8956 30656 8968
rect 27172 8928 30656 8956
rect 26201 8925 26213 8928
rect 26155 8919 26213 8925
rect 25682 8848 25688 8900
rect 25740 8888 25746 8900
rect 26068 8888 26096 8919
rect 25740 8860 26096 8888
rect 25740 8848 25746 8860
rect 26326 8848 26332 8900
rect 26384 8888 26390 8900
rect 26605 8891 26663 8897
rect 26605 8888 26617 8891
rect 26384 8860 26617 8888
rect 26384 8848 26390 8860
rect 26605 8857 26617 8860
rect 26651 8857 26663 8891
rect 26605 8851 26663 8857
rect 26694 8848 26700 8900
rect 26752 8888 26758 8900
rect 26789 8891 26847 8897
rect 26789 8888 26801 8891
rect 26752 8860 26801 8888
rect 26752 8848 26758 8860
rect 26789 8857 26801 8860
rect 26835 8857 26847 8891
rect 26789 8851 26847 8857
rect 21591 8792 22048 8820
rect 21591 8789 21603 8792
rect 21545 8783 21603 8789
rect 22370 8780 22376 8832
rect 22428 8820 22434 8832
rect 24302 8820 24308 8832
rect 22428 8792 24308 8820
rect 22428 8780 22434 8792
rect 24302 8780 24308 8792
rect 24360 8780 24366 8832
rect 24394 8780 24400 8832
rect 24452 8820 24458 8832
rect 24578 8820 24584 8832
rect 24452 8792 24584 8820
rect 24452 8780 24458 8792
rect 24578 8780 24584 8792
rect 24636 8780 24642 8832
rect 25038 8780 25044 8832
rect 25096 8780 25102 8832
rect 25133 8823 25191 8829
rect 25133 8789 25145 8823
rect 25179 8820 25191 8823
rect 25222 8820 25228 8832
rect 25179 8792 25228 8820
rect 25179 8789 25191 8792
rect 25133 8783 25191 8789
rect 25222 8780 25228 8792
rect 25280 8780 25286 8832
rect 26050 8780 26056 8832
rect 26108 8820 26114 8832
rect 27172 8820 27200 8928
rect 30650 8916 30656 8928
rect 30708 8956 30714 8968
rect 31036 8965 31064 8996
rect 30883 8959 30941 8965
rect 30883 8956 30895 8959
rect 30708 8928 30895 8956
rect 30708 8916 30714 8928
rect 30883 8925 30895 8928
rect 30929 8925 30941 8959
rect 30883 8919 30941 8925
rect 31021 8959 31079 8965
rect 31021 8925 31033 8959
rect 31067 8925 31079 8959
rect 31021 8919 31079 8925
rect 31118 8959 31176 8965
rect 31118 8925 31130 8959
rect 31164 8956 31176 8959
rect 31220 8956 31248 8996
rect 32490 8984 32496 8996
rect 32548 8984 32554 9036
rect 31164 8928 31248 8956
rect 31297 8959 31355 8965
rect 31164 8925 31176 8928
rect 31118 8919 31176 8925
rect 31297 8925 31309 8959
rect 31343 8956 31355 8959
rect 31478 8956 31484 8968
rect 31343 8928 31484 8956
rect 31343 8925 31355 8928
rect 31297 8919 31355 8925
rect 31478 8916 31484 8928
rect 31536 8916 31542 8968
rect 27700 8891 27758 8897
rect 27700 8857 27712 8891
rect 27746 8888 27758 8891
rect 27890 8888 27896 8900
rect 27746 8860 27896 8888
rect 27746 8857 27758 8860
rect 27700 8851 27758 8857
rect 27890 8848 27896 8860
rect 27948 8848 27954 8900
rect 47762 8888 47768 8900
rect 47723 8860 47768 8888
rect 47762 8848 47768 8860
rect 47820 8848 47826 8900
rect 26108 8792 27200 8820
rect 26108 8780 26114 8792
rect 27246 8780 27252 8832
rect 27304 8820 27310 8832
rect 28813 8823 28871 8829
rect 28813 8820 28825 8823
rect 27304 8792 28825 8820
rect 27304 8780 27310 8792
rect 28813 8789 28825 8792
rect 28859 8789 28871 8823
rect 30650 8820 30656 8832
rect 30611 8792 30656 8820
rect 28813 8783 28871 8789
rect 30650 8780 30656 8792
rect 30708 8780 30714 8832
rect 1104 8730 48852 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 48852 8730
rect 1104 8656 48852 8678
rect 6886 8588 23520 8616
rect 2225 8551 2283 8557
rect 2225 8517 2237 8551
rect 2271 8548 2283 8551
rect 6886 8548 6914 8588
rect 2271 8520 6914 8548
rect 22088 8551 22146 8557
rect 2271 8517 2283 8520
rect 2225 8511 2283 8517
rect 22088 8517 22100 8551
rect 22134 8548 22146 8551
rect 22738 8548 22744 8560
rect 22134 8520 22744 8548
rect 22134 8517 22146 8520
rect 22088 8511 22146 8517
rect 22738 8508 22744 8520
rect 22796 8508 22802 8560
rect 23492 8548 23520 8588
rect 23566 8576 23572 8628
rect 23624 8616 23630 8628
rect 24029 8619 24087 8625
rect 24029 8616 24041 8619
rect 23624 8588 24041 8616
rect 23624 8576 23630 8588
rect 24029 8585 24041 8588
rect 24075 8616 24087 8619
rect 24075 8588 24348 8616
rect 24075 8585 24087 8588
rect 24029 8579 24087 8585
rect 24210 8548 24216 8560
rect 23492 8520 24216 8548
rect 24210 8508 24216 8520
rect 24268 8508 24274 8560
rect 24320 8548 24348 8588
rect 24394 8576 24400 8628
rect 24452 8616 24458 8628
rect 24452 8588 24497 8616
rect 24452 8576 24458 8588
rect 24762 8576 24768 8628
rect 24820 8616 24826 8628
rect 25685 8619 25743 8625
rect 25685 8616 25697 8619
rect 24820 8588 25697 8616
rect 24820 8576 24826 8588
rect 25685 8585 25697 8588
rect 25731 8585 25743 8619
rect 25685 8579 25743 8585
rect 27614 8576 27620 8628
rect 27672 8616 27678 8628
rect 27890 8616 27896 8628
rect 27672 8588 27752 8616
rect 27851 8588 27896 8616
rect 27672 8576 27678 8588
rect 24489 8551 24547 8557
rect 24320 8520 24440 8548
rect 1854 8480 1860 8492
rect 1815 8452 1860 8480
rect 1854 8440 1860 8452
rect 1912 8440 1918 8492
rect 17586 8480 17592 8492
rect 17547 8452 17592 8480
rect 17586 8440 17592 8452
rect 17644 8440 17650 8492
rect 17856 8483 17914 8489
rect 17856 8449 17868 8483
rect 17902 8480 17914 8483
rect 19242 8480 19248 8492
rect 17902 8452 19248 8480
rect 17902 8449 17914 8452
rect 17856 8443 17914 8449
rect 19242 8440 19248 8452
rect 19300 8440 19306 8492
rect 19334 8372 19340 8424
rect 19392 8412 19398 8424
rect 19429 8415 19487 8421
rect 19429 8412 19441 8415
rect 19392 8384 19441 8412
rect 19392 8372 19398 8384
rect 19429 8381 19441 8384
rect 19475 8381 19487 8415
rect 19429 8375 19487 8381
rect 19613 8415 19671 8421
rect 19613 8381 19625 8415
rect 19659 8381 19671 8415
rect 21266 8412 21272 8424
rect 21227 8384 21272 8412
rect 19613 8375 19671 8381
rect 18966 8276 18972 8288
rect 18927 8248 18972 8276
rect 18966 8236 18972 8248
rect 19024 8236 19030 8288
rect 19334 8236 19340 8288
rect 19392 8276 19398 8288
rect 19628 8276 19656 8375
rect 21266 8372 21272 8384
rect 21324 8372 21330 8424
rect 21818 8412 21824 8424
rect 21779 8384 21824 8412
rect 21818 8372 21824 8384
rect 21876 8372 21882 8424
rect 24412 8412 24440 8520
rect 24489 8517 24501 8551
rect 24535 8548 24547 8551
rect 24854 8548 24860 8560
rect 24535 8520 24860 8548
rect 24535 8517 24547 8520
rect 24489 8511 24547 8517
rect 24854 8508 24860 8520
rect 24912 8548 24918 8560
rect 24912 8520 25544 8548
rect 24912 8508 24918 8520
rect 25130 8440 25136 8492
rect 25188 8480 25194 8492
rect 25516 8489 25544 8520
rect 25225 8483 25283 8489
rect 25225 8480 25237 8483
rect 25188 8452 25237 8480
rect 25188 8440 25194 8452
rect 25225 8449 25237 8452
rect 25271 8449 25283 8483
rect 25225 8443 25283 8449
rect 25501 8483 25559 8489
rect 25501 8449 25513 8483
rect 25547 8449 25559 8483
rect 27154 8480 27160 8492
rect 27115 8452 27160 8480
rect 25501 8443 25559 8449
rect 27154 8440 27160 8452
rect 27212 8440 27218 8492
rect 27341 8483 27399 8489
rect 27341 8449 27353 8483
rect 27387 8480 27399 8483
rect 27614 8480 27620 8492
rect 27387 8452 27620 8480
rect 27387 8449 27399 8452
rect 27341 8443 27399 8449
rect 27614 8440 27620 8452
rect 27672 8440 27678 8492
rect 27724 8489 27752 8588
rect 27890 8576 27896 8588
rect 27948 8576 27954 8628
rect 29454 8576 29460 8628
rect 29512 8576 29518 8628
rect 31570 8616 31576 8628
rect 31531 8588 31576 8616
rect 31570 8576 31576 8588
rect 31628 8576 31634 8628
rect 32490 8616 32496 8628
rect 32451 8588 32496 8616
rect 32490 8576 32496 8588
rect 32548 8576 32554 8628
rect 29472 8495 29500 8576
rect 30460 8551 30518 8557
rect 29748 8520 30374 8548
rect 29454 8489 29512 8495
rect 29748 8492 29776 8520
rect 27709 8483 27767 8489
rect 27709 8449 27721 8483
rect 27755 8449 27767 8483
rect 27709 8443 27767 8449
rect 29365 8483 29423 8489
rect 29365 8449 29377 8483
rect 29411 8449 29423 8483
rect 29454 8455 29466 8489
rect 29500 8455 29512 8489
rect 29454 8449 29512 8455
rect 29549 8486 29607 8492
rect 29549 8452 29561 8486
rect 29595 8452 29607 8486
rect 29730 8480 29736 8492
rect 29691 8452 29736 8480
rect 29365 8443 29423 8449
rect 29549 8446 29607 8452
rect 24412 8384 24532 8412
rect 24504 8344 24532 8384
rect 24578 8372 24584 8424
rect 24636 8412 24642 8424
rect 25314 8412 25320 8424
rect 24636 8384 24681 8412
rect 25275 8384 25320 8412
rect 24636 8372 24642 8384
rect 25314 8372 25320 8384
rect 25372 8372 25378 8424
rect 27246 8372 27252 8424
rect 27304 8412 27310 8424
rect 27433 8415 27491 8421
rect 27433 8412 27445 8415
rect 27304 8384 27445 8412
rect 27304 8372 27310 8384
rect 27433 8381 27445 8384
rect 27479 8381 27491 8415
rect 27433 8375 27491 8381
rect 27522 8372 27528 8424
rect 27580 8412 27586 8424
rect 27580 8384 27625 8412
rect 27580 8372 27586 8384
rect 24946 8344 24952 8356
rect 24504 8316 24952 8344
rect 24946 8304 24952 8316
rect 25004 8304 25010 8356
rect 25056 8316 25360 8344
rect 23198 8276 23204 8288
rect 19392 8248 19656 8276
rect 23111 8248 23204 8276
rect 19392 8236 19398 8248
rect 23198 8236 23204 8248
rect 23256 8276 23262 8288
rect 25056 8276 25084 8316
rect 25332 8285 25360 8316
rect 26050 8304 26056 8356
rect 26108 8344 26114 8356
rect 29380 8344 29408 8443
rect 29564 8356 29592 8446
rect 29730 8440 29736 8452
rect 29788 8440 29794 8492
rect 30190 8480 30196 8492
rect 30151 8452 30196 8480
rect 30190 8440 30196 8452
rect 30248 8440 30254 8492
rect 30346 8480 30374 8520
rect 30460 8517 30472 8551
rect 30506 8548 30518 8551
rect 30650 8548 30656 8560
rect 30506 8520 30656 8548
rect 30506 8517 30518 8520
rect 30460 8511 30518 8517
rect 30650 8508 30656 8520
rect 30708 8508 30714 8560
rect 31478 8480 31484 8492
rect 30346 8452 31484 8480
rect 31478 8440 31484 8452
rect 31536 8440 31542 8492
rect 32122 8480 32128 8492
rect 32083 8452 32128 8480
rect 32122 8440 32128 8452
rect 32180 8440 32186 8492
rect 32309 8483 32367 8489
rect 32309 8449 32321 8483
rect 32355 8449 32367 8483
rect 47854 8480 47860 8492
rect 47815 8452 47860 8480
rect 32309 8443 32367 8449
rect 31570 8372 31576 8424
rect 31628 8412 31634 8424
rect 32324 8412 32352 8443
rect 47854 8440 47860 8452
rect 47912 8440 47918 8492
rect 31628 8384 32352 8412
rect 31628 8372 31634 8384
rect 26108 8316 29408 8344
rect 26108 8304 26114 8316
rect 29546 8304 29552 8356
rect 29604 8304 29610 8356
rect 33042 8304 33048 8356
rect 33100 8344 33106 8356
rect 48041 8347 48099 8353
rect 48041 8344 48053 8347
rect 33100 8316 48053 8344
rect 33100 8304 33106 8316
rect 48041 8313 48053 8316
rect 48087 8313 48099 8347
rect 48041 8307 48099 8313
rect 23256 8248 25084 8276
rect 25317 8279 25375 8285
rect 23256 8236 23262 8248
rect 25317 8245 25329 8279
rect 25363 8245 25375 8279
rect 25317 8239 25375 8245
rect 25406 8236 25412 8288
rect 25464 8276 25470 8288
rect 25958 8276 25964 8288
rect 25464 8248 25964 8276
rect 25464 8236 25470 8248
rect 25958 8236 25964 8248
rect 26016 8276 26022 8288
rect 26234 8276 26240 8288
rect 26016 8248 26240 8276
rect 26016 8236 26022 8248
rect 26234 8236 26240 8248
rect 26292 8236 26298 8288
rect 29086 8276 29092 8288
rect 29047 8248 29092 8276
rect 29086 8236 29092 8248
rect 29144 8236 29150 8288
rect 29178 8236 29184 8288
rect 29236 8276 29242 8288
rect 38010 8276 38016 8288
rect 29236 8248 38016 8276
rect 29236 8236 29242 8248
rect 38010 8236 38016 8248
rect 38068 8236 38074 8288
rect 1104 8186 48852 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 48852 8186
rect 1104 8112 48852 8134
rect 6886 8044 19840 8072
rect 2133 7939 2191 7945
rect 2133 7905 2145 7939
rect 2179 7936 2191 7939
rect 6886 7936 6914 8044
rect 18782 7964 18788 8016
rect 18840 8004 18846 8016
rect 19812 8004 19840 8044
rect 21266 8032 21272 8084
rect 21324 8072 21330 8084
rect 29178 8072 29184 8084
rect 21324 8044 29184 8072
rect 21324 8032 21330 8044
rect 29178 8032 29184 8044
rect 29236 8032 29242 8084
rect 29546 8032 29552 8084
rect 29604 8072 29610 8084
rect 30009 8075 30067 8081
rect 30009 8072 30021 8075
rect 29604 8044 30021 8072
rect 29604 8032 29610 8044
rect 30009 8041 30021 8044
rect 30055 8041 30067 8075
rect 30009 8035 30067 8041
rect 30098 8032 30104 8084
rect 30156 8072 30162 8084
rect 32122 8072 32128 8084
rect 30156 8044 32128 8072
rect 30156 8032 30162 8044
rect 32122 8032 32128 8044
rect 32180 8032 32186 8084
rect 45646 8072 45652 8084
rect 41386 8044 45652 8072
rect 21450 8004 21456 8016
rect 18840 7976 19748 8004
rect 19812 7976 21456 8004
rect 18840 7964 18846 7976
rect 18966 7936 18972 7948
rect 2179 7908 6914 7936
rect 18524 7908 18972 7936
rect 2179 7905 2191 7908
rect 2133 7899 2191 7905
rect 18046 7828 18052 7880
rect 18104 7868 18110 7880
rect 18524 7877 18552 7908
rect 18966 7896 18972 7908
rect 19024 7936 19030 7948
rect 19720 7945 19748 7976
rect 21450 7964 21456 7976
rect 21508 7964 21514 8016
rect 22094 7964 22100 8016
rect 22152 8004 22158 8016
rect 22152 7976 22197 8004
rect 22152 7964 22158 7976
rect 26234 7964 26240 8016
rect 26292 8004 26298 8016
rect 26605 8007 26663 8013
rect 26605 8004 26617 8007
rect 26292 7976 26617 8004
rect 26292 7964 26298 7976
rect 26605 7973 26617 7976
rect 26651 7973 26663 8007
rect 41386 8004 41414 8044
rect 45646 8032 45652 8044
rect 45704 8032 45710 8084
rect 26605 7967 26663 7973
rect 27540 7976 41414 8004
rect 19245 7939 19303 7945
rect 19245 7936 19257 7939
rect 19024 7908 19257 7936
rect 19024 7896 19030 7908
rect 19245 7905 19257 7908
rect 19291 7905 19303 7939
rect 19245 7899 19303 7905
rect 19705 7939 19763 7945
rect 19705 7905 19717 7939
rect 19751 7905 19763 7939
rect 19705 7899 19763 7905
rect 22741 7939 22799 7945
rect 22741 7905 22753 7939
rect 22787 7936 22799 7939
rect 23658 7936 23664 7948
rect 22787 7908 23664 7936
rect 22787 7905 22799 7908
rect 22741 7899 22799 7905
rect 23658 7896 23664 7908
rect 23716 7936 23722 7948
rect 24578 7936 24584 7948
rect 23716 7908 24584 7936
rect 23716 7896 23722 7908
rect 24578 7896 24584 7908
rect 24636 7896 24642 7948
rect 18325 7871 18383 7877
rect 18325 7868 18337 7871
rect 18104 7840 18337 7868
rect 18104 7828 18110 7840
rect 18325 7837 18337 7840
rect 18371 7837 18383 7871
rect 18325 7831 18383 7837
rect 18509 7871 18567 7877
rect 18509 7837 18521 7871
rect 18555 7837 18567 7871
rect 18509 7831 18567 7837
rect 22557 7871 22615 7877
rect 22557 7837 22569 7871
rect 22603 7868 22615 7871
rect 23198 7868 23204 7880
rect 22603 7840 23204 7868
rect 22603 7837 22615 7840
rect 22557 7831 22615 7837
rect 23198 7828 23204 7840
rect 23256 7828 23262 7880
rect 23474 7828 23480 7880
rect 23532 7868 23538 7880
rect 24394 7868 24400 7880
rect 23532 7840 24400 7868
rect 23532 7828 23538 7840
rect 24394 7828 24400 7840
rect 24452 7868 24458 7880
rect 25225 7871 25283 7877
rect 25225 7868 25237 7871
rect 24452 7840 25237 7868
rect 24452 7828 24458 7840
rect 25225 7837 25237 7840
rect 25271 7868 25283 7871
rect 27430 7868 27436 7880
rect 25271 7840 27436 7868
rect 25271 7837 25283 7840
rect 25225 7831 25283 7837
rect 27430 7828 27436 7840
rect 27488 7828 27494 7880
rect 1854 7800 1860 7812
rect 1815 7772 1860 7800
rect 1854 7760 1860 7772
rect 1912 7760 1918 7812
rect 18598 7760 18604 7812
rect 18656 7800 18662 7812
rect 25498 7809 25504 7812
rect 19429 7803 19487 7809
rect 19429 7800 19441 7803
rect 18656 7772 19441 7800
rect 18656 7760 18662 7772
rect 19429 7769 19441 7772
rect 19475 7769 19487 7803
rect 25492 7800 25504 7809
rect 19429 7763 19487 7769
rect 22066 7772 22692 7800
rect 25459 7772 25504 7800
rect 18690 7732 18696 7744
rect 18651 7704 18696 7732
rect 18690 7692 18696 7704
rect 18748 7692 18754 7744
rect 20530 7692 20536 7744
rect 20588 7732 20594 7744
rect 22066 7732 22094 7772
rect 22462 7732 22468 7744
rect 20588 7704 22094 7732
rect 22423 7704 22468 7732
rect 20588 7692 20594 7704
rect 22462 7692 22468 7704
rect 22520 7692 22526 7744
rect 22664 7732 22692 7772
rect 25492 7763 25504 7772
rect 25498 7760 25504 7763
rect 25556 7760 25562 7812
rect 27540 7800 27568 7976
rect 30469 7939 30527 7945
rect 30469 7905 30481 7939
rect 30515 7936 30527 7939
rect 31570 7936 31576 7948
rect 30515 7908 31576 7936
rect 30515 7905 30527 7908
rect 30469 7899 30527 7905
rect 31570 7896 31576 7908
rect 31628 7896 31634 7948
rect 31849 7939 31907 7945
rect 31849 7905 31861 7939
rect 31895 7905 31907 7939
rect 31849 7899 31907 7905
rect 29641 7871 29699 7877
rect 29641 7837 29653 7871
rect 29687 7868 29699 7871
rect 30098 7868 30104 7880
rect 29687 7840 30104 7868
rect 29687 7837 29699 7840
rect 29641 7831 29699 7837
rect 30098 7828 30104 7840
rect 30156 7828 30162 7880
rect 26528 7772 27568 7800
rect 29825 7803 29883 7809
rect 26528 7732 26556 7772
rect 29825 7769 29837 7803
rect 29871 7800 29883 7803
rect 30282 7800 30288 7812
rect 29871 7772 30288 7800
rect 29871 7769 29883 7772
rect 29825 7763 29883 7769
rect 30282 7760 30288 7772
rect 30340 7760 30346 7812
rect 30653 7803 30711 7809
rect 30653 7769 30665 7803
rect 30699 7800 30711 7803
rect 30926 7800 30932 7812
rect 30699 7772 30932 7800
rect 30699 7769 30711 7772
rect 30653 7763 30711 7769
rect 30926 7760 30932 7772
rect 30984 7760 30990 7812
rect 22664 7704 26556 7732
rect 29638 7692 29644 7744
rect 29696 7732 29702 7744
rect 31864 7732 31892 7899
rect 46290 7868 46296 7880
rect 46251 7840 46296 7868
rect 46290 7828 46296 7840
rect 46348 7828 46354 7880
rect 46477 7803 46535 7809
rect 46477 7769 46489 7803
rect 46523 7800 46535 7803
rect 46750 7800 46756 7812
rect 46523 7772 46756 7800
rect 46523 7769 46535 7772
rect 46477 7763 46535 7769
rect 46750 7760 46756 7772
rect 46808 7760 46814 7812
rect 48130 7800 48136 7812
rect 48091 7772 48136 7800
rect 48130 7760 48136 7772
rect 48188 7760 48194 7812
rect 29696 7704 31892 7732
rect 29696 7692 29702 7704
rect 1104 7642 48852 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 48852 7642
rect 1104 7568 48852 7590
rect 18509 7531 18567 7537
rect 18509 7497 18521 7531
rect 18555 7528 18567 7531
rect 18598 7528 18604 7540
rect 18555 7500 18604 7528
rect 18555 7497 18567 7500
rect 18509 7491 18567 7497
rect 18598 7488 18604 7500
rect 18656 7488 18662 7540
rect 19242 7488 19248 7540
rect 19300 7528 19306 7540
rect 19337 7531 19395 7537
rect 19337 7528 19349 7531
rect 19300 7500 19349 7528
rect 19300 7488 19306 7500
rect 19337 7497 19349 7500
rect 19383 7497 19395 7531
rect 19978 7528 19984 7540
rect 19337 7491 19395 7497
rect 19720 7500 19984 7528
rect 18690 7420 18696 7472
rect 18748 7460 18754 7472
rect 18748 7432 19334 7460
rect 18748 7420 18754 7432
rect 17954 7352 17960 7404
rect 18012 7392 18018 7404
rect 18414 7392 18420 7404
rect 18012 7364 18420 7392
rect 18012 7352 18018 7364
rect 18414 7352 18420 7364
rect 18472 7352 18478 7404
rect 19306 7324 19334 7432
rect 19610 7392 19616 7404
rect 19571 7364 19616 7392
rect 19610 7352 19616 7364
rect 19668 7352 19674 7404
rect 19720 7401 19748 7500
rect 19978 7488 19984 7500
rect 20036 7488 20042 7540
rect 24854 7528 24860 7540
rect 22066 7500 24716 7528
rect 24815 7500 24860 7528
rect 19718 7395 19776 7401
rect 19718 7361 19730 7395
rect 19764 7361 19776 7395
rect 19718 7355 19776 7361
rect 19818 7395 19876 7401
rect 19818 7361 19830 7395
rect 19864 7392 19876 7395
rect 19981 7395 20039 7401
rect 19864 7364 19932 7392
rect 19864 7361 19876 7364
rect 19818 7355 19876 7361
rect 19904 7324 19932 7364
rect 19981 7361 19993 7395
rect 20027 7392 20039 7395
rect 22066 7392 22094 7500
rect 24688 7460 24716 7500
rect 24854 7488 24860 7500
rect 24912 7488 24918 7540
rect 27798 7488 27804 7540
rect 27856 7528 27862 7540
rect 28074 7528 28080 7540
rect 27856 7500 28080 7528
rect 27856 7488 27862 7500
rect 28074 7488 28080 7500
rect 28132 7488 28138 7540
rect 29730 7528 29736 7540
rect 29012 7500 29736 7528
rect 29012 7460 29040 7500
rect 29730 7488 29736 7500
rect 29788 7488 29794 7540
rect 30926 7528 30932 7540
rect 30887 7500 30932 7528
rect 30926 7488 30932 7500
rect 30984 7488 30990 7540
rect 46750 7528 46756 7540
rect 46711 7500 46756 7528
rect 46750 7488 46756 7500
rect 46808 7488 46814 7540
rect 24688 7432 29040 7460
rect 29086 7420 29092 7472
rect 29144 7460 29150 7472
rect 29242 7463 29300 7469
rect 29242 7460 29254 7463
rect 29144 7432 29254 7460
rect 29144 7420 29150 7432
rect 29242 7429 29254 7432
rect 29288 7429 29300 7463
rect 29242 7423 29300 7429
rect 46290 7420 46296 7472
rect 46348 7460 46354 7472
rect 46348 7432 47808 7460
rect 46348 7420 46354 7432
rect 23474 7392 23480 7404
rect 20027 7364 22094 7392
rect 23435 7364 23480 7392
rect 20027 7361 20039 7364
rect 19981 7355 20039 7361
rect 23474 7352 23480 7364
rect 23532 7352 23538 7404
rect 23744 7395 23802 7401
rect 23744 7361 23756 7395
rect 23790 7392 23802 7395
rect 25222 7392 25228 7404
rect 23790 7364 25228 7392
rect 23790 7361 23802 7364
rect 23744 7355 23802 7361
rect 25222 7352 25228 7364
rect 25280 7352 25286 7404
rect 28353 7395 28411 7401
rect 28353 7361 28365 7395
rect 28399 7392 28411 7395
rect 30837 7395 30895 7401
rect 30837 7392 30849 7395
rect 28399 7364 30849 7392
rect 28399 7361 28411 7364
rect 28353 7355 28411 7361
rect 30837 7361 30849 7364
rect 30883 7392 30895 7395
rect 32582 7392 32588 7404
rect 30883 7364 32588 7392
rect 30883 7361 30895 7364
rect 30837 7355 30895 7361
rect 32582 7352 32588 7364
rect 32640 7352 32646 7404
rect 45554 7352 45560 7404
rect 45612 7392 45618 7404
rect 47780 7401 47808 7432
rect 46661 7395 46719 7401
rect 46661 7392 46673 7395
rect 45612 7364 46673 7392
rect 45612 7352 45618 7364
rect 46661 7361 46673 7364
rect 46707 7361 46719 7395
rect 46661 7355 46719 7361
rect 47765 7395 47823 7401
rect 47765 7361 47777 7395
rect 47811 7361 47823 7395
rect 47765 7355 47823 7361
rect 19306 7296 19932 7324
rect 27430 7284 27436 7336
rect 27488 7324 27494 7336
rect 28997 7327 29055 7333
rect 28997 7324 29009 7327
rect 27488 7296 29009 7324
rect 27488 7284 27494 7296
rect 28997 7293 29009 7296
rect 29043 7293 29055 7327
rect 28997 7287 29055 7293
rect 19058 7216 19064 7268
rect 19116 7256 19122 7268
rect 20346 7256 20352 7268
rect 19116 7228 20352 7256
rect 19116 7216 19122 7228
rect 20346 7216 20352 7228
rect 20404 7216 20410 7268
rect 2038 7148 2044 7200
rect 2096 7188 2102 7200
rect 2317 7191 2375 7197
rect 2317 7188 2329 7191
rect 2096 7160 2329 7188
rect 2096 7148 2102 7160
rect 2317 7157 2329 7160
rect 2363 7157 2375 7191
rect 2317 7151 2375 7157
rect 28445 7191 28503 7197
rect 28445 7157 28457 7191
rect 28491 7188 28503 7191
rect 29730 7188 29736 7200
rect 28491 7160 29736 7188
rect 28491 7157 28503 7160
rect 28445 7151 28503 7157
rect 29730 7148 29736 7160
rect 29788 7148 29794 7200
rect 30282 7148 30288 7200
rect 30340 7188 30346 7200
rect 30377 7191 30435 7197
rect 30377 7188 30389 7191
rect 30340 7160 30389 7188
rect 30340 7148 30346 7160
rect 30377 7157 30389 7160
rect 30423 7157 30435 7191
rect 30377 7151 30435 7157
rect 1104 7098 48852 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 48852 7098
rect 1104 7024 48852 7046
rect 19334 6944 19340 6996
rect 19392 6984 19398 6996
rect 19429 6987 19487 6993
rect 19429 6984 19441 6987
rect 19392 6956 19441 6984
rect 19392 6944 19398 6956
rect 19429 6953 19441 6956
rect 19475 6953 19487 6987
rect 19429 6947 19487 6953
rect 30282 6916 30288 6928
rect 29564 6888 30288 6916
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 29564 6857 29592 6888
rect 30282 6876 30288 6888
rect 30340 6876 30346 6928
rect 29549 6851 29607 6857
rect 3476 6820 26740 6848
rect 3476 6808 3482 6820
rect 2961 6783 3019 6789
rect 2961 6749 2973 6783
rect 3007 6780 3019 6783
rect 17218 6780 17224 6792
rect 3007 6752 17224 6780
rect 3007 6749 3019 6752
rect 2961 6743 3019 6749
rect 17218 6740 17224 6752
rect 17276 6780 17282 6792
rect 17494 6780 17500 6792
rect 17276 6752 17500 6780
rect 17276 6740 17282 6752
rect 17494 6740 17500 6752
rect 17552 6740 17558 6792
rect 18414 6740 18420 6792
rect 18472 6780 18478 6792
rect 19337 6783 19395 6789
rect 19337 6780 19349 6783
rect 18472 6752 19349 6780
rect 18472 6740 18478 6752
rect 19337 6749 19349 6752
rect 19383 6749 19395 6783
rect 19337 6743 19395 6749
rect 19610 6740 19616 6792
rect 19668 6780 19674 6792
rect 21085 6783 21143 6789
rect 21085 6780 21097 6783
rect 19668 6752 21097 6780
rect 19668 6740 19674 6752
rect 21085 6749 21097 6752
rect 21131 6780 21143 6783
rect 22462 6780 22468 6792
rect 21131 6752 22468 6780
rect 21131 6749 21143 6752
rect 21085 6743 21143 6749
rect 22462 6740 22468 6752
rect 22520 6740 22526 6792
rect 20898 6712 20904 6724
rect 20859 6684 20904 6712
rect 20898 6672 20904 6684
rect 20956 6672 20962 6724
rect 26712 6712 26740 6820
rect 29549 6817 29561 6851
rect 29595 6817 29607 6851
rect 29730 6848 29736 6860
rect 29691 6820 29736 6848
rect 29549 6811 29607 6817
rect 29730 6808 29736 6820
rect 29788 6808 29794 6860
rect 30929 6851 30987 6857
rect 30929 6817 30941 6851
rect 30975 6817 30987 6851
rect 30929 6811 30987 6817
rect 30944 6712 30972 6811
rect 44910 6808 44916 6860
rect 44968 6848 44974 6860
rect 45649 6851 45707 6857
rect 45649 6848 45661 6851
rect 44968 6820 45661 6848
rect 44968 6808 44974 6820
rect 45649 6817 45661 6820
rect 45695 6817 45707 6851
rect 46842 6848 46848 6860
rect 46803 6820 46848 6848
rect 45649 6811 45707 6817
rect 46842 6808 46848 6820
rect 46900 6808 46906 6860
rect 26712 6684 30972 6712
rect 45833 6715 45891 6721
rect 45833 6681 45845 6715
rect 45879 6712 45891 6715
rect 45922 6712 45928 6724
rect 45879 6684 45928 6712
rect 45879 6681 45891 6684
rect 45833 6675 45891 6681
rect 45922 6672 45928 6684
rect 45980 6672 45986 6724
rect 2222 6604 2228 6656
rect 2280 6644 2286 6656
rect 3053 6647 3111 6653
rect 3053 6644 3065 6647
rect 2280 6616 3065 6644
rect 2280 6604 2286 6616
rect 3053 6613 3065 6616
rect 3099 6613 3111 6647
rect 3053 6607 3111 6613
rect 19426 6604 19432 6656
rect 19484 6644 19490 6656
rect 20162 6644 20168 6656
rect 19484 6616 20168 6644
rect 19484 6604 19490 6616
rect 20162 6604 20168 6616
rect 20220 6604 20226 6656
rect 21082 6604 21088 6656
rect 21140 6644 21146 6656
rect 21269 6647 21327 6653
rect 21269 6644 21281 6647
rect 21140 6616 21281 6644
rect 21140 6604 21146 6616
rect 21269 6613 21281 6616
rect 21315 6613 21327 6647
rect 21269 6607 21327 6613
rect 1104 6554 48852 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 48852 6554
rect 1104 6480 48852 6502
rect 20898 6440 20904 6452
rect 20811 6412 20904 6440
rect 2222 6372 2228 6384
rect 2183 6344 2228 6372
rect 2222 6332 2228 6344
rect 2280 6332 2286 6384
rect 20824 6381 20852 6412
rect 20898 6400 20904 6412
rect 20956 6440 20962 6452
rect 45922 6440 45928 6452
rect 20956 6412 24164 6440
rect 45883 6412 45928 6440
rect 20956 6400 20962 6412
rect 24136 6384 24164 6412
rect 45922 6400 45928 6412
rect 45980 6400 45986 6452
rect 20809 6375 20867 6381
rect 20809 6341 20821 6375
rect 20855 6341 20867 6375
rect 20990 6372 20996 6384
rect 20951 6344 20996 6372
rect 20809 6335 20867 6341
rect 20990 6332 20996 6344
rect 21048 6372 21054 6384
rect 22002 6372 22008 6384
rect 21048 6344 22008 6372
rect 21048 6332 21054 6344
rect 22002 6332 22008 6344
rect 22060 6332 22066 6384
rect 24118 6332 24124 6384
rect 24176 6372 24182 6384
rect 27617 6375 27675 6381
rect 27617 6372 27629 6375
rect 24176 6344 27629 6372
rect 24176 6332 24182 6344
rect 27617 6341 27629 6344
rect 27663 6372 27675 6375
rect 28626 6372 28632 6384
rect 27663 6344 28632 6372
rect 27663 6341 27675 6344
rect 27617 6335 27675 6341
rect 28626 6332 28632 6344
rect 28684 6332 28690 6384
rect 2038 6304 2044 6316
rect 1999 6276 2044 6304
rect 2038 6264 2044 6276
rect 2096 6264 2102 6316
rect 23566 6264 23572 6316
rect 23624 6304 23630 6316
rect 23661 6307 23719 6313
rect 23661 6304 23673 6307
rect 23624 6276 23673 6304
rect 23624 6264 23630 6276
rect 23661 6273 23673 6276
rect 23707 6273 23719 6307
rect 23661 6267 23719 6273
rect 23753 6307 23811 6313
rect 23753 6273 23765 6307
rect 23799 6273 23811 6307
rect 23753 6267 23811 6273
rect 2774 6236 2780 6248
rect 2735 6208 2780 6236
rect 2774 6196 2780 6208
rect 2832 6196 2838 6248
rect 23768 6236 23796 6267
rect 23842 6264 23848 6316
rect 23900 6304 23906 6316
rect 23900 6276 23945 6304
rect 23900 6264 23906 6276
rect 24026 6264 24032 6316
rect 24084 6304 24090 6316
rect 24084 6276 24129 6304
rect 24084 6264 24090 6276
rect 24486 6264 24492 6316
rect 24544 6304 24550 6316
rect 27798 6304 27804 6316
rect 24544 6276 27804 6304
rect 24544 6264 24550 6276
rect 27798 6264 27804 6276
rect 27856 6264 27862 6316
rect 29914 6264 29920 6316
rect 29972 6304 29978 6316
rect 35618 6304 35624 6316
rect 29972 6276 35624 6304
rect 29972 6264 29978 6276
rect 35618 6264 35624 6276
rect 35676 6264 35682 6316
rect 45830 6304 45836 6316
rect 45791 6276 45836 6304
rect 45830 6264 45836 6276
rect 45888 6264 45894 6316
rect 24210 6236 24216 6248
rect 23768 6208 24216 6236
rect 24210 6196 24216 6208
rect 24268 6196 24274 6248
rect 2406 6128 2412 6180
rect 2464 6168 2470 6180
rect 2682 6168 2688 6180
rect 2464 6140 2688 6168
rect 2464 6128 2470 6140
rect 2682 6128 2688 6140
rect 2740 6168 2746 6180
rect 39482 6168 39488 6180
rect 2740 6140 39488 6168
rect 2740 6128 2746 6140
rect 39482 6128 39488 6140
rect 39540 6128 39546 6180
rect 1578 6100 1584 6112
rect 1539 6072 1584 6100
rect 1578 6060 1584 6072
rect 1636 6060 1642 6112
rect 21177 6103 21235 6109
rect 21177 6069 21189 6103
rect 21223 6100 21235 6103
rect 22922 6100 22928 6112
rect 21223 6072 22928 6100
rect 21223 6069 21235 6072
rect 21177 6063 21235 6069
rect 22922 6060 22928 6072
rect 22980 6060 22986 6112
rect 23382 6100 23388 6112
rect 23343 6072 23388 6100
rect 23382 6060 23388 6072
rect 23440 6060 23446 6112
rect 27985 6103 28043 6109
rect 27985 6069 27997 6103
rect 28031 6100 28043 6103
rect 28166 6100 28172 6112
rect 28031 6072 28172 6100
rect 28031 6069 28043 6072
rect 27985 6063 28043 6069
rect 28166 6060 28172 6072
rect 28224 6060 28230 6112
rect 46290 6060 46296 6112
rect 46348 6100 46354 6112
rect 47765 6103 47823 6109
rect 47765 6100 47777 6103
rect 46348 6072 47777 6100
rect 46348 6060 46354 6072
rect 47765 6069 47777 6072
rect 47811 6069 47823 6103
rect 47765 6063 47823 6069
rect 1104 6010 48852 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 48852 6010
rect 1104 5936 48852 5958
rect 6886 5868 26924 5896
rect 2314 5760 2320 5772
rect 2227 5732 2320 5760
rect 1762 5692 1768 5704
rect 1723 5664 1768 5692
rect 1762 5652 1768 5664
rect 1820 5652 1826 5704
rect 2240 5701 2268 5732
rect 2314 5720 2320 5732
rect 2372 5760 2378 5772
rect 6886 5760 6914 5868
rect 22002 5828 22008 5840
rect 21963 5800 22008 5828
rect 22002 5788 22008 5800
rect 22060 5788 22066 5840
rect 24210 5828 24216 5840
rect 22848 5800 24216 5828
rect 2372 5732 6914 5760
rect 2372 5720 2378 5732
rect 21634 5720 21640 5772
rect 21692 5760 21698 5772
rect 22848 5760 22876 5800
rect 24210 5788 24216 5800
rect 24268 5788 24274 5840
rect 25774 5828 25780 5840
rect 25735 5800 25780 5828
rect 25774 5788 25780 5800
rect 25832 5788 25838 5840
rect 24026 5760 24032 5772
rect 21692 5732 22876 5760
rect 21692 5720 21698 5732
rect 2225 5695 2283 5701
rect 2225 5661 2237 5695
rect 2271 5661 2283 5695
rect 2225 5655 2283 5661
rect 2682 5652 2688 5704
rect 2740 5692 2746 5704
rect 2869 5695 2927 5701
rect 2869 5692 2881 5695
rect 2740 5664 2881 5692
rect 2740 5652 2746 5664
rect 2869 5661 2881 5664
rect 2915 5661 2927 5695
rect 2869 5655 2927 5661
rect 20625 5695 20683 5701
rect 20625 5661 20637 5695
rect 20671 5692 20683 5695
rect 21818 5692 21824 5704
rect 20671 5664 21824 5692
rect 20671 5661 20683 5664
rect 20625 5655 20683 5661
rect 21818 5652 21824 5664
rect 21876 5652 21882 5704
rect 22278 5652 22284 5704
rect 22336 5692 22342 5704
rect 22848 5701 22876 5732
rect 23124 5732 24032 5760
rect 23124 5704 23152 5732
rect 24026 5720 24032 5732
rect 24084 5720 24090 5772
rect 24394 5760 24400 5772
rect 24355 5732 24400 5760
rect 24394 5720 24400 5732
rect 24452 5720 24458 5772
rect 22695 5695 22753 5701
rect 22695 5692 22707 5695
rect 22336 5664 22707 5692
rect 22336 5652 22342 5664
rect 22695 5661 22707 5664
rect 22741 5661 22753 5695
rect 22695 5655 22753 5661
rect 22833 5695 22891 5701
rect 22833 5661 22845 5695
rect 22879 5661 22891 5695
rect 22833 5655 22891 5661
rect 22922 5652 22928 5704
rect 22980 5692 22986 5704
rect 22980 5664 23025 5692
rect 22980 5652 22986 5664
rect 23106 5652 23112 5704
rect 23164 5692 23170 5704
rect 23164 5664 23257 5692
rect 23164 5652 23170 5664
rect 23382 5652 23388 5704
rect 23440 5692 23446 5704
rect 24653 5695 24711 5701
rect 24653 5692 24665 5695
rect 23440 5664 24665 5692
rect 23440 5652 23446 5664
rect 24653 5661 24665 5664
rect 24699 5661 24711 5695
rect 26896 5692 26924 5868
rect 27798 5856 27804 5908
rect 27856 5896 27862 5908
rect 28537 5899 28595 5905
rect 28537 5896 28549 5899
rect 27856 5868 28549 5896
rect 27856 5856 27862 5868
rect 28537 5865 28549 5868
rect 28583 5865 28595 5899
rect 45462 5896 45468 5908
rect 28537 5859 28595 5865
rect 31726 5868 45468 5896
rect 27154 5760 27160 5772
rect 27115 5732 27160 5760
rect 27154 5720 27160 5732
rect 27212 5720 27218 5772
rect 31726 5692 31754 5868
rect 45462 5856 45468 5868
rect 45520 5856 45526 5908
rect 46290 5760 46296 5772
rect 46251 5732 46296 5760
rect 46290 5720 46296 5732
rect 46348 5720 46354 5772
rect 26896 5664 31754 5692
rect 24653 5655 24711 5661
rect 20892 5627 20950 5633
rect 20892 5593 20904 5627
rect 20938 5624 20950 5627
rect 22465 5627 22523 5633
rect 22465 5624 22477 5627
rect 20938 5596 22477 5624
rect 20938 5593 20950 5596
rect 20892 5587 20950 5593
rect 22465 5593 22477 5596
rect 22511 5593 22523 5627
rect 22465 5587 22523 5593
rect 24394 5584 24400 5636
rect 24452 5624 24458 5636
rect 27154 5624 27160 5636
rect 24452 5596 27160 5624
rect 24452 5584 24458 5596
rect 27154 5584 27160 5596
rect 27212 5584 27218 5636
rect 27424 5627 27482 5633
rect 27424 5593 27436 5627
rect 27470 5624 27482 5627
rect 27706 5624 27712 5636
rect 27470 5596 27712 5624
rect 27470 5593 27482 5596
rect 27424 5587 27482 5593
rect 27706 5584 27712 5596
rect 27764 5584 27770 5636
rect 46477 5627 46535 5633
rect 46477 5593 46489 5627
rect 46523 5624 46535 5627
rect 46934 5624 46940 5636
rect 46523 5596 46940 5624
rect 46523 5593 46535 5596
rect 46477 5587 46535 5593
rect 46934 5584 46940 5596
rect 46992 5584 46998 5636
rect 48130 5624 48136 5636
rect 48091 5596 48136 5624
rect 48130 5584 48136 5596
rect 48188 5584 48194 5636
rect 1946 5516 1952 5568
rect 2004 5556 2010 5568
rect 2317 5559 2375 5565
rect 2317 5556 2329 5559
rect 2004 5528 2329 5556
rect 2004 5516 2010 5528
rect 2317 5525 2329 5528
rect 2363 5525 2375 5559
rect 2958 5556 2964 5568
rect 2919 5528 2964 5556
rect 2317 5519 2375 5525
rect 2958 5516 2964 5528
rect 3016 5516 3022 5568
rect 1104 5466 48852 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 48852 5466
rect 1104 5392 48852 5414
rect 3418 5312 3424 5364
rect 3476 5352 3482 5364
rect 18138 5352 18144 5364
rect 3476 5324 18144 5352
rect 3476 5312 3482 5324
rect 18138 5312 18144 5324
rect 18196 5312 18202 5364
rect 22462 5312 22468 5364
rect 22520 5352 22526 5364
rect 23201 5355 23259 5361
rect 23201 5352 23213 5355
rect 22520 5324 23213 5352
rect 22520 5312 22526 5324
rect 23201 5321 23213 5324
rect 23247 5321 23259 5355
rect 23201 5315 23259 5321
rect 23842 5312 23848 5364
rect 23900 5352 23906 5364
rect 24029 5355 24087 5361
rect 24029 5352 24041 5355
rect 23900 5324 24041 5352
rect 23900 5312 23906 5324
rect 24029 5321 24041 5324
rect 24075 5321 24087 5355
rect 27706 5352 27712 5364
rect 27667 5324 27712 5352
rect 24029 5315 24087 5321
rect 27706 5312 27712 5324
rect 27764 5312 27770 5364
rect 39298 5312 39304 5364
rect 39356 5352 39362 5364
rect 46658 5352 46664 5364
rect 39356 5324 46664 5352
rect 39356 5312 39362 5324
rect 46658 5312 46664 5324
rect 46716 5312 46722 5364
rect 46934 5352 46940 5364
rect 46895 5324 46940 5352
rect 46934 5312 46940 5324
rect 46992 5312 46998 5364
rect 1946 5284 1952 5296
rect 1907 5256 1952 5284
rect 1946 5244 1952 5256
rect 2004 5244 2010 5296
rect 14734 5244 14740 5296
rect 14792 5284 14798 5296
rect 19242 5284 19248 5296
rect 14792 5256 19248 5284
rect 14792 5244 14798 5256
rect 19242 5244 19248 5256
rect 19300 5244 19306 5296
rect 20625 5287 20683 5293
rect 20625 5253 20637 5287
rect 20671 5284 20683 5287
rect 22066 5287 22124 5293
rect 22066 5284 22078 5287
rect 20671 5256 22078 5284
rect 20671 5253 20683 5256
rect 20625 5247 20683 5253
rect 22066 5253 22078 5256
rect 22112 5253 22124 5287
rect 22066 5247 22124 5253
rect 23661 5287 23719 5293
rect 23661 5253 23673 5287
rect 23707 5284 23719 5287
rect 24118 5284 24124 5296
rect 23707 5256 24124 5284
rect 23707 5253 23719 5256
rect 23661 5247 23719 5253
rect 24118 5244 24124 5256
rect 24176 5244 24182 5296
rect 24210 5244 24216 5296
rect 24268 5284 24274 5296
rect 28994 5284 29000 5296
rect 24268 5256 29000 5284
rect 24268 5244 24274 5256
rect 1578 5176 1584 5228
rect 1636 5216 1642 5228
rect 1765 5219 1823 5225
rect 1765 5216 1777 5219
rect 1636 5188 1777 5216
rect 1636 5176 1642 5188
rect 1765 5185 1777 5188
rect 1811 5185 1823 5219
rect 1765 5179 1823 5185
rect 19334 5176 19340 5228
rect 19392 5216 19398 5228
rect 20855 5219 20913 5225
rect 20855 5216 20867 5219
rect 19392 5188 20867 5216
rect 19392 5176 19398 5188
rect 20855 5185 20867 5188
rect 20901 5185 20913 5219
rect 20855 5179 20913 5185
rect 20993 5219 21051 5225
rect 20993 5185 21005 5219
rect 21039 5185 21051 5219
rect 20993 5179 21051 5185
rect 2774 5148 2780 5160
rect 2735 5120 2780 5148
rect 2774 5108 2780 5120
rect 2832 5108 2838 5160
rect 21008 5080 21036 5179
rect 21082 5176 21088 5228
rect 21140 5222 21164 5228
rect 21152 5188 21164 5222
rect 21140 5182 21164 5188
rect 21269 5219 21327 5225
rect 21269 5185 21281 5219
rect 21315 5185 21327 5219
rect 21818 5216 21824 5228
rect 21779 5188 21824 5216
rect 21140 5176 21146 5182
rect 21269 5179 21327 5185
rect 21284 5148 21312 5179
rect 21818 5176 21824 5188
rect 21876 5176 21882 5228
rect 23106 5216 23112 5228
rect 21928 5188 23112 5216
rect 21928 5148 21956 5188
rect 23106 5176 23112 5188
rect 23164 5176 23170 5228
rect 23845 5219 23903 5225
rect 23845 5185 23857 5219
rect 23891 5216 23903 5219
rect 25774 5216 25780 5228
rect 23891 5188 25780 5216
rect 23891 5185 23903 5188
rect 23845 5179 23903 5185
rect 25774 5176 25780 5188
rect 25832 5176 25838 5228
rect 28092 5225 28120 5256
rect 28994 5244 29000 5256
rect 29052 5244 29058 5296
rect 27985 5219 28043 5225
rect 27985 5185 27997 5219
rect 28031 5185 28043 5219
rect 27985 5179 28043 5185
rect 28077 5219 28135 5225
rect 28077 5185 28089 5219
rect 28123 5185 28135 5219
rect 28077 5179 28135 5185
rect 21284 5120 21956 5148
rect 28000 5148 28028 5179
rect 28166 5176 28172 5228
rect 28224 5216 28230 5228
rect 28353 5219 28411 5225
rect 28224 5188 28269 5216
rect 28224 5176 28230 5188
rect 28353 5185 28365 5219
rect 28399 5216 28411 5219
rect 28718 5216 28724 5228
rect 28399 5188 28724 5216
rect 28399 5185 28411 5188
rect 28353 5179 28411 5185
rect 28718 5176 28724 5188
rect 28776 5176 28782 5228
rect 46842 5216 46848 5228
rect 46803 5188 46848 5216
rect 46842 5176 46848 5188
rect 46900 5176 46906 5228
rect 47854 5216 47860 5228
rect 47815 5188 47860 5216
rect 47854 5176 47860 5188
rect 47912 5176 47918 5228
rect 38746 5148 38752 5160
rect 28000 5120 38752 5148
rect 38746 5108 38752 5120
rect 38804 5108 38810 5160
rect 21634 5080 21640 5092
rect 21008 5052 21640 5080
rect 21634 5040 21640 5052
rect 21692 5040 21698 5092
rect 24026 5040 24032 5092
rect 24084 5080 24090 5092
rect 28718 5080 28724 5092
rect 24084 5052 28724 5080
rect 24084 5040 24090 5052
rect 28718 5040 28724 5052
rect 28776 5040 28782 5092
rect 29822 5040 29828 5092
rect 29880 5080 29886 5092
rect 48041 5083 48099 5089
rect 48041 5080 48053 5083
rect 29880 5052 48053 5080
rect 29880 5040 29886 5052
rect 48041 5049 48053 5052
rect 48087 5049 48099 5083
rect 48041 5043 48099 5049
rect 1104 4922 48852 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 48852 4922
rect 1104 4848 48852 4870
rect 17218 4700 17224 4752
rect 17276 4740 17282 4752
rect 46842 4740 46848 4752
rect 17276 4712 46848 4740
rect 17276 4700 17282 4712
rect 46842 4700 46848 4712
rect 46900 4700 46906 4752
rect 1397 4675 1455 4681
rect 1397 4641 1409 4675
rect 1443 4672 1455 4675
rect 1762 4672 1768 4684
rect 1443 4644 1768 4672
rect 1443 4641 1455 4644
rect 1397 4635 1455 4641
rect 1762 4632 1768 4644
rect 1820 4632 1826 4684
rect 2774 4672 2780 4684
rect 2735 4644 2780 4672
rect 2774 4632 2780 4644
rect 2832 4632 2838 4684
rect 30926 4672 30932 4684
rect 30887 4644 30932 4672
rect 30926 4632 30932 4644
rect 30984 4632 30990 4684
rect 6178 4564 6184 4616
rect 6236 4604 6242 4616
rect 6457 4607 6515 4613
rect 6457 4604 6469 4607
rect 6236 4576 6469 4604
rect 6236 4564 6242 4576
rect 6457 4573 6469 4576
rect 6503 4573 6515 4607
rect 6457 4567 6515 4573
rect 13170 4564 13176 4616
rect 13228 4604 13234 4616
rect 13357 4607 13415 4613
rect 13357 4604 13369 4607
rect 13228 4576 13369 4604
rect 13228 4564 13234 4576
rect 13357 4573 13369 4576
rect 13403 4573 13415 4607
rect 13357 4567 13415 4573
rect 30285 4607 30343 4613
rect 30285 4573 30297 4607
rect 30331 4573 30343 4607
rect 41966 4604 41972 4616
rect 41927 4576 41972 4604
rect 30285 4567 30343 4573
rect 1581 4539 1639 4545
rect 1581 4505 1593 4539
rect 1627 4536 1639 4539
rect 2958 4536 2964 4548
rect 1627 4508 2964 4536
rect 1627 4505 1639 4508
rect 1581 4499 1639 4505
rect 2958 4496 2964 4508
rect 3016 4496 3022 4548
rect 30300 4468 30328 4567
rect 41966 4564 41972 4576
rect 42024 4564 42030 4616
rect 45833 4607 45891 4613
rect 45833 4573 45845 4607
rect 45879 4604 45891 4607
rect 46293 4607 46351 4613
rect 46293 4604 46305 4607
rect 45879 4576 46305 4604
rect 45879 4573 45891 4576
rect 45833 4567 45891 4573
rect 46293 4573 46305 4576
rect 46339 4573 46351 4607
rect 46293 4567 46351 4573
rect 30469 4539 30527 4545
rect 30469 4505 30481 4539
rect 30515 4536 30527 4539
rect 30650 4536 30656 4548
rect 30515 4508 30656 4536
rect 30515 4505 30527 4508
rect 30469 4499 30527 4505
rect 30650 4496 30656 4508
rect 30708 4496 30714 4548
rect 46477 4539 46535 4545
rect 46477 4505 46489 4539
rect 46523 4536 46535 4539
rect 46934 4536 46940 4548
rect 46523 4508 46940 4536
rect 46523 4505 46535 4508
rect 46477 4499 46535 4505
rect 46934 4496 46940 4508
rect 46992 4496 46998 4548
rect 48133 4539 48191 4545
rect 48133 4505 48145 4539
rect 48179 4536 48191 4539
rect 48314 4536 48320 4548
rect 48179 4508 48320 4536
rect 48179 4505 48191 4508
rect 48133 4499 48191 4505
rect 48314 4496 48320 4508
rect 48372 4496 48378 4548
rect 30374 4468 30380 4480
rect 30300 4440 30380 4468
rect 30374 4428 30380 4440
rect 30432 4428 30438 4480
rect 1104 4378 48852 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 48852 4378
rect 1104 4304 48852 4326
rect 29472 4236 30788 4264
rect 22005 4199 22063 4205
rect 22005 4196 22017 4199
rect 6932 4168 7144 4196
rect 1578 4128 1584 4140
rect 1539 4100 1584 4128
rect 1578 4088 1584 4100
rect 1636 4088 1642 4140
rect 2225 4131 2283 4137
rect 2225 4097 2237 4131
rect 2271 4097 2283 4131
rect 3050 4128 3056 4140
rect 3011 4100 3056 4128
rect 2225 4091 2283 4097
rect 2240 3992 2268 4091
rect 3050 4088 3056 4100
rect 3108 4088 3114 4140
rect 6365 4131 6423 4137
rect 6365 4097 6377 4131
rect 6411 4128 6423 4131
rect 6932 4128 6960 4168
rect 6411 4100 6960 4128
rect 7009 4131 7067 4137
rect 6411 4097 6423 4100
rect 6365 4091 6423 4097
rect 7009 4097 7021 4131
rect 7055 4097 7067 4131
rect 7116 4128 7144 4168
rect 21836 4168 22017 4196
rect 12250 4128 12256 4140
rect 7116 4100 12256 4128
rect 7009 4091 7067 4097
rect 7024 4060 7052 4091
rect 12250 4088 12256 4100
rect 12308 4088 12314 4140
rect 13170 4128 13176 4140
rect 13131 4100 13176 4128
rect 13170 4088 13176 4100
rect 13228 4088 13234 4140
rect 16758 4088 16764 4140
rect 16816 4128 16822 4140
rect 20901 4131 20959 4137
rect 20901 4128 20913 4131
rect 16816 4100 20913 4128
rect 16816 4088 16822 4100
rect 20901 4097 20913 4100
rect 20947 4097 20959 4131
rect 20901 4091 20959 4097
rect 20993 4131 21051 4137
rect 20993 4097 21005 4131
rect 21039 4128 21051 4131
rect 21836 4128 21864 4168
rect 22005 4165 22017 4168
rect 22051 4165 22063 4199
rect 22005 4159 22063 4165
rect 21039 4100 21864 4128
rect 21039 4097 21051 4100
rect 20993 4091 21051 4097
rect 26234 4088 26240 4140
rect 26292 4128 26298 4140
rect 26602 4128 26608 4140
rect 26292 4100 26608 4128
rect 26292 4088 26298 4100
rect 26602 4088 26608 4100
rect 26660 4088 26666 4140
rect 7024 4032 13032 4060
rect 11606 3992 11612 4004
rect 2240 3964 11612 3992
rect 11606 3952 11612 3964
rect 11664 3952 11670 4004
rect 11974 3952 11980 4004
rect 12032 3992 12038 4004
rect 12713 3995 12771 4001
rect 12713 3992 12725 3995
rect 12032 3964 12725 3992
rect 12032 3952 12038 3964
rect 12713 3961 12725 3964
rect 12759 3961 12771 3995
rect 13004 3992 13032 4032
rect 13078 4020 13084 4072
rect 13136 4060 13142 4072
rect 13357 4063 13415 4069
rect 13357 4060 13369 4063
rect 13136 4032 13369 4060
rect 13136 4020 13142 4032
rect 13357 4029 13369 4032
rect 13403 4029 13415 4063
rect 13357 4023 13415 4029
rect 13538 4020 13544 4072
rect 13596 4060 13602 4072
rect 13633 4063 13691 4069
rect 13633 4060 13645 4063
rect 13596 4032 13645 4060
rect 13596 4020 13602 4032
rect 13633 4029 13645 4032
rect 13679 4029 13691 4063
rect 13633 4023 13691 4029
rect 16206 4020 16212 4072
rect 16264 4060 16270 4072
rect 20806 4060 20812 4072
rect 16264 4032 20812 4060
rect 16264 4020 16270 4032
rect 20806 4020 20812 4032
rect 20864 4020 20870 4072
rect 21174 4020 21180 4072
rect 21232 4060 21238 4072
rect 21821 4063 21879 4069
rect 21821 4060 21833 4063
rect 21232 4032 21833 4060
rect 21232 4020 21238 4032
rect 21821 4029 21833 4032
rect 21867 4029 21879 4063
rect 22281 4063 22339 4069
rect 22281 4060 22293 4063
rect 21821 4023 21879 4029
rect 21928 4032 22293 4060
rect 15286 3992 15292 4004
rect 13004 3964 15292 3992
rect 12713 3955 12771 3961
rect 15286 3952 15292 3964
rect 15344 3952 15350 4004
rect 20346 3952 20352 4004
rect 20404 3992 20410 4004
rect 20404 3964 20576 3992
rect 20404 3952 20410 3964
rect 1673 3927 1731 3933
rect 1673 3893 1685 3927
rect 1719 3924 1731 3927
rect 1946 3924 1952 3936
rect 1719 3896 1952 3924
rect 1719 3893 1731 3896
rect 1673 3887 1731 3893
rect 1946 3884 1952 3896
rect 2004 3884 2010 3936
rect 2314 3924 2320 3936
rect 2275 3896 2320 3924
rect 2314 3884 2320 3896
rect 2372 3884 2378 3936
rect 3142 3924 3148 3936
rect 3103 3896 3148 3924
rect 3142 3884 3148 3896
rect 3200 3884 3206 3936
rect 3878 3924 3884 3936
rect 3839 3896 3884 3924
rect 3878 3884 3884 3896
rect 3936 3884 3942 3936
rect 6457 3927 6515 3933
rect 6457 3893 6469 3927
rect 6503 3924 6515 3927
rect 6546 3924 6552 3936
rect 6503 3896 6552 3924
rect 6503 3893 6515 3896
rect 6457 3887 6515 3893
rect 6546 3884 6552 3896
rect 6604 3884 6610 3936
rect 7098 3924 7104 3936
rect 7059 3896 7104 3924
rect 7098 3884 7104 3896
rect 7156 3884 7162 3936
rect 11698 3884 11704 3936
rect 11756 3924 11762 3936
rect 12069 3927 12127 3933
rect 12069 3924 12081 3927
rect 11756 3896 12081 3924
rect 11756 3884 11762 3896
rect 12069 3893 12081 3896
rect 12115 3893 12127 3927
rect 12069 3887 12127 3893
rect 12618 3884 12624 3936
rect 12676 3924 12682 3936
rect 17126 3924 17132 3936
rect 12676 3896 17132 3924
rect 12676 3884 12682 3896
rect 17126 3884 17132 3896
rect 17184 3924 17190 3936
rect 17402 3924 17408 3936
rect 17184 3896 17408 3924
rect 17184 3884 17190 3896
rect 17402 3884 17408 3896
rect 17460 3884 17466 3936
rect 20162 3884 20168 3936
rect 20220 3924 20226 3936
rect 20441 3927 20499 3933
rect 20441 3924 20453 3927
rect 20220 3896 20453 3924
rect 20220 3884 20226 3896
rect 20441 3893 20453 3896
rect 20487 3893 20499 3927
rect 20548 3924 20576 3964
rect 21266 3952 21272 4004
rect 21324 3992 21330 4004
rect 21928 3992 21956 4032
rect 22281 4029 22293 4032
rect 22327 4029 22339 4063
rect 22281 4023 22339 4029
rect 22370 4020 22376 4072
rect 22428 4060 22434 4072
rect 29472 4060 29500 4236
rect 30484 4168 30696 4196
rect 29546 4088 29552 4140
rect 29604 4128 29610 4140
rect 29641 4131 29699 4137
rect 29641 4128 29653 4131
rect 29604 4100 29653 4128
rect 29604 4088 29610 4100
rect 29641 4097 29653 4100
rect 29687 4097 29699 4131
rect 29641 4091 29699 4097
rect 29730 4088 29736 4140
rect 29788 4128 29794 4140
rect 30484 4128 30512 4168
rect 29788 4100 30512 4128
rect 30561 4131 30619 4137
rect 29788 4088 29794 4100
rect 30561 4097 30573 4131
rect 30607 4097 30619 4131
rect 30561 4091 30619 4097
rect 30576 4060 30604 4091
rect 22428 4032 29500 4060
rect 29564 4032 30604 4060
rect 22428 4020 22434 4032
rect 21324 3964 21956 3992
rect 21324 3952 21330 3964
rect 22002 3952 22008 4004
rect 22060 3992 22066 4004
rect 29564 3992 29592 4032
rect 22060 3964 29592 3992
rect 30668 3992 30696 4168
rect 30760 4128 30788 4236
rect 46750 4156 46756 4208
rect 46808 4196 46814 4208
rect 47949 4199 48007 4205
rect 47949 4196 47961 4199
rect 46808 4168 47961 4196
rect 46808 4156 46814 4168
rect 47949 4165 47961 4168
rect 47995 4165 48007 4199
rect 47949 4159 48007 4165
rect 36357 4131 36415 4137
rect 36357 4128 36369 4131
rect 30760 4100 36369 4128
rect 36357 4097 36369 4100
rect 36403 4097 36415 4131
rect 36357 4091 36415 4097
rect 36446 4088 36452 4140
rect 36504 4128 36510 4140
rect 38013 4131 38071 4137
rect 38013 4128 38025 4131
rect 36504 4100 38025 4128
rect 36504 4088 36510 4100
rect 38013 4097 38025 4100
rect 38059 4097 38071 4131
rect 39482 4128 39488 4140
rect 39443 4100 39488 4128
rect 38013 4091 38071 4097
rect 39482 4088 39488 4100
rect 39540 4088 39546 4140
rect 42426 4128 42432 4140
rect 42387 4100 42432 4128
rect 42426 4088 42432 4100
rect 42484 4088 42490 4140
rect 44177 4131 44235 4137
rect 44177 4097 44189 4131
rect 44223 4128 44235 4131
rect 45554 4128 45560 4140
rect 44223 4100 45560 4128
rect 44223 4097 44235 4100
rect 44177 4091 44235 4097
rect 45554 4088 45560 4100
rect 45612 4088 45618 4140
rect 45830 4128 45836 4140
rect 45791 4100 45836 4128
rect 45830 4088 45836 4100
rect 45888 4088 45894 4140
rect 46842 4128 46848 4140
rect 46803 4100 46848 4128
rect 46842 4088 46848 4100
rect 46900 4088 46906 4140
rect 46934 4088 46940 4140
rect 46992 4128 46998 4140
rect 46992 4100 47037 4128
rect 46992 4088 46998 4100
rect 42444 4060 42472 4088
rect 42444 4032 44772 4060
rect 40770 3992 40776 4004
rect 30668 3964 40776 3992
rect 22060 3952 22066 3964
rect 40770 3952 40776 3964
rect 40828 3952 40834 4004
rect 43717 3995 43775 4001
rect 43717 3961 43729 3995
rect 43763 3992 43775 3995
rect 44634 3992 44640 4004
rect 43763 3964 44640 3992
rect 43763 3961 43775 3964
rect 43717 3955 43775 3961
rect 44634 3952 44640 3964
rect 44692 3952 44698 4004
rect 29546 3924 29552 3936
rect 20548 3896 29552 3924
rect 20441 3887 20499 3893
rect 29546 3884 29552 3896
rect 29604 3884 29610 3936
rect 29733 3927 29791 3933
rect 29733 3893 29745 3927
rect 29779 3924 29791 3927
rect 30558 3924 30564 3936
rect 29779 3896 30564 3924
rect 29779 3893 29791 3896
rect 29733 3887 29791 3893
rect 30558 3884 30564 3896
rect 30616 3884 30622 3936
rect 30650 3884 30656 3936
rect 30708 3924 30714 3936
rect 31386 3924 31392 3936
rect 30708 3896 30753 3924
rect 31347 3896 31392 3924
rect 30708 3884 30714 3896
rect 31386 3884 31392 3896
rect 31444 3884 31450 3936
rect 32766 3884 32772 3936
rect 32824 3924 32830 3936
rect 32953 3927 33011 3933
rect 32953 3924 32965 3927
rect 32824 3896 32965 3924
rect 32824 3884 32830 3896
rect 32953 3893 32965 3896
rect 32999 3893 33011 3927
rect 32953 3887 33011 3893
rect 36170 3884 36176 3936
rect 36228 3924 36234 3936
rect 36449 3927 36507 3933
rect 36449 3924 36461 3927
rect 36228 3896 36461 3924
rect 36228 3884 36234 3896
rect 36449 3893 36461 3896
rect 36495 3893 36507 3927
rect 36449 3887 36507 3893
rect 37918 3884 37924 3936
rect 37976 3924 37982 3936
rect 38105 3927 38163 3933
rect 38105 3924 38117 3927
rect 37976 3896 38117 3924
rect 37976 3884 37982 3896
rect 38105 3893 38117 3896
rect 38151 3893 38163 3927
rect 38105 3887 38163 3893
rect 39577 3927 39635 3933
rect 39577 3893 39589 3927
rect 39623 3924 39635 3927
rect 40218 3924 40224 3936
rect 39623 3896 40224 3924
rect 39623 3893 39635 3896
rect 39577 3887 39635 3893
rect 40218 3884 40224 3896
rect 40276 3884 40282 3936
rect 41414 3884 41420 3936
rect 41472 3924 41478 3936
rect 41693 3927 41751 3933
rect 41693 3924 41705 3927
rect 41472 3896 41705 3924
rect 41472 3884 41478 3896
rect 41693 3893 41705 3896
rect 41739 3893 41751 3927
rect 41693 3887 41751 3893
rect 42521 3927 42579 3933
rect 42521 3893 42533 3927
rect 42567 3924 42579 3927
rect 42610 3924 42616 3936
rect 42567 3896 42616 3924
rect 42567 3893 42579 3896
rect 42521 3887 42579 3893
rect 42610 3884 42616 3896
rect 42668 3884 42674 3936
rect 43990 3884 43996 3936
rect 44048 3924 44054 3936
rect 44269 3927 44327 3933
rect 44269 3924 44281 3927
rect 44048 3896 44281 3924
rect 44048 3884 44054 3896
rect 44269 3893 44281 3896
rect 44315 3893 44327 3927
rect 44744 3924 44772 4032
rect 44818 4020 44824 4072
rect 44876 4060 44882 4072
rect 48133 4063 48191 4069
rect 48133 4060 48145 4063
rect 44876 4032 48145 4060
rect 44876 4020 44882 4032
rect 48133 4029 48145 4032
rect 48179 4029 48191 4063
rect 48133 4023 48191 4029
rect 46290 3992 46296 4004
rect 45112 3964 46296 3992
rect 45112 3924 45140 3964
rect 46290 3952 46296 3964
rect 46348 3952 46354 4004
rect 45370 3924 45376 3936
rect 44744 3896 45140 3924
rect 45331 3896 45376 3924
rect 44269 3887 44327 3893
rect 45370 3884 45376 3896
rect 45428 3884 45434 3936
rect 45925 3927 45983 3933
rect 45925 3893 45937 3927
rect 45971 3924 45983 3927
rect 46198 3924 46204 3936
rect 45971 3896 46204 3924
rect 45971 3893 45983 3896
rect 45925 3887 45983 3893
rect 46198 3884 46204 3896
rect 46256 3884 46262 3936
rect 1104 3834 48852 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 48852 3834
rect 1104 3760 48852 3782
rect 3878 3720 3884 3732
rect 1412 3692 3884 3720
rect 1412 3593 1440 3692
rect 3878 3680 3884 3692
rect 3936 3680 3942 3732
rect 9030 3680 9036 3732
rect 9088 3720 9094 3732
rect 9088 3692 32168 3720
rect 9088 3680 9094 3692
rect 2314 3652 2320 3664
rect 1596 3624 2320 3652
rect 1596 3593 1624 3624
rect 2314 3612 2320 3624
rect 2372 3612 2378 3664
rect 3234 3612 3240 3664
rect 3292 3652 3298 3664
rect 3292 3624 4292 3652
rect 3292 3612 3298 3624
rect 1397 3587 1455 3593
rect 1397 3553 1409 3587
rect 1443 3553 1455 3587
rect 1397 3547 1455 3553
rect 1581 3587 1639 3593
rect 1581 3553 1593 3587
rect 1627 3553 1639 3587
rect 1854 3584 1860 3596
rect 1815 3556 1860 3584
rect 1581 3547 1639 3553
rect 1854 3544 1860 3556
rect 1912 3544 1918 3596
rect 3142 3544 3148 3596
rect 3200 3584 3206 3596
rect 4264 3593 4292 3624
rect 5810 3612 5816 3664
rect 5868 3652 5874 3664
rect 5868 3624 7236 3652
rect 5868 3612 5874 3624
rect 3973 3587 4031 3593
rect 3973 3584 3985 3587
rect 3200 3556 3985 3584
rect 3200 3544 3206 3556
rect 3973 3553 3985 3556
rect 4019 3553 4031 3587
rect 3973 3547 4031 3553
rect 4249 3587 4307 3593
rect 4249 3553 4261 3587
rect 4295 3553 4307 3587
rect 6178 3584 6184 3596
rect 6139 3556 6184 3584
rect 4249 3547 4307 3553
rect 6178 3544 6184 3556
rect 6236 3544 6242 3596
rect 6365 3587 6423 3593
rect 6365 3553 6377 3587
rect 6411 3584 6423 3587
rect 7098 3584 7104 3596
rect 6411 3556 7104 3584
rect 6411 3553 6423 3556
rect 6365 3547 6423 3553
rect 7098 3544 7104 3556
rect 7156 3544 7162 3596
rect 7208 3593 7236 3624
rect 10318 3612 10324 3664
rect 10376 3652 10382 3664
rect 12894 3652 12900 3664
rect 10376 3624 12900 3652
rect 10376 3612 10382 3624
rect 12894 3612 12900 3624
rect 12952 3612 12958 3664
rect 13078 3652 13084 3664
rect 13039 3624 13084 3652
rect 13078 3612 13084 3624
rect 13136 3612 13142 3664
rect 13170 3612 13176 3664
rect 13228 3652 13234 3664
rect 13228 3624 16252 3652
rect 13228 3612 13234 3624
rect 7193 3587 7251 3593
rect 7193 3553 7205 3587
rect 7239 3553 7251 3587
rect 12618 3584 12624 3596
rect 7193 3547 7251 3553
rect 11716 3556 12624 3584
rect 3786 3516 3792 3528
rect 3747 3488 3792 3516
rect 3786 3476 3792 3488
rect 3844 3476 3850 3528
rect 11606 3516 11612 3528
rect 11519 3488 11612 3516
rect 11606 3476 11612 3488
rect 11664 3516 11670 3528
rect 11716 3516 11744 3556
rect 12618 3544 12624 3556
rect 12676 3544 12682 3596
rect 16114 3584 16120 3596
rect 12912 3556 16120 3584
rect 12250 3516 12256 3528
rect 11664 3488 11744 3516
rect 12163 3488 12256 3516
rect 11664 3476 11670 3488
rect 12250 3476 12256 3488
rect 12308 3516 12314 3528
rect 12912 3516 12940 3556
rect 16114 3544 16120 3556
rect 16172 3544 16178 3596
rect 16224 3584 16252 3624
rect 18506 3612 18512 3664
rect 18564 3652 18570 3664
rect 30282 3652 30288 3664
rect 18564 3624 30288 3652
rect 18564 3612 18570 3624
rect 30282 3612 30288 3624
rect 30340 3612 30346 3664
rect 31386 3652 31392 3664
rect 30392 3624 31392 3652
rect 20162 3584 20168 3596
rect 16224 3556 20024 3584
rect 20123 3556 20168 3584
rect 12308 3488 12940 3516
rect 12308 3476 12314 3488
rect 12986 3476 12992 3528
rect 13044 3516 13050 3528
rect 13044 3488 13089 3516
rect 13044 3476 13050 3488
rect 14274 3476 14280 3528
rect 14332 3516 14338 3528
rect 14645 3519 14703 3525
rect 14645 3516 14657 3519
rect 14332 3488 14657 3516
rect 14332 3476 14338 3488
rect 14645 3485 14657 3488
rect 14691 3485 14703 3519
rect 14645 3479 14703 3485
rect 15105 3519 15163 3525
rect 15105 3485 15117 3519
rect 15151 3516 15163 3519
rect 15194 3516 15200 3528
rect 15151 3488 15200 3516
rect 15151 3485 15163 3488
rect 15105 3479 15163 3485
rect 15194 3476 15200 3488
rect 15252 3516 15258 3528
rect 15654 3516 15660 3528
rect 15252 3488 15660 3516
rect 15252 3476 15258 3488
rect 15654 3476 15660 3488
rect 15712 3516 15718 3528
rect 17589 3519 17647 3525
rect 17589 3516 17601 3519
rect 15712 3488 17601 3516
rect 15712 3476 15718 3488
rect 17589 3485 17601 3488
rect 17635 3485 17647 3519
rect 17589 3479 17647 3485
rect 17678 3476 17684 3528
rect 17736 3476 17742 3528
rect 17770 3476 17776 3528
rect 17828 3516 17834 3528
rect 18417 3519 18475 3525
rect 18417 3516 18429 3519
rect 17828 3488 18429 3516
rect 17828 3476 17834 3488
rect 18417 3485 18429 3488
rect 18463 3485 18475 3519
rect 18417 3479 18475 3485
rect 2590 3408 2596 3460
rect 2648 3448 2654 3460
rect 17696 3448 17724 3476
rect 2648 3420 17724 3448
rect 19996 3448 20024 3556
rect 20162 3544 20168 3556
rect 20220 3544 20226 3596
rect 20346 3584 20352 3596
rect 20307 3556 20352 3584
rect 20346 3544 20352 3556
rect 20404 3544 20410 3596
rect 20622 3584 20628 3596
rect 20583 3556 20628 3584
rect 20622 3544 20628 3556
rect 20680 3544 20686 3596
rect 20806 3544 20812 3596
rect 20864 3584 20870 3596
rect 21910 3584 21916 3596
rect 20864 3556 21916 3584
rect 20864 3544 20870 3556
rect 21910 3544 21916 3556
rect 21968 3544 21974 3596
rect 26053 3587 26111 3593
rect 22066 3556 23336 3584
rect 22066 3448 22094 3556
rect 22738 3516 22744 3528
rect 22699 3488 22744 3516
rect 22738 3476 22744 3488
rect 22796 3476 22802 3528
rect 23201 3519 23259 3525
rect 23201 3516 23213 3519
rect 22848 3488 23213 3516
rect 19996 3420 22094 3448
rect 2648 3408 2654 3420
rect 1578 3340 1584 3392
rect 1636 3380 1642 3392
rect 11606 3380 11612 3392
rect 1636 3352 11612 3380
rect 1636 3340 1642 3352
rect 11606 3340 11612 3352
rect 11664 3340 11670 3392
rect 11701 3383 11759 3389
rect 11701 3349 11713 3383
rect 11747 3380 11759 3383
rect 11882 3380 11888 3392
rect 11747 3352 11888 3380
rect 11747 3349 11759 3352
rect 11701 3343 11759 3349
rect 11882 3340 11888 3352
rect 11940 3340 11946 3392
rect 12158 3340 12164 3392
rect 12216 3380 12222 3392
rect 12345 3383 12403 3389
rect 12345 3380 12357 3383
rect 12216 3352 12357 3380
rect 12216 3340 12222 3352
rect 12345 3349 12357 3352
rect 12391 3349 12403 3383
rect 12345 3343 12403 3349
rect 14458 3340 14464 3392
rect 14516 3380 14522 3392
rect 15197 3383 15255 3389
rect 15197 3380 15209 3383
rect 14516 3352 15209 3380
rect 14516 3340 14522 3352
rect 15197 3349 15209 3352
rect 15243 3349 15255 3383
rect 15197 3343 15255 3349
rect 17681 3383 17739 3389
rect 17681 3349 17693 3383
rect 17727 3380 17739 3383
rect 17954 3380 17960 3392
rect 17727 3352 17960 3380
rect 17727 3349 17739 3352
rect 17681 3343 17739 3349
rect 17954 3340 17960 3352
rect 18012 3340 18018 3392
rect 18230 3340 18236 3392
rect 18288 3380 18294 3392
rect 22848 3380 22876 3488
rect 23201 3485 23213 3488
rect 23247 3485 23259 3519
rect 23201 3479 23259 3485
rect 23308 3448 23336 3556
rect 26053 3553 26065 3587
rect 26099 3584 26111 3587
rect 26234 3584 26240 3596
rect 26099 3556 26240 3584
rect 26099 3553 26111 3556
rect 26053 3547 26111 3553
rect 26234 3544 26240 3556
rect 26292 3544 26298 3596
rect 26418 3584 26424 3596
rect 26379 3556 26424 3584
rect 26418 3544 26424 3556
rect 26476 3544 26482 3596
rect 25866 3516 25872 3528
rect 25827 3488 25872 3516
rect 25866 3476 25872 3488
rect 25924 3476 25930 3528
rect 28994 3516 29000 3528
rect 28955 3488 29000 3516
rect 28994 3476 29000 3488
rect 29052 3476 29058 3528
rect 29549 3519 29607 3525
rect 29549 3485 29561 3519
rect 29595 3516 29607 3519
rect 29730 3516 29736 3528
rect 29595 3488 29736 3516
rect 29595 3485 29607 3488
rect 29549 3479 29607 3485
rect 29454 3448 29460 3460
rect 23308 3420 29460 3448
rect 29454 3408 29460 3420
rect 29512 3408 29518 3460
rect 18288 3352 22876 3380
rect 23293 3383 23351 3389
rect 18288 3340 18294 3352
rect 23293 3349 23305 3383
rect 23339 3380 23351 3383
rect 23658 3380 23664 3392
rect 23339 3352 23664 3380
rect 23339 3349 23351 3352
rect 23293 3343 23351 3349
rect 23658 3340 23664 3352
rect 23716 3340 23722 3392
rect 23750 3340 23756 3392
rect 23808 3380 23814 3392
rect 29564 3380 29592 3479
rect 29730 3476 29736 3488
rect 29788 3476 29794 3528
rect 30392 3525 30420 3624
rect 31386 3612 31392 3624
rect 31444 3612 31450 3664
rect 31570 3584 31576 3596
rect 31531 3556 31576 3584
rect 31570 3544 31576 3556
rect 31628 3544 31634 3596
rect 30377 3519 30435 3525
rect 30377 3485 30389 3519
rect 30423 3485 30435 3519
rect 32140 3516 32168 3692
rect 32214 3680 32220 3732
rect 32272 3720 32278 3732
rect 33962 3720 33968 3732
rect 32272 3692 33968 3720
rect 32272 3680 32278 3692
rect 33962 3680 33968 3692
rect 34020 3680 34026 3732
rect 37366 3680 37372 3732
rect 37424 3720 37430 3732
rect 39574 3720 39580 3732
rect 37424 3692 39580 3720
rect 37424 3680 37430 3692
rect 39574 3680 39580 3692
rect 39632 3680 39638 3732
rect 32306 3612 32312 3664
rect 32364 3652 32370 3664
rect 42426 3652 42432 3664
rect 32364 3624 42432 3652
rect 32364 3612 32370 3624
rect 42426 3612 42432 3624
rect 42484 3612 42490 3664
rect 47486 3652 47492 3664
rect 45020 3624 47492 3652
rect 36170 3584 36176 3596
rect 32324 3556 33824 3584
rect 36131 3556 36176 3584
rect 32324 3516 32352 3556
rect 32140 3488 32352 3516
rect 33137 3519 33195 3525
rect 30377 3479 30435 3485
rect 33137 3485 33149 3519
rect 33183 3485 33195 3519
rect 33137 3479 33195 3485
rect 30558 3448 30564 3460
rect 30519 3420 30564 3448
rect 30558 3408 30564 3420
rect 30616 3408 30622 3460
rect 33152 3448 33180 3479
rect 32416 3420 33180 3448
rect 33796 3448 33824 3556
rect 36170 3544 36176 3556
rect 36228 3544 36234 3596
rect 36722 3584 36728 3596
rect 36683 3556 36728 3584
rect 36722 3544 36728 3556
rect 36780 3544 36786 3596
rect 41414 3584 41420 3596
rect 41375 3556 41420 3584
rect 41414 3544 41420 3556
rect 41472 3544 41478 3596
rect 41874 3584 41880 3596
rect 41835 3556 41880 3584
rect 41874 3544 41880 3556
rect 41932 3544 41938 3596
rect 35986 3516 35992 3528
rect 35947 3488 35992 3516
rect 35986 3476 35992 3488
rect 36044 3476 36050 3528
rect 37734 3476 37740 3528
rect 37792 3516 37798 3528
rect 38933 3519 38991 3525
rect 38933 3516 38945 3519
rect 37792 3488 38945 3516
rect 37792 3476 37798 3488
rect 38933 3485 38945 3488
rect 38979 3485 38991 3519
rect 40770 3516 40776 3528
rect 40731 3488 40776 3516
rect 38933 3479 38991 3485
rect 40770 3476 40776 3488
rect 40828 3476 40834 3528
rect 43806 3476 43812 3528
rect 43864 3516 43870 3528
rect 45020 3525 45048 3624
rect 47486 3612 47492 3624
rect 47544 3612 47550 3664
rect 45370 3544 45376 3596
rect 45428 3584 45434 3596
rect 46017 3587 46075 3593
rect 46017 3584 46029 3587
rect 45428 3556 46029 3584
rect 45428 3544 45434 3556
rect 46017 3553 46029 3556
rect 46063 3553 46075 3587
rect 46198 3584 46204 3596
rect 46159 3556 46204 3584
rect 46017 3547 46075 3553
rect 46198 3544 46204 3556
rect 46256 3544 46262 3596
rect 46474 3584 46480 3596
rect 46435 3556 46480 3584
rect 46474 3544 46480 3556
rect 46532 3544 46538 3596
rect 43993 3519 44051 3525
rect 43993 3516 44005 3519
rect 43864 3488 44005 3516
rect 43864 3476 43870 3488
rect 43993 3485 44005 3488
rect 44039 3485 44051 3519
rect 43993 3479 44051 3485
rect 45005 3519 45063 3525
rect 45005 3485 45017 3519
rect 45051 3485 45063 3519
rect 45005 3479 45063 3485
rect 39942 3448 39948 3460
rect 33796 3420 39948 3448
rect 23808 3352 29592 3380
rect 29641 3383 29699 3389
rect 23808 3340 23814 3352
rect 29641 3349 29653 3383
rect 29687 3380 29699 3383
rect 29914 3380 29920 3392
rect 29687 3352 29920 3380
rect 29687 3349 29699 3352
rect 29641 3343 29699 3349
rect 29914 3340 29920 3352
rect 29972 3340 29978 3392
rect 30006 3340 30012 3392
rect 30064 3380 30070 3392
rect 32416 3380 32444 3420
rect 39942 3408 39948 3420
rect 40000 3408 40006 3460
rect 30064 3352 32444 3380
rect 30064 3340 30070 3352
rect 32950 3340 32956 3392
rect 33008 3380 33014 3392
rect 33229 3383 33287 3389
rect 33229 3380 33241 3383
rect 33008 3352 33241 3380
rect 33008 3340 33014 3352
rect 33229 3349 33241 3352
rect 33275 3349 33287 3383
rect 33229 3343 33287 3349
rect 40034 3340 40040 3392
rect 40092 3380 40098 3392
rect 40129 3383 40187 3389
rect 40129 3380 40141 3383
rect 40092 3352 40141 3380
rect 40092 3340 40098 3352
rect 40129 3349 40141 3352
rect 40175 3349 40187 3383
rect 40788 3380 40816 3476
rect 40865 3451 40923 3457
rect 40865 3417 40877 3451
rect 40911 3448 40923 3451
rect 41601 3451 41659 3457
rect 41601 3448 41613 3451
rect 40911 3420 41613 3448
rect 40911 3417 40923 3420
rect 40865 3411 40923 3417
rect 41601 3417 41613 3420
rect 41647 3417 41659 3451
rect 46382 3448 46388 3460
rect 41601 3411 41659 3417
rect 41708 3420 46388 3448
rect 41708 3380 41736 3420
rect 46382 3408 46388 3420
rect 46440 3408 46446 3460
rect 40788 3352 41736 3380
rect 45097 3383 45155 3389
rect 40129 3343 40187 3349
rect 45097 3349 45109 3383
rect 45143 3380 45155 3383
rect 45186 3380 45192 3392
rect 45143 3352 45192 3380
rect 45143 3349 45155 3352
rect 45097 3343 45155 3349
rect 45186 3340 45192 3352
rect 45244 3340 45250 3392
rect 1104 3290 48852 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 48852 3290
rect 1104 3216 48852 3238
rect 3050 3136 3056 3188
rect 3108 3176 3114 3188
rect 19978 3176 19984 3188
rect 3108 3148 19984 3176
rect 3108 3136 3114 3148
rect 19978 3136 19984 3148
rect 20036 3136 20042 3188
rect 20165 3179 20223 3185
rect 20165 3145 20177 3179
rect 20211 3176 20223 3179
rect 20346 3176 20352 3188
rect 20211 3148 20352 3176
rect 20211 3145 20223 3148
rect 20165 3139 20223 3145
rect 20346 3136 20352 3148
rect 20404 3136 20410 3188
rect 20714 3136 20720 3188
rect 20772 3176 20778 3188
rect 22462 3176 22468 3188
rect 20772 3148 22468 3176
rect 20772 3136 20778 3148
rect 22462 3136 22468 3148
rect 22520 3136 22526 3188
rect 22646 3136 22652 3188
rect 22704 3176 22710 3188
rect 30006 3176 30012 3188
rect 22704 3148 30012 3176
rect 22704 3136 22710 3148
rect 30006 3136 30012 3148
rect 30064 3136 30070 3188
rect 34974 3176 34980 3188
rect 31726 3148 34980 3176
rect 1946 3108 1952 3120
rect 1907 3080 1952 3108
rect 1946 3068 1952 3080
rect 2004 3068 2010 3120
rect 6546 3108 6552 3120
rect 6507 3080 6552 3108
rect 6546 3068 6552 3080
rect 6604 3068 6610 3120
rect 12158 3108 12164 3120
rect 12119 3080 12164 3108
rect 12158 3068 12164 3080
rect 12216 3068 12222 3120
rect 14458 3108 14464 3120
rect 14419 3080 14464 3108
rect 14458 3068 14464 3080
rect 14516 3068 14522 3120
rect 17954 3108 17960 3120
rect 17915 3080 17960 3108
rect 17954 3068 17960 3080
rect 18012 3068 18018 3120
rect 20254 3108 20260 3120
rect 20088 3080 20260 3108
rect 3786 3000 3792 3052
rect 3844 3040 3850 3052
rect 4249 3043 4307 3049
rect 4249 3040 4261 3043
rect 3844 3012 4261 3040
rect 3844 3000 3850 3012
rect 4249 3009 4261 3012
rect 4295 3009 4307 3043
rect 4249 3003 4307 3009
rect 8386 3000 8392 3052
rect 8444 3040 8450 3052
rect 8665 3043 8723 3049
rect 8665 3040 8677 3043
rect 8444 3012 8677 3040
rect 8444 3000 8450 3012
rect 8665 3009 8677 3012
rect 8711 3009 8723 3043
rect 11974 3040 11980 3052
rect 11935 3012 11980 3040
rect 8665 3003 8723 3009
rect 11974 3000 11980 3012
rect 12032 3000 12038 3052
rect 14274 3040 14280 3052
rect 14235 3012 14280 3040
rect 14274 3000 14280 3012
rect 14332 3000 14338 3052
rect 17770 3040 17776 3052
rect 17731 3012 17776 3040
rect 17770 3000 17776 3012
rect 17828 3000 17834 3052
rect 20088 3049 20116 3080
rect 20254 3068 20260 3080
rect 20312 3108 20318 3120
rect 23658 3108 23664 3120
rect 20312 3080 22508 3108
rect 23619 3080 23664 3108
rect 20312 3068 20318 3080
rect 20073 3043 20131 3049
rect 20073 3009 20085 3043
rect 20119 3009 20131 3043
rect 21174 3040 21180 3052
rect 21135 3012 21180 3040
rect 20073 3003 20131 3009
rect 21174 3000 21180 3012
rect 21232 3000 21238 3052
rect 1765 2975 1823 2981
rect 1765 2941 1777 2975
rect 1811 2972 1823 2975
rect 2958 2972 2964 2984
rect 1811 2944 2964 2972
rect 1811 2941 1823 2944
rect 1765 2935 1823 2941
rect 2958 2932 2964 2944
rect 3016 2932 3022 2984
rect 3145 2975 3203 2981
rect 3145 2941 3157 2975
rect 3191 2941 3203 2975
rect 3145 2935 3203 2941
rect 5445 2975 5503 2981
rect 5445 2941 5457 2975
rect 5491 2972 5503 2975
rect 6365 2975 6423 2981
rect 6365 2972 6377 2975
rect 5491 2944 6377 2972
rect 5491 2941 5503 2944
rect 5445 2935 5503 2941
rect 6365 2941 6377 2944
rect 6411 2941 6423 2975
rect 6365 2935 6423 2941
rect 6825 2975 6883 2981
rect 6825 2941 6837 2975
rect 6871 2941 6883 2975
rect 12894 2972 12900 2984
rect 12855 2944 12900 2972
rect 6825 2935 6883 2941
rect 1302 2864 1308 2916
rect 1360 2904 1366 2916
rect 3160 2904 3188 2935
rect 1360 2876 3188 2904
rect 1360 2864 1366 2876
rect 5166 2864 5172 2916
rect 5224 2904 5230 2916
rect 6840 2904 6868 2935
rect 12894 2932 12900 2944
rect 12952 2932 12958 2984
rect 15470 2972 15476 2984
rect 15431 2944 15476 2972
rect 15470 2932 15476 2944
rect 15528 2932 15534 2984
rect 18046 2932 18052 2984
rect 18104 2972 18110 2984
rect 18233 2975 18291 2981
rect 18233 2972 18245 2975
rect 18104 2944 18245 2972
rect 18104 2932 18110 2944
rect 18233 2941 18245 2944
rect 18279 2941 18291 2975
rect 22370 2972 22376 2984
rect 18233 2935 18291 2941
rect 21376 2944 22376 2972
rect 8846 2904 8852 2916
rect 5224 2876 6868 2904
rect 8807 2876 8852 2904
rect 5224 2864 5230 2876
rect 8846 2864 8852 2876
rect 8904 2864 8910 2916
rect 10962 2864 10968 2916
rect 11020 2904 11026 2916
rect 17310 2904 17316 2916
rect 11020 2876 17316 2904
rect 11020 2864 11026 2876
rect 17310 2864 17316 2876
rect 17368 2864 17374 2916
rect 17402 2864 17408 2916
rect 17460 2904 17466 2916
rect 21174 2904 21180 2916
rect 17460 2876 21180 2904
rect 17460 2864 17466 2876
rect 21174 2864 21180 2876
rect 21232 2864 21238 2916
rect 11606 2796 11612 2848
rect 11664 2836 11670 2848
rect 15194 2836 15200 2848
rect 11664 2808 15200 2836
rect 11664 2796 11670 2808
rect 15194 2796 15200 2808
rect 15252 2796 15258 2848
rect 17494 2796 17500 2848
rect 17552 2836 17558 2848
rect 21376 2836 21404 2944
rect 22370 2932 22376 2944
rect 22428 2932 22434 2984
rect 22480 2972 22508 3080
rect 23658 3068 23664 3080
rect 23716 3068 23722 3120
rect 29914 3108 29920 3120
rect 29875 3080 29920 3108
rect 29914 3068 29920 3080
rect 29972 3068 29978 3120
rect 22738 3000 22744 3052
rect 22796 3040 22802 3052
rect 23477 3043 23535 3049
rect 23477 3040 23489 3043
rect 22796 3012 23489 3040
rect 22796 3000 22802 3012
rect 23477 3009 23489 3012
rect 23523 3009 23535 3043
rect 23477 3003 23535 3009
rect 25866 3000 25872 3052
rect 25924 3040 25930 3052
rect 26053 3043 26111 3049
rect 26053 3040 26065 3043
rect 25924 3012 26065 3040
rect 25924 3000 25930 3012
rect 26053 3009 26065 3012
rect 26099 3009 26111 3043
rect 26053 3003 26111 3009
rect 28994 3000 29000 3052
rect 29052 3040 29058 3052
rect 29733 3043 29791 3049
rect 29733 3040 29745 3043
rect 29052 3012 29745 3040
rect 29052 3000 29058 3012
rect 29733 3009 29745 3012
rect 29779 3009 29791 3043
rect 29733 3003 29791 3009
rect 23750 2972 23756 2984
rect 22480 2944 23756 2972
rect 23750 2932 23756 2944
rect 23808 2932 23814 2984
rect 23842 2932 23848 2984
rect 23900 2972 23906 2984
rect 23937 2975 23995 2981
rect 23937 2972 23949 2975
rect 23900 2944 23949 2972
rect 23900 2932 23906 2944
rect 23937 2941 23949 2944
rect 23983 2941 23995 2975
rect 30282 2972 30288 2984
rect 30243 2944 30288 2972
rect 23937 2935 23995 2941
rect 30282 2932 30288 2944
rect 30340 2932 30346 2984
rect 31726 2972 31754 3148
rect 34974 3136 34980 3148
rect 35032 3136 35038 3188
rect 35268 3148 45554 3176
rect 32950 3108 32956 3120
rect 32911 3080 32956 3108
rect 32950 3068 32956 3080
rect 33008 3068 33014 3120
rect 35069 3111 35127 3117
rect 35069 3077 35081 3111
rect 35115 3108 35127 3111
rect 35268 3108 35296 3148
rect 35115 3080 35296 3108
rect 35115 3077 35127 3080
rect 35069 3071 35127 3077
rect 35342 3068 35348 3120
rect 35400 3108 35406 3120
rect 35805 3111 35863 3117
rect 35805 3108 35817 3111
rect 35400 3080 35817 3108
rect 35400 3068 35406 3080
rect 35805 3077 35817 3080
rect 35851 3077 35863 3111
rect 37918 3108 37924 3120
rect 37879 3080 37924 3108
rect 35805 3071 35863 3077
rect 37918 3068 37924 3080
rect 37976 3068 37982 3120
rect 40218 3108 40224 3120
rect 40179 3080 40224 3108
rect 40218 3068 40224 3080
rect 40276 3068 40282 3120
rect 43990 3108 43996 3120
rect 43951 3080 43996 3108
rect 43990 3068 43996 3080
rect 44048 3068 44054 3120
rect 45526 3108 45554 3148
rect 45646 3136 45652 3188
rect 45704 3176 45710 3188
rect 46293 3179 46351 3185
rect 46293 3176 46305 3179
rect 45704 3148 46305 3176
rect 45704 3136 45710 3148
rect 46293 3145 46305 3148
rect 46339 3145 46351 3179
rect 46293 3139 46351 3145
rect 47118 3108 47124 3120
rect 45526 3080 47124 3108
rect 47118 3068 47124 3080
rect 47176 3068 47182 3120
rect 32766 3040 32772 3052
rect 32727 3012 32772 3040
rect 32766 3000 32772 3012
rect 32824 3000 32830 3052
rect 35986 3000 35992 3052
rect 36044 3040 36050 3052
rect 36449 3043 36507 3049
rect 36449 3040 36461 3043
rect 36044 3012 36461 3040
rect 36044 3000 36050 3012
rect 36449 3009 36461 3012
rect 36495 3009 36507 3043
rect 37734 3040 37740 3052
rect 37695 3012 37740 3040
rect 36449 3003 36507 3009
rect 37734 3000 37740 3012
rect 37792 3000 37798 3052
rect 40034 3040 40040 3052
rect 39995 3012 40040 3040
rect 40034 3000 40040 3012
rect 40092 3000 40098 3052
rect 42981 3043 43039 3049
rect 42981 3009 42993 3043
rect 43027 3040 43039 3043
rect 43162 3040 43168 3052
rect 43027 3012 43168 3040
rect 43027 3009 43039 3012
rect 42981 3003 43039 3009
rect 43162 3000 43168 3012
rect 43220 3000 43226 3052
rect 43806 3040 43812 3052
rect 43767 3012 43812 3040
rect 43806 3000 43812 3012
rect 43864 3000 43870 3052
rect 45738 3000 45744 3052
rect 45796 3040 45802 3052
rect 46201 3043 46259 3049
rect 46201 3040 46213 3043
rect 45796 3012 46213 3040
rect 45796 3000 45802 3012
rect 46201 3009 46213 3012
rect 46247 3009 46259 3043
rect 46201 3003 46259 3009
rect 47857 3043 47915 3049
rect 47857 3009 47869 3043
rect 47903 3040 47915 3043
rect 49602 3040 49608 3052
rect 47903 3012 49608 3040
rect 47903 3009 47915 3012
rect 47857 3003 47915 3009
rect 49602 3000 49608 3012
rect 49660 3000 49666 3052
rect 33502 2972 33508 2984
rect 30392 2944 31754 2972
rect 33463 2944 33508 2972
rect 21450 2864 21456 2916
rect 21508 2904 21514 2916
rect 30392 2904 30420 2944
rect 33502 2932 33508 2944
rect 33560 2932 33566 2984
rect 35434 2972 35440 2984
rect 35395 2944 35440 2972
rect 35434 2932 35440 2944
rect 35492 2932 35498 2984
rect 39577 2975 39635 2981
rect 39577 2941 39589 2975
rect 39623 2972 39635 2975
rect 39942 2972 39948 2984
rect 39623 2944 39948 2972
rect 39623 2941 39635 2944
rect 39577 2935 39635 2941
rect 39942 2932 39948 2944
rect 40000 2932 40006 2984
rect 41230 2972 41236 2984
rect 41191 2944 41236 2972
rect 41230 2932 41236 2944
rect 41288 2932 41294 2984
rect 44450 2972 44456 2984
rect 44411 2944 44456 2972
rect 44450 2932 44456 2944
rect 44508 2932 44514 2984
rect 34054 2904 34060 2916
rect 21508 2876 30420 2904
rect 30484 2876 34060 2904
rect 21508 2864 21514 2876
rect 17552 2808 21404 2836
rect 17552 2796 17558 2808
rect 22462 2796 22468 2848
rect 22520 2836 22526 2848
rect 30484 2836 30512 2876
rect 34054 2864 34060 2876
rect 34112 2864 34118 2916
rect 34238 2864 34244 2916
rect 34296 2904 34302 2916
rect 34296 2876 35572 2904
rect 34296 2864 34302 2876
rect 22520 2808 30512 2836
rect 22520 2796 22526 2808
rect 34514 2796 34520 2848
rect 34572 2836 34578 2848
rect 35207 2839 35265 2845
rect 35207 2836 35219 2839
rect 34572 2808 35219 2836
rect 34572 2796 34578 2808
rect 35207 2805 35219 2808
rect 35253 2805 35265 2839
rect 35207 2799 35265 2805
rect 35342 2796 35348 2848
rect 35400 2836 35406 2848
rect 35544 2836 35572 2876
rect 35618 2864 35624 2916
rect 35676 2904 35682 2916
rect 48041 2907 48099 2913
rect 48041 2904 48053 2907
rect 35676 2876 48053 2904
rect 35676 2864 35682 2876
rect 48041 2873 48053 2876
rect 48087 2873 48099 2907
rect 48041 2867 48099 2873
rect 43073 2839 43131 2845
rect 43073 2836 43085 2839
rect 35400 2808 35445 2836
rect 35544 2808 43085 2836
rect 35400 2796 35406 2808
rect 43073 2805 43085 2808
rect 43119 2805 43131 2839
rect 43073 2799 43131 2805
rect 1104 2746 48852 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 48852 2746
rect 1104 2672 48852 2694
rect 2958 2592 2964 2644
rect 3016 2632 3022 2644
rect 3053 2635 3111 2641
rect 3053 2632 3065 2635
rect 3016 2604 3065 2632
rect 3016 2592 3022 2604
rect 3053 2601 3065 2604
rect 3099 2601 3111 2635
rect 3053 2595 3111 2601
rect 9171 2635 9229 2641
rect 9171 2601 9183 2635
rect 9217 2632 9229 2635
rect 20257 2635 20315 2641
rect 9217 2604 16574 2632
rect 9217 2601 9229 2604
rect 9171 2595 9229 2601
rect 1581 2567 1639 2573
rect 1581 2533 1593 2567
rect 1627 2564 1639 2567
rect 14734 2564 14740 2576
rect 1627 2536 12020 2564
rect 14695 2536 14740 2564
rect 1627 2533 1639 2536
rect 1581 2527 1639 2533
rect 11698 2496 11704 2508
rect 11659 2468 11704 2496
rect 11698 2456 11704 2468
rect 11756 2456 11762 2508
rect 11882 2496 11888 2508
rect 11843 2468 11888 2496
rect 11882 2456 11888 2468
rect 11940 2456 11946 2508
rect 11992 2496 12020 2536
rect 14734 2524 14740 2536
rect 14792 2524 14798 2576
rect 16546 2564 16574 2604
rect 20257 2601 20269 2635
rect 20303 2632 20315 2635
rect 20438 2632 20444 2644
rect 20303 2604 20444 2632
rect 20303 2601 20315 2604
rect 20257 2595 20315 2601
rect 20438 2592 20444 2604
rect 20496 2592 20502 2644
rect 22554 2592 22560 2644
rect 22612 2632 22618 2644
rect 22833 2635 22891 2641
rect 22833 2632 22845 2635
rect 22612 2604 22845 2632
rect 22612 2592 22618 2604
rect 22833 2601 22845 2604
rect 22879 2601 22891 2635
rect 22833 2595 22891 2601
rect 23385 2635 23443 2641
rect 23385 2601 23397 2635
rect 23431 2632 23443 2635
rect 23566 2632 23572 2644
rect 23431 2604 23572 2632
rect 23431 2601 23443 2604
rect 23385 2595 23443 2601
rect 23566 2592 23572 2604
rect 23624 2592 23630 2644
rect 26326 2592 26332 2644
rect 26384 2632 26390 2644
rect 27341 2635 27399 2641
rect 27341 2632 27353 2635
rect 26384 2604 27353 2632
rect 26384 2592 26390 2604
rect 27341 2601 27353 2604
rect 27387 2601 27399 2635
rect 27341 2595 27399 2601
rect 28074 2592 28080 2644
rect 28132 2632 28138 2644
rect 28132 2604 30420 2632
rect 28132 2592 28138 2604
rect 19334 2564 19340 2576
rect 16546 2536 19340 2564
rect 19334 2524 19340 2536
rect 19392 2524 19398 2576
rect 24673 2567 24731 2573
rect 24673 2533 24685 2567
rect 24719 2564 24731 2567
rect 28902 2564 28908 2576
rect 24719 2536 28908 2564
rect 24719 2533 24731 2536
rect 24673 2527 24731 2533
rect 28902 2524 28908 2536
rect 28960 2524 28966 2576
rect 30392 2564 30420 2604
rect 30466 2592 30472 2644
rect 30524 2632 30530 2644
rect 46382 2632 46388 2644
rect 30524 2604 46388 2632
rect 30524 2592 30530 2604
rect 46382 2592 46388 2604
rect 46440 2592 46446 2644
rect 33137 2567 33195 2573
rect 33137 2564 33149 2567
rect 30392 2536 33149 2564
rect 33137 2533 33149 2536
rect 33183 2533 33195 2567
rect 33137 2527 33195 2533
rect 33965 2567 34023 2573
rect 33965 2533 33977 2567
rect 34011 2564 34023 2567
rect 34514 2564 34520 2576
rect 34011 2536 34520 2564
rect 34011 2533 34023 2536
rect 33965 2527 34023 2533
rect 34514 2524 34520 2536
rect 34572 2524 34578 2576
rect 34885 2567 34943 2573
rect 34885 2533 34897 2567
rect 34931 2564 34943 2567
rect 35434 2564 35440 2576
rect 34931 2536 35440 2564
rect 34931 2533 34943 2536
rect 34885 2527 34943 2533
rect 35434 2524 35440 2536
rect 35492 2524 35498 2576
rect 38746 2564 38752 2576
rect 38707 2536 38752 2564
rect 38746 2524 38752 2536
rect 38804 2524 38810 2576
rect 19426 2496 19432 2508
rect 11992 2468 19432 2496
rect 19426 2456 19432 2468
rect 19484 2456 19490 2508
rect 20530 2456 20536 2508
rect 20588 2496 20594 2508
rect 25501 2499 25559 2505
rect 25501 2496 25513 2499
rect 20588 2468 25513 2496
rect 20588 2456 20594 2468
rect 25501 2465 25513 2468
rect 25547 2465 25559 2499
rect 25501 2459 25559 2465
rect 30374 2456 30380 2508
rect 30432 2496 30438 2508
rect 30469 2499 30527 2505
rect 30469 2496 30481 2499
rect 30432 2468 30481 2496
rect 30432 2456 30438 2468
rect 30469 2465 30481 2468
rect 30515 2465 30527 2499
rect 30469 2459 30527 2465
rect 41966 2456 41972 2508
rect 42024 2496 42030 2508
rect 42429 2499 42487 2505
rect 42429 2496 42441 2499
rect 42024 2468 42441 2496
rect 42024 2456 42030 2468
rect 42429 2465 42441 2468
rect 42475 2465 42487 2499
rect 42610 2496 42616 2508
rect 42571 2468 42616 2496
rect 42429 2459 42487 2465
rect 42610 2456 42616 2468
rect 42668 2456 42674 2508
rect 42702 2456 42708 2508
rect 42760 2496 42766 2508
rect 42889 2499 42947 2505
rect 42889 2496 42901 2499
rect 42760 2468 42901 2496
rect 42760 2456 42766 2468
rect 42889 2465 42901 2468
rect 42935 2465 42947 2499
rect 42889 2459 42947 2465
rect 44634 2456 44640 2508
rect 44692 2496 44698 2508
rect 45005 2499 45063 2505
rect 45005 2496 45017 2499
rect 44692 2468 45017 2496
rect 44692 2456 44698 2468
rect 45005 2465 45017 2468
rect 45051 2465 45063 2499
rect 45186 2496 45192 2508
rect 45147 2468 45192 2496
rect 45005 2459 45063 2465
rect 45186 2456 45192 2468
rect 45244 2456 45250 2508
rect 45370 2456 45376 2508
rect 45428 2496 45434 2508
rect 45557 2499 45615 2505
rect 45557 2496 45569 2499
rect 45428 2468 45569 2496
rect 45428 2456 45434 2468
rect 45557 2465 45569 2468
rect 45603 2465 45615 2499
rect 45557 2459 45615 2465
rect 1394 2428 1400 2440
rect 1355 2400 1400 2428
rect 1394 2388 1400 2400
rect 1452 2388 1458 2440
rect 1946 2388 1952 2440
rect 2004 2428 2010 2440
rect 2133 2431 2191 2437
rect 2133 2428 2145 2431
rect 2004 2400 2145 2428
rect 2004 2388 2010 2400
rect 2133 2397 2145 2400
rect 2179 2397 2191 2431
rect 2133 2391 2191 2397
rect 7098 2388 7104 2440
rect 7156 2428 7162 2440
rect 7193 2431 7251 2437
rect 7193 2428 7205 2431
rect 7156 2400 7205 2428
rect 7156 2388 7162 2400
rect 7193 2397 7205 2400
rect 7239 2397 7251 2431
rect 7466 2428 7472 2440
rect 7427 2400 7472 2428
rect 7193 2391 7251 2397
rect 7466 2388 7472 2400
rect 7524 2388 7530 2440
rect 7742 2388 7748 2440
rect 7800 2428 7806 2440
rect 8941 2431 8999 2437
rect 8941 2428 8953 2431
rect 7800 2400 8953 2428
rect 7800 2388 7806 2400
rect 8941 2397 8953 2400
rect 8987 2397 8999 2431
rect 8941 2391 8999 2397
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 10229 2431 10287 2437
rect 10229 2428 10241 2431
rect 9732 2400 10241 2428
rect 9732 2388 9738 2400
rect 10229 2397 10241 2400
rect 10275 2397 10287 2431
rect 10229 2391 10287 2397
rect 13648 2400 16574 2428
rect 4522 2320 4528 2372
rect 4580 2360 4586 2372
rect 4709 2363 4767 2369
rect 4709 2360 4721 2363
rect 4580 2332 4721 2360
rect 4580 2320 4586 2332
rect 4709 2329 4721 2332
rect 4755 2329 4767 2363
rect 4709 2323 4767 2329
rect 4816 2332 11744 2360
rect 2317 2295 2375 2301
rect 2317 2261 2329 2295
rect 2363 2292 2375 2295
rect 4816 2292 4844 2332
rect 4982 2292 4988 2304
rect 2363 2264 4844 2292
rect 4943 2264 4988 2292
rect 2363 2261 2375 2264
rect 2317 2255 2375 2261
rect 4982 2252 4988 2264
rect 5040 2252 5046 2304
rect 10410 2292 10416 2304
rect 10371 2264 10416 2292
rect 10410 2252 10416 2264
rect 10468 2252 10474 2304
rect 11716 2292 11744 2332
rect 12250 2320 12256 2372
rect 12308 2360 12314 2372
rect 13541 2363 13599 2369
rect 13541 2360 13553 2363
rect 12308 2332 13553 2360
rect 12308 2320 12314 2332
rect 13541 2329 13553 2332
rect 13587 2329 13599 2363
rect 13541 2323 13599 2329
rect 13648 2292 13676 2400
rect 14182 2320 14188 2372
rect 14240 2360 14246 2372
rect 14553 2363 14611 2369
rect 14553 2360 14565 2363
rect 14240 2332 14565 2360
rect 14240 2320 14246 2332
rect 14553 2329 14565 2332
rect 14599 2329 14611 2363
rect 16546 2360 16574 2400
rect 17402 2388 17408 2440
rect 17460 2428 17466 2440
rect 17497 2431 17555 2437
rect 17497 2428 17509 2431
rect 17460 2400 17509 2428
rect 17460 2388 17466 2400
rect 17497 2397 17509 2400
rect 17543 2397 17555 2431
rect 17770 2428 17776 2440
rect 17731 2400 17776 2428
rect 17497 2391 17555 2397
rect 17770 2388 17776 2400
rect 17828 2388 17834 2440
rect 19978 2388 19984 2440
rect 20036 2428 20042 2440
rect 20073 2431 20131 2437
rect 20073 2428 20085 2431
rect 20036 2400 20085 2428
rect 20036 2388 20042 2400
rect 20073 2397 20085 2400
rect 20119 2397 20131 2431
rect 20073 2391 20131 2397
rect 20456 2400 22876 2428
rect 20456 2360 20484 2400
rect 16546 2332 20484 2360
rect 14553 2323 14611 2329
rect 22554 2320 22560 2372
rect 22612 2360 22618 2372
rect 22741 2363 22799 2369
rect 22741 2360 22753 2363
rect 22612 2332 22753 2360
rect 22612 2320 22618 2332
rect 22741 2329 22753 2332
rect 22787 2329 22799 2363
rect 22848 2360 22876 2400
rect 23198 2388 23204 2440
rect 23256 2428 23262 2440
rect 23569 2431 23627 2437
rect 23569 2428 23581 2431
rect 23256 2400 23581 2428
rect 23256 2388 23262 2400
rect 23569 2397 23581 2400
rect 23615 2397 23627 2431
rect 24394 2428 24400 2440
rect 23569 2391 23627 2397
rect 23676 2400 24400 2428
rect 23676 2360 23704 2400
rect 24394 2388 24400 2400
rect 24452 2388 24458 2440
rect 27062 2388 27068 2440
rect 27120 2428 27126 2440
rect 27157 2431 27215 2437
rect 27157 2428 27169 2431
rect 27120 2400 27169 2428
rect 27120 2388 27126 2400
rect 27157 2397 27169 2400
rect 27203 2397 27215 2431
rect 27157 2391 27215 2397
rect 32858 2388 32864 2440
rect 32916 2428 32922 2440
rect 32953 2431 33011 2437
rect 32953 2428 32965 2431
rect 32916 2400 32965 2428
rect 32916 2388 32922 2400
rect 32953 2397 32965 2400
rect 32999 2397 33011 2431
rect 34146 2428 34152 2440
rect 34107 2400 34152 2428
rect 32953 2391 33011 2397
rect 34146 2388 34152 2400
rect 34204 2388 34210 2440
rect 34790 2388 34796 2440
rect 34848 2428 34854 2440
rect 35069 2431 35127 2437
rect 35069 2428 35081 2431
rect 34848 2400 35081 2428
rect 34848 2388 34854 2400
rect 35069 2397 35081 2400
rect 35115 2397 35127 2431
rect 35069 2391 35127 2397
rect 38654 2388 38660 2440
rect 38712 2428 38718 2440
rect 38933 2431 38991 2437
rect 38933 2428 38945 2431
rect 38712 2400 38945 2428
rect 38712 2388 38718 2400
rect 38933 2397 38945 2400
rect 38979 2397 38991 2431
rect 38933 2391 38991 2397
rect 24486 2360 24492 2372
rect 22848 2332 23704 2360
rect 24447 2332 24492 2360
rect 22741 2323 22799 2329
rect 24486 2320 24492 2332
rect 24544 2320 24550 2372
rect 25130 2320 25136 2372
rect 25188 2360 25194 2372
rect 25317 2363 25375 2369
rect 25317 2360 25329 2363
rect 25188 2332 25329 2360
rect 25188 2320 25194 2332
rect 25317 2329 25329 2332
rect 25363 2329 25375 2363
rect 25317 2323 25375 2329
rect 26206 2332 27476 2360
rect 11716 2264 13676 2292
rect 20070 2252 20076 2304
rect 20128 2292 20134 2304
rect 26206 2292 26234 2332
rect 20128 2264 26234 2292
rect 27448 2292 27476 2332
rect 27706 2320 27712 2372
rect 27764 2360 27770 2372
rect 27985 2363 28043 2369
rect 27985 2360 27997 2363
rect 27764 2332 27997 2360
rect 27764 2320 27770 2332
rect 27985 2329 27997 2332
rect 28031 2329 28043 2363
rect 27985 2323 28043 2329
rect 36078 2320 36084 2372
rect 36136 2360 36142 2372
rect 36265 2363 36323 2369
rect 36265 2360 36277 2363
rect 36136 2332 36277 2360
rect 36136 2320 36142 2332
rect 36265 2329 36277 2332
rect 36311 2329 36323 2363
rect 47762 2360 47768 2372
rect 47723 2332 47768 2360
rect 36265 2323 36323 2329
rect 47762 2320 47768 2332
rect 47820 2320 47826 2372
rect 28077 2295 28135 2301
rect 28077 2292 28089 2295
rect 27448 2264 28089 2292
rect 20128 2252 20134 2264
rect 28077 2261 28089 2264
rect 28123 2261 28135 2295
rect 28077 2255 28135 2261
rect 28166 2252 28172 2304
rect 28224 2292 28230 2304
rect 36357 2295 36415 2301
rect 36357 2292 36369 2295
rect 28224 2264 36369 2292
rect 28224 2252 28230 2264
rect 36357 2261 36369 2264
rect 36403 2261 36415 2295
rect 47854 2292 47860 2304
rect 47815 2264 47860 2292
rect 36357 2255 36415 2261
rect 47854 2252 47860 2264
rect 47912 2252 47918 2304
rect 1104 2202 48852 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 48852 2202
rect 1104 2128 48852 2150
rect 3418 1980 3424 2032
rect 3476 2020 3482 2032
rect 39022 2020 39028 2032
rect 3476 1992 39028 2020
rect 3476 1980 3482 1992
rect 39022 1980 39028 1992
rect 39080 1980 39086 2032
rect 7466 1912 7472 1964
rect 7524 1952 7530 1964
rect 22278 1952 22284 1964
rect 7524 1924 22284 1952
rect 7524 1912 7530 1924
rect 22278 1912 22284 1924
rect 22336 1912 22342 1964
rect 23934 1912 23940 1964
rect 23992 1952 23998 1964
rect 47854 1952 47860 1964
rect 23992 1924 47860 1952
rect 23992 1912 23998 1924
rect 47854 1912 47860 1924
rect 47912 1912 47918 1964
rect 4982 1844 4988 1896
rect 5040 1884 5046 1896
rect 28442 1884 28448 1896
rect 5040 1856 28448 1884
rect 5040 1844 5046 1856
rect 28442 1844 28448 1856
rect 28500 1844 28506 1896
rect 17770 1776 17776 1828
rect 17828 1816 17834 1828
rect 35342 1816 35348 1828
rect 17828 1788 35348 1816
rect 17828 1776 17834 1788
rect 35342 1776 35348 1788
rect 35400 1776 35406 1828
<< via1 >>
rect 3424 49852 3476 49904
rect 8208 49852 8260 49904
rect 43996 49716 44048 49768
rect 46756 49716 46808 49768
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 1308 49240 1360 49292
rect 5816 49240 5868 49292
rect 10324 49240 10376 49292
rect 12348 49240 12400 49292
rect 18052 49240 18104 49292
rect 22008 49283 22060 49292
rect 22008 49249 22017 49283
rect 22017 49249 22051 49283
rect 22051 49249 22060 49283
rect 22008 49240 22060 49249
rect 24216 49240 24268 49292
rect 27620 49283 27672 49292
rect 27620 49249 27629 49283
rect 27629 49249 27663 49283
rect 27663 49249 27672 49283
rect 27620 49240 27672 49249
rect 43168 49283 43220 49292
rect 43168 49249 43177 49283
rect 43177 49249 43211 49283
rect 43211 49249 43220 49283
rect 43168 49240 43220 49249
rect 48320 49240 48372 49292
rect 3608 49172 3660 49224
rect 6552 49215 6604 49224
rect 6552 49181 6561 49215
rect 6561 49181 6595 49215
rect 6595 49181 6604 49215
rect 6552 49172 6604 49181
rect 7472 49215 7524 49224
rect 7472 49181 7481 49215
rect 7481 49181 7515 49215
rect 7515 49181 7524 49215
rect 7472 49172 7524 49181
rect 14188 49172 14240 49224
rect 16580 49172 16632 49224
rect 19340 49215 19392 49224
rect 2596 49104 2648 49156
rect 4620 49147 4672 49156
rect 4620 49113 4629 49147
rect 4629 49113 4663 49147
rect 4663 49113 4672 49147
rect 4620 49104 4672 49113
rect 5172 49147 5224 49156
rect 5172 49113 5181 49147
rect 5181 49113 5215 49147
rect 5215 49113 5224 49147
rect 5172 49104 5224 49113
rect 11704 49147 11756 49156
rect 11704 49113 11713 49147
rect 11713 49113 11747 49147
rect 11747 49113 11756 49147
rect 11704 49104 11756 49113
rect 19340 49181 19349 49215
rect 19349 49181 19383 49215
rect 19383 49181 19392 49215
rect 19340 49172 19392 49181
rect 20168 49215 20220 49224
rect 20168 49181 20177 49215
rect 20177 49181 20211 49215
rect 20211 49181 20220 49215
rect 20168 49172 20220 49181
rect 22284 49215 22336 49224
rect 22284 49181 22293 49215
rect 22293 49181 22327 49215
rect 22327 49181 22336 49215
rect 22284 49172 22336 49181
rect 23848 49215 23900 49224
rect 23848 49181 23857 49215
rect 23857 49181 23891 49215
rect 23891 49181 23900 49215
rect 23848 49172 23900 49181
rect 24676 49215 24728 49224
rect 24676 49181 24685 49215
rect 24685 49181 24719 49215
rect 24719 49181 24728 49215
rect 24676 49172 24728 49181
rect 26424 49215 26476 49224
rect 26424 49181 26433 49215
rect 26433 49181 26467 49215
rect 26467 49181 26476 49215
rect 26424 49172 26476 49181
rect 26976 49215 27028 49224
rect 26976 49181 26985 49215
rect 26985 49181 27019 49215
rect 27019 49181 27028 49215
rect 26976 49172 27028 49181
rect 29000 49172 29052 49224
rect 24492 49104 24544 49156
rect 27160 49147 27212 49156
rect 27160 49113 27169 49147
rect 27169 49113 27203 49147
rect 27203 49113 27212 49147
rect 27160 49104 27212 49113
rect 29736 49104 29788 49156
rect 33508 49172 33560 49224
rect 34888 49172 34940 49224
rect 36268 49215 36320 49224
rect 36268 49181 36277 49215
rect 36277 49181 36311 49215
rect 36311 49181 36320 49215
rect 36268 49172 36320 49181
rect 38108 49215 38160 49224
rect 38108 49181 38117 49215
rect 38117 49181 38151 49215
rect 38151 49181 38160 49215
rect 38108 49172 38160 49181
rect 40776 49215 40828 49224
rect 40776 49181 40785 49215
rect 40785 49181 40819 49215
rect 40819 49181 40828 49215
rect 40776 49172 40828 49181
rect 41604 49215 41656 49224
rect 41604 49181 41613 49215
rect 41613 49181 41647 49215
rect 41647 49181 41656 49215
rect 41604 49172 41656 49181
rect 42432 49215 42484 49224
rect 42432 49181 42441 49215
rect 42441 49181 42475 49215
rect 42475 49181 42484 49215
rect 42432 49172 42484 49181
rect 47768 49215 47820 49224
rect 41420 49104 41472 49156
rect 3976 49036 4028 49088
rect 5264 49079 5316 49088
rect 5264 49045 5273 49079
rect 5273 49045 5307 49079
rect 5307 49045 5316 49079
rect 5264 49036 5316 49045
rect 6736 49079 6788 49088
rect 6736 49045 6745 49079
rect 6745 49045 6779 49079
rect 6779 49045 6788 49079
rect 6736 49036 6788 49045
rect 10140 49079 10192 49088
rect 10140 49045 10149 49079
rect 10149 49045 10183 49079
rect 10183 49045 10192 49079
rect 10140 49036 10192 49045
rect 15016 49079 15068 49088
rect 15016 49045 15025 49079
rect 15025 49045 15059 49079
rect 15059 49045 15068 49079
rect 15016 49036 15068 49045
rect 17224 49079 17276 49088
rect 17224 49045 17233 49079
rect 17233 49045 17267 49079
rect 17267 49045 17276 49079
rect 17224 49036 17276 49045
rect 20076 49036 20128 49088
rect 20260 49079 20312 49088
rect 20260 49045 20269 49079
rect 20269 49045 20303 49079
rect 20303 49045 20312 49079
rect 20260 49036 20312 49045
rect 29276 49036 29328 49088
rect 32128 49079 32180 49088
rect 32128 49045 32137 49079
rect 32137 49045 32171 49079
rect 32171 49045 32180 49079
rect 32128 49036 32180 49045
rect 38292 49079 38344 49088
rect 38292 49045 38301 49079
rect 38301 49045 38335 49079
rect 38335 49045 38344 49079
rect 38292 49036 38344 49045
rect 40868 49079 40920 49088
rect 40868 49045 40877 49079
rect 40877 49045 40911 49079
rect 40911 49045 40920 49079
rect 40868 49036 40920 49045
rect 41604 49036 41656 49088
rect 47768 49181 47777 49215
rect 47777 49181 47811 49215
rect 47811 49181 47820 49215
rect 47768 49172 47820 49181
rect 45744 49104 45796 49156
rect 45284 49036 45336 49088
rect 47124 49036 47176 49088
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 24676 48832 24728 48884
rect 30012 48832 30064 48884
rect 20 48764 72 48816
rect 664 48696 716 48748
rect 3884 48764 3936 48816
rect 1492 48628 1544 48680
rect 3148 48671 3200 48680
rect 3148 48637 3157 48671
rect 3157 48637 3191 48671
rect 3191 48637 3200 48671
rect 3148 48628 3200 48637
rect 4068 48628 4120 48680
rect 4160 48671 4212 48680
rect 4160 48637 4169 48671
rect 4169 48637 4203 48671
rect 4203 48637 4212 48671
rect 4896 48764 4948 48816
rect 7472 48764 7524 48816
rect 8208 48764 8260 48816
rect 4160 48628 4212 48637
rect 5540 48628 5592 48680
rect 6920 48671 6972 48680
rect 6920 48637 6929 48671
rect 6929 48637 6963 48671
rect 6963 48637 6972 48671
rect 7196 48671 7248 48680
rect 6920 48628 6972 48637
rect 7196 48637 7205 48671
rect 7205 48637 7239 48671
rect 7239 48637 7248 48671
rect 7196 48628 7248 48637
rect 9128 48671 9180 48680
rect 9128 48637 9137 48671
rect 9137 48637 9171 48671
rect 9171 48637 9180 48671
rect 9128 48628 9180 48637
rect 10232 48628 10284 48680
rect 13820 48764 13872 48816
rect 11612 48739 11664 48748
rect 11612 48705 11621 48739
rect 11621 48705 11655 48739
rect 11655 48705 11664 48739
rect 11612 48696 11664 48705
rect 12348 48739 12400 48748
rect 12348 48705 12357 48739
rect 12357 48705 12391 48739
rect 12391 48705 12400 48739
rect 12348 48696 12400 48705
rect 19432 48764 19484 48816
rect 31944 48764 31996 48816
rect 25412 48696 25464 48748
rect 26424 48696 26476 48748
rect 29736 48739 29788 48748
rect 29736 48705 29745 48739
rect 29745 48705 29779 48739
rect 29779 48705 29788 48739
rect 29736 48696 29788 48705
rect 32128 48739 32180 48748
rect 32128 48705 32137 48739
rect 32137 48705 32171 48739
rect 32171 48705 32180 48739
rect 32128 48696 32180 48705
rect 34888 48739 34940 48748
rect 34888 48705 34897 48739
rect 34897 48705 34931 48739
rect 34931 48705 34940 48739
rect 34888 48696 34940 48705
rect 42340 48696 42392 48748
rect 46296 48832 46348 48884
rect 44456 48764 44508 48816
rect 48964 48764 49016 48816
rect 46756 48739 46808 48748
rect 46756 48705 46765 48739
rect 46765 48705 46799 48739
rect 46799 48705 46808 48739
rect 46756 48696 46808 48705
rect 12532 48671 12584 48680
rect 12532 48637 12541 48671
rect 12541 48637 12575 48671
rect 12575 48637 12584 48671
rect 12532 48628 12584 48637
rect 12624 48628 12676 48680
rect 16856 48671 16908 48680
rect 16856 48637 16865 48671
rect 16865 48637 16899 48671
rect 16899 48637 16908 48671
rect 16856 48628 16908 48637
rect 16948 48628 17000 48680
rect 19524 48628 19576 48680
rect 20628 48628 20680 48680
rect 22744 48671 22796 48680
rect 22744 48637 22753 48671
rect 22753 48637 22787 48671
rect 22787 48637 22796 48671
rect 22744 48628 22796 48637
rect 23480 48671 23532 48680
rect 23480 48637 23489 48671
rect 23489 48637 23523 48671
rect 23523 48637 23532 48671
rect 23480 48628 23532 48637
rect 26516 48628 26568 48680
rect 27620 48671 27672 48680
rect 27620 48637 27629 48671
rect 27629 48637 27663 48671
rect 27663 48637 27672 48671
rect 27620 48628 27672 48637
rect 27896 48671 27948 48680
rect 27896 48637 27905 48671
rect 27905 48637 27939 48671
rect 27939 48637 27948 48671
rect 27896 48628 27948 48637
rect 30564 48628 30616 48680
rect 32312 48671 32364 48680
rect 32312 48637 32321 48671
rect 32321 48637 32355 48671
rect 32355 48637 32364 48671
rect 32312 48628 32364 48637
rect 32864 48671 32916 48680
rect 32864 48637 32873 48671
rect 32873 48637 32907 48671
rect 32907 48637 32916 48671
rect 32864 48628 32916 48637
rect 36084 48671 36136 48680
rect 30748 48560 30800 48612
rect 5632 48535 5684 48544
rect 5632 48501 5641 48535
rect 5641 48501 5675 48535
rect 5675 48501 5684 48535
rect 5632 48492 5684 48501
rect 11796 48535 11848 48544
rect 11796 48501 11805 48535
rect 11805 48501 11839 48535
rect 11839 48501 11848 48535
rect 11796 48492 11848 48501
rect 14832 48535 14884 48544
rect 14832 48501 14841 48535
rect 14841 48501 14875 48535
rect 14875 48501 14884 48535
rect 14832 48492 14884 48501
rect 27528 48492 27580 48544
rect 36084 48637 36093 48671
rect 36093 48637 36127 48671
rect 36127 48637 36136 48671
rect 36084 48628 36136 48637
rect 39488 48671 39540 48680
rect 39488 48637 39497 48671
rect 39497 48637 39531 48671
rect 39531 48637 39540 48671
rect 39488 48628 39540 48637
rect 40040 48671 40092 48680
rect 40040 48637 40049 48671
rect 40049 48637 40083 48671
rect 40083 48637 40092 48671
rect 40040 48628 40092 48637
rect 44456 48671 44508 48680
rect 44456 48637 44465 48671
rect 44465 48637 44499 48671
rect 44499 48637 44508 48671
rect 44456 48628 44508 48637
rect 44640 48671 44692 48680
rect 44640 48637 44649 48671
rect 44649 48637 44683 48671
rect 44683 48637 44692 48671
rect 44640 48628 44692 48637
rect 45836 48671 45888 48680
rect 45836 48637 45845 48671
rect 45845 48637 45879 48671
rect 45879 48637 45888 48671
rect 45836 48628 45888 48637
rect 35992 48492 36044 48544
rect 37648 48492 37700 48544
rect 38568 48492 38620 48544
rect 41788 48492 41840 48544
rect 42800 48492 42852 48544
rect 43904 48535 43956 48544
rect 43904 48501 43913 48535
rect 43913 48501 43947 48535
rect 43947 48501 43956 48535
rect 43904 48492 43956 48501
rect 46940 48535 46992 48544
rect 46940 48501 46949 48535
rect 46949 48501 46983 48535
rect 46983 48501 46992 48535
rect 46940 48492 46992 48501
rect 47216 48492 47268 48544
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 3148 48288 3200 48340
rect 6920 48288 6972 48340
rect 9128 48288 9180 48340
rect 16856 48331 16908 48340
rect 16856 48297 16865 48331
rect 16865 48297 16899 48331
rect 16899 48297 16908 48331
rect 16856 48288 16908 48297
rect 39488 48288 39540 48340
rect 44640 48288 44692 48340
rect 1952 48220 2004 48272
rect 5172 48220 5224 48272
rect 9680 48220 9732 48272
rect 2780 48195 2832 48204
rect 2780 48161 2789 48195
rect 2789 48161 2823 48195
rect 2823 48161 2832 48195
rect 2780 48152 2832 48161
rect 5816 48152 5868 48204
rect 10140 48195 10192 48204
rect 10140 48161 10149 48195
rect 10149 48161 10183 48195
rect 10183 48161 10192 48195
rect 10140 48152 10192 48161
rect 11704 48220 11756 48272
rect 19432 48263 19484 48272
rect 14924 48195 14976 48204
rect 14924 48161 14933 48195
rect 14933 48161 14967 48195
rect 14967 48161 14976 48195
rect 14924 48152 14976 48161
rect 1400 48127 1452 48136
rect 1400 48093 1409 48127
rect 1409 48093 1443 48127
rect 1443 48093 1452 48127
rect 1400 48084 1452 48093
rect 7012 48127 7064 48136
rect 7012 48093 7021 48127
rect 7021 48093 7055 48127
rect 7055 48093 7064 48127
rect 7012 48084 7064 48093
rect 7380 48084 7432 48136
rect 13084 48127 13136 48136
rect 13084 48093 13093 48127
rect 13093 48093 13127 48127
rect 13127 48093 13136 48127
rect 13084 48084 13136 48093
rect 14464 48127 14516 48136
rect 14464 48093 14473 48127
rect 14473 48093 14507 48127
rect 14507 48093 14516 48127
rect 14464 48084 14516 48093
rect 1584 48059 1636 48068
rect 1584 48025 1593 48059
rect 1593 48025 1627 48059
rect 1627 48025 1636 48059
rect 1584 48016 1636 48025
rect 6184 48016 6236 48068
rect 3792 47948 3844 48000
rect 10876 48016 10928 48068
rect 14372 48016 14424 48068
rect 6644 47948 6696 48000
rect 10508 47948 10560 48000
rect 14924 47948 14976 48000
rect 19432 48229 19441 48263
rect 19441 48229 19475 48263
rect 19475 48229 19484 48263
rect 19432 48220 19484 48229
rect 19984 48220 20036 48272
rect 17592 48152 17644 48204
rect 22100 48152 22152 48204
rect 22560 48195 22612 48204
rect 22560 48161 22569 48195
rect 22569 48161 22603 48195
rect 22603 48161 22612 48195
rect 22560 48152 22612 48161
rect 23848 48152 23900 48204
rect 24584 48152 24636 48204
rect 22008 48059 22060 48068
rect 22008 48025 22017 48059
rect 22017 48025 22051 48059
rect 22051 48025 22060 48059
rect 22008 48016 22060 48025
rect 22100 48016 22152 48068
rect 24308 48084 24360 48136
rect 24216 48016 24268 48068
rect 24676 48016 24728 48068
rect 28080 48152 28132 48204
rect 28356 48195 28408 48204
rect 28356 48161 28365 48195
rect 28365 48161 28399 48195
rect 28399 48161 28408 48195
rect 28356 48152 28408 48161
rect 26516 48084 26568 48136
rect 27896 48016 27948 48068
rect 28172 48016 28224 48068
rect 29828 48152 29880 48204
rect 29920 48152 29972 48204
rect 30932 48152 30984 48204
rect 36268 48152 36320 48204
rect 36728 48195 36780 48204
rect 36728 48161 36737 48195
rect 36737 48161 36771 48195
rect 36771 48161 36780 48195
rect 36728 48152 36780 48161
rect 37280 48220 37332 48272
rect 41236 48220 41288 48272
rect 42432 48220 42484 48272
rect 41420 48152 41472 48204
rect 41788 48195 41840 48204
rect 41788 48161 41797 48195
rect 41797 48161 41831 48195
rect 41831 48161 41840 48195
rect 41788 48152 41840 48161
rect 42524 48195 42576 48204
rect 42524 48161 42533 48195
rect 42533 48161 42567 48195
rect 42567 48161 42576 48195
rect 42524 48152 42576 48161
rect 46296 48195 46348 48204
rect 46296 48161 46305 48195
rect 46305 48161 46339 48195
rect 46339 48161 46348 48195
rect 46296 48152 46348 48161
rect 46848 48195 46900 48204
rect 46848 48161 46857 48195
rect 46857 48161 46891 48195
rect 46891 48161 46900 48195
rect 46848 48152 46900 48161
rect 31852 48127 31904 48136
rect 31852 48093 31861 48127
rect 31861 48093 31895 48127
rect 31895 48093 31904 48127
rect 31852 48084 31904 48093
rect 35808 48084 35860 48136
rect 44088 48127 44140 48136
rect 29736 48059 29788 48068
rect 29736 48025 29745 48059
rect 29745 48025 29779 48059
rect 29779 48025 29788 48059
rect 29736 48016 29788 48025
rect 29828 48016 29880 48068
rect 31760 48016 31812 48068
rect 32036 48059 32088 48068
rect 32036 48025 32045 48059
rect 32045 48025 32079 48059
rect 32079 48025 32088 48059
rect 32036 48016 32088 48025
rect 36544 48016 36596 48068
rect 35900 47948 35952 48000
rect 36452 47948 36504 48000
rect 44088 48093 44097 48127
rect 44097 48093 44131 48127
rect 44131 48093 44140 48127
rect 44088 48084 44140 48093
rect 45652 48127 45704 48136
rect 41788 48016 41840 48068
rect 45652 48093 45661 48127
rect 45661 48093 45695 48127
rect 45695 48093 45704 48127
rect 45652 48084 45704 48093
rect 47676 48016 47728 48068
rect 44180 47948 44232 48000
rect 44364 47948 44416 48000
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 1584 47744 1636 47796
rect 4160 47787 4212 47796
rect 4160 47753 4169 47787
rect 4169 47753 4203 47787
rect 4203 47753 4212 47787
rect 4160 47744 4212 47753
rect 5448 47744 5500 47796
rect 10232 47787 10284 47796
rect 2596 47719 2648 47728
rect 2596 47685 2605 47719
rect 2605 47685 2639 47719
rect 2639 47685 2648 47719
rect 2596 47676 2648 47685
rect 2688 47676 2740 47728
rect 1860 47651 1912 47660
rect 1860 47617 1869 47651
rect 1869 47617 1903 47651
rect 1903 47617 1912 47651
rect 1860 47608 1912 47617
rect 2504 47651 2556 47660
rect 2504 47617 2513 47651
rect 2513 47617 2547 47651
rect 2547 47617 2556 47651
rect 2504 47608 2556 47617
rect 3148 47651 3200 47660
rect 3148 47617 3157 47651
rect 3157 47617 3191 47651
rect 3191 47617 3200 47651
rect 3148 47608 3200 47617
rect 4068 47651 4120 47660
rect 4068 47617 4077 47651
rect 4077 47617 4111 47651
rect 4111 47617 4120 47651
rect 4068 47608 4120 47617
rect 6644 47676 6696 47728
rect 7380 47651 7432 47660
rect 2412 47472 2464 47524
rect 4804 47472 4856 47524
rect 7380 47617 7389 47651
rect 7389 47617 7423 47651
rect 7423 47617 7432 47651
rect 7380 47608 7432 47617
rect 6828 47540 6880 47592
rect 7840 47583 7892 47592
rect 7840 47549 7849 47583
rect 7849 47549 7883 47583
rect 7883 47549 7892 47583
rect 7840 47540 7892 47549
rect 9956 47472 10008 47524
rect 10232 47753 10241 47787
rect 10241 47753 10275 47787
rect 10275 47753 10284 47787
rect 10232 47744 10284 47753
rect 10876 47787 10928 47796
rect 10876 47753 10885 47787
rect 10885 47753 10919 47787
rect 10919 47753 10928 47787
rect 10876 47744 10928 47753
rect 12532 47744 12584 47796
rect 14372 47787 14424 47796
rect 14372 47753 14381 47787
rect 14381 47753 14415 47787
rect 14415 47753 14424 47787
rect 14372 47744 14424 47753
rect 14924 47744 14976 47796
rect 18512 47744 18564 47796
rect 19432 47744 19484 47796
rect 22008 47744 22060 47796
rect 22744 47744 22796 47796
rect 24216 47787 24268 47796
rect 24216 47753 24225 47787
rect 24225 47753 24259 47787
rect 24259 47753 24268 47787
rect 24216 47744 24268 47753
rect 24308 47744 24360 47796
rect 26148 47744 26200 47796
rect 27160 47744 27212 47796
rect 27620 47744 27672 47796
rect 28080 47744 28132 47796
rect 30380 47744 30432 47796
rect 30564 47787 30616 47796
rect 30564 47753 30573 47787
rect 30573 47753 30607 47787
rect 30607 47753 30616 47787
rect 30564 47744 30616 47753
rect 32036 47744 32088 47796
rect 32312 47744 32364 47796
rect 35992 47744 36044 47796
rect 36544 47787 36596 47796
rect 36544 47753 36553 47787
rect 36553 47753 36587 47787
rect 36587 47753 36596 47787
rect 36544 47744 36596 47753
rect 41788 47787 41840 47796
rect 41788 47753 41797 47787
rect 41797 47753 41831 47787
rect 41831 47753 41840 47787
rect 41788 47744 41840 47753
rect 13176 47676 13228 47728
rect 19984 47676 20036 47728
rect 10784 47651 10836 47660
rect 10784 47617 10793 47651
rect 10793 47617 10827 47651
rect 10827 47617 10836 47651
rect 10784 47608 10836 47617
rect 10968 47608 11020 47660
rect 13268 47651 13320 47660
rect 10508 47540 10560 47592
rect 12348 47583 12400 47592
rect 12348 47549 12357 47583
rect 12357 47549 12391 47583
rect 12391 47549 12400 47583
rect 12348 47540 12400 47549
rect 13268 47617 13277 47651
rect 13277 47617 13311 47651
rect 13311 47617 13320 47651
rect 13268 47608 13320 47617
rect 14464 47608 14516 47660
rect 15844 47608 15896 47660
rect 18052 47608 18104 47660
rect 22836 47651 22888 47660
rect 22836 47617 22845 47651
rect 22845 47617 22879 47651
rect 22879 47617 22888 47651
rect 22836 47608 22888 47617
rect 23664 47608 23716 47660
rect 24676 47608 24728 47660
rect 24952 47651 25004 47660
rect 24952 47617 24961 47651
rect 24961 47617 24995 47651
rect 24995 47617 25004 47651
rect 24952 47608 25004 47617
rect 26056 47608 26108 47660
rect 27252 47651 27304 47660
rect 23112 47540 23164 47592
rect 25872 47540 25924 47592
rect 25964 47540 26016 47592
rect 27252 47617 27261 47651
rect 27261 47617 27295 47651
rect 27295 47617 27304 47651
rect 27252 47608 27304 47617
rect 28172 47651 28224 47660
rect 28172 47617 28181 47651
rect 28181 47617 28215 47651
rect 28215 47617 28224 47651
rect 28172 47608 28224 47617
rect 31116 47651 31168 47660
rect 27988 47540 28040 47592
rect 28540 47540 28592 47592
rect 4988 47447 5040 47456
rect 4988 47413 4997 47447
rect 4997 47413 5031 47447
rect 5031 47413 5040 47447
rect 4988 47404 5040 47413
rect 6184 47404 6236 47456
rect 22100 47404 22152 47456
rect 25964 47404 26016 47456
rect 26148 47404 26200 47456
rect 27252 47404 27304 47456
rect 31116 47617 31125 47651
rect 31125 47617 31159 47651
rect 31159 47617 31168 47651
rect 31116 47608 31168 47617
rect 32128 47651 32180 47660
rect 32128 47617 32137 47651
rect 32137 47617 32171 47651
rect 32171 47617 32180 47651
rect 32128 47608 32180 47617
rect 33508 47651 33560 47660
rect 33508 47617 33517 47651
rect 33517 47617 33551 47651
rect 33551 47617 33560 47651
rect 33508 47608 33560 47617
rect 35808 47651 35860 47660
rect 35808 47617 35817 47651
rect 35817 47617 35851 47651
rect 35851 47617 35860 47651
rect 35808 47608 35860 47617
rect 36452 47651 36504 47660
rect 36452 47617 36461 47651
rect 36461 47617 36495 47651
rect 36495 47617 36504 47651
rect 36452 47608 36504 47617
rect 41696 47651 41748 47660
rect 41696 47617 41705 47651
rect 41705 47617 41739 47651
rect 41739 47617 41748 47651
rect 41696 47608 41748 47617
rect 45468 47744 45520 47796
rect 44364 47676 44416 47728
rect 31760 47540 31812 47592
rect 32496 47540 32548 47592
rect 34704 47583 34756 47592
rect 34704 47549 34713 47583
rect 34713 47549 34747 47583
rect 34747 47549 34756 47583
rect 34704 47540 34756 47549
rect 43996 47583 44048 47592
rect 43996 47549 44005 47583
rect 44005 47549 44039 47583
rect 44039 47549 44048 47583
rect 43996 47540 44048 47549
rect 30564 47472 30616 47524
rect 45652 47676 45704 47728
rect 47860 47651 47912 47660
rect 47860 47617 47869 47651
rect 47869 47617 47903 47651
rect 47903 47617 47912 47651
rect 47860 47608 47912 47617
rect 44732 47583 44784 47592
rect 44732 47549 44741 47583
rect 44741 47549 44775 47583
rect 44775 47549 44784 47583
rect 44732 47540 44784 47549
rect 45100 47540 45152 47592
rect 45192 47583 45244 47592
rect 45192 47549 45201 47583
rect 45201 47549 45235 47583
rect 45235 47549 45244 47583
rect 45192 47540 45244 47549
rect 48044 47447 48096 47456
rect 48044 47413 48053 47447
rect 48053 47413 48087 47447
rect 48087 47413 48096 47447
rect 48044 47404 48096 47413
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 1400 47200 1452 47252
rect 3976 47243 4028 47252
rect 3976 47209 3985 47243
rect 3985 47209 4019 47243
rect 4019 47209 4028 47243
rect 3976 47200 4028 47209
rect 18512 47200 18564 47252
rect 24308 47200 24360 47252
rect 25412 47243 25464 47252
rect 25412 47209 25421 47243
rect 25421 47209 25455 47243
rect 25455 47209 25464 47243
rect 25412 47200 25464 47209
rect 26056 47243 26108 47252
rect 26056 47209 26065 47243
rect 26065 47209 26099 47243
rect 26099 47209 26108 47243
rect 26056 47200 26108 47209
rect 26976 47200 27028 47252
rect 27896 47243 27948 47252
rect 27896 47209 27905 47243
rect 27905 47209 27939 47243
rect 27939 47209 27948 47243
rect 27896 47200 27948 47209
rect 27988 47200 28040 47252
rect 12348 47132 12400 47184
rect 29736 47200 29788 47252
rect 31852 47200 31904 47252
rect 45100 47243 45152 47252
rect 45100 47209 45109 47243
rect 45109 47209 45143 47243
rect 45143 47209 45152 47243
rect 45100 47200 45152 47209
rect 45744 47243 45796 47252
rect 45744 47209 45753 47243
rect 45753 47209 45787 47243
rect 45787 47209 45796 47243
rect 45744 47200 45796 47209
rect 4804 47107 4856 47116
rect 4804 47073 4813 47107
rect 4813 47073 4847 47107
rect 4847 47073 4856 47107
rect 4804 47064 4856 47073
rect 4988 47107 5040 47116
rect 4988 47073 4997 47107
rect 4997 47073 5031 47107
rect 5031 47073 5040 47107
rect 4988 47064 5040 47073
rect 5540 47107 5592 47116
rect 5540 47073 5549 47107
rect 5549 47073 5583 47107
rect 5583 47073 5592 47107
rect 5540 47064 5592 47073
rect 2228 47039 2280 47048
rect 2228 47005 2237 47039
rect 2237 47005 2271 47039
rect 2271 47005 2280 47039
rect 2228 46996 2280 47005
rect 2688 46996 2740 47048
rect 2872 46996 2924 47048
rect 6184 46996 6236 47048
rect 10508 47039 10560 47048
rect 1584 46860 1636 46912
rect 10508 47005 10517 47039
rect 10517 47005 10551 47039
rect 10551 47005 10560 47039
rect 10508 46996 10560 47005
rect 10784 47064 10836 47116
rect 35808 47132 35860 47184
rect 45652 47132 45704 47184
rect 24952 46996 25004 47048
rect 25596 47039 25648 47048
rect 25596 47005 25605 47039
rect 25605 47005 25639 47039
rect 25639 47005 25648 47039
rect 25596 46996 25648 47005
rect 26240 47039 26292 47048
rect 26240 47005 26249 47039
rect 26249 47005 26283 47039
rect 26283 47005 26292 47039
rect 26240 46996 26292 47005
rect 10968 46928 11020 46980
rect 12256 46928 12308 46980
rect 28540 47107 28592 47116
rect 28540 47073 28549 47107
rect 28549 47073 28583 47107
rect 28583 47073 28592 47107
rect 28540 47064 28592 47073
rect 43168 47064 43220 47116
rect 49608 47132 49660 47184
rect 46664 47064 46716 47116
rect 45192 46996 45244 47048
rect 45652 47039 45704 47048
rect 45652 47005 45661 47039
rect 45661 47005 45695 47039
rect 45695 47005 45704 47039
rect 45652 46996 45704 47005
rect 32128 46928 32180 46980
rect 42800 46971 42852 46980
rect 42800 46937 42809 46971
rect 42809 46937 42843 46971
rect 42843 46937 42852 46971
rect 42800 46928 42852 46937
rect 44272 46928 44324 46980
rect 46480 46971 46532 46980
rect 46480 46937 46489 46971
rect 46489 46937 46523 46971
rect 46523 46937 46532 46971
rect 46480 46928 46532 46937
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 10968 46656 11020 46708
rect 13176 46699 13228 46708
rect 2872 46588 2924 46640
rect 13176 46665 13185 46699
rect 13185 46665 13219 46699
rect 13219 46665 13228 46699
rect 13176 46656 13228 46665
rect 9956 46520 10008 46572
rect 15936 46520 15988 46572
rect 1952 46495 2004 46504
rect 1952 46461 1961 46495
rect 1961 46461 1995 46495
rect 1995 46461 2004 46495
rect 1952 46452 2004 46461
rect 2780 46495 2832 46504
rect 2780 46461 2789 46495
rect 2789 46461 2823 46495
rect 2823 46461 2832 46495
rect 2780 46452 2832 46461
rect 10692 46384 10744 46436
rect 38660 46656 38712 46708
rect 47676 46699 47728 46708
rect 47676 46665 47685 46699
rect 47685 46665 47719 46699
rect 47719 46665 47728 46699
rect 47676 46656 47728 46665
rect 22836 46588 22888 46640
rect 43168 46563 43220 46572
rect 43168 46529 43177 46563
rect 43177 46529 43211 46563
rect 43211 46529 43220 46563
rect 43168 46520 43220 46529
rect 44272 46520 44324 46572
rect 44456 46520 44508 46572
rect 1400 46316 1452 46368
rect 38476 46452 38528 46504
rect 38660 46495 38712 46504
rect 38660 46461 38669 46495
rect 38669 46461 38703 46495
rect 38703 46461 38712 46495
rect 38660 46452 38712 46461
rect 45100 46452 45152 46504
rect 45376 46495 45428 46504
rect 45376 46461 45385 46495
rect 45385 46461 45419 46495
rect 45419 46461 45428 46495
rect 45376 46452 45428 46461
rect 46848 46495 46900 46504
rect 46848 46461 46857 46495
rect 46857 46461 46891 46495
rect 46891 46461 46900 46495
rect 46848 46452 46900 46461
rect 38660 46316 38712 46368
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 38476 46155 38528 46164
rect 38476 46121 38485 46155
rect 38485 46121 38519 46155
rect 38519 46121 38528 46155
rect 38476 46112 38528 46121
rect 44732 46112 44784 46164
rect 45376 46112 45428 46164
rect 1400 46019 1452 46028
rect 1400 45985 1409 46019
rect 1409 45985 1443 46019
rect 1443 45985 1452 46019
rect 1400 45976 1452 45985
rect 1584 46019 1636 46028
rect 1584 45985 1593 46019
rect 1593 45985 1627 46019
rect 1627 45985 1636 46019
rect 1584 45976 1636 45985
rect 2780 46019 2832 46028
rect 2780 45985 2789 46019
rect 2789 45985 2823 46019
rect 2823 45985 2832 46019
rect 2780 45976 2832 45985
rect 48136 46019 48188 46028
rect 48136 45985 48145 46019
rect 48145 45985 48179 46019
rect 48179 45985 48188 46019
rect 48136 45976 48188 45985
rect 10968 45908 11020 45960
rect 41696 45908 41748 45960
rect 45192 45951 45244 45960
rect 45192 45917 45201 45951
rect 45201 45917 45235 45951
rect 45235 45917 45244 45951
rect 45192 45908 45244 45917
rect 46296 45951 46348 45960
rect 46296 45917 46305 45951
rect 46305 45917 46339 45951
rect 46339 45917 46348 45951
rect 46296 45908 46348 45917
rect 7472 45840 7524 45892
rect 22100 45840 22152 45892
rect 47032 45840 47084 45892
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 22100 45568 22152 45620
rect 22836 45568 22888 45620
rect 47032 45500 47084 45552
rect 1400 45475 1452 45484
rect 1400 45441 1409 45475
rect 1409 45441 1443 45475
rect 1443 45441 1452 45475
rect 1400 45432 1452 45441
rect 2228 45475 2280 45484
rect 2228 45441 2237 45475
rect 2237 45441 2271 45475
rect 2271 45441 2280 45475
rect 2228 45432 2280 45441
rect 12992 45432 13044 45484
rect 47768 45432 47820 45484
rect 2412 45364 2464 45416
rect 2596 45364 2648 45416
rect 45100 45407 45152 45416
rect 45100 45373 45109 45407
rect 45109 45373 45143 45407
rect 45143 45373 45152 45407
rect 45100 45364 45152 45373
rect 45284 45364 45336 45416
rect 46296 45364 46348 45416
rect 46480 45364 46532 45416
rect 2412 45271 2464 45280
rect 2412 45237 2421 45271
rect 2421 45237 2455 45271
rect 2455 45237 2464 45271
rect 2412 45228 2464 45237
rect 19432 45228 19484 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 1952 45024 2004 45076
rect 45468 45024 45520 45076
rect 32128 44888 32180 44940
rect 37280 44888 37332 44940
rect 48136 44931 48188 44940
rect 48136 44897 48145 44931
rect 48145 44897 48179 44931
rect 48179 44897 48188 44931
rect 48136 44888 48188 44897
rect 1400 44863 1452 44872
rect 1400 44829 1409 44863
rect 1409 44829 1443 44863
rect 1443 44829 1452 44863
rect 1400 44820 1452 44829
rect 2228 44820 2280 44872
rect 2044 44752 2096 44804
rect 16764 44820 16816 44872
rect 46296 44863 46348 44872
rect 46296 44829 46305 44863
rect 46305 44829 46339 44863
rect 46339 44829 46348 44863
rect 46296 44820 46348 44829
rect 1676 44684 1728 44736
rect 47676 44752 47728 44804
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 47676 44523 47728 44532
rect 47676 44489 47685 44523
rect 47685 44489 47719 44523
rect 47719 44489 47728 44523
rect 47676 44480 47728 44489
rect 2044 44387 2096 44396
rect 2044 44353 2053 44387
rect 2053 44353 2087 44387
rect 2087 44353 2096 44387
rect 2044 44344 2096 44353
rect 46296 44344 46348 44396
rect 47584 44387 47636 44396
rect 47584 44353 47593 44387
rect 47593 44353 47627 44387
rect 47627 44353 47636 44387
rect 47584 44344 47636 44353
rect 2964 44276 3016 44328
rect 3056 44319 3108 44328
rect 3056 44285 3065 44319
rect 3065 44285 3099 44319
rect 3099 44285 3108 44319
rect 3056 44276 3108 44285
rect 17224 44140 17276 44192
rect 26148 44140 26200 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 2964 43979 3016 43988
rect 2964 43945 2973 43979
rect 2973 43945 3007 43979
rect 3007 43945 3016 43979
rect 2964 43936 3016 43945
rect 1400 43775 1452 43784
rect 1400 43741 1409 43775
rect 1409 43741 1443 43775
rect 1443 43741 1452 43775
rect 1400 43732 1452 43741
rect 3332 43732 3384 43784
rect 36084 43732 36136 43784
rect 47308 43775 47360 43784
rect 47308 43741 47317 43775
rect 47317 43741 47351 43775
rect 47351 43741 47360 43775
rect 47308 43732 47360 43741
rect 47492 43732 47544 43784
rect 1768 43664 1820 43716
rect 36544 43707 36596 43716
rect 36544 43673 36553 43707
rect 36553 43673 36587 43707
rect 36587 43673 36596 43707
rect 36544 43664 36596 43673
rect 46848 43664 46900 43716
rect 47400 43639 47452 43648
rect 47400 43605 47409 43639
rect 47409 43605 47443 43639
rect 47443 43605 47452 43639
rect 47400 43596 47452 43605
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 36544 43435 36596 43444
rect 36544 43401 36553 43435
rect 36553 43401 36587 43435
rect 36587 43401 36596 43435
rect 36544 43392 36596 43401
rect 36452 43299 36504 43308
rect 36452 43265 36461 43299
rect 36461 43265 36495 43299
rect 36495 43265 36504 43299
rect 36452 43256 36504 43265
rect 47860 43299 47912 43308
rect 47860 43265 47869 43299
rect 47869 43265 47903 43299
rect 47903 43265 47912 43299
rect 47860 43256 47912 43265
rect 47676 43052 47728 43104
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 47400 42712 47452 42764
rect 48136 42755 48188 42764
rect 48136 42721 48145 42755
rect 48145 42721 48179 42755
rect 48179 42721 48188 42755
rect 48136 42712 48188 42721
rect 47492 42576 47544 42628
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 47952 42211 48004 42220
rect 47952 42177 47961 42211
rect 47961 42177 47995 42211
rect 47995 42177 48004 42211
rect 47952 42168 48004 42177
rect 28448 42032 28500 42084
rect 1400 41964 1452 42016
rect 46296 41964 46348 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 1400 41667 1452 41676
rect 1400 41633 1409 41667
rect 1409 41633 1443 41667
rect 1443 41633 1452 41667
rect 1400 41624 1452 41633
rect 1860 41667 1912 41676
rect 1860 41633 1869 41667
rect 1869 41633 1903 41667
rect 1903 41633 1912 41667
rect 1860 41624 1912 41633
rect 46296 41667 46348 41676
rect 46296 41633 46305 41667
rect 46305 41633 46339 41667
rect 46339 41633 46348 41667
rect 46296 41624 46348 41633
rect 1584 41531 1636 41540
rect 1584 41497 1593 41531
rect 1593 41497 1627 41531
rect 1627 41497 1636 41531
rect 1584 41488 1636 41497
rect 46480 41531 46532 41540
rect 46480 41497 46489 41531
rect 46489 41497 46523 41531
rect 46523 41497 46532 41531
rect 46480 41488 46532 41497
rect 48136 41531 48188 41540
rect 48136 41497 48145 41531
rect 48145 41497 48179 41531
rect 48179 41497 48188 41531
rect 48136 41488 48188 41497
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 1584 41216 1636 41268
rect 46480 41216 46532 41268
rect 1400 41123 1452 41132
rect 1400 41089 1409 41123
rect 1409 41089 1443 41123
rect 1443 41089 1452 41123
rect 1400 41080 1452 41089
rect 2320 41080 2372 41132
rect 41696 41080 41748 41132
rect 46664 41080 46716 41132
rect 47860 41123 47912 41132
rect 47860 41089 47869 41123
rect 47869 41089 47903 41123
rect 47903 41089 47912 41123
rect 47860 41080 47912 41089
rect 1952 40876 2004 40928
rect 48228 40876 48280 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 47032 40536 47084 40588
rect 1860 40443 1912 40452
rect 1860 40409 1869 40443
rect 1869 40409 1903 40443
rect 1903 40409 1912 40443
rect 1860 40400 1912 40409
rect 3700 40400 3752 40452
rect 47676 40400 47728 40452
rect 48136 40443 48188 40452
rect 48136 40409 48145 40443
rect 48145 40409 48179 40443
rect 48179 40409 48188 40443
rect 48136 40400 48188 40409
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 47032 40035 47084 40044
rect 47032 40001 47041 40035
rect 47041 40001 47075 40035
rect 47075 40001 47084 40035
rect 47032 39992 47084 40001
rect 45652 39924 45704 39976
rect 47676 40035 47728 40044
rect 47676 40001 47685 40035
rect 47685 40001 47719 40035
rect 47719 40001 47728 40035
rect 47676 39992 47728 40001
rect 1400 39788 1452 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 1400 39491 1452 39500
rect 1400 39457 1409 39491
rect 1409 39457 1443 39491
rect 1443 39457 1452 39491
rect 1400 39448 1452 39457
rect 2780 39491 2832 39500
rect 2780 39457 2789 39491
rect 2789 39457 2823 39491
rect 2823 39457 2832 39491
rect 2780 39448 2832 39457
rect 24400 39448 24452 39500
rect 6644 39380 6696 39432
rect 7472 39423 7524 39432
rect 7472 39389 7481 39423
rect 7481 39389 7515 39423
rect 7515 39389 7524 39423
rect 7472 39380 7524 39389
rect 24492 39380 24544 39432
rect 2136 39312 2188 39364
rect 24952 39380 25004 39432
rect 46848 39380 46900 39432
rect 26332 39312 26384 39364
rect 32220 39312 32272 39364
rect 6828 39244 6880 39296
rect 24492 39244 24544 39296
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 2136 39083 2188 39092
rect 2136 39049 2145 39083
rect 2145 39049 2179 39083
rect 2179 39049 2188 39083
rect 2136 39040 2188 39049
rect 6828 39015 6880 39024
rect 6828 38981 6837 39015
rect 6837 38981 6871 39015
rect 6871 38981 6880 39015
rect 6828 38972 6880 38981
rect 20536 38972 20588 39024
rect 1400 38904 1452 38956
rect 6644 38947 6696 38956
rect 6644 38913 6653 38947
rect 6653 38913 6687 38947
rect 6687 38913 6696 38947
rect 6644 38904 6696 38913
rect 20904 38947 20956 38956
rect 20904 38913 20913 38947
rect 20913 38913 20947 38947
rect 20947 38913 20956 38947
rect 20904 38904 20956 38913
rect 24032 38904 24084 38956
rect 5540 38836 5592 38888
rect 23940 38879 23992 38888
rect 23940 38845 23949 38879
rect 23949 38845 23983 38879
rect 23983 38845 23992 38879
rect 23940 38836 23992 38845
rect 21088 38700 21140 38752
rect 25044 38700 25096 38752
rect 47768 38743 47820 38752
rect 47768 38709 47777 38743
rect 47777 38709 47811 38743
rect 47811 38709 47820 38743
rect 47768 38700 47820 38709
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 20812 38428 20864 38480
rect 5632 38360 5684 38412
rect 21456 38360 21508 38412
rect 47768 38360 47820 38412
rect 48136 38403 48188 38412
rect 48136 38369 48145 38403
rect 48145 38369 48179 38403
rect 48179 38369 48188 38403
rect 48136 38360 48188 38369
rect 21272 38292 21324 38344
rect 21548 38335 21600 38344
rect 21548 38301 21557 38335
rect 21557 38301 21591 38335
rect 21591 38301 21600 38335
rect 21548 38292 21600 38301
rect 23940 38292 23992 38344
rect 22744 38156 22796 38208
rect 24492 38292 24544 38344
rect 26700 38224 26752 38276
rect 46940 38224 46992 38276
rect 24768 38156 24820 38208
rect 25780 38199 25832 38208
rect 25780 38165 25789 38199
rect 25789 38165 25823 38199
rect 25823 38165 25832 38199
rect 25780 38156 25832 38165
rect 27988 38156 28040 38208
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 20904 37952 20956 38004
rect 24032 37995 24084 38004
rect 24032 37961 24041 37995
rect 24041 37961 24075 37995
rect 24075 37961 24084 37995
rect 24032 37952 24084 37961
rect 24400 37952 24452 38004
rect 26332 37995 26384 38004
rect 26332 37961 26341 37995
rect 26341 37961 26375 37995
rect 26375 37961 26384 37995
rect 26332 37952 26384 37961
rect 19340 37859 19392 37868
rect 19340 37825 19349 37859
rect 19349 37825 19383 37859
rect 19383 37825 19392 37859
rect 19340 37816 19392 37825
rect 20536 37816 20588 37868
rect 1400 37791 1452 37800
rect 1400 37757 1409 37791
rect 1409 37757 1443 37791
rect 1443 37757 1452 37791
rect 1400 37748 1452 37757
rect 19800 37748 19852 37800
rect 20812 37748 20864 37800
rect 21088 37859 21140 37868
rect 21088 37825 21097 37859
rect 21097 37825 21131 37859
rect 21131 37825 21140 37859
rect 21088 37816 21140 37825
rect 21272 37859 21324 37868
rect 21272 37825 21281 37859
rect 21281 37825 21315 37859
rect 21315 37825 21324 37859
rect 21272 37816 21324 37825
rect 22376 37816 22428 37868
rect 17776 37680 17828 37732
rect 20996 37680 21048 37732
rect 22468 37791 22520 37800
rect 22468 37757 22477 37791
rect 22477 37757 22511 37791
rect 22511 37757 22520 37791
rect 22468 37748 22520 37757
rect 24308 37859 24360 37868
rect 24308 37825 24317 37859
rect 24317 37825 24351 37859
rect 24351 37825 24360 37859
rect 24308 37816 24360 37825
rect 24952 37816 25004 37868
rect 25136 37859 25188 37868
rect 25136 37825 25145 37859
rect 25145 37825 25179 37859
rect 25179 37825 25188 37859
rect 25136 37816 25188 37825
rect 25964 37859 26016 37868
rect 24124 37680 24176 37732
rect 25964 37825 25973 37859
rect 25973 37825 26007 37859
rect 26007 37825 26016 37859
rect 25964 37816 26016 37825
rect 26056 37748 26108 37800
rect 40868 37952 40920 38004
rect 46940 37995 46992 38004
rect 46940 37961 46949 37995
rect 46949 37961 46983 37995
rect 46983 37961 46992 37995
rect 46940 37952 46992 37961
rect 29552 37884 29604 37936
rect 29920 37927 29972 37936
rect 29920 37893 29929 37927
rect 29929 37893 29963 37927
rect 29963 37893 29972 37927
rect 29920 37884 29972 37893
rect 31116 37884 31168 37936
rect 47952 37927 48004 37936
rect 47952 37893 47961 37927
rect 47961 37893 47995 37927
rect 47995 37893 48004 37927
rect 47952 37884 48004 37893
rect 27804 37859 27856 37868
rect 27804 37825 27838 37859
rect 27838 37825 27856 37859
rect 27804 37816 27856 37825
rect 46572 37816 46624 37868
rect 47032 37748 47084 37800
rect 47216 37748 47268 37800
rect 19708 37655 19760 37664
rect 19708 37621 19717 37655
rect 19717 37621 19751 37655
rect 19751 37621 19760 37655
rect 19708 37612 19760 37621
rect 20904 37612 20956 37664
rect 28172 37612 28224 37664
rect 30104 37655 30156 37664
rect 30104 37621 30113 37655
rect 30113 37621 30147 37655
rect 30147 37621 30156 37655
rect 30104 37612 30156 37621
rect 30288 37655 30340 37664
rect 30288 37621 30297 37655
rect 30297 37621 30331 37655
rect 30331 37621 30340 37655
rect 30288 37612 30340 37621
rect 47400 37612 47452 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 19340 37408 19392 37460
rect 20076 37408 20128 37460
rect 20352 37408 20404 37460
rect 20076 37272 20128 37324
rect 17776 37204 17828 37256
rect 1860 37179 1912 37188
rect 1860 37145 1869 37179
rect 1869 37145 1903 37179
rect 1903 37145 1912 37179
rect 1860 37136 1912 37145
rect 2044 37179 2096 37188
rect 2044 37145 2053 37179
rect 2053 37145 2087 37179
rect 2087 37145 2096 37179
rect 2044 37136 2096 37145
rect 18144 37068 18196 37120
rect 19708 37136 19760 37188
rect 19800 37136 19852 37188
rect 20628 37204 20680 37256
rect 21548 37408 21600 37460
rect 25964 37408 26016 37460
rect 26700 37451 26752 37460
rect 26700 37417 26709 37451
rect 26709 37417 26743 37451
rect 26743 37417 26752 37451
rect 26700 37408 26752 37417
rect 30196 37408 30248 37460
rect 47216 37408 47268 37460
rect 47676 37408 47728 37460
rect 24124 37340 24176 37392
rect 27988 37340 28040 37392
rect 25504 37315 25556 37324
rect 25504 37281 25513 37315
rect 25513 37281 25547 37315
rect 25547 37281 25556 37315
rect 25504 37272 25556 37281
rect 20904 37204 20956 37256
rect 26516 37204 26568 37256
rect 27252 37272 27304 37324
rect 28356 37315 28408 37324
rect 28356 37281 28365 37315
rect 28365 37281 28399 37315
rect 28399 37281 28408 37315
rect 28356 37272 28408 37281
rect 34612 37272 34664 37324
rect 46848 37272 46900 37324
rect 20996 37136 21048 37188
rect 19340 37068 19392 37120
rect 19984 37111 20036 37120
rect 19984 37077 19993 37111
rect 19993 37077 20027 37111
rect 20027 37077 20036 37111
rect 19984 37068 20036 37077
rect 25780 37136 25832 37188
rect 27344 37247 27396 37256
rect 27344 37213 27353 37247
rect 27353 37213 27387 37247
rect 27387 37213 27396 37247
rect 27344 37204 27396 37213
rect 27712 37204 27764 37256
rect 29552 37247 29604 37256
rect 29552 37213 29561 37247
rect 29561 37213 29595 37247
rect 29595 37213 29604 37247
rect 29552 37204 29604 37213
rect 47676 37247 47728 37256
rect 47676 37213 47685 37247
rect 47685 37213 47719 37247
rect 47719 37213 47728 37247
rect 47676 37204 47728 37213
rect 29184 37136 29236 37188
rect 29828 37179 29880 37188
rect 29828 37145 29862 37179
rect 29862 37145 29880 37179
rect 29828 37136 29880 37145
rect 31116 37136 31168 37188
rect 32220 37179 32272 37188
rect 22376 37068 22428 37120
rect 23296 37068 23348 37120
rect 26700 37068 26752 37120
rect 26792 37068 26844 37120
rect 28080 37068 28132 37120
rect 30104 37068 30156 37120
rect 32220 37145 32229 37179
rect 32229 37145 32263 37179
rect 32263 37145 32272 37179
rect 32220 37136 32272 37145
rect 32588 37111 32640 37120
rect 32588 37077 32597 37111
rect 32597 37077 32631 37111
rect 32631 37077 32640 37111
rect 32588 37068 32640 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 21456 36864 21508 36916
rect 25136 36864 25188 36916
rect 25228 36864 25280 36916
rect 27344 36864 27396 36916
rect 29184 36907 29236 36916
rect 2044 36796 2096 36848
rect 24584 36796 24636 36848
rect 25044 36839 25096 36848
rect 25044 36805 25053 36839
rect 25053 36805 25087 36839
rect 25087 36805 25096 36839
rect 25044 36796 25096 36805
rect 26792 36796 26844 36848
rect 29184 36873 29193 36907
rect 29193 36873 29227 36907
rect 29227 36873 29236 36907
rect 29184 36864 29236 36873
rect 18144 36728 18196 36780
rect 18052 36703 18104 36712
rect 18052 36669 18061 36703
rect 18061 36669 18095 36703
rect 18095 36669 18104 36703
rect 18052 36660 18104 36669
rect 20536 36728 20588 36780
rect 21824 36771 21876 36780
rect 21824 36737 21833 36771
rect 21833 36737 21867 36771
rect 21867 36737 21876 36771
rect 21824 36728 21876 36737
rect 21916 36728 21968 36780
rect 26240 36771 26292 36780
rect 21272 36660 21324 36712
rect 25504 36660 25556 36712
rect 26240 36737 26249 36771
rect 26249 36737 26283 36771
rect 26283 36737 26292 36771
rect 27988 36771 28040 36780
rect 26240 36728 26292 36737
rect 27988 36737 27997 36771
rect 27997 36737 28031 36771
rect 28031 36737 28040 36771
rect 27988 36728 28040 36737
rect 28264 36728 28316 36780
rect 27896 36660 27948 36712
rect 27620 36592 27672 36644
rect 28356 36660 28408 36712
rect 29552 36728 29604 36780
rect 30012 36771 30064 36780
rect 30012 36737 30046 36771
rect 30046 36737 30064 36771
rect 30012 36728 30064 36737
rect 31944 36728 31996 36780
rect 47584 36771 47636 36780
rect 47584 36737 47593 36771
rect 47593 36737 47627 36771
rect 47627 36737 47636 36771
rect 47584 36728 47636 36737
rect 32128 36703 32180 36712
rect 32128 36669 32137 36703
rect 32137 36669 32171 36703
rect 32171 36669 32180 36703
rect 32128 36660 32180 36669
rect 1952 36524 2004 36576
rect 19984 36524 20036 36576
rect 20812 36567 20864 36576
rect 20812 36533 20821 36567
rect 20821 36533 20855 36567
rect 20855 36533 20864 36567
rect 20812 36524 20864 36533
rect 24952 36524 25004 36576
rect 25228 36524 25280 36576
rect 28356 36524 28408 36576
rect 30380 36524 30432 36576
rect 33508 36567 33560 36576
rect 33508 36533 33517 36567
rect 33517 36533 33551 36567
rect 33551 36533 33560 36567
rect 33508 36524 33560 36533
rect 46480 36524 46532 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 21824 36320 21876 36372
rect 24584 36320 24636 36372
rect 27804 36320 27856 36372
rect 29828 36363 29880 36372
rect 29828 36329 29837 36363
rect 29837 36329 29871 36363
rect 29871 36329 29880 36363
rect 29828 36320 29880 36329
rect 30196 36320 30248 36372
rect 31944 36363 31996 36372
rect 31944 36329 31953 36363
rect 31953 36329 31987 36363
rect 31987 36329 31996 36363
rect 31944 36320 31996 36329
rect 2596 36184 2648 36236
rect 3424 36116 3476 36168
rect 20628 36227 20680 36236
rect 20628 36193 20637 36227
rect 20637 36193 20671 36227
rect 20671 36193 20680 36227
rect 20628 36184 20680 36193
rect 22468 36184 22520 36236
rect 22652 36184 22704 36236
rect 24768 36227 24820 36236
rect 24768 36193 24777 36227
rect 24777 36193 24811 36227
rect 24811 36193 24820 36227
rect 24768 36184 24820 36193
rect 24400 36116 24452 36168
rect 27252 36184 27304 36236
rect 30104 36227 30156 36236
rect 26608 36159 26660 36168
rect 26608 36125 26617 36159
rect 26617 36125 26651 36159
rect 26651 36125 26660 36159
rect 26608 36116 26660 36125
rect 27896 36116 27948 36168
rect 30104 36193 30113 36227
rect 30113 36193 30147 36227
rect 30147 36193 30156 36227
rect 30104 36184 30156 36193
rect 30288 36227 30340 36236
rect 30288 36193 30297 36227
rect 30297 36193 30331 36227
rect 30331 36193 30340 36227
rect 30288 36184 30340 36193
rect 28356 36159 28408 36168
rect 28356 36125 28365 36159
rect 28365 36125 28399 36159
rect 28399 36125 28408 36159
rect 28356 36116 28408 36125
rect 28540 36159 28592 36168
rect 28540 36125 28549 36159
rect 28549 36125 28583 36159
rect 28583 36125 28592 36159
rect 28540 36116 28592 36125
rect 29920 36116 29972 36168
rect 30564 36116 30616 36168
rect 19156 36048 19208 36100
rect 19340 36048 19392 36100
rect 2872 36023 2924 36032
rect 2872 35989 2881 36023
rect 2881 35989 2915 36023
rect 2915 35989 2924 36023
rect 2872 35980 2924 35989
rect 18236 35980 18288 36032
rect 20720 36048 20772 36100
rect 20996 36048 21048 36100
rect 24860 36048 24912 36100
rect 30840 36252 30892 36304
rect 31668 36184 31720 36236
rect 32588 36184 32640 36236
rect 32036 36116 32088 36168
rect 47676 36252 47728 36304
rect 46480 36227 46532 36236
rect 46480 36193 46489 36227
rect 46489 36193 46523 36227
rect 46523 36193 46532 36227
rect 46480 36184 46532 36193
rect 48136 36227 48188 36236
rect 48136 36193 48145 36227
rect 48145 36193 48179 36227
rect 48179 36193 48188 36227
rect 48136 36184 48188 36193
rect 33508 36116 33560 36168
rect 31116 36048 31168 36100
rect 21456 35980 21508 36032
rect 21916 35980 21968 36032
rect 22468 35980 22520 36032
rect 22744 35980 22796 36032
rect 23572 35980 23624 36032
rect 25320 35980 25372 36032
rect 27344 35980 27396 36032
rect 28264 35980 28316 36032
rect 30840 35980 30892 36032
rect 31392 36023 31444 36032
rect 31392 35989 31401 36023
rect 31401 35989 31435 36023
rect 31435 35989 31444 36023
rect 31392 35980 31444 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 20720 35776 20772 35828
rect 21272 35776 21324 35828
rect 24860 35776 24912 35828
rect 25044 35776 25096 35828
rect 2872 35708 2924 35760
rect 18052 35708 18104 35760
rect 1952 35683 2004 35692
rect 1952 35649 1961 35683
rect 1961 35649 1995 35683
rect 1995 35649 2004 35683
rect 1952 35640 2004 35649
rect 19708 35708 19760 35760
rect 18236 35640 18288 35692
rect 20260 35640 20312 35692
rect 20812 35708 20864 35760
rect 27068 35776 27120 35828
rect 2780 35615 2832 35624
rect 2780 35581 2789 35615
rect 2789 35581 2823 35615
rect 2823 35581 2832 35615
rect 2780 35572 2832 35581
rect 19156 35572 19208 35624
rect 19616 35572 19668 35624
rect 20996 35640 21048 35692
rect 22468 35683 22520 35692
rect 22468 35649 22477 35683
rect 22477 35649 22511 35683
rect 22511 35649 22520 35683
rect 22468 35640 22520 35649
rect 22836 35640 22888 35692
rect 24216 35640 24268 35692
rect 24308 35640 24360 35692
rect 25228 35683 25280 35692
rect 22652 35615 22704 35624
rect 22652 35581 22661 35615
rect 22661 35581 22695 35615
rect 22695 35581 22704 35615
rect 22652 35572 22704 35581
rect 24400 35572 24452 35624
rect 25228 35649 25237 35683
rect 25237 35649 25271 35683
rect 25271 35649 25280 35683
rect 25228 35640 25280 35649
rect 26240 35683 26292 35692
rect 26240 35649 26249 35683
rect 26249 35649 26283 35683
rect 26283 35649 26292 35683
rect 26240 35640 26292 35649
rect 20076 35504 20128 35556
rect 25504 35504 25556 35556
rect 27344 35683 27396 35692
rect 27344 35649 27353 35683
rect 27353 35649 27387 35683
rect 27387 35649 27396 35683
rect 27344 35640 27396 35649
rect 27620 35708 27672 35760
rect 27712 35708 27764 35760
rect 28540 35708 28592 35760
rect 28172 35640 28224 35692
rect 29000 35683 29052 35692
rect 29000 35649 29009 35683
rect 29009 35649 29043 35683
rect 29043 35649 29052 35683
rect 29000 35640 29052 35649
rect 30012 35776 30064 35828
rect 29920 35708 29972 35760
rect 29368 35640 29420 35692
rect 32036 35708 32088 35760
rect 47952 35751 48004 35760
rect 47952 35717 47961 35751
rect 47961 35717 47995 35751
rect 47995 35717 48004 35751
rect 47952 35708 48004 35717
rect 30380 35683 30432 35692
rect 30380 35649 30389 35683
rect 30389 35649 30423 35683
rect 30423 35649 30432 35683
rect 30380 35640 30432 35649
rect 31392 35640 31444 35692
rect 32220 35640 32272 35692
rect 45652 35640 45704 35692
rect 30104 35572 30156 35624
rect 32128 35615 32180 35624
rect 32128 35581 32137 35615
rect 32137 35581 32171 35615
rect 32171 35581 32180 35615
rect 32128 35572 32180 35581
rect 19524 35479 19576 35488
rect 19524 35445 19533 35479
rect 19533 35445 19567 35479
rect 19567 35445 19576 35479
rect 19524 35436 19576 35445
rect 19708 35436 19760 35488
rect 20628 35436 20680 35488
rect 30564 35504 30616 35556
rect 45836 35504 45888 35556
rect 29460 35479 29512 35488
rect 29460 35445 29469 35479
rect 29469 35445 29503 35479
rect 29503 35445 29512 35479
rect 29460 35436 29512 35445
rect 33508 35479 33560 35488
rect 33508 35445 33517 35479
rect 33517 35445 33551 35479
rect 33551 35445 33560 35479
rect 33508 35436 33560 35445
rect 46296 35479 46348 35488
rect 46296 35445 46305 35479
rect 46305 35445 46339 35479
rect 46339 35445 46348 35479
rect 46296 35436 46348 35445
rect 46480 35436 46532 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 19340 35232 19392 35284
rect 20996 35275 21048 35284
rect 20996 35241 21005 35275
rect 21005 35241 21039 35275
rect 21039 35241 21048 35275
rect 20996 35232 21048 35241
rect 25044 35232 25096 35284
rect 25504 35275 25556 35284
rect 25504 35241 25513 35275
rect 25513 35241 25547 35275
rect 25547 35241 25556 35275
rect 25504 35232 25556 35241
rect 29460 35232 29512 35284
rect 30288 35232 30340 35284
rect 32220 35232 32272 35284
rect 1768 35164 1820 35216
rect 2596 35164 2648 35216
rect 19616 35164 19668 35216
rect 24216 35164 24268 35216
rect 20076 35139 20128 35148
rect 1768 35028 1820 35080
rect 20076 35105 20085 35139
rect 20085 35105 20119 35139
rect 20119 35105 20128 35139
rect 20076 35096 20128 35105
rect 24492 35139 24544 35148
rect 24492 35105 24501 35139
rect 24501 35105 24535 35139
rect 24535 35105 24544 35139
rect 24492 35096 24544 35105
rect 24308 35028 24360 35080
rect 24676 35071 24728 35080
rect 24676 35037 24685 35071
rect 24685 35037 24719 35071
rect 24719 35037 24728 35071
rect 24676 35028 24728 35037
rect 29368 35164 29420 35216
rect 28724 35028 28776 35080
rect 30472 35028 30524 35080
rect 1860 35003 1912 35012
rect 1860 34969 1869 35003
rect 1869 34969 1903 35003
rect 1903 34969 1912 35003
rect 1860 34960 1912 34969
rect 19524 34960 19576 35012
rect 20904 35003 20956 35012
rect 20076 34892 20128 34944
rect 20904 34969 20913 35003
rect 20913 34969 20947 35003
rect 20947 34969 20956 35003
rect 20904 34960 20956 34969
rect 22652 34960 22704 35012
rect 24124 34960 24176 35012
rect 31116 35096 31168 35148
rect 33508 35096 33560 35148
rect 46296 35139 46348 35148
rect 46296 35105 46305 35139
rect 46305 35105 46339 35139
rect 46339 35105 46348 35139
rect 46296 35096 46348 35105
rect 46480 35139 46532 35148
rect 46480 35105 46489 35139
rect 46489 35105 46523 35139
rect 46523 35105 46532 35139
rect 46480 35096 46532 35105
rect 48136 35139 48188 35148
rect 48136 35105 48145 35139
rect 48145 35105 48179 35139
rect 48179 35105 48188 35139
rect 48136 35096 48188 35105
rect 30748 35028 30800 35080
rect 31576 35028 31628 35080
rect 32036 35028 32088 35080
rect 21272 34892 21324 34944
rect 24860 34935 24912 34944
rect 24860 34901 24869 34935
rect 24869 34901 24903 34935
rect 24903 34901 24912 34935
rect 24860 34892 24912 34901
rect 25596 34892 25648 34944
rect 30840 34960 30892 35012
rect 31668 34960 31720 35012
rect 32680 35028 32732 35080
rect 31208 34892 31260 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 23572 34731 23624 34740
rect 23572 34697 23581 34731
rect 23581 34697 23615 34731
rect 23615 34697 23624 34731
rect 23572 34688 23624 34697
rect 24492 34688 24544 34740
rect 28724 34731 28776 34740
rect 28724 34697 28733 34731
rect 28733 34697 28767 34731
rect 28767 34697 28776 34731
rect 28724 34688 28776 34697
rect 31116 34688 31168 34740
rect 32036 34688 32088 34740
rect 32680 34731 32732 34740
rect 32680 34697 32689 34731
rect 32689 34697 32723 34731
rect 32723 34697 32732 34731
rect 32680 34688 32732 34697
rect 2412 34620 2464 34672
rect 1768 34595 1820 34604
rect 1768 34561 1777 34595
rect 1777 34561 1811 34595
rect 1811 34561 1820 34595
rect 1768 34552 1820 34561
rect 19432 34552 19484 34604
rect 20352 34595 20404 34604
rect 2780 34527 2832 34536
rect 2780 34493 2789 34527
rect 2789 34493 2823 34527
rect 2823 34493 2832 34527
rect 2780 34484 2832 34493
rect 20352 34561 20361 34595
rect 20361 34561 20395 34595
rect 20395 34561 20404 34595
rect 20352 34552 20404 34561
rect 20536 34595 20588 34604
rect 20536 34561 20545 34595
rect 20545 34561 20579 34595
rect 20579 34561 20588 34595
rect 24768 34620 24820 34672
rect 20536 34552 20588 34561
rect 22468 34595 22520 34604
rect 22468 34561 22502 34595
rect 22502 34561 22520 34595
rect 22468 34552 22520 34561
rect 25412 34552 25464 34604
rect 25780 34595 25832 34604
rect 25780 34561 25789 34595
rect 25789 34561 25823 34595
rect 25823 34561 25832 34595
rect 25780 34552 25832 34561
rect 20628 34484 20680 34536
rect 24584 34527 24636 34536
rect 24584 34493 24593 34527
rect 24593 34493 24627 34527
rect 24627 34493 24636 34527
rect 24584 34484 24636 34493
rect 25228 34484 25280 34536
rect 27804 34620 27856 34672
rect 28264 34595 28316 34604
rect 28264 34561 28273 34595
rect 28273 34561 28307 34595
rect 28307 34561 28316 34595
rect 28264 34552 28316 34561
rect 28632 34552 28684 34604
rect 31484 34620 31536 34672
rect 30288 34552 30340 34604
rect 30564 34552 30616 34604
rect 30840 34595 30892 34604
rect 30840 34561 30849 34595
rect 30849 34561 30883 34595
rect 30883 34561 30892 34595
rect 30840 34552 30892 34561
rect 31208 34552 31260 34604
rect 46020 34620 46072 34672
rect 46756 34595 46808 34604
rect 46756 34561 46765 34595
rect 46765 34561 46799 34595
rect 46799 34561 46808 34595
rect 46756 34552 46808 34561
rect 19340 34348 19392 34400
rect 22192 34416 22244 34468
rect 29644 34484 29696 34536
rect 30748 34527 30800 34536
rect 30748 34493 30757 34527
rect 30757 34493 30791 34527
rect 30791 34493 30800 34527
rect 30748 34484 30800 34493
rect 28080 34416 28132 34468
rect 30288 34416 30340 34468
rect 23480 34348 23532 34400
rect 24032 34391 24084 34400
rect 24032 34357 24041 34391
rect 24041 34357 24075 34391
rect 24075 34357 24084 34391
rect 24032 34348 24084 34357
rect 25320 34348 25372 34400
rect 25964 34391 26016 34400
rect 25964 34357 25973 34391
rect 25973 34357 26007 34391
rect 26007 34357 26016 34391
rect 25964 34348 26016 34357
rect 27988 34348 28040 34400
rect 30380 34348 30432 34400
rect 46480 34348 46532 34400
rect 47768 34391 47820 34400
rect 47768 34357 47777 34391
rect 47777 34357 47811 34391
rect 47811 34357 47820 34391
rect 47768 34348 47820 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 20352 34144 20404 34196
rect 22468 34144 22520 34196
rect 24584 34144 24636 34196
rect 19800 34008 19852 34060
rect 20628 34008 20680 34060
rect 25228 34076 25280 34128
rect 25412 34076 25464 34128
rect 21180 34008 21232 34060
rect 20536 33940 20588 33992
rect 24860 34008 24912 34060
rect 19800 33915 19852 33924
rect 19800 33881 19809 33915
rect 19809 33881 19843 33915
rect 19843 33881 19852 33915
rect 19800 33872 19852 33881
rect 20352 33872 20404 33924
rect 24032 33940 24084 33992
rect 24124 33940 24176 33992
rect 1768 33804 1820 33856
rect 20628 33804 20680 33856
rect 22284 33804 22336 33856
rect 22376 33804 22428 33856
rect 22560 33804 22612 33856
rect 24216 33872 24268 33924
rect 24492 33872 24544 33924
rect 25504 33940 25556 33992
rect 25964 33983 26016 33992
rect 25964 33949 25973 33983
rect 25973 33949 26007 33983
rect 26007 33949 26016 33983
rect 25964 33940 26016 33949
rect 28080 34051 28132 34060
rect 28080 34017 28089 34051
rect 28089 34017 28123 34051
rect 28123 34017 28132 34051
rect 28080 34008 28132 34017
rect 29552 34051 29604 34060
rect 29552 34017 29561 34051
rect 29561 34017 29595 34051
rect 29595 34017 29604 34051
rect 29552 34008 29604 34017
rect 32036 34051 32088 34060
rect 32036 34017 32045 34051
rect 32045 34017 32079 34051
rect 32079 34017 32088 34051
rect 32036 34008 32088 34017
rect 47768 34076 47820 34128
rect 46480 34051 46532 34060
rect 46480 34017 46489 34051
rect 46489 34017 46523 34051
rect 46523 34017 46532 34051
rect 46480 34008 46532 34017
rect 48136 34051 48188 34060
rect 48136 34017 48145 34051
rect 48145 34017 48179 34051
rect 48179 34017 48188 34051
rect 48136 34008 48188 34017
rect 23756 33804 23808 33856
rect 26056 33872 26108 33924
rect 26240 33872 26292 33924
rect 25964 33804 26016 33856
rect 27252 33804 27304 33856
rect 28356 33940 28408 33992
rect 30380 33940 30432 33992
rect 31760 33983 31812 33992
rect 31760 33949 31769 33983
rect 31769 33949 31803 33983
rect 31803 33949 31812 33983
rect 31760 33940 31812 33949
rect 29000 33804 29052 33856
rect 30840 33804 30892 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 20536 33643 20588 33652
rect 20536 33609 20545 33643
rect 20545 33609 20579 33643
rect 20579 33609 20588 33643
rect 20536 33600 20588 33609
rect 24124 33600 24176 33652
rect 24768 33600 24820 33652
rect 1768 33507 1820 33516
rect 1768 33473 1777 33507
rect 1777 33473 1811 33507
rect 1811 33473 1820 33507
rect 1768 33464 1820 33473
rect 19340 33532 19392 33584
rect 21088 33464 21140 33516
rect 21640 33464 21692 33516
rect 1952 33439 2004 33448
rect 1952 33405 1961 33439
rect 1961 33405 1995 33439
rect 1995 33405 2004 33439
rect 1952 33396 2004 33405
rect 2780 33439 2832 33448
rect 2780 33405 2789 33439
rect 2789 33405 2823 33439
rect 2823 33405 2832 33439
rect 2780 33396 2832 33405
rect 21180 33439 21232 33448
rect 21180 33405 21189 33439
rect 21189 33405 21223 33439
rect 21223 33405 21232 33439
rect 21180 33396 21232 33405
rect 21916 33396 21968 33448
rect 22284 33507 22336 33516
rect 22284 33473 22293 33507
rect 22293 33473 22327 33507
rect 22327 33473 22336 33507
rect 22560 33532 22612 33584
rect 22284 33464 22336 33473
rect 22928 33507 22980 33516
rect 22928 33473 22937 33507
rect 22937 33473 22971 33507
rect 22971 33473 22980 33507
rect 22928 33464 22980 33473
rect 23480 33532 23532 33584
rect 26056 33600 26108 33652
rect 28356 33643 28408 33652
rect 28356 33609 28365 33643
rect 28365 33609 28399 33643
rect 28399 33609 28408 33643
rect 28356 33600 28408 33609
rect 29552 33600 29604 33652
rect 31760 33532 31812 33584
rect 23940 33464 23992 33516
rect 24216 33464 24268 33516
rect 25412 33464 25464 33516
rect 26424 33507 26476 33516
rect 26424 33473 26433 33507
rect 26433 33473 26467 33507
rect 26467 33473 26476 33507
rect 26424 33464 26476 33473
rect 26976 33507 27028 33516
rect 26976 33473 26985 33507
rect 26985 33473 27019 33507
rect 27019 33473 27028 33507
rect 26976 33464 27028 33473
rect 27068 33464 27120 33516
rect 30564 33464 30616 33516
rect 31024 33507 31076 33516
rect 31024 33473 31033 33507
rect 31033 33473 31067 33507
rect 31067 33473 31076 33507
rect 31024 33464 31076 33473
rect 31944 33464 31996 33516
rect 46020 33464 46072 33516
rect 22376 33396 22428 33448
rect 22560 33396 22612 33448
rect 24584 33396 24636 33448
rect 46204 33439 46256 33448
rect 19892 33260 19944 33312
rect 20444 33260 20496 33312
rect 21364 33260 21416 33312
rect 25320 33328 25372 33380
rect 23296 33260 23348 33312
rect 23572 33260 23624 33312
rect 24400 33260 24452 33312
rect 46204 33405 46213 33439
rect 46213 33405 46247 33439
rect 46247 33405 46256 33439
rect 46204 33396 46256 33405
rect 32864 33260 32916 33312
rect 47768 33303 47820 33312
rect 47768 33269 47777 33303
rect 47777 33269 47811 33303
rect 47811 33269 47820 33303
rect 47768 33260 47820 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 1952 33056 2004 33108
rect 19984 33056 20036 33108
rect 20444 33056 20496 33108
rect 22928 33056 22980 33108
rect 23848 33056 23900 33108
rect 20996 32988 21048 33040
rect 15200 32920 15252 32972
rect 19984 32920 20036 32972
rect 20352 32963 20404 32972
rect 20352 32929 20361 32963
rect 20361 32929 20395 32963
rect 20395 32929 20404 32963
rect 20352 32920 20404 32929
rect 24216 32988 24268 33040
rect 1952 32852 2004 32904
rect 2136 32852 2188 32904
rect 2412 32852 2464 32904
rect 2688 32895 2740 32904
rect 2688 32861 2697 32895
rect 2697 32861 2731 32895
rect 2731 32861 2740 32895
rect 2688 32852 2740 32861
rect 15568 32895 15620 32904
rect 15568 32861 15577 32895
rect 15577 32861 15611 32895
rect 15611 32861 15620 32895
rect 15568 32852 15620 32861
rect 20076 32852 20128 32904
rect 22008 32920 22060 32972
rect 20536 32895 20588 32904
rect 20536 32861 20545 32895
rect 20545 32861 20579 32895
rect 20579 32861 20588 32895
rect 20536 32852 20588 32861
rect 20812 32852 20864 32904
rect 15752 32827 15804 32836
rect 15752 32793 15761 32827
rect 15761 32793 15795 32827
rect 15795 32793 15804 32827
rect 15752 32784 15804 32793
rect 20720 32784 20772 32836
rect 20904 32784 20956 32836
rect 23572 32852 23624 32904
rect 23756 32852 23808 32904
rect 24308 32920 24360 32972
rect 24768 33056 24820 33108
rect 27068 33056 27120 33108
rect 30472 33099 30524 33108
rect 30472 33065 30481 33099
rect 30481 33065 30515 33099
rect 30515 33065 30524 33099
rect 30472 33056 30524 33065
rect 30564 33056 30616 33108
rect 35900 33056 35952 33108
rect 31300 32988 31352 33040
rect 26148 32852 26200 32904
rect 27344 32920 27396 32972
rect 28816 32963 28868 32972
rect 27252 32895 27304 32904
rect 27252 32861 27261 32895
rect 27261 32861 27295 32895
rect 27295 32861 27304 32895
rect 27252 32852 27304 32861
rect 27712 32852 27764 32904
rect 23480 32827 23532 32836
rect 23480 32793 23489 32827
rect 23489 32793 23523 32827
rect 23523 32793 23532 32827
rect 23480 32784 23532 32793
rect 2136 32716 2188 32768
rect 20812 32716 20864 32768
rect 23204 32716 23256 32768
rect 25780 32784 25832 32836
rect 28080 32784 28132 32836
rect 28816 32929 28825 32963
rect 28825 32929 28859 32963
rect 28859 32929 28868 32963
rect 28816 32920 28868 32929
rect 30840 32920 30892 32972
rect 31668 32963 31720 32972
rect 31668 32929 31677 32963
rect 31677 32929 31711 32963
rect 31711 32929 31720 32963
rect 31668 32920 31720 32929
rect 32128 32920 32180 32972
rect 32588 32963 32640 32972
rect 32588 32929 32597 32963
rect 32597 32929 32631 32963
rect 32631 32929 32640 32963
rect 32588 32920 32640 32929
rect 47768 32920 47820 32972
rect 48044 32963 48096 32972
rect 48044 32929 48053 32963
rect 48053 32929 48087 32963
rect 48087 32929 48096 32963
rect 48044 32920 48096 32929
rect 31484 32895 31536 32904
rect 31484 32861 31493 32895
rect 31493 32861 31527 32895
rect 31527 32861 31536 32895
rect 31484 32852 31536 32861
rect 31208 32784 31260 32836
rect 24860 32716 24912 32768
rect 28172 32716 28224 32768
rect 28632 32759 28684 32768
rect 28632 32725 28641 32759
rect 28641 32725 28675 32759
rect 28675 32725 28684 32759
rect 28632 32716 28684 32725
rect 31116 32759 31168 32768
rect 31116 32725 31125 32759
rect 31125 32725 31159 32759
rect 31159 32725 31168 32759
rect 31116 32716 31168 32725
rect 32312 32852 32364 32904
rect 32404 32784 32456 32836
rect 46480 32827 46532 32836
rect 46480 32793 46489 32827
rect 46489 32793 46523 32827
rect 46523 32793 46532 32827
rect 46480 32784 46532 32793
rect 34060 32716 34112 32768
rect 40776 32716 40828 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 15752 32512 15804 32564
rect 19432 32512 19484 32564
rect 23204 32555 23256 32564
rect 23204 32521 23213 32555
rect 23213 32521 23247 32555
rect 23247 32521 23256 32555
rect 23204 32512 23256 32521
rect 23388 32512 23440 32564
rect 23480 32512 23532 32564
rect 24676 32555 24728 32564
rect 24676 32521 24685 32555
rect 24685 32521 24719 32555
rect 24719 32521 24728 32555
rect 24676 32512 24728 32521
rect 28632 32512 28684 32564
rect 28908 32512 28960 32564
rect 2136 32487 2188 32496
rect 2136 32453 2145 32487
rect 2145 32453 2179 32487
rect 2179 32453 2188 32487
rect 2136 32444 2188 32453
rect 1952 32419 2004 32428
rect 1952 32385 1961 32419
rect 1961 32385 1995 32419
rect 1995 32385 2004 32419
rect 1952 32376 2004 32385
rect 12624 32376 12676 32428
rect 18236 32419 18288 32428
rect 18236 32385 18245 32419
rect 18245 32385 18279 32419
rect 18279 32385 18288 32419
rect 18236 32376 18288 32385
rect 18420 32419 18472 32428
rect 18420 32385 18429 32419
rect 18429 32385 18463 32419
rect 18463 32385 18472 32419
rect 18420 32376 18472 32385
rect 21548 32444 21600 32496
rect 22560 32487 22612 32496
rect 22560 32453 22569 32487
rect 22569 32453 22603 32487
rect 22603 32453 22612 32487
rect 22560 32444 22612 32453
rect 22928 32444 22980 32496
rect 20352 32376 20404 32428
rect 2780 32351 2832 32360
rect 2780 32317 2789 32351
rect 2789 32317 2823 32351
rect 2823 32317 2832 32351
rect 2780 32308 2832 32317
rect 20628 32419 20680 32428
rect 20628 32385 20637 32419
rect 20637 32385 20671 32419
rect 20671 32385 20680 32419
rect 20628 32376 20680 32385
rect 20812 32419 20864 32428
rect 20812 32385 20821 32419
rect 20821 32385 20855 32419
rect 20855 32385 20864 32419
rect 20812 32376 20864 32385
rect 21640 32376 21692 32428
rect 22008 32376 22060 32428
rect 24032 32444 24084 32496
rect 30564 32444 30616 32496
rect 31944 32512 31996 32564
rect 32128 32512 32180 32564
rect 32496 32512 32548 32564
rect 32588 32512 32640 32564
rect 33784 32512 33836 32564
rect 36452 32555 36504 32564
rect 32312 32444 32364 32496
rect 36452 32521 36461 32555
rect 36461 32521 36495 32555
rect 36495 32521 36504 32555
rect 36452 32512 36504 32521
rect 39120 32487 39172 32496
rect 1952 32240 2004 32292
rect 18420 32240 18472 32292
rect 22192 32308 22244 32360
rect 15660 32172 15712 32224
rect 16856 32172 16908 32224
rect 17960 32172 18012 32224
rect 19432 32172 19484 32224
rect 19984 32172 20036 32224
rect 20076 32172 20128 32224
rect 22376 32240 22428 32292
rect 23572 32385 23581 32412
rect 23581 32385 23615 32412
rect 23615 32385 23624 32412
rect 23572 32360 23624 32385
rect 23940 32376 23992 32428
rect 24492 32376 24544 32428
rect 26424 32419 26476 32428
rect 23756 32308 23808 32360
rect 24584 32308 24636 32360
rect 26424 32385 26433 32419
rect 26433 32385 26467 32419
rect 26467 32385 26476 32419
rect 26424 32376 26476 32385
rect 26976 32376 27028 32428
rect 27436 32376 27488 32428
rect 27988 32376 28040 32428
rect 39120 32453 39129 32487
rect 39129 32453 39163 32487
rect 39163 32453 39172 32487
rect 39120 32444 39172 32453
rect 32588 32419 32640 32428
rect 32588 32385 32597 32419
rect 32597 32385 32631 32419
rect 32631 32385 32640 32419
rect 32588 32376 32640 32385
rect 28356 32308 28408 32360
rect 28908 32308 28960 32360
rect 31300 32351 31352 32360
rect 31300 32317 31309 32351
rect 31309 32317 31343 32351
rect 31343 32317 31352 32351
rect 31300 32308 31352 32317
rect 26240 32283 26292 32292
rect 26240 32249 26249 32283
rect 26249 32249 26283 32283
rect 26283 32249 26292 32283
rect 26240 32240 26292 32249
rect 28816 32240 28868 32292
rect 31668 32308 31720 32360
rect 32496 32308 32548 32360
rect 36360 32419 36412 32428
rect 36360 32385 36369 32419
rect 36369 32385 36403 32419
rect 36403 32385 36412 32419
rect 36360 32376 36412 32385
rect 46388 32419 46440 32428
rect 46388 32385 46397 32419
rect 46397 32385 46431 32419
rect 46431 32385 46440 32419
rect 46388 32376 46440 32385
rect 37464 32351 37516 32360
rect 21456 32172 21508 32224
rect 22560 32172 22612 32224
rect 22836 32172 22888 32224
rect 23204 32172 23256 32224
rect 23480 32172 23532 32224
rect 24492 32172 24544 32224
rect 25780 32172 25832 32224
rect 28356 32172 28408 32224
rect 32036 32172 32088 32224
rect 37464 32317 37473 32351
rect 37473 32317 37507 32351
rect 37507 32317 37516 32351
rect 37464 32308 37516 32317
rect 46204 32308 46256 32360
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 15568 31968 15620 32020
rect 16856 31968 16908 32020
rect 22192 31968 22244 32020
rect 23020 31968 23072 32020
rect 23940 31968 23992 32020
rect 21180 31943 21232 31952
rect 21180 31909 21189 31943
rect 21189 31909 21223 31943
rect 21223 31909 21232 31943
rect 21180 31900 21232 31909
rect 22376 31943 22428 31952
rect 22376 31909 22385 31943
rect 22385 31909 22419 31943
rect 22419 31909 22428 31943
rect 22376 31900 22428 31909
rect 23572 31900 23624 31952
rect 2780 31832 2832 31884
rect 2872 31875 2924 31884
rect 2872 31841 2881 31875
rect 2881 31841 2915 31875
rect 2915 31841 2924 31875
rect 2872 31832 2924 31841
rect 19340 31832 19392 31884
rect 20812 31832 20864 31884
rect 23296 31832 23348 31884
rect 16580 31764 16632 31816
rect 21824 31764 21876 31816
rect 22284 31764 22336 31816
rect 23480 31807 23532 31816
rect 23480 31773 23489 31807
rect 23489 31773 23523 31807
rect 23523 31773 23532 31807
rect 23480 31764 23532 31773
rect 24124 31764 24176 31816
rect 24860 31807 24912 31816
rect 24860 31773 24869 31807
rect 24869 31773 24903 31807
rect 24903 31773 24912 31807
rect 27436 31968 27488 32020
rect 27712 31968 27764 32020
rect 24860 31764 24912 31773
rect 25228 31764 25280 31816
rect 2044 31696 2096 31748
rect 15660 31696 15712 31748
rect 16856 31696 16908 31748
rect 20076 31739 20128 31748
rect 20076 31705 20110 31739
rect 20110 31705 20128 31739
rect 20076 31696 20128 31705
rect 23020 31696 23072 31748
rect 27344 31900 27396 31952
rect 27344 31807 27396 31816
rect 27344 31773 27353 31807
rect 27353 31773 27387 31807
rect 27387 31773 27396 31807
rect 27344 31764 27396 31773
rect 32036 31900 32088 31952
rect 32404 31943 32456 31952
rect 32404 31909 32413 31943
rect 32413 31909 32447 31943
rect 32447 31909 32456 31943
rect 32404 31900 32456 31909
rect 37464 31968 37516 32020
rect 46480 31968 46532 32020
rect 27712 31807 27764 31816
rect 27712 31773 27721 31807
rect 27721 31773 27755 31807
rect 27755 31773 27764 31807
rect 27712 31764 27764 31773
rect 28172 31807 28224 31816
rect 28172 31773 28181 31807
rect 28181 31773 28215 31807
rect 28215 31773 28224 31807
rect 28172 31764 28224 31773
rect 28356 31807 28408 31816
rect 28356 31773 28365 31807
rect 28365 31773 28399 31807
rect 28399 31773 28408 31807
rect 28356 31764 28408 31773
rect 18512 31671 18564 31680
rect 18512 31637 18521 31671
rect 18521 31637 18555 31671
rect 18555 31637 18564 31671
rect 18512 31628 18564 31637
rect 21732 31628 21784 31680
rect 22192 31628 22244 31680
rect 24492 31628 24544 31680
rect 26608 31696 26660 31748
rect 27252 31696 27304 31748
rect 31116 31764 31168 31816
rect 31760 31807 31812 31816
rect 31760 31773 31769 31807
rect 31769 31773 31803 31807
rect 31803 31773 31812 31807
rect 31760 31764 31812 31773
rect 32128 31696 32180 31748
rect 32956 31764 33008 31816
rect 33232 31832 33284 31884
rect 34060 31832 34112 31884
rect 38568 31875 38620 31884
rect 38568 31841 38577 31875
rect 38577 31841 38611 31875
rect 38611 31841 38620 31875
rect 38568 31832 38620 31841
rect 46572 31832 46624 31884
rect 33600 31807 33652 31816
rect 33600 31773 33609 31807
rect 33609 31773 33643 31807
rect 33643 31773 33652 31807
rect 33600 31764 33652 31773
rect 35900 31764 35952 31816
rect 36360 31764 36412 31816
rect 36636 31764 36688 31816
rect 37188 31807 37240 31816
rect 37188 31773 37197 31807
rect 37197 31773 37231 31807
rect 37231 31773 37240 31807
rect 37188 31764 37240 31773
rect 45468 31764 45520 31816
rect 47400 31764 47452 31816
rect 33784 31739 33836 31748
rect 33784 31705 33793 31739
rect 33793 31705 33827 31739
rect 33827 31705 33836 31739
rect 33784 31696 33836 31705
rect 37372 31739 37424 31748
rect 37372 31705 37381 31739
rect 37381 31705 37415 31739
rect 37415 31705 37424 31739
rect 37372 31696 37424 31705
rect 32956 31628 33008 31680
rect 33048 31628 33100 31680
rect 35808 31628 35860 31680
rect 46204 31628 46256 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 2780 31467 2832 31476
rect 2780 31433 2789 31467
rect 2789 31433 2823 31467
rect 2823 31433 2832 31467
rect 2780 31424 2832 31433
rect 16856 31467 16908 31476
rect 16856 31433 16865 31467
rect 16865 31433 16899 31467
rect 16899 31433 16908 31467
rect 16856 31424 16908 31433
rect 1400 31331 1452 31340
rect 1400 31297 1409 31331
rect 1409 31297 1443 31331
rect 1443 31297 1452 31331
rect 1400 31288 1452 31297
rect 1768 31288 1820 31340
rect 3700 31288 3752 31340
rect 17960 31356 18012 31408
rect 18236 31424 18288 31476
rect 19432 31424 19484 31476
rect 20168 31424 20220 31476
rect 20628 31424 20680 31476
rect 28448 31467 28500 31476
rect 17500 31331 17552 31340
rect 17500 31297 17509 31331
rect 17509 31297 17543 31331
rect 17543 31297 17552 31331
rect 17500 31288 17552 31297
rect 18512 31288 18564 31340
rect 21916 31356 21968 31408
rect 22376 31356 22428 31408
rect 23480 31356 23532 31408
rect 17592 31220 17644 31272
rect 19156 31263 19208 31272
rect 19156 31229 19165 31263
rect 19165 31229 19199 31263
rect 19199 31229 19208 31263
rect 19156 31220 19208 31229
rect 20720 31220 20772 31272
rect 25044 31288 25096 31340
rect 25780 31288 25832 31340
rect 23388 31220 23440 31272
rect 24216 31220 24268 31272
rect 28448 31433 28457 31467
rect 28457 31433 28491 31467
rect 28491 31433 28500 31467
rect 28448 31424 28500 31433
rect 26976 31356 27028 31408
rect 27988 31399 28040 31408
rect 29736 31424 29788 31476
rect 31024 31424 31076 31476
rect 32496 31424 32548 31476
rect 37372 31467 37424 31476
rect 27988 31365 28013 31399
rect 28013 31365 28040 31399
rect 27988 31356 28040 31365
rect 37372 31433 37381 31467
rect 37381 31433 37415 31467
rect 37415 31433 37424 31467
rect 37372 31424 37424 31433
rect 39764 31399 39816 31408
rect 31300 31288 31352 31340
rect 31392 31331 31444 31340
rect 31392 31297 31401 31331
rect 31401 31297 31435 31331
rect 31435 31297 31444 31331
rect 31392 31288 31444 31297
rect 32588 31288 32640 31340
rect 29828 31263 29880 31272
rect 29828 31229 29837 31263
rect 29837 31229 29871 31263
rect 29871 31229 29880 31263
rect 29828 31220 29880 31229
rect 30012 31263 30064 31272
rect 30012 31229 30021 31263
rect 30021 31229 30055 31263
rect 30055 31229 30064 31263
rect 30012 31220 30064 31229
rect 20168 31152 20220 31204
rect 15016 31084 15068 31136
rect 26976 31152 27028 31204
rect 32036 31220 32088 31272
rect 32864 31331 32916 31340
rect 32864 31297 32873 31331
rect 32873 31297 32907 31331
rect 32907 31297 32916 31331
rect 32864 31288 32916 31297
rect 33232 31288 33284 31340
rect 35992 31288 36044 31340
rect 39764 31365 39773 31399
rect 39773 31365 39807 31399
rect 39807 31365 39816 31399
rect 39764 31356 39816 31365
rect 43904 31288 43956 31340
rect 35348 31220 35400 31272
rect 35808 31220 35860 31272
rect 36268 31220 36320 31272
rect 36544 31220 36596 31272
rect 38108 31263 38160 31272
rect 38108 31229 38117 31263
rect 38117 31229 38151 31263
rect 38151 31229 38160 31263
rect 38108 31220 38160 31229
rect 38016 31152 38068 31204
rect 20720 31084 20772 31136
rect 21088 31084 21140 31136
rect 22560 31084 22612 31136
rect 23388 31084 23440 31136
rect 24584 31084 24636 31136
rect 28908 31084 28960 31136
rect 29184 31127 29236 31136
rect 29184 31093 29193 31127
rect 29193 31093 29227 31127
rect 29227 31093 29236 31127
rect 29184 31084 29236 31093
rect 30012 31084 30064 31136
rect 35348 31084 35400 31136
rect 35624 31084 35676 31136
rect 46572 31084 46624 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 2044 30923 2096 30932
rect 2044 30889 2053 30923
rect 2053 30889 2087 30923
rect 2087 30889 2096 30923
rect 2044 30880 2096 30889
rect 17500 30880 17552 30932
rect 20996 30880 21048 30932
rect 21640 30880 21692 30932
rect 27344 30880 27396 30932
rect 29000 30923 29052 30932
rect 29000 30889 29009 30923
rect 29009 30889 29043 30923
rect 29043 30889 29052 30923
rect 29000 30880 29052 30889
rect 31300 30923 31352 30932
rect 31300 30889 31309 30923
rect 31309 30889 31343 30923
rect 31343 30889 31352 30923
rect 31300 30880 31352 30889
rect 38108 30880 38160 30932
rect 18420 30812 18472 30864
rect 16580 30787 16632 30796
rect 16580 30753 16589 30787
rect 16589 30753 16623 30787
rect 16623 30753 16632 30787
rect 16580 30744 16632 30753
rect 17592 30744 17644 30796
rect 21732 30812 21784 30864
rect 22008 30812 22060 30864
rect 19340 30676 19392 30728
rect 19984 30676 20036 30728
rect 16672 30608 16724 30660
rect 18144 30608 18196 30660
rect 19432 30651 19484 30660
rect 19432 30617 19441 30651
rect 19441 30617 19475 30651
rect 19475 30617 19484 30651
rect 19432 30608 19484 30617
rect 17132 30540 17184 30592
rect 20444 30540 20496 30592
rect 21088 30676 21140 30728
rect 21456 30744 21508 30796
rect 21732 30676 21784 30728
rect 22744 30744 22796 30796
rect 28908 30812 28960 30864
rect 29092 30812 29144 30864
rect 24308 30744 24360 30796
rect 21916 30608 21968 30660
rect 24492 30676 24544 30728
rect 27160 30676 27212 30728
rect 22284 30540 22336 30592
rect 23296 30608 23348 30660
rect 24768 30608 24820 30660
rect 29552 30676 29604 30728
rect 29920 30719 29972 30728
rect 29920 30685 29929 30719
rect 29929 30685 29963 30719
rect 29963 30685 29972 30719
rect 29920 30676 29972 30685
rect 30012 30676 30064 30728
rect 36544 30719 36596 30728
rect 36544 30685 36553 30719
rect 36553 30685 36587 30719
rect 36587 30685 36596 30719
rect 36544 30676 36596 30685
rect 36636 30676 36688 30728
rect 45468 30676 45520 30728
rect 22468 30540 22520 30592
rect 22652 30540 22704 30592
rect 23388 30540 23440 30592
rect 28632 30608 28684 30660
rect 35992 30651 36044 30660
rect 35992 30617 36001 30651
rect 36001 30617 36035 30651
rect 36035 30617 36044 30651
rect 35992 30608 36044 30617
rect 36912 30651 36964 30660
rect 36912 30617 36921 30651
rect 36921 30617 36955 30651
rect 36955 30617 36964 30651
rect 36912 30608 36964 30617
rect 46388 30608 46440 30660
rect 36636 30540 36688 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 3424 30336 3476 30388
rect 36912 30336 36964 30388
rect 16672 30311 16724 30320
rect 16672 30277 16681 30311
rect 16681 30277 16715 30311
rect 16715 30277 16724 30311
rect 16672 30268 16724 30277
rect 20536 30268 20588 30320
rect 2412 30200 2464 30252
rect 14832 30200 14884 30252
rect 1860 30132 1912 30184
rect 2228 30132 2280 30184
rect 17132 30243 17184 30252
rect 17132 30209 17146 30243
rect 17146 30209 17180 30243
rect 17180 30209 17184 30243
rect 17132 30200 17184 30209
rect 17500 30200 17552 30252
rect 18420 30200 18472 30252
rect 19708 30243 19760 30252
rect 19708 30209 19717 30243
rect 19717 30209 19751 30243
rect 19751 30209 19760 30243
rect 19708 30200 19760 30209
rect 20812 30268 20864 30320
rect 21180 30268 21232 30320
rect 22284 30268 22336 30320
rect 20904 30243 20956 30252
rect 20904 30209 20913 30243
rect 20913 30209 20947 30243
rect 20947 30209 20956 30243
rect 20904 30200 20956 30209
rect 17040 30064 17092 30116
rect 17592 30064 17644 30116
rect 18144 30107 18196 30116
rect 18144 30073 18153 30107
rect 18153 30073 18187 30107
rect 18187 30073 18196 30107
rect 18144 30064 18196 30073
rect 19156 30064 19208 30116
rect 1400 29996 1452 30048
rect 2228 30039 2280 30048
rect 2228 30005 2237 30039
rect 2237 30005 2271 30039
rect 2271 30005 2280 30039
rect 2228 29996 2280 30005
rect 17776 29996 17828 30048
rect 21916 30200 21968 30252
rect 23940 30200 23992 30252
rect 24584 30200 24636 30252
rect 24860 30243 24912 30252
rect 24860 30209 24869 30243
rect 24869 30209 24903 30243
rect 24903 30209 24912 30243
rect 24860 30200 24912 30209
rect 25596 30243 25648 30252
rect 25596 30209 25605 30243
rect 25605 30209 25639 30243
rect 25639 30209 25648 30243
rect 25596 30200 25648 30209
rect 26424 30200 26476 30252
rect 27436 30243 27488 30252
rect 27436 30209 27445 30243
rect 27445 30209 27479 30243
rect 27479 30209 27488 30243
rect 27436 30200 27488 30209
rect 28908 30243 28960 30252
rect 28908 30209 28917 30243
rect 28917 30209 28951 30243
rect 28951 30209 28960 30243
rect 28908 30200 28960 30209
rect 29184 30200 29236 30252
rect 29920 30243 29972 30252
rect 29920 30209 29929 30243
rect 29929 30209 29963 30243
rect 29963 30209 29972 30243
rect 29920 30200 29972 30209
rect 30012 30200 30064 30252
rect 36544 30200 36596 30252
rect 47952 30243 48004 30252
rect 47952 30209 47961 30243
rect 47961 30209 47995 30243
rect 47995 30209 48004 30243
rect 47952 30200 48004 30209
rect 21732 30132 21784 30184
rect 23296 30175 23348 30184
rect 23296 30141 23305 30175
rect 23305 30141 23339 30175
rect 23339 30141 23348 30175
rect 23296 30132 23348 30141
rect 23388 30175 23440 30184
rect 23388 30141 23397 30175
rect 23397 30141 23431 30175
rect 23431 30141 23440 30175
rect 28632 30175 28684 30184
rect 23388 30132 23440 30141
rect 28632 30141 28641 30175
rect 28641 30141 28675 30175
rect 28675 30141 28684 30175
rect 28632 30132 28684 30141
rect 21548 30064 21600 30116
rect 22008 30064 22060 30116
rect 29368 30132 29420 30184
rect 31208 30064 31260 30116
rect 22652 29996 22704 30048
rect 22744 29996 22796 30048
rect 24952 29996 25004 30048
rect 27344 29996 27396 30048
rect 27988 29996 28040 30048
rect 29000 29996 29052 30048
rect 37464 30039 37516 30048
rect 37464 30005 37473 30039
rect 37473 30005 37507 30039
rect 37507 30005 37516 30039
rect 37464 29996 37516 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 19432 29792 19484 29844
rect 19708 29792 19760 29844
rect 24860 29792 24912 29844
rect 23940 29724 23992 29776
rect 27436 29792 27488 29844
rect 30012 29792 30064 29844
rect 31576 29792 31628 29844
rect 1400 29699 1452 29708
rect 1400 29665 1409 29699
rect 1409 29665 1443 29699
rect 1443 29665 1452 29699
rect 1400 29656 1452 29665
rect 2228 29656 2280 29708
rect 2780 29699 2832 29708
rect 2780 29665 2789 29699
rect 2789 29665 2823 29699
rect 2823 29665 2832 29699
rect 2780 29656 2832 29665
rect 21824 29656 21876 29708
rect 29000 29656 29052 29708
rect 29828 29656 29880 29708
rect 30012 29699 30064 29708
rect 30012 29665 30021 29699
rect 30021 29665 30055 29699
rect 30055 29665 30064 29699
rect 30012 29656 30064 29665
rect 31208 29656 31260 29708
rect 16856 29588 16908 29640
rect 20444 29631 20496 29640
rect 20444 29597 20478 29631
rect 20478 29597 20496 29631
rect 20444 29588 20496 29597
rect 25044 29588 25096 29640
rect 29368 29588 29420 29640
rect 30196 29631 30248 29640
rect 30196 29597 30205 29631
rect 30205 29597 30239 29631
rect 30239 29597 30248 29631
rect 30196 29588 30248 29597
rect 30288 29631 30340 29640
rect 30288 29597 30297 29631
rect 30297 29597 30331 29631
rect 30331 29597 30340 29631
rect 30288 29588 30340 29597
rect 16672 29520 16724 29572
rect 22284 29520 22336 29572
rect 24308 29520 24360 29572
rect 27988 29520 28040 29572
rect 30012 29520 30064 29572
rect 31760 29520 31812 29572
rect 20904 29452 20956 29504
rect 21732 29452 21784 29504
rect 28724 29452 28776 29504
rect 32956 29792 33008 29844
rect 34796 29835 34848 29844
rect 34796 29801 34805 29835
rect 34805 29801 34839 29835
rect 34839 29801 34848 29835
rect 34796 29792 34848 29801
rect 38660 29835 38712 29844
rect 38660 29801 38669 29835
rect 38669 29801 38703 29835
rect 38703 29801 38712 29835
rect 38660 29792 38712 29801
rect 33784 29656 33836 29708
rect 34704 29631 34756 29640
rect 34704 29597 34713 29631
rect 34713 29597 34747 29631
rect 34747 29597 34756 29631
rect 34704 29588 34756 29597
rect 34888 29631 34940 29640
rect 34888 29597 34897 29631
rect 34897 29597 34931 29631
rect 34931 29597 34940 29631
rect 34888 29588 34940 29597
rect 46296 29588 46348 29640
rect 37280 29520 37332 29572
rect 37556 29563 37608 29572
rect 37556 29529 37590 29563
rect 37590 29529 37608 29563
rect 37556 29520 37608 29529
rect 33876 29452 33928 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 16672 29291 16724 29300
rect 16672 29257 16681 29291
rect 16681 29257 16715 29291
rect 16715 29257 16724 29291
rect 16672 29248 16724 29257
rect 22284 29248 22336 29300
rect 24308 29291 24360 29300
rect 24308 29257 24317 29291
rect 24317 29257 24351 29291
rect 24351 29257 24360 29291
rect 24308 29248 24360 29257
rect 29000 29248 29052 29300
rect 29184 29248 29236 29300
rect 8852 29112 8904 29164
rect 17037 29158 17089 29167
rect 17037 29124 17064 29158
rect 17064 29124 17089 29158
rect 17037 29115 17089 29124
rect 22192 29180 22244 29232
rect 17500 29112 17552 29164
rect 17776 29155 17828 29164
rect 17776 29121 17785 29155
rect 17785 29121 17819 29155
rect 17819 29121 17828 29155
rect 17776 29112 17828 29121
rect 19340 29112 19392 29164
rect 22560 29180 22612 29232
rect 29828 29248 29880 29300
rect 30288 29248 30340 29300
rect 31392 29248 31444 29300
rect 32588 29248 32640 29300
rect 46940 29248 46992 29300
rect 47400 29248 47452 29300
rect 3424 28976 3476 29028
rect 15476 28976 15528 29028
rect 22468 29155 22520 29164
rect 22468 29121 22477 29155
rect 22477 29121 22511 29155
rect 22511 29121 22520 29155
rect 22468 29112 22520 29121
rect 23204 29112 23256 29164
rect 23388 29044 23440 29096
rect 24768 29155 24820 29164
rect 24768 29121 24777 29155
rect 24777 29121 24811 29155
rect 24811 29121 24820 29155
rect 24952 29155 25004 29164
rect 24768 29112 24820 29121
rect 24952 29121 24961 29155
rect 24961 29121 24995 29155
rect 24995 29121 25004 29155
rect 24952 29112 25004 29121
rect 28448 29155 28500 29164
rect 28448 29121 28457 29155
rect 28457 29121 28491 29155
rect 28491 29121 28500 29155
rect 28448 29112 28500 29121
rect 28724 29155 28776 29164
rect 28724 29121 28733 29155
rect 28733 29121 28767 29155
rect 28767 29121 28776 29155
rect 28724 29112 28776 29121
rect 30380 29112 30432 29164
rect 34520 29180 34572 29232
rect 34796 29180 34848 29232
rect 22652 28976 22704 29028
rect 25596 29044 25648 29096
rect 35532 29112 35584 29164
rect 37280 29155 37332 29164
rect 34704 29044 34756 29096
rect 37280 29121 37289 29155
rect 37289 29121 37323 29155
rect 37323 29121 37332 29155
rect 37280 29112 37332 29121
rect 46940 29112 46992 29164
rect 37464 29044 37516 29096
rect 38476 29044 38528 29096
rect 39580 29044 39632 29096
rect 29000 28976 29052 29028
rect 29368 28976 29420 29028
rect 2044 28951 2096 28960
rect 2044 28917 2053 28951
rect 2053 28917 2087 28951
rect 2087 28917 2096 28951
rect 2044 28908 2096 28917
rect 29092 28908 29144 28960
rect 29828 28908 29880 28960
rect 34244 28908 34296 28960
rect 34888 28976 34940 29028
rect 46572 28976 46624 29028
rect 34796 28908 34848 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 2044 28568 2096 28620
rect 2780 28611 2832 28620
rect 2780 28577 2789 28611
rect 2789 28577 2823 28611
rect 2823 28577 2832 28611
rect 2780 28568 2832 28577
rect 26424 28704 26476 28756
rect 26608 28704 26660 28756
rect 27988 28747 28040 28756
rect 27988 28713 27997 28747
rect 27997 28713 28031 28747
rect 28031 28713 28040 28747
rect 27988 28704 28040 28713
rect 24676 28636 24728 28688
rect 22836 28568 22888 28620
rect 22008 28500 22060 28552
rect 24676 28543 24728 28552
rect 24676 28509 24685 28543
rect 24685 28509 24719 28543
rect 24719 28509 24728 28543
rect 24676 28500 24728 28509
rect 24860 28543 24912 28552
rect 24860 28509 24869 28543
rect 24869 28509 24903 28543
rect 24903 28509 24912 28543
rect 24860 28500 24912 28509
rect 25228 28500 25280 28552
rect 25780 28568 25832 28620
rect 26424 28568 26476 28620
rect 27160 28568 27212 28620
rect 26332 28500 26384 28552
rect 2320 28432 2372 28484
rect 17316 28432 17368 28484
rect 18328 28432 18380 28484
rect 21180 28432 21232 28484
rect 23388 28432 23440 28484
rect 24584 28432 24636 28484
rect 27436 28432 27488 28484
rect 29000 28636 29052 28688
rect 32220 28704 32272 28756
rect 31760 28636 31812 28688
rect 37464 28636 37516 28688
rect 28540 28432 28592 28484
rect 31852 28432 31904 28484
rect 32956 28500 33008 28552
rect 33876 28543 33928 28552
rect 33876 28509 33885 28543
rect 33885 28509 33919 28543
rect 33919 28509 33928 28543
rect 33876 28500 33928 28509
rect 32680 28432 32732 28484
rect 34152 28543 34204 28552
rect 34152 28509 34161 28543
rect 34161 28509 34195 28543
rect 34195 28509 34204 28543
rect 39304 28568 39356 28620
rect 48136 28611 48188 28620
rect 48136 28577 48145 28611
rect 48145 28577 48179 28611
rect 48179 28577 48188 28611
rect 48136 28568 48188 28577
rect 34152 28500 34204 28509
rect 18696 28364 18748 28416
rect 19340 28407 19392 28416
rect 19340 28373 19349 28407
rect 19349 28373 19383 28407
rect 19383 28373 19392 28407
rect 19340 28364 19392 28373
rect 19984 28364 20036 28416
rect 20352 28364 20404 28416
rect 22284 28407 22336 28416
rect 22284 28373 22293 28407
rect 22293 28373 22327 28407
rect 22327 28373 22336 28407
rect 22284 28364 22336 28373
rect 23664 28364 23716 28416
rect 24400 28407 24452 28416
rect 24400 28373 24409 28407
rect 24409 28373 24443 28407
rect 24443 28373 24452 28407
rect 24400 28364 24452 28373
rect 25228 28364 25280 28416
rect 31576 28407 31628 28416
rect 31576 28373 31585 28407
rect 31585 28373 31619 28407
rect 31619 28373 31628 28407
rect 31576 28364 31628 28373
rect 33600 28364 33652 28416
rect 34796 28432 34848 28484
rect 38660 28500 38712 28552
rect 39028 28543 39080 28552
rect 39028 28509 39037 28543
rect 39037 28509 39071 28543
rect 39071 28509 39080 28543
rect 39028 28500 39080 28509
rect 46112 28500 46164 28552
rect 36636 28475 36688 28484
rect 36636 28441 36645 28475
rect 36645 28441 36679 28475
rect 36679 28441 36688 28475
rect 36636 28432 36688 28441
rect 39856 28432 39908 28484
rect 46480 28475 46532 28484
rect 46480 28441 46489 28475
rect 46489 28441 46523 28475
rect 46523 28441 46532 28475
rect 46480 28432 46532 28441
rect 37372 28364 37424 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 2320 28203 2372 28212
rect 2320 28169 2329 28203
rect 2329 28169 2363 28203
rect 2363 28169 2372 28203
rect 2320 28160 2372 28169
rect 18328 28160 18380 28212
rect 20812 28160 20864 28212
rect 2872 28024 2924 28076
rect 3148 28024 3200 28076
rect 12624 28067 12676 28076
rect 12624 28033 12633 28067
rect 12633 28033 12667 28067
rect 12667 28033 12676 28067
rect 12624 28024 12676 28033
rect 19521 28067 19573 28076
rect 1676 27956 1728 28008
rect 2320 27956 2372 28008
rect 16856 27956 16908 28008
rect 12716 27863 12768 27872
rect 12716 27829 12725 27863
rect 12725 27829 12759 27863
rect 12759 27829 12768 27863
rect 12716 27820 12768 27829
rect 18236 27820 18288 27872
rect 19521 28033 19530 28067
rect 19530 28033 19564 28067
rect 19564 28033 19573 28067
rect 19521 28024 19573 28033
rect 20076 28024 20128 28076
rect 21088 28024 21140 28076
rect 21456 28024 21508 28076
rect 22560 28067 22612 28076
rect 22560 28033 22569 28067
rect 22569 28033 22603 28067
rect 22603 28033 22612 28067
rect 22560 28024 22612 28033
rect 19800 27888 19852 27940
rect 19616 27820 19668 27872
rect 21272 27956 21324 28008
rect 23480 28024 23532 28076
rect 23940 28092 23992 28144
rect 24400 28092 24452 28144
rect 25780 28160 25832 28212
rect 24032 28067 24084 28076
rect 24032 28033 24041 28067
rect 24041 28033 24075 28067
rect 24075 28033 24084 28067
rect 24032 28024 24084 28033
rect 25044 28067 25096 28076
rect 25044 28033 25053 28067
rect 25053 28033 25087 28067
rect 25087 28033 25096 28067
rect 25044 28024 25096 28033
rect 28540 28024 28592 28076
rect 29552 28024 29604 28076
rect 31576 28024 31628 28076
rect 32312 28067 32364 28076
rect 32312 28033 32321 28067
rect 32321 28033 32355 28067
rect 32355 28033 32364 28067
rect 32312 28024 32364 28033
rect 24768 27956 24820 28008
rect 29460 27956 29512 28008
rect 21088 27888 21140 27940
rect 23664 27888 23716 27940
rect 31852 27888 31904 27940
rect 31944 27888 31996 27940
rect 34704 28092 34756 28144
rect 33876 28024 33928 28076
rect 36636 28160 36688 28212
rect 37556 28203 37608 28212
rect 37556 28169 37565 28203
rect 37565 28169 37599 28203
rect 37599 28169 37608 28203
rect 37556 28160 37608 28169
rect 35532 28092 35584 28144
rect 35992 28024 36044 28076
rect 37464 28067 37516 28076
rect 37464 28033 37473 28067
rect 37473 28033 37507 28067
rect 37507 28033 37516 28067
rect 37464 28024 37516 28033
rect 38476 28024 38528 28076
rect 47860 28067 47912 28076
rect 47860 28033 47869 28067
rect 47869 28033 47903 28067
rect 47903 28033 47912 28067
rect 47860 28024 47912 28033
rect 44732 27956 44784 28008
rect 45560 27956 45612 28008
rect 46020 27999 46072 28008
rect 46020 27965 46029 27999
rect 46029 27965 46063 27999
rect 46063 27965 46072 27999
rect 46020 27956 46072 27965
rect 19984 27820 20036 27872
rect 22744 27820 22796 27872
rect 23940 27820 23992 27872
rect 27436 27820 27488 27872
rect 29644 27820 29696 27872
rect 32128 27863 32180 27872
rect 32128 27829 32137 27863
rect 32137 27829 32171 27863
rect 32171 27829 32180 27863
rect 32128 27820 32180 27829
rect 33232 27820 33284 27872
rect 39028 27820 39080 27872
rect 47676 27820 47728 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 7012 27548 7064 27600
rect 15752 27548 15804 27600
rect 17316 27591 17368 27600
rect 17316 27557 17325 27591
rect 17325 27557 17359 27591
rect 17359 27557 17368 27591
rect 17316 27548 17368 27557
rect 18512 27548 18564 27600
rect 19800 27616 19852 27668
rect 20812 27591 20864 27600
rect 20812 27557 20821 27591
rect 20821 27557 20855 27591
rect 20855 27557 20864 27591
rect 20812 27548 20864 27557
rect 21732 27548 21784 27600
rect 2596 27480 2648 27532
rect 2964 27480 3016 27532
rect 1768 27455 1820 27464
rect 1768 27421 1777 27455
rect 1777 27421 1811 27455
rect 1811 27421 1820 27455
rect 1768 27412 1820 27421
rect 3056 27455 3108 27464
rect 3056 27421 3065 27455
rect 3065 27421 3099 27455
rect 3099 27421 3108 27455
rect 3056 27412 3108 27421
rect 18420 27455 18472 27464
rect 18420 27421 18429 27455
rect 18429 27421 18463 27455
rect 18463 27421 18472 27455
rect 18420 27412 18472 27421
rect 18512 27455 18564 27464
rect 18512 27421 18521 27455
rect 18521 27421 18555 27455
rect 18555 27421 18564 27455
rect 18696 27455 18748 27464
rect 18512 27412 18564 27421
rect 18696 27421 18705 27455
rect 18705 27421 18739 27455
rect 18739 27421 18748 27455
rect 18696 27412 18748 27421
rect 19432 27455 19484 27464
rect 2596 27344 2648 27396
rect 12256 27344 12308 27396
rect 1952 27276 2004 27328
rect 8300 27276 8352 27328
rect 16580 27276 16632 27328
rect 16856 27344 16908 27396
rect 19432 27421 19441 27455
rect 19441 27421 19475 27455
rect 19475 27421 19484 27455
rect 19432 27412 19484 27421
rect 21180 27412 21232 27464
rect 21456 27412 21508 27464
rect 24032 27616 24084 27668
rect 29552 27659 29604 27668
rect 29552 27625 29561 27659
rect 29561 27625 29595 27659
rect 29595 27625 29604 27659
rect 29552 27616 29604 27625
rect 25964 27548 26016 27600
rect 26056 27548 26108 27600
rect 32312 27616 32364 27668
rect 33232 27659 33284 27668
rect 33232 27625 33241 27659
rect 33241 27625 33275 27659
rect 33275 27625 33284 27659
rect 33232 27616 33284 27625
rect 22560 27480 22612 27532
rect 19248 27276 19300 27328
rect 21272 27344 21324 27396
rect 24676 27412 24728 27464
rect 24584 27387 24636 27396
rect 21916 27276 21968 27328
rect 24584 27353 24593 27387
rect 24593 27353 24627 27387
rect 24627 27353 24636 27387
rect 24584 27344 24636 27353
rect 25228 27276 25280 27328
rect 26148 27455 26200 27464
rect 26148 27421 26157 27455
rect 26157 27421 26191 27455
rect 26191 27421 26200 27455
rect 26148 27412 26200 27421
rect 29460 27480 29512 27532
rect 27712 27344 27764 27396
rect 28448 27344 28500 27396
rect 28724 27344 28776 27396
rect 32220 27548 32272 27600
rect 32772 27548 32824 27600
rect 45560 27591 45612 27600
rect 29644 27412 29696 27464
rect 30196 27412 30248 27464
rect 32128 27412 32180 27464
rect 28172 27319 28224 27328
rect 28172 27285 28181 27319
rect 28181 27285 28215 27319
rect 28215 27285 28224 27319
rect 28172 27276 28224 27285
rect 31944 27344 31996 27396
rect 28908 27276 28960 27328
rect 32680 27412 32732 27464
rect 35808 27412 35860 27464
rect 39672 27480 39724 27532
rect 45560 27557 45569 27591
rect 45569 27557 45603 27591
rect 45603 27557 45612 27591
rect 45560 27548 45612 27557
rect 46296 27523 46348 27532
rect 46296 27489 46305 27523
rect 46305 27489 46339 27523
rect 46339 27489 46348 27523
rect 46296 27480 46348 27489
rect 46572 27480 46624 27532
rect 48228 27480 48280 27532
rect 37096 27412 37148 27464
rect 32588 27344 32640 27396
rect 34060 27387 34112 27396
rect 34060 27353 34069 27387
rect 34069 27353 34103 27387
rect 34103 27353 34112 27387
rect 34060 27344 34112 27353
rect 35164 27387 35216 27396
rect 35164 27353 35173 27387
rect 35173 27353 35207 27387
rect 35207 27353 35216 27387
rect 35164 27344 35216 27353
rect 35624 27344 35676 27396
rect 37280 27344 37332 27396
rect 35532 27319 35584 27328
rect 35532 27285 35541 27319
rect 35541 27285 35575 27319
rect 35575 27285 35584 27319
rect 35532 27276 35584 27285
rect 38476 27412 38528 27464
rect 45468 27455 45520 27464
rect 45468 27421 45477 27455
rect 45477 27421 45511 27455
rect 45511 27421 45520 27455
rect 45468 27412 45520 27421
rect 41696 27387 41748 27396
rect 41696 27353 41705 27387
rect 41705 27353 41739 27387
rect 41739 27353 41748 27387
rect 41696 27344 41748 27353
rect 37464 27276 37516 27328
rect 48044 27276 48096 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 2136 27072 2188 27124
rect 26148 27115 26200 27124
rect 1952 27047 2004 27056
rect 1952 27013 1961 27047
rect 1961 27013 1995 27047
rect 1995 27013 2004 27047
rect 1952 27004 2004 27013
rect 12716 27004 12768 27056
rect 16580 27004 16632 27056
rect 1768 26979 1820 26988
rect 1768 26945 1777 26979
rect 1777 26945 1811 26979
rect 1811 26945 1820 26979
rect 1768 26936 1820 26945
rect 15752 26979 15804 26988
rect 15752 26945 15761 26979
rect 15761 26945 15795 26979
rect 15795 26945 15804 26979
rect 15752 26936 15804 26945
rect 16120 26936 16172 26988
rect 19340 27004 19392 27056
rect 21088 27047 21140 27056
rect 21088 27013 21097 27047
rect 21097 27013 21131 27047
rect 21131 27013 21140 27047
rect 21088 27004 21140 27013
rect 21272 27047 21324 27056
rect 21272 27013 21281 27047
rect 21281 27013 21315 27047
rect 21315 27013 21324 27047
rect 21272 27004 21324 27013
rect 18236 26979 18288 26988
rect 2780 26911 2832 26920
rect 2780 26877 2789 26911
rect 2789 26877 2823 26911
rect 2823 26877 2832 26911
rect 2780 26868 2832 26877
rect 11796 26911 11848 26920
rect 11796 26877 11805 26911
rect 11805 26877 11839 26911
rect 11839 26877 11848 26911
rect 11796 26868 11848 26877
rect 11060 26800 11112 26852
rect 16580 26868 16632 26920
rect 17040 26911 17092 26920
rect 17040 26877 17049 26911
rect 17049 26877 17083 26911
rect 17083 26877 17092 26911
rect 17040 26868 17092 26877
rect 18236 26945 18245 26979
rect 18245 26945 18279 26979
rect 18279 26945 18288 26979
rect 18236 26936 18288 26945
rect 19892 26936 19944 26988
rect 20352 26936 20404 26988
rect 15844 26775 15896 26784
rect 15844 26741 15853 26775
rect 15853 26741 15887 26775
rect 15887 26741 15896 26775
rect 15844 26732 15896 26741
rect 21916 26936 21968 26988
rect 22468 26936 22520 26988
rect 25044 27004 25096 27056
rect 26148 27081 26157 27115
rect 26157 27081 26191 27115
rect 26191 27081 26200 27115
rect 26148 27072 26200 27081
rect 28172 27072 28224 27124
rect 33784 27072 33836 27124
rect 35624 27072 35676 27124
rect 37004 27072 37056 27124
rect 37280 27115 37332 27124
rect 37280 27081 37289 27115
rect 37289 27081 37323 27115
rect 37323 27081 37332 27115
rect 37280 27072 37332 27081
rect 37464 27072 37516 27124
rect 23940 26936 23992 26988
rect 24676 26936 24728 26988
rect 25964 26979 26016 26988
rect 25964 26945 25973 26979
rect 25973 26945 26007 26979
rect 26007 26945 26016 26979
rect 27160 26979 27212 26988
rect 25964 26936 26016 26945
rect 27160 26945 27169 26979
rect 27169 26945 27203 26979
rect 27203 26945 27212 26979
rect 27160 26936 27212 26945
rect 28080 26979 28132 26988
rect 28080 26945 28089 26979
rect 28089 26945 28123 26979
rect 28123 26945 28132 26979
rect 28080 26936 28132 26945
rect 28448 26979 28500 26988
rect 28448 26945 28457 26979
rect 28457 26945 28491 26979
rect 28491 26945 28500 26979
rect 28448 26936 28500 26945
rect 29368 26936 29420 26988
rect 24860 26868 24912 26920
rect 26240 26868 26292 26920
rect 28908 26868 28960 26920
rect 30288 26936 30340 26988
rect 30472 26936 30524 26988
rect 34520 27004 34572 27056
rect 35808 27004 35860 27056
rect 36084 27004 36136 27056
rect 34704 26936 34756 26988
rect 30748 26868 30800 26920
rect 34520 26868 34572 26920
rect 35164 26868 35216 26920
rect 35532 26936 35584 26988
rect 36268 26936 36320 26988
rect 36820 27004 36872 27056
rect 45836 27072 45888 27124
rect 46480 27072 46532 27124
rect 37924 26979 37976 26988
rect 25228 26843 25280 26852
rect 25228 26809 25237 26843
rect 25237 26809 25271 26843
rect 25271 26809 25280 26843
rect 25228 26800 25280 26809
rect 33232 26800 33284 26852
rect 26240 26732 26292 26784
rect 26700 26732 26752 26784
rect 28080 26732 28132 26784
rect 28724 26732 28776 26784
rect 29736 26775 29788 26784
rect 29736 26741 29745 26775
rect 29745 26741 29779 26775
rect 29779 26741 29788 26775
rect 29736 26732 29788 26741
rect 30472 26732 30524 26784
rect 35348 26800 35400 26852
rect 36820 26868 36872 26920
rect 37004 26868 37056 26920
rect 37464 26868 37516 26920
rect 37924 26945 37933 26979
rect 37933 26945 37967 26979
rect 37967 26945 37976 26979
rect 37924 26936 37976 26945
rect 38476 26936 38528 26988
rect 46388 26936 46440 26988
rect 38108 26868 38160 26920
rect 39396 26911 39448 26920
rect 37740 26800 37792 26852
rect 39396 26877 39405 26911
rect 39405 26877 39439 26911
rect 39439 26877 39448 26911
rect 39396 26868 39448 26877
rect 48504 26868 48556 26920
rect 34428 26732 34480 26784
rect 36452 26732 36504 26784
rect 40040 26732 40092 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 2964 26528 3016 26580
rect 11796 26528 11848 26580
rect 19248 26571 19300 26580
rect 19248 26537 19257 26571
rect 19257 26537 19291 26571
rect 19291 26537 19300 26571
rect 19248 26528 19300 26537
rect 19432 26528 19484 26580
rect 3056 26460 3108 26512
rect 2780 26435 2832 26444
rect 2780 26401 2789 26435
rect 2789 26401 2823 26435
rect 2823 26401 2832 26435
rect 2780 26392 2832 26401
rect 17316 26460 17368 26512
rect 20076 26460 20128 26512
rect 22836 26528 22888 26580
rect 23204 26528 23256 26580
rect 24860 26528 24912 26580
rect 25044 26528 25096 26580
rect 26056 26571 26108 26580
rect 26056 26537 26065 26571
rect 26065 26537 26099 26571
rect 26099 26537 26108 26571
rect 26056 26528 26108 26537
rect 15844 26435 15896 26444
rect 15844 26401 15853 26435
rect 15853 26401 15887 26435
rect 15887 26401 15896 26435
rect 15844 26392 15896 26401
rect 17040 26392 17092 26444
rect 18236 26367 18288 26376
rect 18236 26333 18245 26367
rect 18245 26333 18279 26367
rect 18279 26333 18288 26367
rect 18236 26324 18288 26333
rect 18328 26324 18380 26376
rect 18512 26324 18564 26376
rect 19248 26324 19300 26376
rect 2780 26256 2832 26308
rect 17776 26256 17828 26308
rect 19524 26367 19576 26376
rect 19524 26333 19533 26367
rect 19533 26333 19567 26367
rect 19567 26333 19576 26367
rect 19524 26324 19576 26333
rect 20168 26392 20220 26444
rect 19708 26367 19760 26376
rect 19708 26333 19717 26367
rect 19717 26333 19751 26367
rect 19751 26333 19760 26367
rect 19708 26324 19760 26333
rect 19984 26324 20036 26376
rect 23572 26460 23624 26512
rect 26148 26460 26200 26512
rect 22284 26392 22336 26444
rect 22468 26367 22520 26376
rect 22468 26333 22477 26367
rect 22477 26333 22511 26367
rect 22511 26333 22520 26367
rect 22468 26324 22520 26333
rect 24124 26392 24176 26444
rect 27712 26528 27764 26580
rect 27804 26528 27856 26580
rect 28632 26528 28684 26580
rect 29460 26528 29512 26580
rect 26424 26460 26476 26512
rect 30104 26460 30156 26512
rect 32680 26528 32732 26580
rect 35532 26528 35584 26580
rect 37096 26528 37148 26580
rect 39396 26528 39448 26580
rect 35072 26460 35124 26512
rect 30012 26392 30064 26444
rect 30196 26435 30248 26444
rect 30196 26401 30205 26435
rect 30205 26401 30239 26435
rect 30239 26401 30248 26435
rect 30196 26392 30248 26401
rect 21916 26256 21968 26308
rect 22744 26299 22796 26308
rect 22744 26265 22778 26299
rect 22778 26265 22796 26299
rect 22744 26256 22796 26265
rect 22836 26256 22888 26308
rect 29736 26324 29788 26376
rect 32772 26392 32824 26444
rect 32956 26392 33008 26444
rect 34520 26392 34572 26444
rect 34704 26435 34756 26444
rect 34704 26401 34713 26435
rect 34713 26401 34747 26435
rect 34747 26401 34756 26435
rect 34704 26392 34756 26401
rect 25136 26256 25188 26308
rect 26148 26256 26200 26308
rect 26240 26256 26292 26308
rect 33876 26367 33928 26376
rect 33876 26333 33885 26367
rect 33885 26333 33919 26367
rect 33919 26333 33928 26367
rect 35348 26460 35400 26512
rect 33876 26324 33928 26333
rect 33784 26256 33836 26308
rect 35164 26364 35216 26376
rect 39672 26392 39724 26444
rect 40040 26435 40092 26444
rect 40040 26401 40049 26435
rect 40049 26401 40083 26435
rect 40083 26401 40092 26435
rect 40040 26392 40092 26401
rect 35164 26330 35173 26364
rect 35173 26330 35207 26364
rect 35207 26330 35216 26364
rect 35164 26324 35216 26330
rect 35808 26324 35860 26376
rect 36268 26324 36320 26376
rect 36452 26324 36504 26376
rect 37004 26324 37056 26376
rect 37464 26324 37516 26376
rect 38476 26324 38528 26376
rect 47492 26528 47544 26580
rect 45560 26460 45612 26512
rect 41512 26324 41564 26376
rect 46940 26324 46992 26376
rect 48136 26367 48188 26376
rect 48136 26333 48145 26367
rect 48145 26333 48179 26367
rect 48179 26333 48188 26367
rect 48136 26324 48188 26333
rect 41696 26299 41748 26308
rect 41696 26265 41705 26299
rect 41705 26265 41739 26299
rect 41739 26265 41748 26299
rect 41696 26256 41748 26265
rect 17592 26188 17644 26240
rect 25780 26188 25832 26240
rect 29736 26188 29788 26240
rect 31300 26188 31352 26240
rect 34704 26188 34756 26240
rect 35532 26188 35584 26240
rect 47308 26256 47360 26308
rect 47032 26188 47084 26240
rect 47860 26188 47912 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 2780 26027 2832 26036
rect 2780 25993 2789 26027
rect 2789 25993 2823 26027
rect 2823 25993 2832 26027
rect 2780 25984 2832 25993
rect 11796 25984 11848 26036
rect 47032 25984 47084 26036
rect 5264 25916 5316 25968
rect 23296 25916 23348 25968
rect 23480 25916 23532 25968
rect 29644 25959 29696 25968
rect 29644 25925 29653 25959
rect 29653 25925 29687 25959
rect 29687 25925 29696 25959
rect 29644 25916 29696 25925
rect 1400 25891 1452 25900
rect 1400 25857 1409 25891
rect 1409 25857 1443 25891
rect 1443 25857 1452 25891
rect 1400 25848 1452 25857
rect 2136 25848 2188 25900
rect 1676 25823 1728 25832
rect 1676 25789 1685 25823
rect 1685 25789 1719 25823
rect 1719 25789 1728 25823
rect 1676 25780 1728 25789
rect 16028 25848 16080 25900
rect 16212 25848 16264 25900
rect 16580 25848 16632 25900
rect 20352 25891 20404 25900
rect 20352 25857 20361 25891
rect 20361 25857 20395 25891
rect 20395 25857 20404 25891
rect 20352 25848 20404 25857
rect 20536 25891 20588 25900
rect 20536 25857 20545 25891
rect 20545 25857 20579 25891
rect 20579 25857 20588 25891
rect 20536 25848 20588 25857
rect 23388 25891 23440 25900
rect 23388 25857 23397 25891
rect 23397 25857 23431 25891
rect 23431 25857 23440 25891
rect 23388 25848 23440 25857
rect 24584 25848 24636 25900
rect 24952 25848 25004 25900
rect 29736 25848 29788 25900
rect 30288 25916 30340 25968
rect 30748 25959 30800 25968
rect 30748 25925 30757 25959
rect 30757 25925 30791 25959
rect 30791 25925 30800 25959
rect 30748 25916 30800 25925
rect 34060 25916 34112 25968
rect 35808 25916 35860 25968
rect 36084 25916 36136 25968
rect 17040 25780 17092 25832
rect 2504 25712 2556 25764
rect 30104 25780 30156 25832
rect 30288 25780 30340 25832
rect 32956 25848 33008 25900
rect 33140 25848 33192 25900
rect 33321 25891 33373 25900
rect 33321 25857 33330 25891
rect 33330 25857 33364 25891
rect 33364 25857 33373 25891
rect 33321 25848 33373 25857
rect 32772 25780 32824 25832
rect 33784 25848 33836 25900
rect 36636 25916 36688 25968
rect 45560 25916 45612 25968
rect 34520 25780 34572 25832
rect 35440 25780 35492 25832
rect 36544 25894 36596 25900
rect 36544 25860 36553 25894
rect 36553 25860 36587 25894
rect 36587 25860 36596 25894
rect 36544 25848 36596 25860
rect 36820 25848 36872 25900
rect 37004 25848 37056 25900
rect 42340 25848 42392 25900
rect 36636 25780 36688 25832
rect 36912 25780 36964 25832
rect 45744 25780 45796 25832
rect 46848 25823 46900 25832
rect 46848 25789 46857 25823
rect 46857 25789 46891 25823
rect 46891 25789 46900 25823
rect 46848 25780 46900 25789
rect 47492 25780 47544 25832
rect 47768 25780 47820 25832
rect 17224 25712 17276 25764
rect 15660 25644 15712 25696
rect 16212 25644 16264 25696
rect 21088 25712 21140 25764
rect 29000 25712 29052 25764
rect 30472 25712 30524 25764
rect 24860 25644 24912 25696
rect 25596 25644 25648 25696
rect 29736 25644 29788 25696
rect 33508 25644 33560 25696
rect 34520 25644 34572 25696
rect 34796 25644 34848 25696
rect 36360 25644 36412 25696
rect 47768 25687 47820 25696
rect 47768 25653 47777 25687
rect 47777 25653 47811 25687
rect 47811 25653 47820 25687
rect 47768 25644 47820 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 1676 25440 1728 25492
rect 2504 25372 2556 25424
rect 2872 25372 2924 25424
rect 11888 25440 11940 25492
rect 20168 25440 20220 25492
rect 20720 25483 20772 25492
rect 20720 25449 20729 25483
rect 20729 25449 20763 25483
rect 20763 25449 20772 25483
rect 20720 25440 20772 25449
rect 20904 25440 20956 25492
rect 18788 25304 18840 25356
rect 16580 25279 16632 25288
rect 16580 25245 16589 25279
rect 16589 25245 16623 25279
rect 16623 25245 16632 25279
rect 16580 25236 16632 25245
rect 17592 25279 17644 25288
rect 17592 25245 17601 25279
rect 17601 25245 17635 25279
rect 17635 25245 17644 25279
rect 17592 25236 17644 25245
rect 20076 25304 20128 25356
rect 20628 25304 20680 25356
rect 20812 25347 20864 25356
rect 20812 25313 20821 25347
rect 20821 25313 20855 25347
rect 20855 25313 20864 25347
rect 20812 25304 20864 25313
rect 19800 25236 19852 25288
rect 6828 25168 6880 25220
rect 16028 25168 16080 25220
rect 19340 25168 19392 25220
rect 20720 25211 20772 25220
rect 20720 25177 20729 25211
rect 20729 25177 20763 25211
rect 20763 25177 20772 25211
rect 20720 25168 20772 25177
rect 17408 25100 17460 25152
rect 20260 25100 20312 25152
rect 25596 25440 25648 25492
rect 25780 25440 25832 25492
rect 35532 25440 35584 25492
rect 35808 25483 35860 25492
rect 35808 25449 35817 25483
rect 35817 25449 35851 25483
rect 35851 25449 35860 25483
rect 35808 25440 35860 25449
rect 45744 25483 45796 25492
rect 21088 25372 21140 25424
rect 34520 25372 34572 25424
rect 24492 25304 24544 25356
rect 23296 25236 23348 25288
rect 26424 25304 26476 25356
rect 29000 25347 29052 25356
rect 29000 25313 29009 25347
rect 29009 25313 29043 25347
rect 29043 25313 29052 25347
rect 29000 25304 29052 25313
rect 30012 25304 30064 25356
rect 25688 25279 25740 25288
rect 25688 25245 25697 25279
rect 25697 25245 25731 25279
rect 25731 25245 25740 25279
rect 25688 25236 25740 25245
rect 26056 25236 26108 25288
rect 30472 25279 30524 25288
rect 30472 25245 30481 25279
rect 30481 25245 30515 25279
rect 30515 25245 30524 25279
rect 30472 25236 30524 25245
rect 27620 25168 27672 25220
rect 25596 25100 25648 25152
rect 26240 25100 26292 25152
rect 30012 25100 30064 25152
rect 30472 25100 30524 25152
rect 30840 25168 30892 25220
rect 31392 25211 31444 25220
rect 31392 25177 31401 25211
rect 31401 25177 31435 25211
rect 31435 25177 31444 25211
rect 31392 25168 31444 25177
rect 32128 25168 32180 25220
rect 33324 25168 33376 25220
rect 33600 25279 33652 25288
rect 33600 25245 33609 25279
rect 33609 25245 33643 25279
rect 33643 25245 33652 25279
rect 33600 25236 33652 25245
rect 33784 25279 33836 25288
rect 33784 25245 33793 25279
rect 33793 25245 33827 25279
rect 33827 25245 33836 25279
rect 36268 25279 36320 25288
rect 33784 25236 33836 25245
rect 36268 25245 36277 25279
rect 36277 25245 36311 25279
rect 36311 25245 36320 25279
rect 36268 25236 36320 25245
rect 36360 25236 36412 25288
rect 40500 25236 40552 25288
rect 45744 25449 45753 25483
rect 45753 25449 45787 25483
rect 45787 25449 45796 25483
rect 45744 25440 45796 25449
rect 47032 25440 47084 25492
rect 47860 25483 47912 25492
rect 40684 25372 40736 25424
rect 47400 25372 47452 25424
rect 47860 25449 47869 25483
rect 47869 25449 47903 25483
rect 47903 25449 47912 25483
rect 47860 25440 47912 25449
rect 41604 25236 41656 25288
rect 46204 25236 46256 25288
rect 46388 25236 46440 25288
rect 35440 25211 35492 25220
rect 35440 25177 35449 25211
rect 35449 25177 35483 25211
rect 35483 25177 35492 25211
rect 35440 25168 35492 25177
rect 34796 25100 34848 25152
rect 35808 25168 35860 25220
rect 37280 25100 37332 25152
rect 37648 25143 37700 25152
rect 37648 25109 37657 25143
rect 37657 25109 37691 25143
rect 37691 25109 37700 25143
rect 37648 25100 37700 25109
rect 40132 25143 40184 25152
rect 40132 25109 40141 25143
rect 40141 25109 40175 25143
rect 40175 25109 40184 25143
rect 40132 25100 40184 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 20536 24896 20588 24948
rect 20720 24896 20772 24948
rect 27988 24896 28040 24948
rect 29092 24896 29144 24948
rect 32772 24939 32824 24948
rect 32772 24905 32781 24939
rect 32781 24905 32815 24939
rect 32815 24905 32824 24939
rect 32772 24896 32824 24905
rect 2136 24803 2188 24812
rect 2136 24769 2145 24803
rect 2145 24769 2179 24803
rect 2179 24769 2188 24803
rect 2136 24760 2188 24769
rect 15660 24760 15712 24812
rect 16580 24760 16632 24812
rect 17500 24760 17552 24812
rect 17868 24760 17920 24812
rect 18788 24803 18840 24812
rect 18788 24769 18797 24803
rect 18797 24769 18831 24803
rect 18831 24769 18840 24803
rect 18788 24760 18840 24769
rect 20076 24828 20128 24880
rect 20260 24828 20312 24880
rect 20812 24828 20864 24880
rect 19984 24803 20036 24812
rect 1860 24692 1912 24744
rect 17316 24692 17368 24744
rect 19984 24769 19993 24803
rect 19993 24769 20027 24803
rect 20027 24769 20036 24803
rect 19984 24760 20036 24769
rect 20628 24803 20680 24812
rect 20628 24769 20637 24803
rect 20637 24769 20671 24803
rect 20671 24769 20680 24803
rect 20628 24760 20680 24769
rect 20720 24760 20772 24812
rect 21824 24760 21876 24812
rect 28448 24828 28500 24880
rect 30012 24828 30064 24880
rect 32220 24828 32272 24880
rect 33784 24896 33836 24948
rect 35900 24896 35952 24948
rect 40684 24896 40736 24948
rect 33508 24871 33560 24880
rect 33508 24837 33542 24871
rect 33542 24837 33560 24871
rect 33508 24828 33560 24837
rect 35532 24828 35584 24880
rect 36912 24828 36964 24880
rect 6736 24624 6788 24676
rect 19708 24624 19760 24676
rect 21088 24692 21140 24744
rect 23020 24803 23072 24812
rect 23020 24769 23029 24803
rect 23029 24769 23063 24803
rect 23063 24769 23072 24803
rect 23480 24803 23532 24812
rect 23020 24760 23072 24769
rect 23480 24769 23489 24803
rect 23489 24769 23523 24803
rect 23523 24769 23532 24803
rect 23480 24760 23532 24769
rect 25044 24760 25096 24812
rect 25228 24803 25280 24812
rect 25228 24769 25262 24803
rect 25262 24769 25280 24803
rect 27988 24803 28040 24812
rect 25228 24760 25280 24769
rect 27988 24769 27997 24803
rect 27997 24769 28031 24803
rect 28031 24769 28040 24803
rect 27988 24760 28040 24769
rect 23572 24692 23624 24744
rect 28540 24692 28592 24744
rect 29000 24692 29052 24744
rect 29644 24760 29696 24812
rect 30472 24803 30524 24812
rect 30472 24769 30506 24803
rect 30506 24769 30524 24803
rect 30472 24760 30524 24769
rect 30840 24760 30892 24812
rect 32404 24803 32456 24812
rect 32404 24769 32413 24803
rect 32413 24769 32447 24803
rect 32447 24769 32456 24803
rect 32404 24760 32456 24769
rect 33324 24760 33376 24812
rect 30104 24692 30156 24744
rect 30196 24735 30248 24744
rect 30196 24701 30205 24735
rect 30205 24701 30239 24735
rect 30239 24701 30248 24735
rect 30196 24692 30248 24701
rect 32680 24692 32732 24744
rect 34520 24760 34572 24812
rect 41052 24828 41104 24880
rect 40132 24760 40184 24812
rect 40224 24760 40276 24812
rect 41972 24760 42024 24812
rect 42432 24803 42484 24812
rect 1952 24556 2004 24608
rect 20260 24556 20312 24608
rect 21456 24556 21508 24608
rect 22560 24599 22612 24608
rect 22560 24565 22569 24599
rect 22569 24565 22603 24599
rect 22603 24565 22612 24599
rect 22560 24556 22612 24565
rect 22652 24556 22704 24608
rect 23388 24556 23440 24608
rect 23572 24599 23624 24608
rect 23572 24565 23581 24599
rect 23581 24565 23615 24599
rect 23615 24565 23624 24599
rect 23572 24556 23624 24565
rect 24676 24556 24728 24608
rect 26608 24556 26660 24608
rect 27252 24556 27304 24608
rect 28356 24556 28408 24608
rect 29368 24556 29420 24608
rect 29644 24624 29696 24676
rect 34704 24692 34756 24744
rect 36268 24692 36320 24744
rect 42432 24769 42441 24803
rect 42441 24769 42475 24803
rect 42475 24769 42484 24803
rect 42432 24760 42484 24769
rect 45192 24760 45244 24812
rect 47492 24760 47544 24812
rect 47860 24803 47912 24812
rect 47860 24769 47869 24803
rect 47869 24769 47903 24803
rect 47903 24769 47912 24803
rect 47860 24760 47912 24769
rect 31208 24556 31260 24608
rect 31392 24556 31444 24608
rect 38292 24624 38344 24676
rect 35348 24556 35400 24608
rect 39396 24556 39448 24608
rect 43444 24624 43496 24676
rect 41144 24556 41196 24608
rect 42340 24556 42392 24608
rect 46480 24556 46532 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 2320 24352 2372 24404
rect 1400 24191 1452 24200
rect 1400 24157 1409 24191
rect 1409 24157 1443 24191
rect 1443 24157 1452 24191
rect 1400 24148 1452 24157
rect 1676 24191 1728 24200
rect 1676 24157 1685 24191
rect 1685 24157 1719 24191
rect 1719 24157 1728 24191
rect 1676 24148 1728 24157
rect 1768 24148 1820 24200
rect 15752 24191 15804 24200
rect 15752 24157 15761 24191
rect 15761 24157 15795 24191
rect 15795 24157 15804 24191
rect 15752 24148 15804 24157
rect 19340 24284 19392 24336
rect 20352 24352 20404 24404
rect 20996 24352 21048 24404
rect 21180 24352 21232 24404
rect 21364 24352 21416 24404
rect 27988 24352 28040 24404
rect 28540 24395 28592 24404
rect 28540 24361 28549 24395
rect 28549 24361 28583 24395
rect 28583 24361 28592 24395
rect 28540 24352 28592 24361
rect 29092 24352 29144 24404
rect 36636 24352 36688 24404
rect 38752 24352 38804 24404
rect 41420 24352 41472 24404
rect 41972 24395 42024 24404
rect 20720 24284 20772 24336
rect 23388 24284 23440 24336
rect 25320 24284 25372 24336
rect 27436 24327 27488 24336
rect 27436 24293 27445 24327
rect 27445 24293 27479 24327
rect 27479 24293 27488 24327
rect 27436 24284 27488 24293
rect 17592 24216 17644 24268
rect 17868 24259 17920 24268
rect 17868 24225 17877 24259
rect 17877 24225 17911 24259
rect 17911 24225 17920 24259
rect 17868 24216 17920 24225
rect 19800 24259 19852 24268
rect 19800 24225 19809 24259
rect 19809 24225 19843 24259
rect 19843 24225 19852 24259
rect 19800 24216 19852 24225
rect 19892 24216 19944 24268
rect 20812 24259 20864 24268
rect 20812 24225 20821 24259
rect 20821 24225 20855 24259
rect 20855 24225 20864 24259
rect 20812 24216 20864 24225
rect 21916 24259 21968 24268
rect 21916 24225 21925 24259
rect 21925 24225 21959 24259
rect 21959 24225 21968 24259
rect 21916 24216 21968 24225
rect 27528 24259 27580 24268
rect 27528 24225 27537 24259
rect 27537 24225 27571 24259
rect 27571 24225 27580 24259
rect 27528 24216 27580 24225
rect 28356 24216 28408 24268
rect 16304 24055 16356 24064
rect 16304 24021 16313 24055
rect 16313 24021 16347 24055
rect 16347 24021 16356 24055
rect 16304 24012 16356 24021
rect 19340 24148 19392 24200
rect 20076 24148 20128 24200
rect 20904 24191 20956 24200
rect 20904 24157 20913 24191
rect 20913 24157 20947 24191
rect 20947 24157 20956 24191
rect 20904 24148 20956 24157
rect 18052 24080 18104 24132
rect 19432 24080 19484 24132
rect 20628 24123 20680 24132
rect 20628 24089 20637 24123
rect 20637 24089 20671 24123
rect 20671 24089 20680 24123
rect 20628 24080 20680 24089
rect 16948 24012 17000 24064
rect 21824 24148 21876 24200
rect 22560 24148 22612 24200
rect 24492 24191 24544 24200
rect 24492 24157 24501 24191
rect 24501 24157 24535 24191
rect 24535 24157 24544 24191
rect 24492 24148 24544 24157
rect 24676 24191 24728 24200
rect 24676 24157 24685 24191
rect 24685 24157 24719 24191
rect 24719 24157 24728 24191
rect 24676 24148 24728 24157
rect 25044 24148 25096 24200
rect 28264 24148 28316 24200
rect 28448 24148 28500 24200
rect 30104 24284 30156 24336
rect 29276 24216 29328 24268
rect 30564 24216 30616 24268
rect 32128 24284 32180 24336
rect 35716 24284 35768 24336
rect 40224 24284 40276 24336
rect 40500 24327 40552 24336
rect 40500 24293 40509 24327
rect 40509 24293 40543 24327
rect 40543 24293 40552 24327
rect 40500 24284 40552 24293
rect 40960 24327 41012 24336
rect 40960 24293 40969 24327
rect 40969 24293 41003 24327
rect 41003 24293 41012 24327
rect 40960 24284 41012 24293
rect 41972 24361 41981 24395
rect 41981 24361 42015 24395
rect 42015 24361 42024 24395
rect 41972 24352 42024 24361
rect 42064 24352 42116 24404
rect 43352 24284 43404 24336
rect 48044 24352 48096 24404
rect 32680 24216 32732 24268
rect 34704 24259 34756 24268
rect 34704 24225 34713 24259
rect 34713 24225 34747 24259
rect 34747 24225 34756 24259
rect 34704 24216 34756 24225
rect 25596 24123 25648 24132
rect 25596 24089 25630 24123
rect 25630 24089 25648 24123
rect 25596 24080 25648 24089
rect 23020 24012 23072 24064
rect 24308 24012 24360 24064
rect 25136 24012 25188 24064
rect 25320 24012 25372 24064
rect 27528 24080 27580 24132
rect 28080 24080 28132 24132
rect 26884 24012 26936 24064
rect 27712 24012 27764 24064
rect 29092 24080 29144 24132
rect 29552 24123 29604 24132
rect 29552 24089 29561 24123
rect 29561 24089 29595 24123
rect 29595 24089 29604 24123
rect 29552 24080 29604 24089
rect 30840 24123 30892 24132
rect 30840 24089 30849 24123
rect 30849 24089 30883 24123
rect 30883 24089 30892 24123
rect 30840 24080 30892 24089
rect 30932 24080 30984 24132
rect 31668 24123 31720 24132
rect 31668 24089 31677 24123
rect 31677 24089 31711 24123
rect 31711 24089 31720 24123
rect 31668 24080 31720 24089
rect 31852 24080 31904 24132
rect 29276 24012 29328 24064
rect 30472 24012 30524 24064
rect 32220 24148 32272 24200
rect 34796 24148 34848 24200
rect 35440 24148 35492 24200
rect 40868 24216 40920 24268
rect 41052 24216 41104 24268
rect 42156 24216 42208 24268
rect 47768 24284 47820 24336
rect 37372 24148 37424 24200
rect 37648 24148 37700 24200
rect 38108 24191 38160 24200
rect 38108 24157 38117 24191
rect 38117 24157 38151 24191
rect 38151 24157 38160 24191
rect 38108 24148 38160 24157
rect 39764 24148 39816 24200
rect 39856 24148 39908 24200
rect 41144 24191 41196 24200
rect 41144 24157 41153 24191
rect 41153 24157 41187 24191
rect 41187 24157 41196 24191
rect 41144 24148 41196 24157
rect 46480 24259 46532 24268
rect 46480 24225 46489 24259
rect 46489 24225 46523 24259
rect 46523 24225 46532 24259
rect 46480 24216 46532 24225
rect 48136 24259 48188 24268
rect 48136 24225 48145 24259
rect 48145 24225 48179 24259
rect 48179 24225 48188 24259
rect 48136 24216 48188 24225
rect 42892 24148 42944 24200
rect 43168 24191 43220 24200
rect 43168 24157 43177 24191
rect 43177 24157 43211 24191
rect 43211 24157 43220 24191
rect 43168 24148 43220 24157
rect 43352 24191 43404 24200
rect 43352 24157 43361 24191
rect 43361 24157 43395 24191
rect 43395 24157 43404 24191
rect 43352 24148 43404 24157
rect 43444 24148 43496 24200
rect 32864 24080 32916 24132
rect 40592 24080 40644 24132
rect 41420 24080 41472 24132
rect 42248 24080 42300 24132
rect 34796 24012 34848 24064
rect 36084 24055 36136 24064
rect 36084 24021 36093 24055
rect 36093 24021 36127 24055
rect 36127 24021 36136 24055
rect 36084 24012 36136 24021
rect 37280 24055 37332 24064
rect 37280 24021 37289 24055
rect 37289 24021 37323 24055
rect 37323 24021 37332 24055
rect 37280 24012 37332 24021
rect 37924 24012 37976 24064
rect 38844 24012 38896 24064
rect 39672 24012 39724 24064
rect 41788 24055 41840 24064
rect 41788 24021 41813 24055
rect 41813 24021 41840 24055
rect 41788 24012 41840 24021
rect 43260 24012 43312 24064
rect 47676 24080 47728 24132
rect 43812 24055 43864 24064
rect 43812 24021 43821 24055
rect 43821 24021 43855 24055
rect 43855 24021 43864 24055
rect 43812 24012 43864 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 15568 23808 15620 23860
rect 17316 23808 17368 23860
rect 20904 23808 20956 23860
rect 21088 23851 21140 23860
rect 21088 23817 21097 23851
rect 21097 23817 21131 23851
rect 21131 23817 21140 23851
rect 21088 23808 21140 23817
rect 25228 23808 25280 23860
rect 1952 23783 2004 23792
rect 1952 23749 1961 23783
rect 1961 23749 1995 23783
rect 1995 23749 2004 23783
rect 1952 23740 2004 23749
rect 15936 23783 15988 23792
rect 15936 23749 15945 23783
rect 15945 23749 15979 23783
rect 15979 23749 15988 23783
rect 15936 23740 15988 23749
rect 16028 23740 16080 23792
rect 1768 23715 1820 23724
rect 1768 23681 1777 23715
rect 1777 23681 1811 23715
rect 1811 23681 1820 23715
rect 1768 23672 1820 23681
rect 15660 23715 15712 23724
rect 15660 23681 15669 23715
rect 15669 23681 15703 23715
rect 15703 23681 15712 23715
rect 15660 23672 15712 23681
rect 15752 23672 15804 23724
rect 20352 23740 20404 23792
rect 25136 23740 25188 23792
rect 19892 23672 19944 23724
rect 1492 23604 1544 23656
rect 1952 23604 2004 23656
rect 2780 23647 2832 23656
rect 2780 23613 2789 23647
rect 2789 23613 2823 23647
rect 2823 23613 2832 23647
rect 2780 23604 2832 23613
rect 16488 23604 16540 23656
rect 17132 23647 17184 23656
rect 17132 23613 17141 23647
rect 17141 23613 17175 23647
rect 17175 23613 17184 23647
rect 17132 23604 17184 23613
rect 17500 23647 17552 23656
rect 17500 23613 17509 23647
rect 17509 23613 17543 23647
rect 17543 23613 17552 23647
rect 17500 23604 17552 23613
rect 19340 23604 19392 23656
rect 1676 23536 1728 23588
rect 19432 23536 19484 23588
rect 19708 23604 19760 23656
rect 20260 23672 20312 23724
rect 20720 23672 20772 23724
rect 20996 23672 21048 23724
rect 21916 23672 21968 23724
rect 23204 23672 23256 23724
rect 24308 23715 24360 23724
rect 24308 23681 24317 23715
rect 24317 23681 24351 23715
rect 24351 23681 24360 23715
rect 24308 23672 24360 23681
rect 23480 23604 23532 23656
rect 24676 23672 24728 23724
rect 25228 23715 25280 23724
rect 25228 23681 25237 23715
rect 25237 23681 25271 23715
rect 25271 23681 25280 23715
rect 25228 23672 25280 23681
rect 26240 23808 26292 23860
rect 26424 23851 26476 23860
rect 26424 23817 26433 23851
rect 26433 23817 26467 23851
rect 26467 23817 26476 23851
rect 26424 23808 26476 23817
rect 28080 23808 28132 23860
rect 29000 23808 29052 23860
rect 25780 23740 25832 23792
rect 26056 23715 26108 23724
rect 26056 23681 26065 23715
rect 26065 23681 26099 23715
rect 26099 23681 26108 23715
rect 26056 23672 26108 23681
rect 26884 23672 26936 23724
rect 28172 23715 28224 23724
rect 28172 23681 28181 23715
rect 28181 23681 28215 23715
rect 28215 23681 28224 23715
rect 28172 23672 28224 23681
rect 28540 23715 28592 23724
rect 28540 23681 28549 23715
rect 28549 23681 28583 23715
rect 28583 23681 28592 23715
rect 28540 23672 28592 23681
rect 30012 23740 30064 23792
rect 29368 23715 29420 23724
rect 29368 23681 29377 23715
rect 29377 23681 29411 23715
rect 29411 23681 29420 23715
rect 29368 23672 29420 23681
rect 29552 23715 29604 23724
rect 29552 23681 29561 23715
rect 29561 23681 29595 23715
rect 29595 23681 29604 23715
rect 31668 23740 31720 23792
rect 32864 23740 32916 23792
rect 33600 23808 33652 23860
rect 35808 23808 35860 23860
rect 38844 23851 38896 23860
rect 35716 23783 35768 23792
rect 35716 23749 35725 23783
rect 35725 23749 35759 23783
rect 35759 23749 35768 23783
rect 35716 23740 35768 23749
rect 36084 23740 36136 23792
rect 37280 23783 37332 23792
rect 37280 23749 37289 23783
rect 37289 23749 37323 23783
rect 37323 23749 37332 23783
rect 38844 23817 38853 23851
rect 38853 23817 38887 23851
rect 38887 23817 38896 23851
rect 38844 23808 38896 23817
rect 40868 23808 40920 23860
rect 37280 23740 37332 23749
rect 38384 23740 38436 23792
rect 30288 23715 30340 23724
rect 29552 23672 29604 23681
rect 30288 23681 30297 23715
rect 30297 23681 30331 23715
rect 30331 23681 30340 23715
rect 30288 23672 30340 23681
rect 32404 23672 32456 23724
rect 33048 23672 33100 23724
rect 35992 23672 36044 23724
rect 42340 23740 42392 23792
rect 42524 23808 42576 23860
rect 42984 23740 43036 23792
rect 43812 23740 43864 23792
rect 47952 23783 48004 23792
rect 47952 23749 47961 23783
rect 47961 23749 47995 23783
rect 47995 23749 48004 23783
rect 47952 23740 48004 23749
rect 27160 23604 27212 23656
rect 28080 23647 28132 23656
rect 28080 23613 28089 23647
rect 28089 23613 28123 23647
rect 28123 23613 28132 23647
rect 28080 23604 28132 23613
rect 21456 23536 21508 23588
rect 29000 23604 29052 23656
rect 29092 23604 29144 23656
rect 38568 23672 38620 23724
rect 39672 23715 39724 23724
rect 36544 23604 36596 23656
rect 39028 23647 39080 23656
rect 39028 23613 39037 23647
rect 39037 23613 39071 23647
rect 39071 23613 39080 23647
rect 39672 23681 39681 23715
rect 39681 23681 39715 23715
rect 39715 23681 39724 23715
rect 39672 23672 39724 23681
rect 40408 23672 40460 23724
rect 40592 23715 40644 23724
rect 40592 23681 40601 23715
rect 40601 23681 40635 23715
rect 40635 23681 40644 23715
rect 40592 23672 40644 23681
rect 39028 23604 39080 23613
rect 39856 23604 39908 23656
rect 40868 23672 40920 23724
rect 40960 23604 41012 23656
rect 41512 23604 41564 23656
rect 44456 23672 44508 23724
rect 41788 23647 41840 23656
rect 41788 23613 41797 23647
rect 41797 23613 41831 23647
rect 41831 23613 41840 23647
rect 41788 23604 41840 23613
rect 42432 23604 42484 23656
rect 1492 23468 1544 23520
rect 1860 23468 1912 23520
rect 3516 23468 3568 23520
rect 17868 23468 17920 23520
rect 19892 23511 19944 23520
rect 19892 23477 19901 23511
rect 19901 23477 19935 23511
rect 19935 23477 19944 23511
rect 19892 23468 19944 23477
rect 20076 23468 20128 23520
rect 29736 23579 29788 23588
rect 23756 23511 23808 23520
rect 23756 23477 23765 23511
rect 23765 23477 23799 23511
rect 23799 23477 23808 23511
rect 24400 23511 24452 23520
rect 23756 23468 23808 23477
rect 24400 23477 24409 23511
rect 24409 23477 24443 23511
rect 24443 23477 24452 23511
rect 24400 23468 24452 23477
rect 28448 23511 28500 23520
rect 28448 23477 28457 23511
rect 28457 23477 28491 23511
rect 28491 23477 28500 23511
rect 28448 23468 28500 23477
rect 29736 23545 29745 23579
rect 29745 23545 29779 23579
rect 29779 23545 29788 23579
rect 29736 23536 29788 23545
rect 30012 23536 30064 23588
rect 42800 23536 42852 23588
rect 30104 23468 30156 23520
rect 30564 23468 30616 23520
rect 36452 23511 36504 23520
rect 36452 23477 36461 23511
rect 36461 23477 36495 23511
rect 36495 23477 36504 23511
rect 36452 23468 36504 23477
rect 37464 23511 37516 23520
rect 37464 23477 37473 23511
rect 37473 23477 37507 23511
rect 37507 23477 37516 23511
rect 37464 23468 37516 23477
rect 37648 23511 37700 23520
rect 37648 23477 37657 23511
rect 37657 23477 37691 23511
rect 37691 23477 37700 23511
rect 37648 23468 37700 23477
rect 38476 23511 38528 23520
rect 38476 23477 38485 23511
rect 38485 23477 38519 23511
rect 38519 23477 38528 23511
rect 38476 23468 38528 23477
rect 38752 23468 38804 23520
rect 39672 23468 39724 23520
rect 41144 23468 41196 23520
rect 43904 23604 43956 23656
rect 47492 23604 47544 23656
rect 43996 23536 44048 23588
rect 44180 23468 44232 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 17592 23307 17644 23316
rect 17592 23273 17601 23307
rect 17601 23273 17635 23307
rect 17635 23273 17644 23307
rect 17592 23264 17644 23273
rect 18052 23264 18104 23316
rect 19708 23264 19760 23316
rect 20076 23264 20128 23316
rect 20260 23264 20312 23316
rect 20628 23264 20680 23316
rect 22652 23264 22704 23316
rect 23112 23264 23164 23316
rect 19892 23196 19944 23248
rect 28264 23196 28316 23248
rect 28724 23196 28776 23248
rect 19340 23128 19392 23180
rect 20628 23128 20680 23180
rect 30472 23264 30524 23316
rect 32496 23264 32548 23316
rect 33048 23264 33100 23316
rect 33324 23264 33376 23316
rect 35992 23264 36044 23316
rect 36544 23264 36596 23316
rect 38476 23264 38528 23316
rect 40500 23264 40552 23316
rect 40868 23264 40920 23316
rect 30012 23196 30064 23248
rect 30288 23196 30340 23248
rect 30932 23196 30984 23248
rect 16856 23060 16908 23112
rect 20168 23103 20220 23112
rect 16304 22992 16356 23044
rect 16764 22992 16816 23044
rect 20168 23069 20177 23103
rect 20177 23069 20211 23103
rect 20211 23069 20220 23103
rect 20168 23060 20220 23069
rect 20996 23060 21048 23112
rect 22928 23060 22980 23112
rect 23756 23060 23808 23112
rect 29552 23128 29604 23180
rect 35440 23128 35492 23180
rect 36176 23196 36228 23248
rect 36452 23128 36504 23180
rect 37648 23128 37700 23180
rect 29460 23060 29512 23112
rect 31944 23060 31996 23112
rect 34796 23060 34848 23112
rect 35808 23060 35860 23112
rect 19432 22992 19484 23044
rect 23296 23035 23348 23044
rect 23296 23001 23305 23035
rect 23305 23001 23339 23035
rect 23339 23001 23348 23035
rect 23296 22992 23348 23001
rect 24584 22992 24636 23044
rect 27804 22992 27856 23044
rect 31116 22992 31168 23044
rect 32036 22992 32088 23044
rect 18604 22924 18656 22976
rect 24952 22924 25004 22976
rect 27344 22924 27396 22976
rect 27712 22924 27764 22976
rect 28724 22924 28776 22976
rect 31392 22924 31444 22976
rect 32680 22924 32732 22976
rect 35716 22924 35768 22976
rect 36268 23060 36320 23112
rect 37556 23060 37608 23112
rect 38108 23196 38160 23248
rect 38476 23171 38528 23180
rect 38476 23137 38485 23171
rect 38485 23137 38519 23171
rect 38519 23137 38528 23171
rect 38476 23128 38528 23137
rect 39028 23196 39080 23248
rect 39764 23060 39816 23112
rect 40592 23128 40644 23180
rect 42156 23264 42208 23316
rect 45928 23264 45980 23316
rect 46940 23264 46992 23316
rect 42340 23171 42392 23180
rect 38108 22992 38160 23044
rect 41604 23103 41656 23112
rect 41604 23069 41613 23103
rect 41613 23069 41647 23103
rect 41647 23069 41656 23103
rect 41604 23060 41656 23069
rect 42340 23137 42349 23171
rect 42349 23137 42383 23171
rect 42383 23137 42392 23171
rect 42340 23128 42392 23137
rect 43996 23128 44048 23180
rect 42616 23103 42668 23112
rect 42616 23069 42625 23103
rect 42625 23069 42659 23103
rect 42659 23069 42668 23103
rect 42616 23060 42668 23069
rect 43352 23060 43404 23112
rect 42432 22992 42484 23044
rect 42892 22992 42944 23044
rect 45008 23060 45060 23112
rect 36176 22967 36228 22976
rect 36176 22933 36185 22967
rect 36185 22933 36219 22967
rect 36219 22933 36228 22967
rect 36176 22924 36228 22933
rect 37556 22967 37608 22976
rect 37556 22933 37565 22967
rect 37565 22933 37599 22967
rect 37599 22933 37608 22967
rect 37556 22924 37608 22933
rect 41972 22924 42024 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 17132 22720 17184 22772
rect 2044 22695 2096 22704
rect 2044 22661 2053 22695
rect 2053 22661 2087 22695
rect 2087 22661 2096 22695
rect 2044 22652 2096 22661
rect 18696 22720 18748 22772
rect 20536 22720 20588 22772
rect 24400 22720 24452 22772
rect 27804 22763 27856 22772
rect 27804 22729 27813 22763
rect 27813 22729 27847 22763
rect 27847 22729 27856 22763
rect 27804 22720 27856 22729
rect 18972 22652 19024 22704
rect 1860 22627 1912 22636
rect 1860 22593 1869 22627
rect 1869 22593 1903 22627
rect 1903 22593 1912 22627
rect 1860 22584 1912 22593
rect 3424 22627 3476 22636
rect 3424 22593 3433 22627
rect 3433 22593 3467 22627
rect 3467 22593 3476 22627
rect 3424 22584 3476 22593
rect 16580 22584 16632 22636
rect 13820 22516 13872 22568
rect 15200 22448 15252 22500
rect 18328 22584 18380 22636
rect 18512 22627 18564 22636
rect 18512 22593 18535 22627
rect 18535 22593 18564 22627
rect 18512 22584 18564 22593
rect 18696 22630 18748 22636
rect 18696 22596 18705 22630
rect 18705 22596 18739 22630
rect 18739 22596 18748 22630
rect 18880 22627 18932 22636
rect 18696 22584 18748 22596
rect 18880 22593 18889 22627
rect 18889 22593 18923 22627
rect 18923 22593 18932 22627
rect 18880 22584 18932 22593
rect 19248 22584 19300 22636
rect 19524 22584 19576 22636
rect 19892 22627 19944 22636
rect 19892 22593 19901 22627
rect 19901 22593 19935 22627
rect 19935 22593 19944 22627
rect 19892 22584 19944 22593
rect 18144 22516 18196 22568
rect 19432 22516 19484 22568
rect 18512 22448 18564 22500
rect 23572 22652 23624 22704
rect 24492 22652 24544 22704
rect 23204 22491 23256 22500
rect 23204 22457 23213 22491
rect 23213 22457 23247 22491
rect 23247 22457 23256 22491
rect 23204 22448 23256 22457
rect 23664 22584 23716 22636
rect 24860 22627 24912 22636
rect 24860 22593 24869 22627
rect 24869 22593 24903 22627
rect 24903 22593 24912 22627
rect 24860 22584 24912 22593
rect 25412 22652 25464 22704
rect 28080 22652 28132 22704
rect 25136 22584 25188 22636
rect 25688 22584 25740 22636
rect 27712 22584 27764 22636
rect 28724 22627 28776 22636
rect 28724 22593 28733 22627
rect 28733 22593 28767 22627
rect 28767 22593 28776 22627
rect 28724 22584 28776 22593
rect 29552 22584 29604 22636
rect 30932 22584 30984 22636
rect 31484 22652 31536 22704
rect 31392 22627 31444 22636
rect 31392 22593 31401 22627
rect 31401 22593 31435 22627
rect 31435 22593 31444 22627
rect 32864 22720 32916 22772
rect 33416 22720 33468 22772
rect 31668 22652 31720 22704
rect 31392 22584 31444 22593
rect 32496 22627 32548 22636
rect 32496 22593 32505 22627
rect 32505 22593 32539 22627
rect 32539 22593 32548 22627
rect 32496 22584 32548 22593
rect 33140 22652 33192 22704
rect 32680 22627 32732 22636
rect 32680 22593 32689 22627
rect 32689 22593 32723 22627
rect 32723 22593 32732 22627
rect 32680 22584 32732 22593
rect 32864 22627 32916 22636
rect 32864 22593 32873 22627
rect 32873 22593 32907 22627
rect 32907 22593 32916 22627
rect 32864 22584 32916 22593
rect 33324 22584 33376 22636
rect 37280 22720 37332 22772
rect 40316 22763 40368 22772
rect 40316 22729 40325 22763
rect 40325 22729 40359 22763
rect 40359 22729 40368 22763
rect 40316 22720 40368 22729
rect 40500 22763 40552 22772
rect 40500 22729 40509 22763
rect 40509 22729 40543 22763
rect 40543 22729 40552 22763
rect 40500 22720 40552 22729
rect 44456 22720 44508 22772
rect 40868 22652 40920 22704
rect 35808 22627 35860 22636
rect 23572 22516 23624 22568
rect 28632 22448 28684 22500
rect 32404 22516 32456 22568
rect 35808 22593 35817 22627
rect 35817 22593 35851 22627
rect 35851 22593 35860 22627
rect 35808 22584 35860 22593
rect 35992 22627 36044 22636
rect 35992 22593 36001 22627
rect 36001 22593 36035 22627
rect 36035 22593 36044 22627
rect 35992 22584 36044 22593
rect 36176 22584 36228 22636
rect 36820 22584 36872 22636
rect 37096 22516 37148 22568
rect 38384 22627 38436 22636
rect 38384 22593 38393 22627
rect 38393 22593 38427 22627
rect 38427 22593 38436 22627
rect 38384 22584 38436 22593
rect 41604 22652 41656 22704
rect 32128 22448 32180 22500
rect 32496 22448 32548 22500
rect 3516 22423 3568 22432
rect 3516 22389 3525 22423
rect 3525 22389 3559 22423
rect 3559 22389 3568 22423
rect 3516 22380 3568 22389
rect 18236 22423 18288 22432
rect 18236 22389 18245 22423
rect 18245 22389 18279 22423
rect 18279 22389 18288 22423
rect 18236 22380 18288 22389
rect 19340 22380 19392 22432
rect 20076 22380 20128 22432
rect 20536 22380 20588 22432
rect 24952 22380 25004 22432
rect 28080 22380 28132 22432
rect 28356 22380 28408 22432
rect 30932 22423 30984 22432
rect 30932 22389 30941 22423
rect 30941 22389 30975 22423
rect 30975 22389 30984 22423
rect 30932 22380 30984 22389
rect 32220 22423 32272 22432
rect 32220 22389 32229 22423
rect 32229 22389 32263 22423
rect 32263 22389 32272 22423
rect 32220 22380 32272 22389
rect 33324 22423 33376 22432
rect 33324 22389 33333 22423
rect 33333 22389 33367 22423
rect 33367 22389 33376 22423
rect 33324 22380 33376 22389
rect 36084 22448 36136 22500
rect 37464 22448 37516 22500
rect 38476 22516 38528 22568
rect 43076 22584 43128 22636
rect 44088 22584 44140 22636
rect 46848 22584 46900 22636
rect 47952 22627 48004 22636
rect 47952 22593 47961 22627
rect 47961 22593 47995 22627
rect 47995 22593 48004 22627
rect 47952 22584 48004 22593
rect 38108 22491 38160 22500
rect 38108 22457 38117 22491
rect 38117 22457 38151 22491
rect 38151 22457 38160 22491
rect 38108 22448 38160 22457
rect 40868 22448 40920 22500
rect 41328 22516 41380 22568
rect 42432 22516 42484 22568
rect 42616 22559 42668 22568
rect 42616 22525 42625 22559
rect 42625 22525 42659 22559
rect 42659 22525 42668 22559
rect 42616 22516 42668 22525
rect 42340 22448 42392 22500
rect 36176 22423 36228 22432
rect 36176 22389 36185 22423
rect 36185 22389 36219 22423
rect 36219 22389 36228 22423
rect 36176 22380 36228 22389
rect 37372 22423 37424 22432
rect 37372 22389 37381 22423
rect 37381 22389 37415 22423
rect 37415 22389 37424 22423
rect 37372 22380 37424 22389
rect 37648 22423 37700 22432
rect 37648 22389 37657 22423
rect 37657 22389 37691 22423
rect 37691 22389 37700 22423
rect 37648 22380 37700 22389
rect 40684 22423 40736 22432
rect 40684 22389 40693 22423
rect 40693 22389 40727 22423
rect 40727 22389 40736 22423
rect 40684 22380 40736 22389
rect 40960 22380 41012 22432
rect 42432 22423 42484 22432
rect 42432 22389 42441 22423
rect 42441 22389 42475 22423
rect 42475 22389 42484 22423
rect 42432 22380 42484 22389
rect 42524 22380 42576 22432
rect 45468 22380 45520 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 2872 22040 2924 22092
rect 18512 22176 18564 22228
rect 18328 22108 18380 22160
rect 15476 22083 15528 22092
rect 15476 22049 15485 22083
rect 15485 22049 15519 22083
rect 15519 22049 15528 22083
rect 15476 22040 15528 22049
rect 18144 22040 18196 22092
rect 18420 22040 18472 22092
rect 3424 21972 3476 22024
rect 3792 22015 3844 22024
rect 3792 21981 3801 22015
rect 3801 21981 3835 22015
rect 3835 21981 3844 22015
rect 3792 21972 3844 21981
rect 16856 22015 16908 22024
rect 16856 21981 16865 22015
rect 16865 21981 16899 22015
rect 16899 21981 16908 22015
rect 16856 21972 16908 21981
rect 17408 21972 17460 22024
rect 13912 21904 13964 21956
rect 18236 21972 18288 22024
rect 18696 21904 18748 21956
rect 21824 22040 21876 22092
rect 22100 22040 22152 22092
rect 25044 22176 25096 22228
rect 25412 22176 25464 22228
rect 27344 22176 27396 22228
rect 30656 22176 30708 22228
rect 32036 22176 32088 22228
rect 41328 22176 41380 22228
rect 42064 22219 42116 22228
rect 42064 22185 42073 22219
rect 42073 22185 42107 22219
rect 42107 22185 42116 22219
rect 42064 22176 42116 22185
rect 30380 22108 30432 22160
rect 31576 22108 31628 22160
rect 25688 22040 25740 22092
rect 27344 22015 27396 22024
rect 18512 21836 18564 21888
rect 20536 21904 20588 21956
rect 20720 21904 20772 21956
rect 23572 21904 23624 21956
rect 24952 21947 25004 21956
rect 24952 21913 24986 21947
rect 24986 21913 25004 21947
rect 24952 21904 25004 21913
rect 27344 21981 27353 22015
rect 27353 21981 27387 22015
rect 27387 21981 27396 22015
rect 27344 21972 27396 21981
rect 27528 21972 27580 22024
rect 28816 22040 28868 22092
rect 36820 22083 36872 22092
rect 36820 22049 36829 22083
rect 36829 22049 36863 22083
rect 36863 22049 36872 22083
rect 36820 22040 36872 22049
rect 37188 22040 37240 22092
rect 43444 22108 43496 22160
rect 28172 22015 28224 22024
rect 28172 21981 28181 22015
rect 28181 21981 28215 22015
rect 28215 21981 28224 22015
rect 28172 21972 28224 21981
rect 28264 21972 28316 22024
rect 31024 21972 31076 22024
rect 32588 21972 32640 22024
rect 34704 21972 34756 22024
rect 36176 22015 36228 22024
rect 36176 21981 36185 22015
rect 36185 21981 36219 22015
rect 36219 21981 36228 22015
rect 36176 21972 36228 21981
rect 36268 21972 36320 22024
rect 37832 21972 37884 22024
rect 40500 21972 40552 22024
rect 41144 22015 41196 22024
rect 41144 21981 41153 22015
rect 41153 21981 41187 22015
rect 41187 21981 41196 22015
rect 41144 21972 41196 21981
rect 30472 21947 30524 21956
rect 19984 21836 20036 21888
rect 25688 21836 25740 21888
rect 27436 21836 27488 21888
rect 28172 21836 28224 21888
rect 29000 21836 29052 21888
rect 30472 21913 30481 21947
rect 30481 21913 30515 21947
rect 30515 21913 30524 21947
rect 30472 21904 30524 21913
rect 32220 21904 32272 21956
rect 44180 22040 44232 22092
rect 42524 21972 42576 22024
rect 42616 21972 42668 22024
rect 43352 22015 43404 22024
rect 43352 21981 43361 22015
rect 43361 21981 43395 22015
rect 43395 21981 43404 22015
rect 43352 21972 43404 21981
rect 43444 22015 43496 22024
rect 43444 21981 43458 22015
rect 43458 21981 43492 22015
rect 43492 21981 43496 22015
rect 43444 21972 43496 21981
rect 41420 21904 41472 21956
rect 41788 21904 41840 21956
rect 41972 21904 42024 21956
rect 42432 21904 42484 21956
rect 44456 21904 44508 21956
rect 47952 21947 48004 21956
rect 47952 21913 47961 21947
rect 47961 21913 47995 21947
rect 47995 21913 48004 21947
rect 47952 21904 48004 21913
rect 36360 21879 36412 21888
rect 36360 21845 36369 21879
rect 36369 21845 36403 21879
rect 36403 21845 36412 21879
rect 36360 21836 36412 21845
rect 43628 21836 43680 21888
rect 46112 21836 46164 21888
rect 46480 21879 46532 21888
rect 46480 21845 46489 21879
rect 46489 21845 46523 21879
rect 46523 21845 46532 21879
rect 46480 21836 46532 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 3792 21632 3844 21684
rect 13728 21632 13780 21684
rect 13912 21675 13964 21684
rect 13912 21641 13921 21675
rect 13921 21641 13955 21675
rect 13955 21641 13964 21675
rect 13912 21632 13964 21641
rect 3516 21607 3568 21616
rect 3516 21573 3525 21607
rect 3525 21573 3559 21607
rect 3559 21573 3568 21607
rect 3516 21564 3568 21573
rect 24952 21632 25004 21684
rect 2504 21496 2556 21548
rect 16580 21564 16632 21616
rect 18328 21564 18380 21616
rect 18696 21564 18748 21616
rect 19340 21564 19392 21616
rect 30656 21632 30708 21684
rect 30748 21632 30800 21684
rect 31116 21632 31168 21684
rect 33048 21632 33100 21684
rect 36176 21632 36228 21684
rect 36360 21632 36412 21684
rect 13820 21539 13872 21548
rect 13820 21505 13829 21539
rect 13829 21505 13863 21539
rect 13863 21505 13872 21539
rect 13820 21496 13872 21505
rect 14924 21539 14976 21548
rect 14924 21505 14933 21539
rect 14933 21505 14967 21539
rect 14967 21505 14976 21539
rect 14924 21496 14976 21505
rect 17408 21496 17460 21548
rect 5172 21471 5224 21480
rect 5172 21437 5181 21471
rect 5181 21437 5215 21471
rect 5215 21437 5224 21471
rect 5172 21428 5224 21437
rect 15476 21428 15528 21480
rect 21640 21496 21692 21548
rect 21732 21496 21784 21548
rect 21916 21496 21968 21548
rect 13728 21360 13780 21412
rect 18328 21335 18380 21344
rect 18328 21301 18337 21335
rect 18337 21301 18371 21335
rect 18371 21301 18380 21335
rect 18328 21292 18380 21301
rect 20536 21360 20588 21412
rect 23572 21496 23624 21548
rect 24124 21539 24176 21548
rect 24124 21505 24133 21539
rect 24133 21505 24167 21539
rect 24167 21505 24176 21539
rect 25044 21539 25096 21548
rect 24124 21496 24176 21505
rect 25044 21505 25053 21539
rect 25053 21505 25087 21539
rect 25087 21505 25096 21539
rect 25044 21496 25096 21505
rect 25320 21539 25372 21548
rect 25320 21505 25354 21539
rect 25354 21505 25372 21539
rect 25320 21496 25372 21505
rect 27436 21496 27488 21548
rect 28540 21496 28592 21548
rect 28724 21496 28776 21548
rect 29552 21496 29604 21548
rect 30196 21564 30248 21616
rect 30932 21564 30984 21616
rect 32128 21496 32180 21548
rect 38292 21564 38344 21616
rect 33140 21539 33192 21548
rect 33140 21505 33149 21539
rect 33149 21505 33183 21539
rect 33183 21505 33192 21539
rect 33140 21496 33192 21505
rect 33232 21539 33284 21548
rect 33232 21505 33241 21539
rect 33241 21505 33275 21539
rect 33275 21505 33284 21539
rect 33232 21496 33284 21505
rect 33416 21539 33468 21548
rect 33416 21505 33425 21539
rect 33425 21505 33459 21539
rect 33459 21505 33468 21539
rect 33416 21496 33468 21505
rect 37832 21496 37884 21548
rect 40776 21632 40828 21684
rect 42432 21632 42484 21684
rect 46848 21675 46900 21684
rect 46848 21641 46857 21675
rect 46857 21641 46891 21675
rect 46891 21641 46900 21675
rect 46848 21632 46900 21641
rect 41328 21564 41380 21616
rect 23848 21360 23900 21412
rect 23296 21292 23348 21344
rect 23480 21292 23532 21344
rect 26240 21292 26292 21344
rect 27160 21292 27212 21344
rect 32772 21428 32824 21480
rect 38016 21428 38068 21480
rect 40868 21496 40920 21548
rect 40224 21428 40276 21480
rect 43628 21496 43680 21548
rect 45744 21539 45796 21548
rect 45744 21505 45778 21539
rect 45778 21505 45796 21539
rect 45744 21496 45796 21505
rect 35348 21360 35400 21412
rect 37740 21360 37792 21412
rect 40684 21360 40736 21412
rect 29552 21335 29604 21344
rect 29552 21301 29561 21335
rect 29561 21301 29595 21335
rect 29595 21301 29604 21335
rect 29552 21292 29604 21301
rect 31944 21292 31996 21344
rect 34796 21292 34848 21344
rect 37280 21292 37332 21344
rect 37832 21335 37884 21344
rect 37832 21301 37841 21335
rect 37841 21301 37875 21335
rect 37875 21301 37884 21335
rect 37832 21292 37884 21301
rect 38016 21335 38068 21344
rect 38016 21301 38025 21335
rect 38025 21301 38059 21335
rect 38059 21301 38068 21335
rect 38016 21292 38068 21301
rect 38936 21292 38988 21344
rect 40408 21292 40460 21344
rect 40960 21335 41012 21344
rect 40960 21301 40969 21335
rect 40969 21301 41003 21335
rect 41003 21301 41012 21335
rect 40960 21292 41012 21301
rect 41880 21292 41932 21344
rect 44916 21335 44968 21344
rect 44916 21301 44925 21335
rect 44925 21301 44959 21335
rect 44959 21301 44968 21335
rect 44916 21292 44968 21301
rect 47768 21335 47820 21344
rect 47768 21301 47777 21335
rect 47777 21301 47811 21335
rect 47811 21301 47820 21335
rect 47768 21292 47820 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 19340 21088 19392 21140
rect 15660 21020 15712 21072
rect 18052 21020 18104 21072
rect 18880 21020 18932 21072
rect 21916 21131 21968 21140
rect 21916 21097 21925 21131
rect 21925 21097 21959 21131
rect 21959 21097 21968 21131
rect 21916 21088 21968 21097
rect 33048 21088 33100 21140
rect 33140 21088 33192 21140
rect 37556 21088 37608 21140
rect 37740 21131 37792 21140
rect 37740 21097 37749 21131
rect 37749 21097 37783 21131
rect 37783 21097 37792 21131
rect 37740 21088 37792 21097
rect 38292 21088 38344 21140
rect 40132 21088 40184 21140
rect 43444 21088 43496 21140
rect 45744 21088 45796 21140
rect 3424 20952 3476 21004
rect 14924 20927 14976 20936
rect 14924 20893 14933 20927
rect 14933 20893 14967 20927
rect 14967 20893 14976 20927
rect 14924 20884 14976 20893
rect 2412 20748 2464 20800
rect 15660 20816 15712 20868
rect 17408 20884 17460 20936
rect 19984 20952 20036 21004
rect 16212 20859 16264 20868
rect 16212 20825 16221 20859
rect 16221 20825 16255 20859
rect 16255 20825 16264 20859
rect 16212 20816 16264 20825
rect 18328 20859 18380 20868
rect 18328 20825 18337 20859
rect 18337 20825 18371 20859
rect 18371 20825 18380 20859
rect 18328 20816 18380 20825
rect 18972 20816 19024 20868
rect 20536 20884 20588 20936
rect 22100 20927 22152 20936
rect 22100 20893 22109 20927
rect 22109 20893 22143 20927
rect 22143 20893 22152 20927
rect 22284 20927 22336 20936
rect 22100 20884 22152 20893
rect 22284 20893 22293 20927
rect 22293 20893 22327 20927
rect 22327 20893 22336 20927
rect 22284 20884 22336 20893
rect 25320 21020 25372 21072
rect 23388 20995 23440 21004
rect 23388 20961 23397 20995
rect 23397 20961 23431 20995
rect 23431 20961 23440 20995
rect 23388 20952 23440 20961
rect 23572 20952 23624 21004
rect 24124 20952 24176 21004
rect 27160 21020 27212 21072
rect 27528 21020 27580 21072
rect 36176 21020 36228 21072
rect 37924 21020 37976 21072
rect 17408 20748 17460 20800
rect 18696 20791 18748 20800
rect 18696 20757 18705 20791
rect 18705 20757 18739 20791
rect 18739 20757 18748 20791
rect 18696 20748 18748 20757
rect 23020 20816 23072 20868
rect 23296 20859 23348 20868
rect 23296 20825 23305 20859
rect 23305 20825 23339 20859
rect 23339 20825 23348 20859
rect 23296 20816 23348 20825
rect 23112 20748 23164 20800
rect 23848 20816 23900 20868
rect 24860 20884 24912 20936
rect 25412 20927 25464 20936
rect 25412 20893 25421 20927
rect 25421 20893 25455 20927
rect 25455 20893 25464 20927
rect 25412 20884 25464 20893
rect 25596 20884 25648 20936
rect 26148 20927 26200 20936
rect 26148 20893 26157 20927
rect 26157 20893 26191 20927
rect 26191 20893 26200 20927
rect 26148 20884 26200 20893
rect 26424 20884 26476 20936
rect 28356 20927 28408 20936
rect 28356 20893 28365 20927
rect 28365 20893 28399 20927
rect 28399 20893 28408 20927
rect 28356 20884 28408 20893
rect 28540 20927 28592 20936
rect 28540 20893 28549 20927
rect 28549 20893 28583 20927
rect 28583 20893 28592 20927
rect 28540 20884 28592 20893
rect 31760 20952 31812 21004
rect 32772 20995 32824 21004
rect 32772 20961 32781 20995
rect 32781 20961 32815 20995
rect 32815 20961 32824 20995
rect 32772 20952 32824 20961
rect 31300 20884 31352 20936
rect 31668 20927 31720 20936
rect 31668 20893 31677 20927
rect 31677 20893 31711 20927
rect 31711 20893 31720 20927
rect 31668 20884 31720 20893
rect 33324 20884 33376 20936
rect 26240 20816 26292 20868
rect 23572 20748 23624 20800
rect 24952 20748 25004 20800
rect 29000 20748 29052 20800
rect 29920 20816 29972 20868
rect 30380 20816 30432 20868
rect 31208 20816 31260 20868
rect 36268 20952 36320 21004
rect 38016 20952 38068 21004
rect 43352 21020 43404 21072
rect 45376 21020 45428 21072
rect 45468 21020 45520 21072
rect 34796 20884 34848 20936
rect 35348 20884 35400 20936
rect 38108 20927 38160 20936
rect 38108 20893 38117 20927
rect 38117 20893 38151 20927
rect 38151 20893 38160 20927
rect 38108 20884 38160 20893
rect 40408 20884 40460 20936
rect 45008 20952 45060 21004
rect 41880 20927 41932 20936
rect 41880 20893 41889 20927
rect 41889 20893 41923 20927
rect 41923 20893 41932 20927
rect 41880 20884 41932 20893
rect 44088 20927 44140 20936
rect 44088 20893 44097 20927
rect 44097 20893 44131 20927
rect 44131 20893 44140 20927
rect 44088 20884 44140 20893
rect 46848 20952 46900 21004
rect 46940 20995 46992 21004
rect 46940 20961 46949 20995
rect 46949 20961 46983 20995
rect 46983 20961 46992 20995
rect 46940 20952 46992 20961
rect 45373 20924 45425 20933
rect 45373 20890 45400 20924
rect 45400 20890 45425 20924
rect 45373 20881 45425 20890
rect 45652 20927 45704 20936
rect 45652 20893 45661 20927
rect 45661 20893 45695 20927
rect 45695 20893 45704 20927
rect 45652 20884 45704 20893
rect 30748 20748 30800 20800
rect 30932 20791 30984 20800
rect 30932 20757 30941 20791
rect 30941 20757 30975 20791
rect 30975 20757 30984 20791
rect 30932 20748 30984 20757
rect 33140 20748 33192 20800
rect 37372 20791 37424 20800
rect 37372 20757 37381 20791
rect 37381 20757 37415 20791
rect 37415 20757 37424 20791
rect 37372 20748 37424 20757
rect 38016 20791 38068 20800
rect 38016 20757 38025 20791
rect 38025 20757 38059 20791
rect 38059 20757 38068 20791
rect 38016 20748 38068 20757
rect 40224 20816 40276 20868
rect 44916 20816 44968 20868
rect 47676 20816 47728 20868
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 2136 20340 2188 20392
rect 11888 20383 11940 20392
rect 11888 20349 11897 20383
rect 11897 20349 11931 20383
rect 11931 20349 11940 20383
rect 11888 20340 11940 20349
rect 2780 20272 2832 20324
rect 5172 20272 5224 20324
rect 20 20204 72 20256
rect 16212 20544 16264 20596
rect 16580 20544 16632 20596
rect 15200 20408 15252 20460
rect 16580 20408 16632 20460
rect 16672 20451 16724 20460
rect 16672 20417 16681 20451
rect 16681 20417 16715 20451
rect 16715 20417 16724 20451
rect 16672 20408 16724 20417
rect 15936 20383 15988 20392
rect 15936 20349 15945 20383
rect 15945 20349 15979 20383
rect 15979 20349 15988 20383
rect 15936 20340 15988 20349
rect 16764 20340 16816 20392
rect 18788 20544 18840 20596
rect 18972 20544 19024 20596
rect 22100 20544 22152 20596
rect 22560 20476 22612 20528
rect 25136 20544 25188 20596
rect 25320 20544 25372 20596
rect 29736 20544 29788 20596
rect 29920 20587 29972 20596
rect 29920 20553 29929 20587
rect 29929 20553 29963 20587
rect 29963 20553 29972 20587
rect 29920 20544 29972 20553
rect 18880 20408 18932 20460
rect 18696 20340 18748 20392
rect 18972 20340 19024 20392
rect 13820 20272 13872 20324
rect 26148 20476 26200 20528
rect 23480 20408 23532 20460
rect 23572 20408 23624 20460
rect 24952 20408 25004 20460
rect 25136 20408 25188 20460
rect 25688 20408 25740 20460
rect 29460 20476 29512 20528
rect 31668 20544 31720 20596
rect 35624 20544 35676 20596
rect 38016 20544 38068 20596
rect 44088 20544 44140 20596
rect 44456 20587 44508 20596
rect 44456 20553 44465 20587
rect 44465 20553 44499 20587
rect 44499 20553 44508 20587
rect 44456 20544 44508 20553
rect 47676 20587 47728 20596
rect 47676 20553 47685 20587
rect 47685 20553 47719 20587
rect 47719 20553 47728 20587
rect 47676 20544 47728 20553
rect 40132 20519 40184 20528
rect 29552 20408 29604 20460
rect 30196 20451 30248 20460
rect 30196 20417 30205 20451
rect 30205 20417 30239 20451
rect 30239 20417 30248 20451
rect 30196 20408 30248 20417
rect 30380 20451 30432 20460
rect 30380 20417 30389 20451
rect 30389 20417 30423 20451
rect 30423 20417 30432 20451
rect 30380 20408 30432 20417
rect 30564 20451 30616 20460
rect 30564 20417 30573 20451
rect 30573 20417 30607 20451
rect 30607 20417 30616 20451
rect 30564 20408 30616 20417
rect 22928 20383 22980 20392
rect 22928 20349 22937 20383
rect 22937 20349 22971 20383
rect 22971 20349 22980 20383
rect 22928 20340 22980 20349
rect 23112 20383 23164 20392
rect 23112 20349 23121 20383
rect 23121 20349 23155 20383
rect 23155 20349 23164 20383
rect 23112 20340 23164 20349
rect 23296 20340 23348 20392
rect 17592 20204 17644 20256
rect 17960 20247 18012 20256
rect 17960 20213 17969 20247
rect 17969 20213 18003 20247
rect 18003 20213 18012 20247
rect 17960 20204 18012 20213
rect 20536 20272 20588 20324
rect 21916 20272 21968 20324
rect 33140 20340 33192 20392
rect 33968 20383 34020 20392
rect 33968 20349 33977 20383
rect 33977 20349 34011 20383
rect 34011 20349 34020 20383
rect 33968 20340 34020 20349
rect 36176 20340 36228 20392
rect 36544 20451 36596 20460
rect 36544 20417 36553 20451
rect 36553 20417 36587 20451
rect 36587 20417 36596 20451
rect 40132 20485 40141 20519
rect 40141 20485 40175 20519
rect 40175 20485 40184 20519
rect 40132 20476 40184 20485
rect 40868 20476 40920 20528
rect 36544 20408 36596 20417
rect 37280 20340 37332 20392
rect 24492 20272 24544 20324
rect 29276 20272 29328 20324
rect 30564 20272 30616 20324
rect 31484 20272 31536 20324
rect 36544 20272 36596 20324
rect 38108 20340 38160 20392
rect 41328 20408 41380 20460
rect 42156 20408 42208 20460
rect 42708 20408 42760 20460
rect 41788 20340 41840 20392
rect 40500 20272 40552 20324
rect 40960 20272 41012 20324
rect 45192 20408 45244 20460
rect 46480 20408 46532 20460
rect 46848 20451 46900 20460
rect 46848 20417 46857 20451
rect 46857 20417 46891 20451
rect 46891 20417 46900 20451
rect 46848 20408 46900 20417
rect 47308 20408 47360 20460
rect 45652 20340 45704 20392
rect 45376 20272 45428 20324
rect 22100 20204 22152 20256
rect 24308 20204 24360 20256
rect 27344 20204 27396 20256
rect 29736 20204 29788 20256
rect 31300 20204 31352 20256
rect 34152 20204 34204 20256
rect 37096 20204 37148 20256
rect 37464 20204 37516 20256
rect 38384 20204 38436 20256
rect 40868 20204 40920 20256
rect 43168 20204 43220 20256
rect 47032 20204 47084 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 11888 20043 11940 20052
rect 11888 20009 11897 20043
rect 11897 20009 11931 20043
rect 11931 20009 11940 20043
rect 11888 20000 11940 20009
rect 17408 20000 17460 20052
rect 17592 20000 17644 20052
rect 21916 20000 21968 20052
rect 17224 19932 17276 19984
rect 18236 19932 18288 19984
rect 18512 19932 18564 19984
rect 21732 19932 21784 19984
rect 22560 20000 22612 20052
rect 22744 20000 22796 20052
rect 23296 20000 23348 20052
rect 23388 20000 23440 20052
rect 26424 20000 26476 20052
rect 29092 20000 29144 20052
rect 30380 20000 30432 20052
rect 32404 20000 32456 20052
rect 37648 20000 37700 20052
rect 39396 20000 39448 20052
rect 40408 20000 40460 20052
rect 41144 20000 41196 20052
rect 22192 19932 22244 19984
rect 46848 19932 46900 19984
rect 10784 19796 10836 19848
rect 13820 19796 13872 19848
rect 15752 19839 15804 19848
rect 15752 19805 15761 19839
rect 15761 19805 15795 19839
rect 15795 19805 15804 19839
rect 15752 19796 15804 19805
rect 17960 19796 18012 19848
rect 18788 19864 18840 19916
rect 19340 19864 19392 19916
rect 18052 19660 18104 19712
rect 18420 19839 18472 19848
rect 18420 19805 18434 19839
rect 18434 19805 18468 19839
rect 18468 19805 18472 19839
rect 18420 19796 18472 19805
rect 18880 19796 18932 19848
rect 19156 19796 19208 19848
rect 20720 19796 20772 19848
rect 22100 19796 22152 19848
rect 26608 19907 26660 19916
rect 26608 19873 26617 19907
rect 26617 19873 26651 19907
rect 26651 19873 26660 19907
rect 26608 19864 26660 19873
rect 37280 19864 37332 19916
rect 38752 19864 38804 19916
rect 40868 19907 40920 19916
rect 40868 19873 40877 19907
rect 40877 19873 40911 19907
rect 40911 19873 40920 19907
rect 40868 19864 40920 19873
rect 21916 19728 21968 19780
rect 22376 19728 22428 19780
rect 22836 19796 22888 19848
rect 26148 19796 26200 19848
rect 31944 19839 31996 19848
rect 25780 19728 25832 19780
rect 31944 19805 31953 19839
rect 31953 19805 31987 19839
rect 31987 19805 31996 19839
rect 31944 19796 31996 19805
rect 33140 19796 33192 19848
rect 36176 19796 36228 19848
rect 37004 19839 37056 19848
rect 37004 19805 37013 19839
rect 37013 19805 37047 19839
rect 37047 19805 37056 19839
rect 37004 19796 37056 19805
rect 38476 19796 38528 19848
rect 45100 19864 45152 19916
rect 47768 19864 47820 19916
rect 41052 19839 41104 19848
rect 41052 19805 41061 19839
rect 41061 19805 41095 19839
rect 41095 19805 41104 19839
rect 48136 19839 48188 19848
rect 41052 19796 41104 19805
rect 48136 19805 48145 19839
rect 48145 19805 48179 19839
rect 48179 19805 48188 19839
rect 48136 19796 48188 19805
rect 26792 19728 26844 19780
rect 28264 19728 28316 19780
rect 28724 19728 28776 19780
rect 30932 19728 30984 19780
rect 31024 19771 31076 19780
rect 31024 19737 31033 19771
rect 31033 19737 31067 19771
rect 31067 19737 31076 19771
rect 31024 19728 31076 19737
rect 33416 19728 33468 19780
rect 34060 19728 34112 19780
rect 38016 19771 38068 19780
rect 38016 19737 38025 19771
rect 38025 19737 38059 19771
rect 38059 19737 38068 19771
rect 38016 19728 38068 19737
rect 38200 19771 38252 19780
rect 38200 19737 38225 19771
rect 38225 19737 38252 19771
rect 38200 19728 38252 19737
rect 38568 19728 38620 19780
rect 38660 19728 38712 19780
rect 40776 19771 40828 19780
rect 40776 19737 40785 19771
rect 40785 19737 40819 19771
rect 40819 19737 40828 19771
rect 40776 19728 40828 19737
rect 40960 19728 41012 19780
rect 41880 19771 41932 19780
rect 41880 19737 41889 19771
rect 41889 19737 41923 19771
rect 41923 19737 41932 19771
rect 41880 19728 41932 19737
rect 44088 19728 44140 19780
rect 45192 19728 45244 19780
rect 46296 19728 46348 19780
rect 46940 19728 46992 19780
rect 18604 19660 18656 19712
rect 18972 19660 19024 19712
rect 21732 19660 21784 19712
rect 22836 19660 22888 19712
rect 23112 19660 23164 19712
rect 23204 19660 23256 19712
rect 26424 19660 26476 19712
rect 27160 19660 27212 19712
rect 27344 19660 27396 19712
rect 35624 19660 35676 19712
rect 38476 19660 38528 19712
rect 39120 19660 39172 19712
rect 40868 19660 40920 19712
rect 41420 19660 41472 19712
rect 45468 19703 45520 19712
rect 45468 19669 45477 19703
rect 45477 19669 45511 19703
rect 45511 19669 45520 19703
rect 45468 19660 45520 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 17224 19388 17276 19440
rect 2412 19320 2464 19372
rect 12348 19320 12400 19372
rect 17408 19320 17460 19372
rect 17960 19320 18012 19372
rect 18696 19456 18748 19508
rect 22928 19456 22980 19508
rect 26608 19456 26660 19508
rect 29276 19499 29328 19508
rect 29276 19465 29285 19499
rect 29285 19465 29319 19499
rect 29319 19465 29328 19499
rect 29276 19456 29328 19465
rect 29460 19456 29512 19508
rect 33416 19456 33468 19508
rect 38200 19456 38252 19508
rect 39396 19456 39448 19508
rect 40776 19456 40828 19508
rect 41880 19456 41932 19508
rect 46940 19499 46992 19508
rect 46940 19465 46949 19499
rect 46949 19465 46983 19499
rect 46983 19465 46992 19499
rect 46940 19456 46992 19465
rect 18788 19388 18840 19440
rect 34152 19388 34204 19440
rect 35900 19388 35952 19440
rect 38108 19388 38160 19440
rect 18880 19320 18932 19372
rect 19984 19363 20036 19372
rect 19984 19329 19993 19363
rect 19993 19329 20027 19363
rect 20027 19329 20036 19363
rect 19984 19320 20036 19329
rect 22560 19320 22612 19372
rect 23480 19320 23532 19372
rect 25136 19320 25188 19372
rect 26240 19320 26292 19372
rect 26424 19320 26476 19372
rect 26976 19363 27028 19372
rect 26976 19329 26985 19363
rect 26985 19329 27019 19363
rect 27019 19329 27028 19363
rect 26976 19320 27028 19329
rect 27068 19320 27120 19372
rect 22376 19252 22428 19304
rect 22836 19252 22888 19304
rect 23388 19295 23440 19304
rect 23388 19261 23397 19295
rect 23397 19261 23431 19295
rect 23431 19261 23440 19295
rect 23388 19252 23440 19261
rect 25596 19295 25648 19304
rect 25596 19261 25605 19295
rect 25605 19261 25639 19295
rect 25639 19261 25648 19295
rect 25596 19252 25648 19261
rect 26148 19252 26200 19304
rect 26792 19252 26844 19304
rect 29092 19320 29144 19372
rect 31024 19320 31076 19372
rect 33416 19363 33468 19372
rect 33416 19329 33425 19363
rect 33425 19329 33459 19363
rect 33459 19329 33468 19363
rect 33416 19320 33468 19329
rect 33600 19363 33652 19372
rect 33600 19329 33609 19363
rect 33609 19329 33643 19363
rect 33643 19329 33652 19363
rect 33600 19320 33652 19329
rect 34060 19320 34112 19372
rect 33876 19252 33928 19304
rect 37004 19320 37056 19372
rect 38200 19363 38252 19372
rect 38200 19329 38209 19363
rect 38209 19329 38243 19363
rect 38243 19329 38252 19363
rect 38200 19320 38252 19329
rect 38384 19363 38436 19372
rect 38384 19329 38393 19363
rect 38393 19329 38427 19363
rect 38427 19329 38436 19363
rect 38384 19320 38436 19329
rect 39028 19320 39080 19372
rect 39120 19363 39172 19372
rect 39120 19329 39129 19363
rect 39129 19329 39163 19363
rect 39163 19329 39172 19363
rect 41328 19388 41380 19440
rect 39120 19320 39172 19329
rect 40684 19320 40736 19372
rect 40960 19320 41012 19372
rect 41604 19320 41656 19372
rect 43168 19320 43220 19372
rect 44824 19363 44876 19372
rect 44824 19329 44858 19363
rect 44858 19329 44876 19363
rect 44824 19320 44876 19329
rect 45100 19320 45152 19372
rect 47952 19363 48004 19372
rect 47952 19329 47961 19363
rect 47961 19329 47995 19363
rect 47995 19329 48004 19363
rect 47952 19320 48004 19329
rect 37464 19252 37516 19304
rect 38660 19252 38712 19304
rect 43812 19252 43864 19304
rect 44548 19295 44600 19304
rect 44548 19261 44557 19295
rect 44557 19261 44591 19295
rect 44591 19261 44600 19295
rect 44548 19252 44600 19261
rect 22100 19227 22152 19236
rect 22100 19193 22109 19227
rect 22109 19193 22143 19227
rect 22143 19193 22152 19227
rect 22744 19227 22796 19236
rect 22100 19184 22152 19193
rect 22744 19193 22753 19227
rect 22753 19193 22787 19227
rect 22787 19193 22796 19227
rect 22744 19184 22796 19193
rect 33508 19184 33560 19236
rect 37280 19184 37332 19236
rect 41144 19184 41196 19236
rect 41604 19227 41656 19236
rect 41604 19193 41613 19227
rect 41613 19193 41647 19227
rect 41647 19193 41656 19227
rect 41604 19184 41656 19193
rect 1400 19116 1452 19168
rect 2320 19159 2372 19168
rect 2320 19125 2329 19159
rect 2329 19125 2363 19159
rect 2363 19125 2372 19159
rect 2320 19116 2372 19125
rect 17960 19159 18012 19168
rect 17960 19125 17969 19159
rect 17969 19125 18003 19159
rect 18003 19125 18012 19159
rect 17960 19116 18012 19125
rect 19616 19116 19668 19168
rect 22192 19116 22244 19168
rect 25688 19116 25740 19168
rect 31668 19116 31720 19168
rect 33140 19159 33192 19168
rect 33140 19125 33149 19159
rect 33149 19125 33183 19159
rect 33183 19125 33192 19159
rect 33140 19116 33192 19125
rect 33784 19116 33836 19168
rect 38476 19159 38528 19168
rect 38476 19125 38485 19159
rect 38485 19125 38519 19159
rect 38519 19125 38528 19159
rect 38476 19116 38528 19125
rect 38660 19159 38712 19168
rect 38660 19125 38669 19159
rect 38669 19125 38703 19159
rect 38703 19125 38712 19159
rect 38660 19116 38712 19125
rect 41420 19159 41472 19168
rect 41420 19125 41429 19159
rect 41429 19125 41463 19159
rect 41463 19125 41472 19159
rect 42432 19159 42484 19168
rect 41420 19116 41472 19125
rect 42432 19125 42441 19159
rect 42441 19125 42475 19159
rect 42475 19125 42484 19159
rect 42432 19116 42484 19125
rect 45928 19159 45980 19168
rect 45928 19125 45937 19159
rect 45937 19125 45971 19159
rect 45971 19125 45980 19159
rect 45928 19116 45980 19125
rect 48044 19159 48096 19168
rect 48044 19125 48053 19159
rect 48053 19125 48087 19159
rect 48087 19125 48096 19159
rect 48044 19116 48096 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 18420 18912 18472 18964
rect 22560 18912 22612 18964
rect 24124 18912 24176 18964
rect 25780 18912 25832 18964
rect 32312 18912 32364 18964
rect 22192 18844 22244 18896
rect 25044 18844 25096 18896
rect 1400 18819 1452 18828
rect 1400 18785 1409 18819
rect 1409 18785 1443 18819
rect 1443 18785 1452 18819
rect 1400 18776 1452 18785
rect 2320 18776 2372 18828
rect 2780 18819 2832 18828
rect 2780 18785 2789 18819
rect 2789 18785 2823 18819
rect 2823 18785 2832 18819
rect 2780 18776 2832 18785
rect 22376 18819 22428 18828
rect 22376 18785 22385 18819
rect 22385 18785 22419 18819
rect 22419 18785 22428 18819
rect 22376 18776 22428 18785
rect 23112 18819 23164 18828
rect 23112 18785 23121 18819
rect 23121 18785 23155 18819
rect 23155 18785 23164 18819
rect 23112 18776 23164 18785
rect 15752 18708 15804 18760
rect 19340 18751 19392 18760
rect 19340 18717 19349 18751
rect 19349 18717 19383 18751
rect 19383 18717 19392 18751
rect 19340 18708 19392 18717
rect 19616 18751 19668 18760
rect 19616 18717 19650 18751
rect 19650 18717 19668 18751
rect 19616 18708 19668 18717
rect 22100 18751 22152 18760
rect 22100 18717 22109 18751
rect 22109 18717 22143 18751
rect 22143 18717 22152 18751
rect 22100 18708 22152 18717
rect 22744 18708 22796 18760
rect 17960 18640 18012 18692
rect 18236 18640 18288 18692
rect 16672 18572 16724 18624
rect 17408 18572 17460 18624
rect 17868 18572 17920 18624
rect 19892 18640 19944 18692
rect 21088 18640 21140 18692
rect 23480 18708 23532 18760
rect 24768 18751 24820 18760
rect 24768 18717 24777 18751
rect 24777 18717 24811 18751
rect 24811 18717 24820 18751
rect 24768 18708 24820 18717
rect 24952 18708 25004 18760
rect 25320 18751 25372 18760
rect 25320 18717 25329 18751
rect 25329 18717 25363 18751
rect 25363 18717 25372 18751
rect 25320 18708 25372 18717
rect 25688 18708 25740 18760
rect 29736 18751 29788 18760
rect 29736 18717 29745 18751
rect 29745 18717 29779 18751
rect 29779 18717 29788 18751
rect 29736 18708 29788 18717
rect 30840 18708 30892 18760
rect 31760 18708 31812 18760
rect 23848 18640 23900 18692
rect 26792 18683 26844 18692
rect 26792 18649 26801 18683
rect 26801 18649 26835 18683
rect 26835 18649 26844 18683
rect 26792 18640 26844 18649
rect 27896 18640 27948 18692
rect 28356 18640 28408 18692
rect 20628 18572 20680 18624
rect 22192 18572 22244 18624
rect 25412 18572 25464 18624
rect 27436 18572 27488 18624
rect 29000 18640 29052 18692
rect 30932 18640 30984 18692
rect 31668 18640 31720 18692
rect 33508 18844 33560 18896
rect 33048 18776 33100 18828
rect 33508 18708 33560 18760
rect 33784 18751 33836 18760
rect 33784 18717 33793 18751
rect 33793 18717 33827 18751
rect 33827 18717 33836 18751
rect 35900 18912 35952 18964
rect 37372 18912 37424 18964
rect 39028 18912 39080 18964
rect 40776 18912 40828 18964
rect 41512 18912 41564 18964
rect 38752 18819 38804 18828
rect 38752 18785 38761 18819
rect 38761 18785 38795 18819
rect 38795 18785 38804 18819
rect 38752 18776 38804 18785
rect 41052 18887 41104 18896
rect 41052 18853 41061 18887
rect 41061 18853 41095 18887
rect 41095 18853 41104 18887
rect 41052 18844 41104 18853
rect 45376 18844 45428 18896
rect 45468 18844 45520 18896
rect 46112 18844 46164 18896
rect 40776 18776 40828 18828
rect 41236 18776 41288 18828
rect 33784 18708 33836 18717
rect 34060 18708 34112 18760
rect 35992 18708 36044 18760
rect 37924 18751 37976 18760
rect 37924 18717 37933 18751
rect 37933 18717 37967 18751
rect 37967 18717 37976 18751
rect 37924 18708 37976 18717
rect 38016 18751 38068 18760
rect 38016 18717 38025 18751
rect 38025 18717 38059 18751
rect 38059 18717 38068 18751
rect 38016 18708 38068 18717
rect 38660 18708 38712 18760
rect 43076 18776 43128 18828
rect 40224 18683 40276 18692
rect 40224 18649 40233 18683
rect 40233 18649 40267 18683
rect 40267 18649 40276 18683
rect 40224 18640 40276 18649
rect 44548 18708 44600 18760
rect 47032 18776 47084 18828
rect 45652 18751 45704 18760
rect 45652 18717 45661 18751
rect 45661 18717 45695 18751
rect 45695 18717 45704 18751
rect 45652 18708 45704 18717
rect 45744 18708 45796 18760
rect 40684 18572 40736 18624
rect 40776 18572 40828 18624
rect 41328 18572 41380 18624
rect 42156 18572 42208 18624
rect 42432 18640 42484 18692
rect 44088 18683 44140 18692
rect 44088 18649 44097 18683
rect 44097 18649 44131 18683
rect 44131 18649 44140 18683
rect 44088 18640 44140 18649
rect 45928 18640 45980 18692
rect 43260 18572 43312 18624
rect 44456 18615 44508 18624
rect 44456 18581 44465 18615
rect 44465 18581 44499 18615
rect 44499 18581 44508 18615
rect 44456 18572 44508 18581
rect 45008 18615 45060 18624
rect 45008 18581 45017 18615
rect 45017 18581 45051 18615
rect 45051 18581 45060 18615
rect 45008 18572 45060 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 15752 18368 15804 18420
rect 19984 18368 20036 18420
rect 21916 18368 21968 18420
rect 22836 18368 22888 18420
rect 23020 18368 23072 18420
rect 15384 18343 15436 18352
rect 15384 18309 15393 18343
rect 15393 18309 15427 18343
rect 15427 18309 15436 18343
rect 15384 18300 15436 18309
rect 18052 18300 18104 18352
rect 1952 18232 2004 18284
rect 20628 18275 20680 18284
rect 20628 18241 20637 18275
rect 20637 18241 20671 18275
rect 20671 18241 20680 18275
rect 20628 18232 20680 18241
rect 3424 18096 3476 18148
rect 1584 18028 1636 18080
rect 2872 18071 2924 18080
rect 2872 18037 2881 18071
rect 2881 18037 2915 18071
rect 2915 18037 2924 18071
rect 2872 18028 2924 18037
rect 20996 18164 21048 18216
rect 17868 18096 17920 18148
rect 22192 18275 22244 18284
rect 22192 18241 22201 18275
rect 22201 18241 22235 18275
rect 22235 18241 22244 18275
rect 22192 18232 22244 18241
rect 22560 18232 22612 18284
rect 24768 18368 24820 18420
rect 26792 18368 26844 18420
rect 27896 18411 27948 18420
rect 27896 18377 27905 18411
rect 27905 18377 27939 18411
rect 27939 18377 27948 18411
rect 27896 18368 27948 18377
rect 28264 18368 28316 18420
rect 30932 18411 30984 18420
rect 30932 18377 30941 18411
rect 30941 18377 30975 18411
rect 30975 18377 30984 18411
rect 30932 18368 30984 18377
rect 37924 18368 37976 18420
rect 41512 18411 41564 18420
rect 41512 18377 41521 18411
rect 41521 18377 41555 18411
rect 41555 18377 41564 18411
rect 41512 18368 41564 18377
rect 43812 18411 43864 18420
rect 43812 18377 43821 18411
rect 43821 18377 43855 18411
rect 43855 18377 43864 18411
rect 43812 18368 43864 18377
rect 46296 18368 46348 18420
rect 25596 18300 25648 18352
rect 26424 18300 26476 18352
rect 23204 18275 23256 18284
rect 23204 18241 23213 18275
rect 23213 18241 23247 18275
rect 23247 18241 23256 18275
rect 23204 18232 23256 18241
rect 23388 18232 23440 18284
rect 25320 18232 25372 18284
rect 26608 18232 26660 18284
rect 27160 18275 27212 18284
rect 27160 18241 27169 18275
rect 27169 18241 27203 18275
rect 27203 18241 27212 18275
rect 27160 18232 27212 18241
rect 27344 18275 27396 18284
rect 27344 18241 27353 18275
rect 27353 18241 27387 18275
rect 27387 18241 27396 18275
rect 27344 18232 27396 18241
rect 27620 18232 27672 18284
rect 28356 18275 28408 18284
rect 25136 18164 25188 18216
rect 25780 18164 25832 18216
rect 23020 18096 23072 18148
rect 26240 18207 26292 18216
rect 26240 18173 26249 18207
rect 26249 18173 26283 18207
rect 26283 18173 26292 18207
rect 27436 18207 27488 18216
rect 26240 18164 26292 18173
rect 27436 18173 27445 18207
rect 27445 18173 27479 18207
rect 27479 18173 27488 18207
rect 27436 18164 27488 18173
rect 28356 18241 28365 18275
rect 28365 18241 28399 18275
rect 28399 18241 28408 18275
rect 28356 18232 28408 18241
rect 30012 18275 30064 18284
rect 30012 18241 30021 18275
rect 30021 18241 30055 18275
rect 30055 18241 30064 18275
rect 30012 18232 30064 18241
rect 33140 18300 33192 18352
rect 41144 18343 41196 18352
rect 41144 18309 41153 18343
rect 41153 18309 41187 18343
rect 41187 18309 41196 18343
rect 41144 18300 41196 18309
rect 45008 18300 45060 18352
rect 29368 18164 29420 18216
rect 31668 18232 31720 18284
rect 31760 18232 31812 18284
rect 31852 18164 31904 18216
rect 32128 18275 32180 18284
rect 32128 18241 32137 18275
rect 32137 18241 32171 18275
rect 32171 18241 32180 18275
rect 32312 18275 32364 18284
rect 32128 18232 32180 18241
rect 32312 18241 32321 18275
rect 32321 18241 32355 18275
rect 32355 18241 32364 18275
rect 32312 18232 32364 18241
rect 36544 18232 36596 18284
rect 32864 18164 32916 18216
rect 37648 18164 37700 18216
rect 37924 18232 37976 18284
rect 40224 18232 40276 18284
rect 40868 18232 40920 18284
rect 41972 18232 42024 18284
rect 44548 18232 44600 18284
rect 47308 18232 47360 18284
rect 38292 18207 38344 18216
rect 38292 18173 38301 18207
rect 38301 18173 38335 18207
rect 38335 18173 38344 18207
rect 38292 18164 38344 18173
rect 40132 18164 40184 18216
rect 41236 18164 41288 18216
rect 18880 18028 18932 18080
rect 23204 18028 23256 18080
rect 24216 18028 24268 18080
rect 25044 18071 25096 18080
rect 25044 18037 25053 18071
rect 25053 18037 25087 18071
rect 25087 18037 25096 18071
rect 25044 18028 25096 18037
rect 25504 18028 25556 18080
rect 26608 18028 26660 18080
rect 26884 18028 26936 18080
rect 33508 18096 33560 18148
rect 29276 18028 29328 18080
rect 29828 18028 29880 18080
rect 30288 18028 30340 18080
rect 35348 18071 35400 18080
rect 35348 18037 35357 18071
rect 35357 18037 35391 18071
rect 35391 18037 35400 18071
rect 35348 18028 35400 18037
rect 45744 18028 45796 18080
rect 47676 18071 47728 18080
rect 47676 18037 47685 18071
rect 47685 18037 47719 18071
rect 47719 18037 47728 18071
rect 47676 18028 47728 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 15384 17824 15436 17876
rect 16120 17824 16172 17876
rect 2872 17756 2924 17808
rect 20812 17756 20864 17808
rect 1584 17731 1636 17740
rect 1584 17697 1593 17731
rect 1593 17697 1627 17731
rect 1627 17697 1636 17731
rect 1584 17688 1636 17697
rect 2780 17731 2832 17740
rect 2780 17697 2789 17731
rect 2789 17697 2823 17731
rect 2823 17697 2832 17731
rect 2780 17688 2832 17697
rect 20996 17688 21048 17740
rect 22560 17688 22612 17740
rect 23664 17867 23716 17876
rect 23664 17833 23673 17867
rect 23673 17833 23707 17867
rect 23707 17833 23716 17867
rect 23664 17824 23716 17833
rect 25136 17824 25188 17876
rect 26240 17824 26292 17876
rect 28264 17824 28316 17876
rect 29276 17824 29328 17876
rect 29552 17824 29604 17876
rect 31760 17824 31812 17876
rect 32864 17867 32916 17876
rect 32864 17833 32873 17867
rect 32873 17833 32907 17867
rect 32907 17833 32916 17867
rect 32864 17824 32916 17833
rect 33600 17824 33652 17876
rect 38016 17824 38068 17876
rect 41972 17867 42024 17876
rect 41972 17833 41981 17867
rect 41981 17833 42015 17867
rect 42015 17833 42024 17867
rect 41972 17824 42024 17833
rect 44824 17824 44876 17876
rect 23572 17756 23624 17808
rect 26056 17756 26108 17808
rect 29460 17756 29512 17808
rect 39396 17756 39448 17808
rect 45652 17756 45704 17808
rect 15844 17620 15896 17672
rect 20352 17620 20404 17672
rect 23204 17663 23256 17672
rect 16580 17552 16632 17604
rect 17960 17552 18012 17604
rect 20628 17552 20680 17604
rect 20352 17527 20404 17536
rect 20352 17493 20361 17527
rect 20361 17493 20395 17527
rect 20395 17493 20404 17527
rect 20352 17484 20404 17493
rect 22560 17595 22612 17604
rect 22560 17561 22569 17595
rect 22569 17561 22603 17595
rect 22603 17561 22612 17595
rect 22560 17552 22612 17561
rect 22836 17552 22888 17604
rect 23204 17629 23213 17663
rect 23213 17629 23247 17663
rect 23247 17629 23256 17663
rect 23204 17620 23256 17629
rect 23296 17620 23348 17672
rect 24216 17620 24268 17672
rect 25412 17663 25464 17672
rect 25412 17629 25421 17663
rect 25421 17629 25455 17663
rect 25455 17629 25464 17663
rect 25412 17620 25464 17629
rect 25504 17663 25556 17672
rect 25504 17629 25513 17663
rect 25513 17629 25547 17663
rect 25547 17629 25556 17663
rect 25504 17620 25556 17629
rect 25688 17552 25740 17604
rect 25964 17620 26016 17672
rect 27896 17620 27948 17672
rect 28356 17620 28408 17672
rect 29552 17663 29604 17672
rect 29552 17629 29561 17663
rect 29561 17629 29595 17663
rect 29595 17629 29604 17663
rect 29552 17620 29604 17629
rect 32036 17688 32088 17740
rect 26424 17552 26476 17604
rect 29828 17595 29880 17604
rect 29828 17561 29862 17595
rect 29862 17561 29880 17595
rect 22928 17484 22980 17536
rect 23296 17484 23348 17536
rect 25780 17484 25832 17536
rect 29828 17552 29880 17561
rect 29368 17484 29420 17536
rect 31484 17552 31536 17604
rect 34152 17620 34204 17672
rect 37924 17663 37976 17672
rect 37924 17629 37933 17663
rect 37933 17629 37967 17663
rect 37967 17629 37976 17663
rect 37924 17620 37976 17629
rect 38292 17688 38344 17740
rect 40776 17688 40828 17740
rect 40040 17620 40092 17672
rect 40408 17620 40460 17672
rect 41052 17620 41104 17672
rect 44456 17688 44508 17740
rect 42156 17663 42208 17672
rect 42156 17629 42165 17663
rect 42165 17629 42199 17663
rect 42199 17629 42208 17663
rect 42156 17620 42208 17629
rect 43260 17663 43312 17672
rect 43260 17629 43269 17663
rect 43269 17629 43303 17663
rect 43303 17629 43312 17663
rect 43260 17620 43312 17629
rect 46296 17731 46348 17740
rect 46296 17697 46305 17731
rect 46305 17697 46339 17731
rect 46339 17697 46348 17731
rect 46296 17688 46348 17697
rect 47676 17688 47728 17740
rect 48136 17731 48188 17740
rect 48136 17697 48145 17731
rect 48145 17697 48179 17731
rect 48179 17697 48188 17731
rect 48136 17688 48188 17697
rect 32128 17552 32180 17604
rect 33876 17552 33928 17604
rect 35348 17552 35400 17604
rect 37648 17484 37700 17536
rect 41604 17484 41656 17536
rect 41880 17484 41932 17536
rect 45376 17484 45428 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 19064 17280 19116 17332
rect 21732 17280 21784 17332
rect 22284 17280 22336 17332
rect 24492 17280 24544 17332
rect 29368 17280 29420 17332
rect 29828 17323 29880 17332
rect 29828 17289 29837 17323
rect 29837 17289 29871 17323
rect 29871 17289 29880 17323
rect 29828 17280 29880 17289
rect 35992 17323 36044 17332
rect 35992 17289 36001 17323
rect 36001 17289 36035 17323
rect 36035 17289 36044 17323
rect 35992 17280 36044 17289
rect 19984 17212 20036 17264
rect 20260 17212 20312 17264
rect 22376 17212 22428 17264
rect 24676 17212 24728 17264
rect 26240 17255 26292 17264
rect 1860 17187 1912 17196
rect 1860 17153 1869 17187
rect 1869 17153 1903 17187
rect 1903 17153 1912 17187
rect 1860 17144 1912 17153
rect 15936 17187 15988 17196
rect 15936 17153 15945 17187
rect 15945 17153 15979 17187
rect 15979 17153 15988 17187
rect 15936 17144 15988 17153
rect 16672 17187 16724 17196
rect 16672 17153 16681 17187
rect 16681 17153 16715 17187
rect 16715 17153 16724 17187
rect 16672 17144 16724 17153
rect 20628 17144 20680 17196
rect 22928 17187 22980 17196
rect 22928 17153 22937 17187
rect 22937 17153 22971 17187
rect 22971 17153 22980 17187
rect 22928 17144 22980 17153
rect 23848 17144 23900 17196
rect 24308 17144 24360 17196
rect 25412 17144 25464 17196
rect 25780 17144 25832 17196
rect 26240 17221 26249 17255
rect 26249 17221 26283 17255
rect 26283 17221 26292 17255
rect 26240 17212 26292 17221
rect 26792 17212 26844 17264
rect 29276 17212 29328 17264
rect 18328 17119 18380 17128
rect 18328 17085 18337 17119
rect 18337 17085 18371 17119
rect 18371 17085 18380 17119
rect 18328 17076 18380 17085
rect 2136 16940 2188 16992
rect 26424 17076 26476 17128
rect 19340 16940 19392 16992
rect 20260 16940 20312 16992
rect 20352 16983 20404 16992
rect 20352 16949 20361 16983
rect 20361 16949 20395 16983
rect 20395 16949 20404 16983
rect 20352 16940 20404 16949
rect 20904 16940 20956 16992
rect 26884 17008 26936 17060
rect 27896 17144 27948 17196
rect 30840 17212 30892 17264
rect 31852 17212 31904 17264
rect 33048 17212 33100 17264
rect 33876 17255 33928 17264
rect 33876 17221 33885 17255
rect 33885 17221 33919 17255
rect 33919 17221 33928 17255
rect 33876 17212 33928 17221
rect 35532 17212 35584 17264
rect 41052 17212 41104 17264
rect 41788 17212 41840 17264
rect 41972 17212 42024 17264
rect 30288 17187 30340 17196
rect 29920 17076 29972 17128
rect 30288 17153 30297 17187
rect 30297 17153 30331 17187
rect 30331 17153 30340 17187
rect 30288 17144 30340 17153
rect 22560 16940 22612 16992
rect 23664 16940 23716 16992
rect 25596 16983 25648 16992
rect 25596 16949 25605 16983
rect 25605 16949 25639 16983
rect 25639 16949 25648 16983
rect 25596 16940 25648 16949
rect 28540 17008 28592 17060
rect 28632 17008 28684 17060
rect 31300 17144 31352 17196
rect 34152 17144 34204 17196
rect 36176 17144 36228 17196
rect 40040 17187 40092 17196
rect 40040 17153 40049 17187
rect 40049 17153 40083 17187
rect 40083 17153 40092 17187
rect 40040 17144 40092 17153
rect 40500 17144 40552 17196
rect 40776 17187 40828 17196
rect 40776 17153 40785 17187
rect 40785 17153 40819 17187
rect 40819 17153 40828 17187
rect 40776 17144 40828 17153
rect 30840 17076 30892 17128
rect 37648 17076 37700 17128
rect 45836 17280 45888 17332
rect 47584 17187 47636 17196
rect 47584 17153 47593 17187
rect 47593 17153 47627 17187
rect 47627 17153 47636 17187
rect 47584 17144 47636 17153
rect 45836 17076 45888 17128
rect 46848 17119 46900 17128
rect 46848 17085 46857 17119
rect 46857 17085 46891 17119
rect 46891 17085 46900 17119
rect 46848 17076 46900 17085
rect 39396 17008 39448 17060
rect 27988 16983 28040 16992
rect 27988 16949 27997 16983
rect 27997 16949 28031 16983
rect 28031 16949 28040 16983
rect 27988 16940 28040 16949
rect 29736 16940 29788 16992
rect 33876 16940 33928 16992
rect 41420 16940 41472 16992
rect 41604 16983 41656 16992
rect 41604 16949 41613 16983
rect 41613 16949 41647 16983
rect 41647 16949 41656 16983
rect 41604 16940 41656 16949
rect 41788 16983 41840 16992
rect 41788 16949 41797 16983
rect 41797 16949 41831 16983
rect 41831 16949 41840 16983
rect 41788 16940 41840 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 1860 16668 1912 16720
rect 2136 16600 2188 16652
rect 3332 16600 3384 16652
rect 16672 16736 16724 16788
rect 20904 16736 20956 16788
rect 23204 16736 23256 16788
rect 23388 16736 23440 16788
rect 23572 16668 23624 16720
rect 17960 16600 18012 16652
rect 20260 16643 20312 16652
rect 20260 16609 20269 16643
rect 20269 16609 20303 16643
rect 20303 16609 20312 16643
rect 20260 16600 20312 16609
rect 23388 16600 23440 16652
rect 15200 16532 15252 16584
rect 15384 16532 15436 16584
rect 19248 16575 19300 16584
rect 19248 16541 19257 16575
rect 19257 16541 19291 16575
rect 19291 16541 19300 16575
rect 19248 16532 19300 16541
rect 22192 16532 22244 16584
rect 23020 16575 23072 16584
rect 23020 16541 23029 16575
rect 23029 16541 23063 16575
rect 23063 16541 23072 16575
rect 23020 16532 23072 16541
rect 23756 16600 23808 16652
rect 24952 16600 25004 16652
rect 25964 16668 26016 16720
rect 25596 16600 25648 16652
rect 26240 16736 26292 16788
rect 26884 16736 26936 16788
rect 42156 16779 42208 16788
rect 27344 16668 27396 16720
rect 27620 16668 27672 16720
rect 27896 16711 27948 16720
rect 27896 16677 27905 16711
rect 27905 16677 27939 16711
rect 27939 16677 27948 16711
rect 27896 16668 27948 16677
rect 29184 16668 29236 16720
rect 30932 16668 30984 16720
rect 33232 16668 33284 16720
rect 34060 16668 34112 16720
rect 37648 16711 37700 16720
rect 37648 16677 37657 16711
rect 37657 16677 37691 16711
rect 37691 16677 37700 16711
rect 37648 16668 37700 16677
rect 42156 16745 42165 16779
rect 42165 16745 42199 16779
rect 42199 16745 42208 16779
rect 42156 16736 42208 16745
rect 45836 16779 45888 16788
rect 45836 16745 45845 16779
rect 45845 16745 45879 16779
rect 45879 16745 45888 16779
rect 45836 16736 45888 16745
rect 47584 16668 47636 16720
rect 25688 16575 25740 16584
rect 25688 16541 25697 16575
rect 25697 16541 25731 16575
rect 25731 16541 25740 16575
rect 25688 16532 25740 16541
rect 25872 16575 25924 16584
rect 25872 16541 25881 16575
rect 25881 16541 25915 16575
rect 25915 16541 25924 16575
rect 25872 16532 25924 16541
rect 26240 16575 26292 16584
rect 26240 16541 26249 16575
rect 26249 16541 26283 16575
rect 26283 16541 26292 16575
rect 26240 16532 26292 16541
rect 27988 16600 28040 16652
rect 33048 16600 33100 16652
rect 31484 16532 31536 16584
rect 31668 16532 31720 16584
rect 1584 16507 1636 16516
rect 1584 16473 1593 16507
rect 1593 16473 1627 16507
rect 1627 16473 1636 16507
rect 1584 16464 1636 16473
rect 2596 16464 2648 16516
rect 15752 16464 15804 16516
rect 15844 16464 15896 16516
rect 19064 16464 19116 16516
rect 22560 16464 22612 16516
rect 22928 16464 22980 16516
rect 30380 16464 30432 16516
rect 32128 16464 32180 16516
rect 13820 16396 13872 16448
rect 15476 16396 15528 16448
rect 17040 16396 17092 16448
rect 21640 16439 21692 16448
rect 21640 16405 21649 16439
rect 21649 16405 21683 16439
rect 21683 16405 21692 16439
rect 21640 16396 21692 16405
rect 21824 16396 21876 16448
rect 22744 16439 22796 16448
rect 22744 16405 22753 16439
rect 22753 16405 22787 16439
rect 22787 16405 22796 16439
rect 22744 16396 22796 16405
rect 24400 16396 24452 16448
rect 25136 16396 25188 16448
rect 32588 16396 32640 16448
rect 33416 16532 33468 16584
rect 33876 16575 33928 16584
rect 33876 16541 33885 16575
rect 33885 16541 33919 16575
rect 33919 16541 33928 16575
rect 35992 16600 36044 16652
rect 40132 16643 40184 16652
rect 40132 16609 40141 16643
rect 40141 16609 40175 16643
rect 40175 16609 40184 16643
rect 40132 16600 40184 16609
rect 45928 16600 45980 16652
rect 33876 16532 33928 16541
rect 33600 16464 33652 16516
rect 37464 16464 37516 16516
rect 45836 16532 45888 16584
rect 41236 16464 41288 16516
rect 41420 16464 41472 16516
rect 41972 16507 42024 16516
rect 34244 16396 34296 16448
rect 40776 16396 40828 16448
rect 41972 16473 41981 16507
rect 41981 16473 42015 16507
rect 42015 16473 42024 16507
rect 41972 16464 42024 16473
rect 46480 16507 46532 16516
rect 46480 16473 46489 16507
rect 46489 16473 46523 16507
rect 46523 16473 46532 16507
rect 46480 16464 46532 16473
rect 42616 16396 42668 16448
rect 46020 16396 46072 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 1584 16192 1636 16244
rect 20628 16235 20680 16244
rect 1492 16056 1544 16108
rect 13820 16124 13872 16176
rect 15476 16124 15528 16176
rect 16212 16124 16264 16176
rect 17040 16167 17092 16176
rect 17040 16133 17049 16167
rect 17049 16133 17083 16167
rect 17083 16133 17092 16167
rect 17040 16124 17092 16133
rect 20628 16201 20637 16235
rect 20637 16201 20671 16235
rect 20671 16201 20680 16235
rect 20628 16192 20680 16201
rect 21640 16124 21692 16176
rect 23020 16192 23072 16244
rect 24124 16192 24176 16244
rect 24584 16192 24636 16244
rect 32128 16235 32180 16244
rect 32128 16201 32137 16235
rect 32137 16201 32171 16235
rect 32171 16201 32180 16235
rect 32128 16192 32180 16201
rect 35532 16235 35584 16244
rect 35532 16201 35541 16235
rect 35541 16201 35575 16235
rect 35575 16201 35584 16235
rect 35532 16192 35584 16201
rect 40040 16192 40092 16244
rect 41236 16235 41288 16244
rect 41236 16201 41245 16235
rect 41245 16201 41279 16235
rect 41279 16201 41288 16235
rect 41236 16192 41288 16201
rect 46480 16235 46532 16244
rect 46480 16201 46489 16235
rect 46489 16201 46523 16235
rect 46523 16201 46532 16235
rect 46480 16192 46532 16201
rect 19248 16099 19300 16108
rect 19248 16065 19257 16099
rect 19257 16065 19291 16099
rect 19291 16065 19300 16099
rect 19248 16056 19300 16065
rect 20812 16099 20864 16108
rect 20812 16065 20821 16099
rect 20821 16065 20855 16099
rect 20855 16065 20864 16099
rect 20812 16056 20864 16065
rect 21824 16099 21876 16108
rect 21824 16065 21833 16099
rect 21833 16065 21867 16099
rect 21867 16065 21876 16099
rect 21824 16056 21876 16065
rect 30380 16124 30432 16176
rect 296 15988 348 16040
rect 14188 16031 14240 16040
rect 14188 15997 14197 16031
rect 14197 15997 14231 16031
rect 14231 15997 14240 16031
rect 14188 15988 14240 15997
rect 19892 16031 19944 16040
rect 18144 15920 18196 15972
rect 12992 15852 13044 15904
rect 19892 15997 19901 16031
rect 19901 15997 19935 16031
rect 19935 15997 19944 16031
rect 19892 15988 19944 15997
rect 21732 15988 21784 16040
rect 23112 16056 23164 16108
rect 24124 16099 24176 16108
rect 24124 16065 24133 16099
rect 24133 16065 24167 16099
rect 24167 16065 24176 16099
rect 24124 16056 24176 16065
rect 24400 16056 24452 16108
rect 24952 16099 25004 16108
rect 24952 16065 24961 16099
rect 24961 16065 24995 16099
rect 24995 16065 25004 16099
rect 24952 16056 25004 16065
rect 29460 16099 29512 16108
rect 29460 16065 29469 16099
rect 29469 16065 29503 16099
rect 29503 16065 29512 16099
rect 29460 16056 29512 16065
rect 30564 16099 30616 16108
rect 30564 16065 30573 16099
rect 30573 16065 30607 16099
rect 30607 16065 30616 16099
rect 30564 16056 30616 16065
rect 31024 16124 31076 16176
rect 30748 16099 30800 16108
rect 30748 16065 30757 16099
rect 30757 16065 30791 16099
rect 30791 16065 30800 16099
rect 30748 16056 30800 16065
rect 22560 16031 22612 16040
rect 22560 15997 22569 16031
rect 22569 15997 22603 16031
rect 22603 15997 22612 16031
rect 22560 15988 22612 15997
rect 31944 16056 31996 16108
rect 33048 16124 33100 16176
rect 34152 16124 34204 16176
rect 32588 16099 32640 16108
rect 32588 16065 32597 16099
rect 32597 16065 32631 16099
rect 32631 16065 32640 16099
rect 32588 16056 32640 16065
rect 33232 16056 33284 16108
rect 33508 16099 33560 16108
rect 33508 16065 33517 16099
rect 33517 16065 33551 16099
rect 33551 16065 33560 16099
rect 33508 16056 33560 16065
rect 34244 16056 34296 16108
rect 37464 16099 37516 16108
rect 37464 16065 37473 16099
rect 37473 16065 37507 16099
rect 37507 16065 37516 16099
rect 37464 16056 37516 16065
rect 45836 16124 45888 16176
rect 46572 16124 46624 16176
rect 22376 15920 22428 15972
rect 31484 15988 31536 16040
rect 23664 15920 23716 15972
rect 26884 15920 26936 15972
rect 33600 15988 33652 16040
rect 38936 15988 38988 16040
rect 39212 16099 39264 16108
rect 39212 16065 39221 16099
rect 39221 16065 39255 16099
rect 39255 16065 39264 16099
rect 39212 16056 39264 16065
rect 39396 16099 39448 16108
rect 39396 16065 39405 16099
rect 39405 16065 39439 16099
rect 39439 16065 39448 16099
rect 40500 16099 40552 16108
rect 39396 16056 39448 16065
rect 40500 16065 40509 16099
rect 40509 16065 40543 16099
rect 40543 16065 40552 16099
rect 40500 16056 40552 16065
rect 41052 16056 41104 16108
rect 41788 16056 41840 16108
rect 42616 16099 42668 16108
rect 42616 16065 42625 16099
rect 42625 16065 42659 16099
rect 42659 16065 42668 16099
rect 42616 16056 42668 16065
rect 42156 15988 42208 16040
rect 38384 15920 38436 15972
rect 47308 16056 47360 16108
rect 47400 16056 47452 16108
rect 23756 15852 23808 15904
rect 26792 15852 26844 15904
rect 30656 15852 30708 15904
rect 31668 15852 31720 15904
rect 34152 15852 34204 15904
rect 39672 15852 39724 15904
rect 42432 15895 42484 15904
rect 42432 15861 42441 15895
rect 42441 15861 42475 15895
rect 42475 15861 42484 15895
rect 42432 15852 42484 15861
rect 46296 15852 46348 15904
rect 46480 15852 46532 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 4620 15648 4672 15700
rect 14188 15691 14240 15700
rect 14188 15657 14197 15691
rect 14197 15657 14231 15691
rect 14231 15657 14240 15691
rect 14188 15648 14240 15657
rect 15752 15648 15804 15700
rect 17684 15648 17736 15700
rect 19892 15648 19944 15700
rect 20260 15648 20312 15700
rect 30564 15648 30616 15700
rect 31944 15691 31996 15700
rect 23664 15580 23716 15632
rect 24216 15580 24268 15632
rect 26700 15580 26752 15632
rect 17868 15512 17920 15564
rect 18144 15555 18196 15564
rect 18144 15521 18153 15555
rect 18153 15521 18187 15555
rect 18187 15521 18196 15555
rect 18144 15512 18196 15521
rect 20996 15512 21048 15564
rect 21640 15512 21692 15564
rect 22284 15512 22336 15564
rect 24952 15512 25004 15564
rect 13268 15444 13320 15496
rect 14096 15487 14148 15496
rect 14096 15453 14105 15487
rect 14105 15453 14139 15487
rect 14139 15453 14148 15487
rect 14096 15444 14148 15453
rect 15384 15487 15436 15496
rect 15384 15453 15393 15487
rect 15393 15453 15427 15487
rect 15427 15453 15436 15487
rect 15384 15444 15436 15453
rect 16580 15444 16632 15496
rect 19248 15444 19300 15496
rect 16580 15308 16632 15360
rect 21456 15376 21508 15428
rect 21824 15419 21876 15428
rect 21824 15385 21833 15419
rect 21833 15385 21867 15419
rect 21867 15385 21876 15419
rect 21824 15376 21876 15385
rect 22560 15444 22612 15496
rect 22744 15487 22796 15496
rect 22744 15453 22778 15487
rect 22778 15453 22796 15487
rect 22744 15444 22796 15453
rect 24400 15487 24452 15496
rect 24400 15453 24409 15487
rect 24409 15453 24443 15487
rect 24443 15453 24452 15487
rect 24400 15444 24452 15453
rect 24584 15487 24636 15496
rect 24584 15453 24593 15487
rect 24593 15453 24627 15487
rect 24627 15453 24636 15487
rect 25780 15512 25832 15564
rect 26148 15512 26200 15564
rect 24584 15444 24636 15453
rect 26240 15444 26292 15496
rect 26884 15376 26936 15428
rect 20260 15308 20312 15360
rect 20352 15351 20404 15360
rect 20352 15317 20361 15351
rect 20361 15317 20395 15351
rect 20395 15317 20404 15351
rect 20352 15308 20404 15317
rect 22192 15308 22244 15360
rect 23204 15308 23256 15360
rect 23848 15351 23900 15360
rect 23848 15317 23857 15351
rect 23857 15317 23891 15351
rect 23891 15317 23900 15351
rect 23848 15308 23900 15317
rect 24584 15308 24636 15360
rect 25780 15308 25832 15360
rect 25964 15351 26016 15360
rect 25964 15317 25973 15351
rect 25973 15317 26007 15351
rect 26007 15317 26016 15351
rect 25964 15308 26016 15317
rect 26424 15351 26476 15360
rect 26424 15317 26433 15351
rect 26433 15317 26467 15351
rect 26467 15317 26476 15351
rect 26424 15308 26476 15317
rect 29552 15444 29604 15496
rect 30564 15487 30616 15496
rect 30564 15453 30573 15487
rect 30573 15453 30607 15487
rect 30607 15453 30616 15487
rect 30564 15444 30616 15453
rect 30656 15444 30708 15496
rect 28264 15376 28316 15428
rect 30104 15376 30156 15428
rect 31944 15657 31953 15691
rect 31953 15657 31987 15691
rect 31987 15657 31996 15691
rect 31944 15648 31996 15657
rect 39212 15648 39264 15700
rect 38936 15580 38988 15632
rect 40132 15512 40184 15564
rect 46296 15555 46348 15564
rect 46296 15521 46305 15555
rect 46305 15521 46339 15555
rect 46339 15521 46348 15555
rect 46296 15512 46348 15521
rect 46480 15555 46532 15564
rect 46480 15521 46489 15555
rect 46489 15521 46523 15555
rect 46523 15521 46532 15555
rect 46480 15512 46532 15521
rect 48136 15555 48188 15564
rect 48136 15521 48145 15555
rect 48145 15521 48179 15555
rect 48179 15521 48188 15555
rect 48136 15512 48188 15521
rect 34704 15419 34756 15428
rect 34704 15385 34713 15419
rect 34713 15385 34747 15419
rect 34747 15385 34756 15419
rect 34704 15376 34756 15385
rect 29000 15351 29052 15360
rect 29000 15317 29009 15351
rect 29009 15317 29043 15351
rect 29043 15317 29052 15351
rect 29000 15308 29052 15317
rect 30656 15308 30708 15360
rect 35716 15376 35768 15428
rect 35348 15308 35400 15360
rect 36728 15308 36780 15360
rect 37188 15444 37240 15496
rect 37924 15419 37976 15428
rect 37924 15385 37933 15419
rect 37933 15385 37967 15419
rect 37967 15385 37976 15419
rect 37924 15376 37976 15385
rect 38844 15419 38896 15428
rect 38844 15385 38853 15419
rect 38853 15385 38887 15419
rect 38887 15385 38896 15419
rect 38844 15376 38896 15385
rect 42432 15444 42484 15496
rect 42708 15376 42760 15428
rect 40500 15308 40552 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 1676 15104 1728 15156
rect 17684 15036 17736 15088
rect 20076 15036 20128 15088
rect 20628 15036 20680 15088
rect 21456 15036 21508 15088
rect 15844 14968 15896 15020
rect 21180 14968 21232 15020
rect 23204 15011 23256 15020
rect 16948 14900 17000 14952
rect 18236 14943 18288 14952
rect 18236 14909 18245 14943
rect 18245 14909 18279 14943
rect 18279 14909 18288 14943
rect 18236 14900 18288 14909
rect 21916 14900 21968 14952
rect 23204 14977 23213 15011
rect 23213 14977 23247 15011
rect 23247 14977 23256 15011
rect 23204 14968 23256 14977
rect 23848 15036 23900 15088
rect 4068 14832 4120 14884
rect 18052 14832 18104 14884
rect 21456 14832 21508 14884
rect 22008 14832 22060 14884
rect 24400 14968 24452 15020
rect 25136 15104 25188 15156
rect 27068 15104 27120 15156
rect 27252 15036 27304 15088
rect 23388 14900 23440 14952
rect 25228 14900 25280 14952
rect 25780 14968 25832 15020
rect 27528 15104 27580 15156
rect 29000 15036 29052 15088
rect 30104 15079 30156 15088
rect 30104 15045 30113 15079
rect 30113 15045 30147 15079
rect 30147 15045 30156 15079
rect 30104 15036 30156 15045
rect 30748 15104 30800 15156
rect 46204 15104 46256 15156
rect 46388 15104 46440 15156
rect 31024 15036 31076 15088
rect 31484 15036 31536 15088
rect 28172 14968 28224 15020
rect 28816 14968 28868 15020
rect 26240 14900 26292 14952
rect 27252 14900 27304 14952
rect 28356 14900 28408 14952
rect 28724 14943 28776 14952
rect 28724 14909 28733 14943
rect 28733 14909 28767 14943
rect 28767 14909 28776 14943
rect 28724 14900 28776 14909
rect 30380 14900 30432 14952
rect 31392 15011 31444 15020
rect 35440 15036 35492 15088
rect 31392 14977 31406 15011
rect 31406 14977 31440 15011
rect 31440 14977 31444 15011
rect 31392 14968 31444 14977
rect 31668 14968 31720 15020
rect 34152 14968 34204 15020
rect 34612 15011 34664 15020
rect 34612 14977 34646 15011
rect 34646 14977 34664 15011
rect 40132 15036 40184 15088
rect 34612 14968 34664 14977
rect 35716 14875 35768 14884
rect 35716 14841 35725 14875
rect 35725 14841 35759 14875
rect 35759 14841 35768 14875
rect 35716 14832 35768 14841
rect 39672 14968 39724 15020
rect 46848 14968 46900 15020
rect 37924 14900 37976 14952
rect 39028 14943 39080 14952
rect 39028 14909 39037 14943
rect 39037 14909 39071 14943
rect 39071 14909 39080 14943
rect 39028 14900 39080 14909
rect 38384 14832 38436 14884
rect 20076 14764 20128 14816
rect 21640 14764 21692 14816
rect 22192 14764 22244 14816
rect 23296 14764 23348 14816
rect 24032 14764 24084 14816
rect 26148 14807 26200 14816
rect 26148 14773 26157 14807
rect 26157 14773 26191 14807
rect 26191 14773 26200 14807
rect 26148 14764 26200 14773
rect 26424 14807 26476 14816
rect 26424 14773 26433 14807
rect 26433 14773 26467 14807
rect 26467 14773 26476 14807
rect 26424 14764 26476 14773
rect 28724 14807 28776 14816
rect 28724 14773 28733 14807
rect 28733 14773 28767 14807
rect 28767 14773 28776 14807
rect 28724 14764 28776 14773
rect 29092 14807 29144 14816
rect 29092 14773 29101 14807
rect 29101 14773 29135 14807
rect 29135 14773 29144 14807
rect 29092 14764 29144 14773
rect 31208 14764 31260 14816
rect 33416 14764 33468 14816
rect 38844 14764 38896 14816
rect 47768 14807 47820 14816
rect 47768 14773 47777 14807
rect 47777 14773 47811 14807
rect 47811 14773 47820 14807
rect 47768 14764 47820 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 16764 14560 16816 14612
rect 17960 14424 18012 14476
rect 18880 14424 18932 14476
rect 21364 14560 21416 14612
rect 25872 14560 25924 14612
rect 26700 14603 26752 14612
rect 26700 14569 26709 14603
rect 26709 14569 26743 14603
rect 26743 14569 26752 14603
rect 26700 14560 26752 14569
rect 20352 14492 20404 14544
rect 21456 14492 21508 14544
rect 21640 14492 21692 14544
rect 23480 14492 23532 14544
rect 29092 14560 29144 14612
rect 31392 14560 31444 14612
rect 34612 14560 34664 14612
rect 22284 14424 22336 14476
rect 23848 14424 23900 14476
rect 26148 14424 26200 14476
rect 1768 14356 1820 14408
rect 16580 14356 16632 14408
rect 17684 14399 17736 14408
rect 17684 14365 17693 14399
rect 17693 14365 17727 14399
rect 17727 14365 17736 14399
rect 17684 14356 17736 14365
rect 21824 14356 21876 14408
rect 22192 14356 22244 14408
rect 23112 14356 23164 14408
rect 25780 14399 25832 14408
rect 18604 14288 18656 14340
rect 20076 14288 20128 14340
rect 21364 14288 21416 14340
rect 25780 14365 25789 14399
rect 25789 14365 25823 14399
rect 25823 14365 25832 14399
rect 25780 14356 25832 14365
rect 25964 14356 26016 14408
rect 26424 14399 26476 14408
rect 26424 14365 26433 14399
rect 26433 14365 26467 14399
rect 26467 14365 26476 14399
rect 26424 14356 26476 14365
rect 26700 14399 26752 14408
rect 26700 14365 26709 14399
rect 26709 14365 26743 14399
rect 26743 14365 26752 14399
rect 26700 14356 26752 14365
rect 27068 14492 27120 14544
rect 27988 14492 28040 14544
rect 28172 14492 28224 14544
rect 31208 14492 31260 14544
rect 33140 14492 33192 14544
rect 33508 14492 33560 14544
rect 34152 14535 34204 14544
rect 34152 14501 34161 14535
rect 34161 14501 34195 14535
rect 34195 14501 34204 14535
rect 34152 14492 34204 14501
rect 27344 14424 27396 14476
rect 29000 14424 29052 14476
rect 31116 14424 31168 14476
rect 34428 14424 34480 14476
rect 37924 14560 37976 14612
rect 27896 14399 27948 14408
rect 26240 14288 26292 14340
rect 27896 14365 27905 14399
rect 27905 14365 27939 14399
rect 27939 14365 27948 14399
rect 27896 14356 27948 14365
rect 28172 14356 28224 14408
rect 28264 14399 28316 14408
rect 28264 14365 28273 14399
rect 28273 14365 28307 14399
rect 28307 14365 28316 14399
rect 28264 14356 28316 14365
rect 29092 14356 29144 14408
rect 34888 14356 34940 14408
rect 37464 14424 37516 14476
rect 44272 14424 44324 14476
rect 47768 14424 47820 14476
rect 35164 14396 35216 14408
rect 35164 14362 35178 14396
rect 35178 14362 35212 14396
rect 35212 14362 35216 14396
rect 35164 14356 35216 14362
rect 35440 14356 35492 14408
rect 36728 14399 36780 14408
rect 36728 14365 36762 14399
rect 36762 14365 36780 14399
rect 36728 14356 36780 14365
rect 38384 14399 38436 14408
rect 38384 14365 38393 14399
rect 38393 14365 38427 14399
rect 38427 14365 38436 14399
rect 38384 14356 38436 14365
rect 30380 14288 30432 14340
rect 22652 14220 22704 14272
rect 22744 14220 22796 14272
rect 23388 14220 23440 14272
rect 24400 14220 24452 14272
rect 27712 14220 27764 14272
rect 28172 14220 28224 14272
rect 31208 14288 31260 14340
rect 33048 14288 33100 14340
rect 38292 14288 38344 14340
rect 33508 14220 33560 14272
rect 34704 14220 34756 14272
rect 35440 14220 35492 14272
rect 38476 14263 38528 14272
rect 38476 14229 38485 14263
rect 38485 14229 38519 14263
rect 38519 14229 38528 14263
rect 38476 14220 38528 14229
rect 46756 14288 46808 14340
rect 48136 14331 48188 14340
rect 48136 14297 48145 14331
rect 48145 14297 48179 14331
rect 48179 14297 48188 14331
rect 48136 14288 48188 14297
rect 47216 14220 47268 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 20076 14059 20128 14068
rect 20076 14025 20085 14059
rect 20085 14025 20119 14059
rect 20119 14025 20128 14059
rect 20076 14016 20128 14025
rect 21180 14059 21232 14068
rect 21180 14025 21189 14059
rect 21189 14025 21223 14059
rect 21223 14025 21232 14059
rect 21180 14016 21232 14025
rect 21824 14016 21876 14068
rect 25964 13948 26016 14000
rect 1768 13923 1820 13932
rect 1768 13889 1777 13923
rect 1777 13889 1811 13923
rect 1811 13889 1820 13923
rect 1768 13880 1820 13889
rect 15844 13880 15896 13932
rect 17684 13923 17736 13932
rect 17684 13889 17693 13923
rect 17693 13889 17727 13923
rect 17727 13889 17736 13923
rect 17684 13880 17736 13889
rect 20260 13923 20312 13932
rect 20260 13889 20269 13923
rect 20269 13889 20303 13923
rect 20303 13889 20312 13923
rect 20260 13880 20312 13889
rect 1952 13855 2004 13864
rect 1952 13821 1961 13855
rect 1961 13821 1995 13855
rect 1995 13821 2004 13855
rect 1952 13812 2004 13821
rect 2780 13855 2832 13864
rect 2780 13821 2789 13855
rect 2789 13821 2823 13855
rect 2823 13821 2832 13855
rect 2780 13812 2832 13821
rect 14096 13812 14148 13864
rect 18052 13855 18104 13864
rect 18052 13821 18061 13855
rect 18061 13821 18095 13855
rect 18095 13821 18104 13855
rect 18052 13812 18104 13821
rect 18420 13812 18472 13864
rect 3056 13744 3108 13796
rect 18144 13744 18196 13796
rect 21640 13880 21692 13932
rect 21916 13880 21968 13932
rect 24308 13880 24360 13932
rect 24400 13923 24452 13932
rect 24400 13889 24409 13923
rect 24409 13889 24443 13923
rect 24443 13889 24452 13923
rect 25320 13923 25372 13932
rect 24400 13880 24452 13889
rect 25320 13889 25329 13923
rect 25329 13889 25363 13923
rect 25363 13889 25372 13923
rect 25320 13880 25372 13889
rect 25780 13880 25832 13932
rect 27988 14016 28040 14068
rect 46756 14059 46808 14068
rect 31576 13948 31628 14000
rect 33140 13948 33192 14000
rect 33508 13991 33560 14000
rect 33508 13957 33517 13991
rect 33517 13957 33551 13991
rect 33551 13957 33560 13991
rect 33508 13948 33560 13957
rect 35348 13948 35400 14000
rect 38476 13991 38528 14000
rect 38476 13957 38485 13991
rect 38485 13957 38519 13991
rect 38519 13957 38528 13991
rect 38476 13948 38528 13957
rect 46756 14025 46765 14059
rect 46765 14025 46799 14059
rect 46799 14025 46808 14059
rect 46756 14016 46808 14025
rect 21456 13812 21508 13864
rect 22284 13855 22336 13864
rect 22284 13821 22293 13855
rect 22293 13821 22327 13855
rect 22327 13821 22336 13855
rect 22284 13812 22336 13821
rect 22008 13744 22060 13796
rect 23480 13744 23532 13796
rect 26240 13812 26292 13864
rect 24584 13787 24636 13796
rect 24584 13753 24593 13787
rect 24593 13753 24627 13787
rect 24627 13753 24636 13787
rect 24584 13744 24636 13753
rect 16856 13676 16908 13728
rect 20536 13676 20588 13728
rect 21180 13676 21232 13728
rect 21364 13676 21416 13728
rect 22560 13676 22612 13728
rect 24952 13676 25004 13728
rect 25504 13719 25556 13728
rect 25504 13685 25513 13719
rect 25513 13685 25547 13719
rect 25547 13685 25556 13719
rect 25504 13676 25556 13685
rect 26700 13744 26752 13796
rect 26148 13676 26200 13728
rect 28356 13812 28408 13864
rect 29092 13855 29144 13864
rect 29092 13821 29101 13855
rect 29101 13821 29135 13855
rect 29135 13821 29144 13855
rect 29092 13812 29144 13821
rect 29828 13812 29880 13864
rect 30380 13855 30432 13864
rect 30380 13821 30389 13855
rect 30389 13821 30423 13855
rect 30423 13821 30432 13855
rect 30380 13812 30432 13821
rect 33324 13880 33376 13932
rect 32220 13812 32272 13864
rect 33048 13855 33100 13864
rect 33048 13821 33057 13855
rect 33057 13821 33091 13855
rect 33091 13821 33100 13855
rect 33048 13812 33100 13821
rect 27988 13744 28040 13796
rect 31024 13744 31076 13796
rect 34520 13880 34572 13932
rect 34428 13812 34480 13864
rect 35256 13880 35308 13932
rect 35440 13923 35492 13932
rect 35440 13889 35449 13923
rect 35449 13889 35483 13923
rect 35483 13889 35492 13923
rect 35440 13880 35492 13889
rect 46204 13880 46256 13932
rect 47860 13923 47912 13932
rect 47860 13889 47869 13923
rect 47869 13889 47903 13923
rect 47903 13889 47912 13923
rect 47860 13880 47912 13889
rect 35808 13855 35860 13864
rect 35808 13821 35817 13855
rect 35817 13821 35851 13855
rect 35851 13821 35860 13855
rect 35808 13812 35860 13821
rect 38844 13812 38896 13864
rect 39948 13855 40000 13864
rect 39948 13821 39957 13855
rect 39957 13821 39991 13855
rect 39991 13821 40000 13855
rect 39948 13812 40000 13821
rect 35624 13744 35676 13796
rect 28724 13676 28776 13728
rect 32496 13676 32548 13728
rect 34520 13676 34572 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 1952 13472 2004 13524
rect 16764 13472 16816 13524
rect 18144 13472 18196 13524
rect 21824 13472 21876 13524
rect 22008 13472 22060 13524
rect 23296 13472 23348 13524
rect 23572 13515 23624 13524
rect 23572 13481 23581 13515
rect 23581 13481 23615 13515
rect 23615 13481 23624 13515
rect 23572 13472 23624 13481
rect 24216 13472 24268 13524
rect 1584 13336 1636 13388
rect 2044 13311 2096 13320
rect 2044 13277 2053 13311
rect 2053 13277 2087 13311
rect 2087 13277 2096 13311
rect 2044 13268 2096 13277
rect 19156 13336 19208 13388
rect 19340 13336 19392 13388
rect 21640 13336 21692 13388
rect 22284 13336 22336 13388
rect 18052 13175 18104 13184
rect 18052 13141 18061 13175
rect 18061 13141 18095 13175
rect 18095 13141 18104 13175
rect 18052 13132 18104 13141
rect 18512 13311 18564 13320
rect 18512 13277 18521 13311
rect 18521 13277 18555 13311
rect 18555 13277 18564 13311
rect 18512 13268 18564 13277
rect 19432 13268 19484 13320
rect 22008 13268 22060 13320
rect 22100 13311 22152 13320
rect 22100 13277 22109 13311
rect 22109 13277 22143 13311
rect 22143 13277 22152 13311
rect 22376 13311 22428 13320
rect 22100 13268 22152 13277
rect 22376 13277 22385 13311
rect 22385 13277 22419 13311
rect 22419 13277 22428 13311
rect 22376 13268 22428 13277
rect 27436 13472 27488 13524
rect 30564 13472 30616 13524
rect 31668 13472 31720 13524
rect 23296 13336 23348 13388
rect 23848 13336 23900 13388
rect 19340 13200 19392 13252
rect 22192 13200 22244 13252
rect 24768 13268 24820 13320
rect 22652 13132 22704 13184
rect 24216 13200 24268 13252
rect 24584 13200 24636 13252
rect 26148 13336 26200 13388
rect 26240 13268 26292 13320
rect 27436 13311 27488 13320
rect 27436 13277 27445 13311
rect 27445 13277 27479 13311
rect 27479 13277 27488 13311
rect 27436 13268 27488 13277
rect 24400 13175 24452 13184
rect 24400 13141 24409 13175
rect 24409 13141 24443 13175
rect 24443 13141 24452 13175
rect 24400 13132 24452 13141
rect 24492 13132 24544 13184
rect 27620 13132 27672 13184
rect 28172 13336 28224 13388
rect 31116 13336 31168 13388
rect 31852 13336 31904 13388
rect 32312 13379 32364 13388
rect 32312 13345 32321 13379
rect 32321 13345 32355 13379
rect 32355 13345 32364 13379
rect 32312 13336 32364 13345
rect 32496 13379 32548 13388
rect 32496 13345 32505 13379
rect 32505 13345 32539 13379
rect 32539 13345 32548 13379
rect 32496 13336 32548 13345
rect 33692 13379 33744 13388
rect 33692 13345 33701 13379
rect 33701 13345 33735 13379
rect 33735 13345 33744 13379
rect 33692 13336 33744 13345
rect 34152 13336 34204 13388
rect 27988 13311 28040 13320
rect 27988 13277 27997 13311
rect 27997 13277 28031 13311
rect 28031 13277 28040 13311
rect 27988 13268 28040 13277
rect 30012 13268 30064 13320
rect 32220 13268 32272 13320
rect 28540 13200 28592 13252
rect 28724 13200 28776 13252
rect 31576 13200 31628 13252
rect 28172 13175 28224 13184
rect 28172 13141 28181 13175
rect 28181 13141 28215 13175
rect 28215 13141 28224 13175
rect 28172 13132 28224 13141
rect 34704 13200 34756 13252
rect 35348 13132 35400 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 1584 12971 1636 12980
rect 1584 12937 1593 12971
rect 1593 12937 1627 12971
rect 1627 12937 1636 12971
rect 1584 12928 1636 12937
rect 2044 12928 2096 12980
rect 18604 12928 18656 12980
rect 21640 12928 21692 12980
rect 24308 12928 24360 12980
rect 27988 12928 28040 12980
rect 28816 12928 28868 12980
rect 16856 12903 16908 12912
rect 16856 12869 16865 12903
rect 16865 12869 16899 12903
rect 16899 12869 16908 12903
rect 16856 12860 16908 12869
rect 18144 12860 18196 12912
rect 1400 12835 1452 12844
rect 1400 12801 1409 12835
rect 1409 12801 1443 12835
rect 1443 12801 1452 12835
rect 1400 12792 1452 12801
rect 19156 12792 19208 12844
rect 3516 12724 3568 12776
rect 16672 12767 16724 12776
rect 16672 12733 16681 12767
rect 16681 12733 16715 12767
rect 16715 12733 16724 12767
rect 16672 12724 16724 12733
rect 18972 12724 19024 12776
rect 21640 12792 21692 12844
rect 22008 12835 22060 12844
rect 22008 12801 22017 12835
rect 22017 12801 22051 12835
rect 22051 12801 22060 12835
rect 22008 12792 22060 12801
rect 25504 12860 25556 12912
rect 29092 12860 29144 12912
rect 22652 12792 22704 12844
rect 26240 12792 26292 12844
rect 28172 12792 28224 12844
rect 32036 12860 32088 12912
rect 34520 12860 34572 12912
rect 31668 12792 31720 12844
rect 32220 12792 32272 12844
rect 34152 12792 34204 12844
rect 20260 12724 20312 12776
rect 21824 12724 21876 12776
rect 22836 12724 22888 12776
rect 24860 12724 24912 12776
rect 25688 12724 25740 12776
rect 26700 12724 26752 12776
rect 20628 12656 20680 12708
rect 20904 12656 20956 12708
rect 19432 12588 19484 12640
rect 19708 12588 19760 12640
rect 20720 12631 20772 12640
rect 20720 12597 20729 12631
rect 20729 12597 20763 12631
rect 20763 12597 20772 12631
rect 20720 12588 20772 12597
rect 23204 12656 23256 12708
rect 24952 12656 25004 12708
rect 32128 12656 32180 12708
rect 24400 12588 24452 12640
rect 24584 12588 24636 12640
rect 25412 12588 25464 12640
rect 26792 12588 26844 12640
rect 27252 12588 27304 12640
rect 27620 12588 27672 12640
rect 28264 12588 28316 12640
rect 32312 12588 32364 12640
rect 35624 12588 35676 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 16672 12384 16724 12436
rect 18512 12384 18564 12436
rect 20720 12384 20772 12436
rect 21640 12427 21692 12436
rect 21640 12393 21649 12427
rect 21649 12393 21683 12427
rect 21683 12393 21692 12427
rect 21640 12384 21692 12393
rect 22928 12427 22980 12436
rect 22928 12393 22937 12427
rect 22937 12393 22971 12427
rect 22971 12393 22980 12427
rect 22928 12384 22980 12393
rect 24584 12384 24636 12436
rect 26240 12384 26292 12436
rect 32220 12384 32272 12436
rect 34704 12427 34756 12436
rect 34704 12393 34713 12427
rect 34713 12393 34747 12427
rect 34747 12393 34756 12427
rect 34704 12384 34756 12393
rect 44732 12384 44784 12436
rect 46848 12384 46900 12436
rect 19248 12316 19300 12368
rect 20352 12316 20404 12368
rect 17960 12180 18012 12232
rect 19156 12180 19208 12232
rect 18052 12112 18104 12164
rect 19708 12112 19760 12164
rect 20352 12112 20404 12164
rect 29276 12316 29328 12368
rect 23572 12248 23624 12300
rect 27344 12248 27396 12300
rect 22100 12223 22152 12232
rect 22100 12189 22109 12223
rect 22109 12189 22143 12223
rect 22143 12189 22152 12223
rect 22100 12180 22152 12189
rect 22376 12180 22428 12232
rect 22836 12223 22888 12232
rect 22836 12189 22845 12223
rect 22845 12189 22879 12223
rect 22879 12189 22888 12223
rect 22836 12180 22888 12189
rect 23296 12180 23348 12232
rect 23756 12180 23808 12232
rect 24952 12180 25004 12232
rect 25320 12155 25372 12164
rect 25320 12121 25329 12155
rect 25329 12121 25363 12155
rect 25363 12121 25372 12155
rect 25320 12112 25372 12121
rect 25504 12223 25556 12232
rect 25504 12189 25513 12223
rect 25513 12189 25547 12223
rect 25547 12189 25556 12223
rect 25504 12180 25556 12189
rect 25780 12180 25832 12232
rect 27620 12180 27672 12232
rect 28632 12180 28684 12232
rect 30840 12180 30892 12232
rect 31576 12223 31628 12232
rect 31576 12189 31585 12223
rect 31585 12189 31619 12223
rect 31619 12189 31628 12223
rect 31576 12180 31628 12189
rect 34428 12248 34480 12300
rect 28264 12112 28316 12164
rect 31300 12112 31352 12164
rect 19340 12044 19392 12096
rect 22376 12044 22428 12096
rect 23388 12087 23440 12096
rect 23388 12053 23397 12087
rect 23397 12053 23431 12087
rect 23431 12053 23440 12087
rect 23388 12044 23440 12053
rect 25688 12044 25740 12096
rect 28172 12044 28224 12096
rect 32312 12180 32364 12232
rect 32680 12180 32732 12232
rect 33324 12180 33376 12232
rect 35808 12248 35860 12300
rect 32128 12112 32180 12164
rect 35532 12180 35584 12232
rect 35900 12223 35952 12232
rect 35900 12189 35909 12223
rect 35909 12189 35943 12223
rect 35943 12189 35952 12223
rect 35900 12180 35952 12189
rect 36176 12180 36228 12232
rect 44824 12112 44876 12164
rect 33140 12044 33192 12096
rect 33324 12087 33376 12096
rect 33324 12053 33333 12087
rect 33333 12053 33367 12087
rect 33367 12053 33376 12087
rect 33324 12044 33376 12053
rect 36084 12087 36136 12096
rect 36084 12053 36093 12087
rect 36093 12053 36127 12087
rect 36127 12053 36136 12087
rect 36084 12044 36136 12053
rect 37188 12044 37240 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 19156 11883 19208 11892
rect 19156 11849 19165 11883
rect 19165 11849 19199 11883
rect 19199 11849 19208 11883
rect 19156 11840 19208 11849
rect 22192 11840 22244 11892
rect 24952 11840 25004 11892
rect 26700 11840 26752 11892
rect 28632 11840 28684 11892
rect 29276 11840 29328 11892
rect 36084 11840 36136 11892
rect 15936 11704 15988 11756
rect 19432 11704 19484 11756
rect 20352 11772 20404 11824
rect 17592 11636 17644 11688
rect 20076 11747 20128 11756
rect 20076 11713 20085 11747
rect 20085 11713 20119 11747
rect 20119 11713 20128 11747
rect 20076 11704 20128 11713
rect 23388 11772 23440 11824
rect 23756 11772 23808 11824
rect 24124 11772 24176 11824
rect 28172 11772 28224 11824
rect 31024 11772 31076 11824
rect 21916 11704 21968 11756
rect 22100 11747 22152 11756
rect 22100 11713 22109 11747
rect 22109 11713 22143 11747
rect 22143 11713 22152 11747
rect 22376 11747 22428 11756
rect 22100 11704 22152 11713
rect 22376 11713 22385 11747
rect 22385 11713 22419 11747
rect 22419 11713 22428 11747
rect 22376 11704 22428 11713
rect 23204 11747 23256 11756
rect 23204 11713 23213 11747
rect 23213 11713 23247 11747
rect 23247 11713 23256 11747
rect 23204 11704 23256 11713
rect 23480 11747 23532 11756
rect 23480 11713 23489 11747
rect 23489 11713 23523 11747
rect 23523 11713 23532 11747
rect 23480 11704 23532 11713
rect 24492 11704 24544 11756
rect 25688 11747 25740 11756
rect 25688 11713 25697 11747
rect 25697 11713 25731 11747
rect 25731 11713 25740 11747
rect 25688 11704 25740 11713
rect 28080 11747 28132 11756
rect 28080 11713 28114 11747
rect 28114 11713 28132 11747
rect 28080 11704 28132 11713
rect 29736 11704 29788 11756
rect 30288 11747 30340 11756
rect 30288 11713 30297 11747
rect 30297 11713 30331 11747
rect 30331 11713 30340 11747
rect 30288 11704 30340 11713
rect 31300 11747 31352 11756
rect 31300 11713 31309 11747
rect 31309 11713 31343 11747
rect 31343 11713 31352 11747
rect 31300 11704 31352 11713
rect 33324 11815 33376 11824
rect 33324 11781 33333 11815
rect 33333 11781 33367 11815
rect 33367 11781 33376 11815
rect 33324 11772 33376 11781
rect 32128 11747 32180 11756
rect 20352 11636 20404 11688
rect 22192 11679 22244 11688
rect 22192 11645 22201 11679
rect 22201 11645 22235 11679
rect 22235 11645 22244 11679
rect 22192 11636 22244 11645
rect 24400 11636 24452 11688
rect 25964 11679 26016 11688
rect 25964 11645 25973 11679
rect 25973 11645 26007 11679
rect 26007 11645 26016 11679
rect 25964 11636 26016 11645
rect 27436 11636 27488 11688
rect 32128 11713 32137 11747
rect 32137 11713 32171 11747
rect 32171 11713 32180 11747
rect 32128 11704 32180 11713
rect 32864 11704 32916 11756
rect 34336 11679 34388 11688
rect 34336 11645 34345 11679
rect 34345 11645 34379 11679
rect 34379 11645 34388 11679
rect 34336 11636 34388 11645
rect 31484 11568 31536 11620
rect 1584 11500 1636 11552
rect 21364 11500 21416 11552
rect 22836 11500 22888 11552
rect 23756 11500 23808 11552
rect 24032 11500 24084 11552
rect 25504 11500 25556 11552
rect 25872 11543 25924 11552
rect 25872 11509 25881 11543
rect 25881 11509 25915 11543
rect 25915 11509 25924 11543
rect 25872 11500 25924 11509
rect 31760 11500 31812 11552
rect 46296 11500 46348 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 20076 11296 20128 11348
rect 22100 11296 22152 11348
rect 23848 11296 23900 11348
rect 24032 11296 24084 11348
rect 28080 11296 28132 11348
rect 28264 11296 28316 11348
rect 46572 11296 46624 11348
rect 1584 11203 1636 11212
rect 1584 11169 1593 11203
rect 1593 11169 1627 11203
rect 1627 11169 1636 11203
rect 1584 11160 1636 11169
rect 2780 11203 2832 11212
rect 2780 11169 2789 11203
rect 2789 11169 2823 11203
rect 2823 11169 2832 11203
rect 2780 11160 2832 11169
rect 23388 11160 23440 11212
rect 27620 11228 27672 11280
rect 32864 11271 32916 11280
rect 32864 11237 32873 11271
rect 32873 11237 32907 11271
rect 32907 11237 32916 11271
rect 32864 11228 32916 11237
rect 19156 11092 19208 11144
rect 21824 11092 21876 11144
rect 23204 11092 23256 11144
rect 26056 11092 26108 11144
rect 27252 11135 27304 11144
rect 27252 11101 27261 11135
rect 27261 11101 27295 11135
rect 27295 11101 27304 11135
rect 27252 11092 27304 11101
rect 27620 11135 27672 11144
rect 2320 11024 2372 11076
rect 19340 11024 19392 11076
rect 21364 11024 21416 11076
rect 23388 11024 23440 11076
rect 24584 11067 24636 11076
rect 24584 11033 24593 11067
rect 24593 11033 24627 11067
rect 24627 11033 24636 11067
rect 24584 11024 24636 11033
rect 24860 11024 24912 11076
rect 25964 11024 26016 11076
rect 27620 11101 27629 11135
rect 27629 11101 27663 11135
rect 27663 11101 27672 11135
rect 27620 11092 27672 11101
rect 28172 11160 28224 11212
rect 46296 11203 46348 11212
rect 46296 11169 46305 11203
rect 46305 11169 46339 11203
rect 46339 11169 46348 11203
rect 46296 11160 46348 11169
rect 27896 11092 27948 11144
rect 30012 11135 30064 11144
rect 30012 11101 30021 11135
rect 30021 11101 30055 11135
rect 30055 11101 30064 11135
rect 30012 11092 30064 11101
rect 31576 11092 31628 11144
rect 31760 11135 31812 11144
rect 31760 11101 31794 11135
rect 31794 11101 31812 11135
rect 31760 11092 31812 11101
rect 27712 11024 27764 11076
rect 28724 11067 28776 11076
rect 28724 11033 28733 11067
rect 28733 11033 28767 11067
rect 28767 11033 28776 11067
rect 28724 11024 28776 11033
rect 30288 11024 30340 11076
rect 35900 11024 35952 11076
rect 46940 11024 46992 11076
rect 48136 11067 48188 11076
rect 48136 11033 48145 11067
rect 48145 11033 48179 11067
rect 48179 11033 48188 11067
rect 48136 11024 48188 11033
rect 18788 10956 18840 11008
rect 23480 10956 23532 11008
rect 25044 10956 25096 11008
rect 29000 10956 29052 11008
rect 30196 10956 30248 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 23388 10795 23440 10804
rect 23388 10761 23397 10795
rect 23397 10761 23431 10795
rect 23431 10761 23440 10795
rect 23388 10752 23440 10761
rect 23848 10752 23900 10804
rect 24860 10752 24912 10804
rect 25688 10752 25740 10804
rect 1400 10659 1452 10668
rect 1400 10625 1409 10659
rect 1409 10625 1443 10659
rect 1443 10625 1452 10659
rect 1400 10616 1452 10625
rect 2320 10659 2372 10668
rect 2320 10625 2329 10659
rect 2329 10625 2363 10659
rect 2363 10625 2372 10659
rect 2320 10616 2372 10625
rect 18788 10659 18840 10668
rect 18788 10625 18797 10659
rect 18797 10625 18831 10659
rect 18831 10625 18840 10659
rect 18788 10616 18840 10625
rect 18972 10659 19024 10668
rect 18972 10625 18981 10659
rect 18981 10625 19015 10659
rect 19015 10625 19024 10659
rect 18972 10616 19024 10625
rect 19432 10616 19484 10668
rect 22836 10659 22888 10668
rect 22836 10625 22845 10659
rect 22845 10625 22879 10659
rect 22879 10625 22888 10659
rect 22836 10616 22888 10625
rect 23020 10659 23072 10668
rect 23020 10625 23029 10659
rect 23029 10625 23063 10659
rect 23063 10625 23072 10659
rect 23020 10616 23072 10625
rect 24216 10684 24268 10736
rect 24492 10684 24544 10736
rect 25964 10684 26016 10736
rect 26516 10752 26568 10804
rect 28724 10752 28776 10804
rect 30564 10752 30616 10804
rect 46940 10795 46992 10804
rect 46940 10761 46949 10795
rect 46949 10761 46983 10795
rect 46983 10761 46992 10795
rect 46940 10752 46992 10761
rect 26700 10684 26752 10736
rect 19524 10548 19576 10600
rect 20260 10548 20312 10600
rect 24584 10616 24636 10668
rect 25044 10616 25096 10668
rect 25136 10659 25188 10668
rect 25136 10625 25145 10659
rect 25145 10625 25179 10659
rect 25179 10625 25188 10659
rect 25136 10616 25188 10625
rect 23664 10548 23716 10600
rect 25412 10616 25464 10668
rect 26332 10659 26384 10668
rect 26332 10625 26341 10659
rect 26341 10625 26375 10659
rect 26375 10625 26384 10659
rect 26332 10616 26384 10625
rect 27068 10616 27120 10668
rect 29828 10616 29880 10668
rect 48044 10684 48096 10736
rect 30196 10659 30248 10668
rect 30196 10625 30202 10659
rect 30202 10625 30236 10659
rect 30236 10625 30248 10659
rect 30196 10616 30248 10625
rect 30380 10616 30432 10668
rect 30564 10616 30616 10668
rect 32588 10659 32640 10668
rect 32588 10625 32597 10659
rect 32597 10625 32631 10659
rect 32631 10625 32640 10659
rect 32588 10616 32640 10625
rect 46388 10616 46440 10668
rect 47860 10659 47912 10668
rect 47860 10625 47869 10659
rect 47869 10625 47903 10659
rect 47903 10625 47912 10659
rect 47860 10616 47912 10625
rect 22744 10480 22796 10532
rect 22928 10480 22980 10532
rect 28632 10548 28684 10600
rect 32956 10548 33008 10600
rect 34612 10591 34664 10600
rect 18512 10455 18564 10464
rect 18512 10421 18521 10455
rect 18521 10421 18555 10455
rect 18555 10421 18564 10455
rect 18512 10412 18564 10421
rect 23480 10412 23532 10464
rect 25504 10455 25556 10464
rect 25504 10421 25513 10455
rect 25513 10421 25547 10455
rect 25547 10421 25556 10455
rect 25504 10412 25556 10421
rect 34612 10557 34621 10591
rect 34621 10557 34655 10591
rect 34655 10557 34664 10591
rect 34612 10548 34664 10557
rect 26516 10412 26568 10464
rect 27160 10412 27212 10464
rect 29828 10455 29880 10464
rect 29828 10421 29837 10455
rect 29837 10421 29871 10455
rect 29871 10421 29880 10455
rect 29828 10412 29880 10421
rect 30932 10412 30984 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 23020 10251 23072 10260
rect 23020 10217 23029 10251
rect 23029 10217 23063 10251
rect 23063 10217 23072 10251
rect 23020 10208 23072 10217
rect 24584 10208 24636 10260
rect 24952 10208 25004 10260
rect 25596 10208 25648 10260
rect 26516 10208 26568 10260
rect 28356 10208 28408 10260
rect 30288 10208 30340 10260
rect 32956 10251 33008 10260
rect 32956 10217 32965 10251
rect 32965 10217 32999 10251
rect 32999 10217 33008 10251
rect 32956 10208 33008 10217
rect 19432 10072 19484 10124
rect 20260 10072 20312 10124
rect 1768 10004 1820 10056
rect 17592 10004 17644 10056
rect 19340 10047 19392 10056
rect 19340 10013 19349 10047
rect 19349 10013 19383 10047
rect 19383 10013 19392 10047
rect 19708 10047 19760 10056
rect 19340 10004 19392 10013
rect 19708 10013 19717 10047
rect 19717 10013 19751 10047
rect 19751 10013 19760 10047
rect 19708 10004 19760 10013
rect 23480 10072 23532 10124
rect 25412 10115 25464 10124
rect 25412 10081 25421 10115
rect 25421 10081 25455 10115
rect 25455 10081 25464 10115
rect 25412 10072 25464 10081
rect 23296 10004 23348 10056
rect 24308 10004 24360 10056
rect 31576 10115 31628 10124
rect 31576 10081 31585 10115
rect 31585 10081 31619 10115
rect 31619 10081 31628 10115
rect 31576 10072 31628 10081
rect 18512 9936 18564 9988
rect 19432 9936 19484 9988
rect 25228 9979 25280 9988
rect 25228 9945 25237 9979
rect 25237 9945 25271 9979
rect 25271 9945 25280 9979
rect 25228 9936 25280 9945
rect 18236 9911 18288 9920
rect 18236 9877 18245 9911
rect 18245 9877 18279 9911
rect 18279 9877 18288 9911
rect 18236 9868 18288 9877
rect 21824 9868 21876 9920
rect 23480 9868 23532 9920
rect 24032 9868 24084 9920
rect 25688 10004 25740 10056
rect 27620 10004 27672 10056
rect 25596 9936 25648 9988
rect 26976 9936 27028 9988
rect 28632 9979 28684 9988
rect 28632 9945 28641 9979
rect 28641 9945 28675 9979
rect 28675 9945 28684 9979
rect 28632 9936 28684 9945
rect 25872 9868 25924 9920
rect 26700 9911 26752 9920
rect 26700 9877 26709 9911
rect 26709 9877 26743 9911
rect 26743 9877 26752 9911
rect 26700 9868 26752 9877
rect 30196 10004 30248 10056
rect 29828 9979 29880 9988
rect 29828 9945 29862 9979
rect 29862 9945 29880 9979
rect 29828 9936 29880 9945
rect 31024 9936 31076 9988
rect 30932 9911 30984 9920
rect 30932 9877 30941 9911
rect 30941 9877 30975 9911
rect 30975 9877 30984 9911
rect 30932 9868 30984 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 18972 9664 19024 9716
rect 3148 9596 3200 9648
rect 18144 9596 18196 9648
rect 19616 9634 19668 9686
rect 21180 9664 21232 9716
rect 22468 9664 22520 9716
rect 23296 9664 23348 9716
rect 1768 9571 1820 9580
rect 1768 9537 1777 9571
rect 1777 9537 1811 9571
rect 1811 9537 1820 9571
rect 1768 9528 1820 9537
rect 17868 9528 17920 9580
rect 18052 9571 18104 9580
rect 18052 9537 18061 9571
rect 18061 9537 18095 9571
rect 18095 9537 18104 9571
rect 18052 9528 18104 9537
rect 18236 9571 18288 9580
rect 18236 9537 18245 9571
rect 18245 9537 18279 9571
rect 18279 9537 18288 9571
rect 18236 9528 18288 9537
rect 19340 9528 19392 9580
rect 20996 9596 21048 9648
rect 22008 9596 22060 9648
rect 24032 9596 24084 9648
rect 2228 9460 2280 9512
rect 2780 9503 2832 9512
rect 2780 9469 2789 9503
rect 2789 9469 2823 9503
rect 2823 9469 2832 9503
rect 2780 9460 2832 9469
rect 19984 9528 20036 9580
rect 20260 9528 20312 9580
rect 22652 9571 22704 9580
rect 22652 9537 22661 9571
rect 22661 9537 22695 9571
rect 22695 9537 22704 9571
rect 22652 9528 22704 9537
rect 22928 9460 22980 9512
rect 23848 9528 23900 9580
rect 25228 9664 25280 9716
rect 25780 9664 25832 9716
rect 25964 9664 26016 9716
rect 26332 9664 26384 9716
rect 31024 9664 31076 9716
rect 31300 9664 31352 9716
rect 31484 9664 31536 9716
rect 26700 9596 26752 9648
rect 27620 9596 27672 9648
rect 25872 9528 25924 9580
rect 26056 9571 26108 9580
rect 26056 9537 26065 9571
rect 26065 9537 26099 9571
rect 26099 9537 26108 9571
rect 26056 9528 26108 9537
rect 26240 9460 26292 9512
rect 27344 9528 27396 9580
rect 27252 9460 27304 9512
rect 30932 9528 30984 9580
rect 32956 9596 33008 9648
rect 32128 9571 32180 9580
rect 19984 9392 20036 9444
rect 20628 9392 20680 9444
rect 26884 9392 26936 9444
rect 32128 9537 32137 9571
rect 32137 9537 32171 9571
rect 32171 9537 32180 9571
rect 32128 9528 32180 9537
rect 17040 9324 17092 9376
rect 19524 9324 19576 9376
rect 21548 9324 21600 9376
rect 23756 9367 23808 9376
rect 23756 9333 23765 9367
rect 23765 9333 23799 9367
rect 23799 9333 23808 9367
rect 23756 9324 23808 9333
rect 24492 9367 24544 9376
rect 24492 9333 24501 9367
rect 24501 9333 24535 9367
rect 24535 9333 24544 9367
rect 24492 9324 24544 9333
rect 24584 9324 24636 9376
rect 26240 9324 26292 9376
rect 26976 9324 27028 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 2228 9163 2280 9172
rect 2228 9129 2237 9163
rect 2237 9129 2271 9163
rect 2271 9129 2280 9163
rect 2228 9120 2280 9129
rect 17408 9120 17460 9172
rect 18236 9052 18288 9104
rect 17040 9027 17092 9036
rect 17040 8993 17049 9027
rect 17049 8993 17083 9027
rect 17083 8993 17092 9027
rect 17040 8984 17092 8993
rect 17316 9027 17368 9036
rect 17316 8993 17325 9027
rect 17325 8993 17359 9027
rect 17359 8993 17368 9027
rect 17316 8984 17368 8993
rect 17592 8984 17644 9036
rect 19524 8959 19576 8968
rect 19524 8925 19558 8959
rect 19558 8925 19576 8959
rect 19524 8916 19576 8925
rect 22468 9120 22520 9172
rect 24492 9120 24544 9172
rect 25136 9120 25188 9172
rect 25872 9120 25924 9172
rect 22100 9052 22152 9104
rect 22652 9052 22704 9104
rect 22744 9095 22796 9104
rect 22744 9061 22753 9095
rect 22753 9061 22787 9095
rect 22787 9061 22796 9095
rect 22744 9052 22796 9061
rect 25044 9052 25096 9104
rect 25228 9052 25280 9104
rect 26884 9120 26936 9172
rect 21548 9027 21600 9036
rect 21548 8993 21557 9027
rect 21557 8993 21591 9027
rect 21591 8993 21600 9027
rect 21548 8984 21600 8993
rect 21916 8984 21968 9036
rect 23204 8984 23256 9036
rect 22192 8959 22244 8968
rect 21824 8848 21876 8900
rect 19340 8780 19392 8832
rect 22192 8925 22201 8959
rect 22201 8925 22235 8959
rect 22235 8925 22244 8959
rect 22192 8916 22244 8925
rect 22376 8959 22428 8968
rect 22376 8925 22385 8959
rect 22385 8925 22419 8959
rect 22419 8925 22428 8959
rect 22376 8916 22428 8925
rect 22468 8916 22520 8968
rect 23572 8959 23624 8968
rect 23572 8925 23581 8959
rect 23581 8925 23615 8959
rect 23615 8925 23624 8959
rect 23572 8916 23624 8925
rect 24032 8984 24084 9036
rect 24308 8984 24360 9036
rect 23848 8959 23900 8968
rect 23848 8925 23857 8959
rect 23857 8925 23891 8959
rect 23891 8925 23900 8959
rect 24400 8959 24452 8968
rect 23848 8916 23900 8925
rect 24400 8925 24409 8959
rect 24409 8925 24443 8959
rect 24443 8925 24452 8959
rect 24400 8916 24452 8925
rect 25780 8959 25832 8968
rect 22652 8848 22704 8900
rect 24860 8848 24912 8900
rect 25780 8925 25789 8959
rect 25789 8925 25823 8959
rect 25823 8925 25832 8959
rect 25780 8916 25832 8925
rect 25872 8959 25924 8968
rect 25872 8925 25881 8959
rect 25881 8925 25915 8959
rect 25915 8925 25924 8959
rect 27068 9052 27120 9104
rect 29460 9052 29512 9104
rect 27436 9027 27488 9036
rect 27436 8993 27445 9027
rect 27445 8993 27479 9027
rect 27479 8993 27488 9027
rect 27436 8984 27488 8993
rect 31300 9052 31352 9104
rect 41696 9052 41748 9104
rect 46848 9052 46900 9104
rect 25872 8916 25924 8925
rect 25688 8848 25740 8900
rect 26332 8848 26384 8900
rect 26700 8848 26752 8900
rect 22376 8780 22428 8832
rect 24308 8780 24360 8832
rect 24400 8780 24452 8832
rect 24584 8780 24636 8832
rect 25044 8780 25096 8832
rect 25228 8780 25280 8832
rect 26056 8780 26108 8832
rect 30656 8916 30708 8968
rect 32496 8984 32548 9036
rect 31484 8916 31536 8968
rect 27896 8848 27948 8900
rect 47768 8891 47820 8900
rect 47768 8857 47777 8891
rect 47777 8857 47811 8891
rect 47811 8857 47820 8891
rect 47768 8848 47820 8857
rect 27252 8780 27304 8832
rect 30656 8823 30708 8832
rect 30656 8789 30665 8823
rect 30665 8789 30699 8823
rect 30699 8789 30708 8823
rect 30656 8780 30708 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 22744 8508 22796 8560
rect 23572 8576 23624 8628
rect 24216 8508 24268 8560
rect 24400 8619 24452 8628
rect 24400 8585 24409 8619
rect 24409 8585 24443 8619
rect 24443 8585 24452 8619
rect 24400 8576 24452 8585
rect 24768 8576 24820 8628
rect 27620 8576 27672 8628
rect 27896 8619 27948 8628
rect 1860 8483 1912 8492
rect 1860 8449 1869 8483
rect 1869 8449 1903 8483
rect 1903 8449 1912 8483
rect 1860 8440 1912 8449
rect 17592 8483 17644 8492
rect 17592 8449 17601 8483
rect 17601 8449 17635 8483
rect 17635 8449 17644 8483
rect 17592 8440 17644 8449
rect 19248 8440 19300 8492
rect 19340 8372 19392 8424
rect 21272 8415 21324 8424
rect 18972 8279 19024 8288
rect 18972 8245 18981 8279
rect 18981 8245 19015 8279
rect 19015 8245 19024 8279
rect 18972 8236 19024 8245
rect 19340 8236 19392 8288
rect 21272 8381 21281 8415
rect 21281 8381 21315 8415
rect 21315 8381 21324 8415
rect 21272 8372 21324 8381
rect 21824 8415 21876 8424
rect 21824 8381 21833 8415
rect 21833 8381 21867 8415
rect 21867 8381 21876 8415
rect 21824 8372 21876 8381
rect 24860 8508 24912 8560
rect 25136 8440 25188 8492
rect 27160 8483 27212 8492
rect 27160 8449 27169 8483
rect 27169 8449 27203 8483
rect 27203 8449 27212 8483
rect 27160 8440 27212 8449
rect 27620 8440 27672 8492
rect 27896 8585 27905 8619
rect 27905 8585 27939 8619
rect 27939 8585 27948 8619
rect 27896 8576 27948 8585
rect 29460 8576 29512 8628
rect 31576 8619 31628 8628
rect 31576 8585 31585 8619
rect 31585 8585 31619 8619
rect 31619 8585 31628 8619
rect 31576 8576 31628 8585
rect 32496 8619 32548 8628
rect 32496 8585 32505 8619
rect 32505 8585 32539 8619
rect 32539 8585 32548 8619
rect 32496 8576 32548 8585
rect 29736 8483 29788 8492
rect 24584 8415 24636 8424
rect 24584 8381 24593 8415
rect 24593 8381 24627 8415
rect 24627 8381 24636 8415
rect 25320 8415 25372 8424
rect 24584 8372 24636 8381
rect 25320 8381 25329 8415
rect 25329 8381 25363 8415
rect 25363 8381 25372 8415
rect 25320 8372 25372 8381
rect 27252 8372 27304 8424
rect 27528 8415 27580 8424
rect 27528 8381 27537 8415
rect 27537 8381 27571 8415
rect 27571 8381 27580 8415
rect 27528 8372 27580 8381
rect 24952 8304 25004 8356
rect 23204 8279 23256 8288
rect 23204 8245 23213 8279
rect 23213 8245 23247 8279
rect 23247 8245 23256 8279
rect 26056 8304 26108 8356
rect 29736 8449 29745 8483
rect 29745 8449 29779 8483
rect 29779 8449 29788 8483
rect 29736 8440 29788 8449
rect 30196 8483 30248 8492
rect 30196 8449 30205 8483
rect 30205 8449 30239 8483
rect 30239 8449 30248 8483
rect 30196 8440 30248 8449
rect 30656 8508 30708 8560
rect 31484 8440 31536 8492
rect 32128 8483 32180 8492
rect 32128 8449 32137 8483
rect 32137 8449 32171 8483
rect 32171 8449 32180 8483
rect 32128 8440 32180 8449
rect 47860 8483 47912 8492
rect 31576 8372 31628 8424
rect 47860 8449 47869 8483
rect 47869 8449 47903 8483
rect 47903 8449 47912 8483
rect 47860 8440 47912 8449
rect 29552 8304 29604 8356
rect 33048 8304 33100 8356
rect 23204 8236 23256 8245
rect 25412 8236 25464 8288
rect 25964 8236 26016 8288
rect 26240 8236 26292 8288
rect 29092 8279 29144 8288
rect 29092 8245 29101 8279
rect 29101 8245 29135 8279
rect 29135 8245 29144 8279
rect 29092 8236 29144 8245
rect 29184 8236 29236 8288
rect 38016 8236 38068 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 18788 7964 18840 8016
rect 21272 8032 21324 8084
rect 29184 8032 29236 8084
rect 29552 8032 29604 8084
rect 30104 8032 30156 8084
rect 32128 8032 32180 8084
rect 18052 7828 18104 7880
rect 18972 7896 19024 7948
rect 21456 7964 21508 8016
rect 22100 8007 22152 8016
rect 22100 7973 22109 8007
rect 22109 7973 22143 8007
rect 22143 7973 22152 8007
rect 22100 7964 22152 7973
rect 26240 7964 26292 8016
rect 45652 8032 45704 8084
rect 23664 7896 23716 7948
rect 24584 7896 24636 7948
rect 23204 7828 23256 7880
rect 23480 7828 23532 7880
rect 24400 7828 24452 7880
rect 27436 7828 27488 7880
rect 1860 7803 1912 7812
rect 1860 7769 1869 7803
rect 1869 7769 1903 7803
rect 1903 7769 1912 7803
rect 1860 7760 1912 7769
rect 18604 7760 18656 7812
rect 25504 7803 25556 7812
rect 18696 7735 18748 7744
rect 18696 7701 18705 7735
rect 18705 7701 18739 7735
rect 18739 7701 18748 7735
rect 18696 7692 18748 7701
rect 20536 7692 20588 7744
rect 22468 7735 22520 7744
rect 22468 7701 22477 7735
rect 22477 7701 22511 7735
rect 22511 7701 22520 7735
rect 22468 7692 22520 7701
rect 25504 7769 25538 7803
rect 25538 7769 25556 7803
rect 25504 7760 25556 7769
rect 31576 7896 31628 7948
rect 30104 7828 30156 7880
rect 30288 7760 30340 7812
rect 30932 7760 30984 7812
rect 29644 7692 29696 7744
rect 46296 7871 46348 7880
rect 46296 7837 46305 7871
rect 46305 7837 46339 7871
rect 46339 7837 46348 7871
rect 46296 7828 46348 7837
rect 46756 7760 46808 7812
rect 48136 7803 48188 7812
rect 48136 7769 48145 7803
rect 48145 7769 48179 7803
rect 48179 7769 48188 7803
rect 48136 7760 48188 7769
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 18604 7488 18656 7540
rect 19248 7488 19300 7540
rect 18696 7420 18748 7472
rect 17960 7352 18012 7404
rect 18420 7395 18472 7404
rect 18420 7361 18429 7395
rect 18429 7361 18463 7395
rect 18463 7361 18472 7395
rect 18420 7352 18472 7361
rect 19616 7395 19668 7404
rect 19616 7361 19625 7395
rect 19625 7361 19659 7395
rect 19659 7361 19668 7395
rect 19616 7352 19668 7361
rect 19984 7488 20036 7540
rect 24860 7531 24912 7540
rect 24860 7497 24869 7531
rect 24869 7497 24903 7531
rect 24903 7497 24912 7531
rect 24860 7488 24912 7497
rect 27804 7488 27856 7540
rect 28080 7488 28132 7540
rect 29736 7488 29788 7540
rect 30932 7531 30984 7540
rect 30932 7497 30941 7531
rect 30941 7497 30975 7531
rect 30975 7497 30984 7531
rect 30932 7488 30984 7497
rect 46756 7531 46808 7540
rect 46756 7497 46765 7531
rect 46765 7497 46799 7531
rect 46799 7497 46808 7531
rect 46756 7488 46808 7497
rect 29092 7420 29144 7472
rect 46296 7420 46348 7472
rect 23480 7395 23532 7404
rect 23480 7361 23489 7395
rect 23489 7361 23523 7395
rect 23523 7361 23532 7395
rect 23480 7352 23532 7361
rect 25228 7352 25280 7404
rect 32588 7352 32640 7404
rect 45560 7352 45612 7404
rect 27436 7284 27488 7336
rect 19064 7216 19116 7268
rect 20352 7216 20404 7268
rect 2044 7148 2096 7200
rect 29736 7148 29788 7200
rect 30288 7148 30340 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 19340 6944 19392 6996
rect 3424 6808 3476 6860
rect 30288 6876 30340 6928
rect 17224 6740 17276 6792
rect 17500 6740 17552 6792
rect 18420 6740 18472 6792
rect 19616 6740 19668 6792
rect 22468 6740 22520 6792
rect 20904 6715 20956 6724
rect 20904 6681 20913 6715
rect 20913 6681 20947 6715
rect 20947 6681 20956 6715
rect 20904 6672 20956 6681
rect 29736 6851 29788 6860
rect 29736 6817 29745 6851
rect 29745 6817 29779 6851
rect 29779 6817 29788 6851
rect 29736 6808 29788 6817
rect 44916 6808 44968 6860
rect 46848 6851 46900 6860
rect 46848 6817 46857 6851
rect 46857 6817 46891 6851
rect 46891 6817 46900 6851
rect 46848 6808 46900 6817
rect 45928 6672 45980 6724
rect 2228 6604 2280 6656
rect 19432 6604 19484 6656
rect 20168 6604 20220 6656
rect 21088 6604 21140 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 2228 6375 2280 6384
rect 2228 6341 2237 6375
rect 2237 6341 2271 6375
rect 2271 6341 2280 6375
rect 2228 6332 2280 6341
rect 20904 6400 20956 6452
rect 45928 6443 45980 6452
rect 45928 6409 45937 6443
rect 45937 6409 45971 6443
rect 45971 6409 45980 6443
rect 45928 6400 45980 6409
rect 20996 6375 21048 6384
rect 20996 6341 21005 6375
rect 21005 6341 21039 6375
rect 21039 6341 21048 6375
rect 20996 6332 21048 6341
rect 22008 6332 22060 6384
rect 24124 6332 24176 6384
rect 28632 6332 28684 6384
rect 2044 6307 2096 6316
rect 2044 6273 2053 6307
rect 2053 6273 2087 6307
rect 2087 6273 2096 6307
rect 2044 6264 2096 6273
rect 23572 6264 23624 6316
rect 2780 6239 2832 6248
rect 2780 6205 2789 6239
rect 2789 6205 2823 6239
rect 2823 6205 2832 6239
rect 2780 6196 2832 6205
rect 23848 6307 23900 6316
rect 23848 6273 23857 6307
rect 23857 6273 23891 6307
rect 23891 6273 23900 6307
rect 23848 6264 23900 6273
rect 24032 6307 24084 6316
rect 24032 6273 24041 6307
rect 24041 6273 24075 6307
rect 24075 6273 24084 6307
rect 24032 6264 24084 6273
rect 24492 6264 24544 6316
rect 27804 6307 27856 6316
rect 27804 6273 27813 6307
rect 27813 6273 27847 6307
rect 27847 6273 27856 6307
rect 27804 6264 27856 6273
rect 29920 6264 29972 6316
rect 35624 6264 35676 6316
rect 45836 6307 45888 6316
rect 45836 6273 45845 6307
rect 45845 6273 45879 6307
rect 45879 6273 45888 6307
rect 45836 6264 45888 6273
rect 24216 6196 24268 6248
rect 2412 6128 2464 6180
rect 2688 6128 2740 6180
rect 39488 6128 39540 6180
rect 1584 6103 1636 6112
rect 1584 6069 1593 6103
rect 1593 6069 1627 6103
rect 1627 6069 1636 6103
rect 1584 6060 1636 6069
rect 22928 6060 22980 6112
rect 23388 6103 23440 6112
rect 23388 6069 23397 6103
rect 23397 6069 23431 6103
rect 23431 6069 23440 6103
rect 23388 6060 23440 6069
rect 28172 6060 28224 6112
rect 46296 6060 46348 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 1768 5695 1820 5704
rect 1768 5661 1777 5695
rect 1777 5661 1811 5695
rect 1811 5661 1820 5695
rect 1768 5652 1820 5661
rect 2320 5720 2372 5772
rect 22008 5831 22060 5840
rect 22008 5797 22017 5831
rect 22017 5797 22051 5831
rect 22051 5797 22060 5831
rect 22008 5788 22060 5797
rect 21640 5720 21692 5772
rect 24216 5788 24268 5840
rect 25780 5831 25832 5840
rect 25780 5797 25789 5831
rect 25789 5797 25823 5831
rect 25823 5797 25832 5831
rect 25780 5788 25832 5797
rect 2688 5652 2740 5704
rect 21824 5652 21876 5704
rect 22284 5652 22336 5704
rect 24032 5720 24084 5772
rect 24400 5763 24452 5772
rect 24400 5729 24409 5763
rect 24409 5729 24443 5763
rect 24443 5729 24452 5763
rect 24400 5720 24452 5729
rect 22928 5695 22980 5704
rect 22928 5661 22937 5695
rect 22937 5661 22971 5695
rect 22971 5661 22980 5695
rect 22928 5652 22980 5661
rect 23112 5695 23164 5704
rect 23112 5661 23121 5695
rect 23121 5661 23155 5695
rect 23155 5661 23164 5695
rect 23112 5652 23164 5661
rect 23388 5652 23440 5704
rect 27804 5856 27856 5908
rect 27160 5763 27212 5772
rect 27160 5729 27169 5763
rect 27169 5729 27203 5763
rect 27203 5729 27212 5763
rect 27160 5720 27212 5729
rect 45468 5856 45520 5908
rect 46296 5763 46348 5772
rect 46296 5729 46305 5763
rect 46305 5729 46339 5763
rect 46339 5729 46348 5763
rect 46296 5720 46348 5729
rect 24400 5584 24452 5636
rect 27160 5584 27212 5636
rect 27712 5584 27764 5636
rect 46940 5584 46992 5636
rect 48136 5627 48188 5636
rect 48136 5593 48145 5627
rect 48145 5593 48179 5627
rect 48179 5593 48188 5627
rect 48136 5584 48188 5593
rect 1952 5516 2004 5568
rect 2964 5559 3016 5568
rect 2964 5525 2973 5559
rect 2973 5525 3007 5559
rect 3007 5525 3016 5559
rect 2964 5516 3016 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 3424 5312 3476 5364
rect 18144 5312 18196 5364
rect 22468 5312 22520 5364
rect 23848 5312 23900 5364
rect 27712 5355 27764 5364
rect 27712 5321 27721 5355
rect 27721 5321 27755 5355
rect 27755 5321 27764 5355
rect 27712 5312 27764 5321
rect 39304 5312 39356 5364
rect 46664 5312 46716 5364
rect 46940 5355 46992 5364
rect 46940 5321 46949 5355
rect 46949 5321 46983 5355
rect 46983 5321 46992 5355
rect 46940 5312 46992 5321
rect 1952 5287 2004 5296
rect 1952 5253 1961 5287
rect 1961 5253 1995 5287
rect 1995 5253 2004 5287
rect 1952 5244 2004 5253
rect 14740 5244 14792 5296
rect 19248 5244 19300 5296
rect 24124 5244 24176 5296
rect 24216 5244 24268 5296
rect 1584 5176 1636 5228
rect 19340 5176 19392 5228
rect 2780 5151 2832 5160
rect 2780 5117 2789 5151
rect 2789 5117 2823 5151
rect 2823 5117 2832 5151
rect 2780 5108 2832 5117
rect 21088 5222 21140 5228
rect 21088 5188 21118 5222
rect 21118 5188 21140 5222
rect 21088 5176 21140 5188
rect 21824 5219 21876 5228
rect 21824 5185 21833 5219
rect 21833 5185 21867 5219
rect 21867 5185 21876 5219
rect 21824 5176 21876 5185
rect 23112 5176 23164 5228
rect 25780 5176 25832 5228
rect 29000 5244 29052 5296
rect 28172 5219 28224 5228
rect 28172 5185 28181 5219
rect 28181 5185 28215 5219
rect 28215 5185 28224 5219
rect 28172 5176 28224 5185
rect 28724 5176 28776 5228
rect 46848 5219 46900 5228
rect 46848 5185 46857 5219
rect 46857 5185 46891 5219
rect 46891 5185 46900 5219
rect 46848 5176 46900 5185
rect 47860 5219 47912 5228
rect 47860 5185 47869 5219
rect 47869 5185 47903 5219
rect 47903 5185 47912 5219
rect 47860 5176 47912 5185
rect 38752 5108 38804 5160
rect 21640 5040 21692 5092
rect 24032 5040 24084 5092
rect 28724 5040 28776 5092
rect 29828 5040 29880 5092
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 17224 4700 17276 4752
rect 46848 4700 46900 4752
rect 1768 4632 1820 4684
rect 2780 4675 2832 4684
rect 2780 4641 2789 4675
rect 2789 4641 2823 4675
rect 2823 4641 2832 4675
rect 2780 4632 2832 4641
rect 30932 4675 30984 4684
rect 30932 4641 30941 4675
rect 30941 4641 30975 4675
rect 30975 4641 30984 4675
rect 30932 4632 30984 4641
rect 6184 4564 6236 4616
rect 13176 4564 13228 4616
rect 41972 4607 42024 4616
rect 2964 4496 3016 4548
rect 41972 4573 41981 4607
rect 41981 4573 42015 4607
rect 42015 4573 42024 4607
rect 41972 4564 42024 4573
rect 30656 4496 30708 4548
rect 46940 4496 46992 4548
rect 48320 4496 48372 4548
rect 30380 4428 30432 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 1584 4131 1636 4140
rect 1584 4097 1593 4131
rect 1593 4097 1627 4131
rect 1627 4097 1636 4131
rect 1584 4088 1636 4097
rect 3056 4131 3108 4140
rect 3056 4097 3065 4131
rect 3065 4097 3099 4131
rect 3099 4097 3108 4131
rect 3056 4088 3108 4097
rect 12256 4088 12308 4140
rect 13176 4131 13228 4140
rect 13176 4097 13185 4131
rect 13185 4097 13219 4131
rect 13219 4097 13228 4131
rect 13176 4088 13228 4097
rect 16764 4088 16816 4140
rect 26240 4088 26292 4140
rect 26608 4088 26660 4140
rect 11612 3952 11664 4004
rect 11980 3952 12032 4004
rect 13084 4020 13136 4072
rect 13544 4020 13596 4072
rect 16212 4020 16264 4072
rect 20812 4020 20864 4072
rect 21180 4020 21232 4072
rect 15292 3952 15344 4004
rect 20352 3952 20404 4004
rect 1952 3884 2004 3936
rect 2320 3927 2372 3936
rect 2320 3893 2329 3927
rect 2329 3893 2363 3927
rect 2363 3893 2372 3927
rect 2320 3884 2372 3893
rect 3148 3927 3200 3936
rect 3148 3893 3157 3927
rect 3157 3893 3191 3927
rect 3191 3893 3200 3927
rect 3148 3884 3200 3893
rect 3884 3927 3936 3936
rect 3884 3893 3893 3927
rect 3893 3893 3927 3927
rect 3927 3893 3936 3927
rect 3884 3884 3936 3893
rect 6552 3884 6604 3936
rect 7104 3927 7156 3936
rect 7104 3893 7113 3927
rect 7113 3893 7147 3927
rect 7147 3893 7156 3927
rect 7104 3884 7156 3893
rect 11704 3884 11756 3936
rect 12624 3884 12676 3936
rect 17132 3884 17184 3936
rect 17408 3884 17460 3936
rect 20168 3884 20220 3936
rect 21272 3952 21324 4004
rect 22376 4020 22428 4072
rect 29552 4088 29604 4140
rect 29736 4088 29788 4140
rect 22008 3952 22060 4004
rect 46756 4156 46808 4208
rect 36452 4088 36504 4140
rect 39488 4131 39540 4140
rect 39488 4097 39497 4131
rect 39497 4097 39531 4131
rect 39531 4097 39540 4131
rect 39488 4088 39540 4097
rect 42432 4131 42484 4140
rect 42432 4097 42441 4131
rect 42441 4097 42475 4131
rect 42475 4097 42484 4131
rect 42432 4088 42484 4097
rect 45560 4088 45612 4140
rect 45836 4131 45888 4140
rect 45836 4097 45845 4131
rect 45845 4097 45879 4131
rect 45879 4097 45888 4131
rect 45836 4088 45888 4097
rect 46848 4131 46900 4140
rect 46848 4097 46857 4131
rect 46857 4097 46891 4131
rect 46891 4097 46900 4131
rect 46848 4088 46900 4097
rect 46940 4131 46992 4140
rect 46940 4097 46949 4131
rect 46949 4097 46983 4131
rect 46983 4097 46992 4131
rect 46940 4088 46992 4097
rect 40776 3952 40828 4004
rect 44640 3952 44692 4004
rect 29552 3884 29604 3936
rect 30564 3884 30616 3936
rect 30656 3927 30708 3936
rect 30656 3893 30665 3927
rect 30665 3893 30699 3927
rect 30699 3893 30708 3927
rect 31392 3927 31444 3936
rect 30656 3884 30708 3893
rect 31392 3893 31401 3927
rect 31401 3893 31435 3927
rect 31435 3893 31444 3927
rect 31392 3884 31444 3893
rect 32772 3884 32824 3936
rect 36176 3884 36228 3936
rect 37924 3884 37976 3936
rect 40224 3884 40276 3936
rect 41420 3884 41472 3936
rect 42616 3884 42668 3936
rect 43996 3884 44048 3936
rect 44824 4020 44876 4072
rect 46296 3952 46348 4004
rect 45376 3927 45428 3936
rect 45376 3893 45385 3927
rect 45385 3893 45419 3927
rect 45419 3893 45428 3927
rect 45376 3884 45428 3893
rect 46204 3884 46256 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 3884 3680 3936 3732
rect 9036 3680 9088 3732
rect 2320 3612 2372 3664
rect 3240 3612 3292 3664
rect 1860 3587 1912 3596
rect 1860 3553 1869 3587
rect 1869 3553 1903 3587
rect 1903 3553 1912 3587
rect 1860 3544 1912 3553
rect 3148 3544 3200 3596
rect 5816 3612 5868 3664
rect 6184 3587 6236 3596
rect 6184 3553 6193 3587
rect 6193 3553 6227 3587
rect 6227 3553 6236 3587
rect 6184 3544 6236 3553
rect 7104 3544 7156 3596
rect 10324 3612 10376 3664
rect 12900 3612 12952 3664
rect 13084 3655 13136 3664
rect 13084 3621 13093 3655
rect 13093 3621 13127 3655
rect 13127 3621 13136 3655
rect 13084 3612 13136 3621
rect 13176 3612 13228 3664
rect 3792 3519 3844 3528
rect 3792 3485 3801 3519
rect 3801 3485 3835 3519
rect 3835 3485 3844 3519
rect 3792 3476 3844 3485
rect 11612 3519 11664 3528
rect 11612 3485 11621 3519
rect 11621 3485 11655 3519
rect 11655 3485 11664 3519
rect 12624 3544 12676 3596
rect 12256 3519 12308 3528
rect 11612 3476 11664 3485
rect 12256 3485 12265 3519
rect 12265 3485 12299 3519
rect 12299 3485 12308 3519
rect 16120 3544 16172 3596
rect 18512 3612 18564 3664
rect 30288 3612 30340 3664
rect 20168 3587 20220 3596
rect 12256 3476 12308 3485
rect 12992 3519 13044 3528
rect 12992 3485 13001 3519
rect 13001 3485 13035 3519
rect 13035 3485 13044 3519
rect 12992 3476 13044 3485
rect 14280 3476 14332 3528
rect 15200 3476 15252 3528
rect 15660 3476 15712 3528
rect 17684 3476 17736 3528
rect 17776 3476 17828 3528
rect 2596 3408 2648 3460
rect 20168 3553 20177 3587
rect 20177 3553 20211 3587
rect 20211 3553 20220 3587
rect 20168 3544 20220 3553
rect 20352 3587 20404 3596
rect 20352 3553 20361 3587
rect 20361 3553 20395 3587
rect 20395 3553 20404 3587
rect 20352 3544 20404 3553
rect 20628 3587 20680 3596
rect 20628 3553 20637 3587
rect 20637 3553 20671 3587
rect 20671 3553 20680 3587
rect 20628 3544 20680 3553
rect 20812 3544 20864 3596
rect 21916 3544 21968 3596
rect 22744 3519 22796 3528
rect 22744 3485 22753 3519
rect 22753 3485 22787 3519
rect 22787 3485 22796 3519
rect 22744 3476 22796 3485
rect 1584 3340 1636 3392
rect 11612 3340 11664 3392
rect 11888 3340 11940 3392
rect 12164 3340 12216 3392
rect 14464 3340 14516 3392
rect 17960 3340 18012 3392
rect 18236 3340 18288 3392
rect 26240 3544 26292 3596
rect 26424 3587 26476 3596
rect 26424 3553 26433 3587
rect 26433 3553 26467 3587
rect 26467 3553 26476 3587
rect 26424 3544 26476 3553
rect 25872 3519 25924 3528
rect 25872 3485 25881 3519
rect 25881 3485 25915 3519
rect 25915 3485 25924 3519
rect 25872 3476 25924 3485
rect 29000 3519 29052 3528
rect 29000 3485 29009 3519
rect 29009 3485 29043 3519
rect 29043 3485 29052 3519
rect 29000 3476 29052 3485
rect 29460 3408 29512 3460
rect 23664 3340 23716 3392
rect 23756 3340 23808 3392
rect 29736 3476 29788 3528
rect 31392 3612 31444 3664
rect 31576 3587 31628 3596
rect 31576 3553 31585 3587
rect 31585 3553 31619 3587
rect 31619 3553 31628 3587
rect 31576 3544 31628 3553
rect 32220 3680 32272 3732
rect 33968 3680 34020 3732
rect 37372 3680 37424 3732
rect 39580 3680 39632 3732
rect 32312 3612 32364 3664
rect 42432 3612 42484 3664
rect 36176 3587 36228 3596
rect 30564 3451 30616 3460
rect 30564 3417 30573 3451
rect 30573 3417 30607 3451
rect 30607 3417 30616 3451
rect 30564 3408 30616 3417
rect 36176 3553 36185 3587
rect 36185 3553 36219 3587
rect 36219 3553 36228 3587
rect 36176 3544 36228 3553
rect 36728 3587 36780 3596
rect 36728 3553 36737 3587
rect 36737 3553 36771 3587
rect 36771 3553 36780 3587
rect 36728 3544 36780 3553
rect 41420 3587 41472 3596
rect 41420 3553 41429 3587
rect 41429 3553 41463 3587
rect 41463 3553 41472 3587
rect 41420 3544 41472 3553
rect 41880 3587 41932 3596
rect 41880 3553 41889 3587
rect 41889 3553 41923 3587
rect 41923 3553 41932 3587
rect 41880 3544 41932 3553
rect 35992 3519 36044 3528
rect 35992 3485 36001 3519
rect 36001 3485 36035 3519
rect 36035 3485 36044 3519
rect 35992 3476 36044 3485
rect 37740 3476 37792 3528
rect 40776 3519 40828 3528
rect 40776 3485 40785 3519
rect 40785 3485 40819 3519
rect 40819 3485 40828 3519
rect 40776 3476 40828 3485
rect 43812 3476 43864 3528
rect 47492 3612 47544 3664
rect 45376 3544 45428 3596
rect 46204 3587 46256 3596
rect 46204 3553 46213 3587
rect 46213 3553 46247 3587
rect 46247 3553 46256 3587
rect 46204 3544 46256 3553
rect 46480 3587 46532 3596
rect 46480 3553 46489 3587
rect 46489 3553 46523 3587
rect 46523 3553 46532 3587
rect 46480 3544 46532 3553
rect 29920 3340 29972 3392
rect 30012 3340 30064 3392
rect 39948 3408 40000 3460
rect 32956 3340 33008 3392
rect 40040 3340 40092 3392
rect 46388 3408 46440 3460
rect 45192 3340 45244 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 3056 3136 3108 3188
rect 19984 3136 20036 3188
rect 20352 3136 20404 3188
rect 20720 3136 20772 3188
rect 22468 3136 22520 3188
rect 22652 3136 22704 3188
rect 30012 3136 30064 3188
rect 1952 3111 2004 3120
rect 1952 3077 1961 3111
rect 1961 3077 1995 3111
rect 1995 3077 2004 3111
rect 1952 3068 2004 3077
rect 6552 3111 6604 3120
rect 6552 3077 6561 3111
rect 6561 3077 6595 3111
rect 6595 3077 6604 3111
rect 6552 3068 6604 3077
rect 12164 3111 12216 3120
rect 12164 3077 12173 3111
rect 12173 3077 12207 3111
rect 12207 3077 12216 3111
rect 12164 3068 12216 3077
rect 14464 3111 14516 3120
rect 14464 3077 14473 3111
rect 14473 3077 14507 3111
rect 14507 3077 14516 3111
rect 14464 3068 14516 3077
rect 17960 3111 18012 3120
rect 17960 3077 17969 3111
rect 17969 3077 18003 3111
rect 18003 3077 18012 3111
rect 17960 3068 18012 3077
rect 3792 3000 3844 3052
rect 8392 3000 8444 3052
rect 11980 3043 12032 3052
rect 11980 3009 11989 3043
rect 11989 3009 12023 3043
rect 12023 3009 12032 3043
rect 11980 3000 12032 3009
rect 14280 3043 14332 3052
rect 14280 3009 14289 3043
rect 14289 3009 14323 3043
rect 14323 3009 14332 3043
rect 14280 3000 14332 3009
rect 17776 3043 17828 3052
rect 17776 3009 17785 3043
rect 17785 3009 17819 3043
rect 17819 3009 17828 3043
rect 17776 3000 17828 3009
rect 20260 3068 20312 3120
rect 23664 3111 23716 3120
rect 21180 3043 21232 3052
rect 21180 3009 21189 3043
rect 21189 3009 21223 3043
rect 21223 3009 21232 3043
rect 21180 3000 21232 3009
rect 2964 2932 3016 2984
rect 12900 2975 12952 2984
rect 1308 2864 1360 2916
rect 5172 2864 5224 2916
rect 12900 2941 12909 2975
rect 12909 2941 12943 2975
rect 12943 2941 12952 2975
rect 12900 2932 12952 2941
rect 15476 2975 15528 2984
rect 15476 2941 15485 2975
rect 15485 2941 15519 2975
rect 15519 2941 15528 2975
rect 15476 2932 15528 2941
rect 18052 2932 18104 2984
rect 8852 2907 8904 2916
rect 8852 2873 8861 2907
rect 8861 2873 8895 2907
rect 8895 2873 8904 2907
rect 8852 2864 8904 2873
rect 10968 2864 11020 2916
rect 17316 2864 17368 2916
rect 17408 2864 17460 2916
rect 21180 2864 21232 2916
rect 11612 2796 11664 2848
rect 15200 2796 15252 2848
rect 17500 2796 17552 2848
rect 22376 2932 22428 2984
rect 23664 3077 23673 3111
rect 23673 3077 23707 3111
rect 23707 3077 23716 3111
rect 23664 3068 23716 3077
rect 29920 3111 29972 3120
rect 29920 3077 29929 3111
rect 29929 3077 29963 3111
rect 29963 3077 29972 3111
rect 29920 3068 29972 3077
rect 22744 3000 22796 3052
rect 25872 3000 25924 3052
rect 29000 3000 29052 3052
rect 23756 2932 23808 2984
rect 23848 2932 23900 2984
rect 30288 2975 30340 2984
rect 30288 2941 30297 2975
rect 30297 2941 30331 2975
rect 30331 2941 30340 2975
rect 30288 2932 30340 2941
rect 34980 3136 35032 3188
rect 32956 3111 33008 3120
rect 32956 3077 32965 3111
rect 32965 3077 32999 3111
rect 32999 3077 33008 3111
rect 32956 3068 33008 3077
rect 35348 3068 35400 3120
rect 37924 3111 37976 3120
rect 37924 3077 37933 3111
rect 37933 3077 37967 3111
rect 37967 3077 37976 3111
rect 37924 3068 37976 3077
rect 40224 3111 40276 3120
rect 40224 3077 40233 3111
rect 40233 3077 40267 3111
rect 40267 3077 40276 3111
rect 40224 3068 40276 3077
rect 43996 3111 44048 3120
rect 43996 3077 44005 3111
rect 44005 3077 44039 3111
rect 44039 3077 44048 3111
rect 43996 3068 44048 3077
rect 45652 3136 45704 3188
rect 47124 3068 47176 3120
rect 32772 3043 32824 3052
rect 32772 3009 32781 3043
rect 32781 3009 32815 3043
rect 32815 3009 32824 3043
rect 32772 3000 32824 3009
rect 35992 3000 36044 3052
rect 37740 3043 37792 3052
rect 37740 3009 37749 3043
rect 37749 3009 37783 3043
rect 37783 3009 37792 3043
rect 37740 3000 37792 3009
rect 40040 3043 40092 3052
rect 40040 3009 40049 3043
rect 40049 3009 40083 3043
rect 40083 3009 40092 3043
rect 40040 3000 40092 3009
rect 43168 3000 43220 3052
rect 43812 3043 43864 3052
rect 43812 3009 43821 3043
rect 43821 3009 43855 3043
rect 43855 3009 43864 3043
rect 43812 3000 43864 3009
rect 45744 3000 45796 3052
rect 49608 3000 49660 3052
rect 33508 2975 33560 2984
rect 21456 2864 21508 2916
rect 33508 2941 33517 2975
rect 33517 2941 33551 2975
rect 33551 2941 33560 2975
rect 33508 2932 33560 2941
rect 35440 2975 35492 2984
rect 35440 2941 35449 2975
rect 35449 2941 35483 2975
rect 35483 2941 35492 2975
rect 35440 2932 35492 2941
rect 39948 2932 40000 2984
rect 41236 2975 41288 2984
rect 41236 2941 41245 2975
rect 41245 2941 41279 2975
rect 41279 2941 41288 2975
rect 41236 2932 41288 2941
rect 44456 2975 44508 2984
rect 44456 2941 44465 2975
rect 44465 2941 44499 2975
rect 44499 2941 44508 2975
rect 44456 2932 44508 2941
rect 22468 2796 22520 2848
rect 34060 2864 34112 2916
rect 34244 2864 34296 2916
rect 34520 2796 34572 2848
rect 35348 2839 35400 2848
rect 35348 2805 35357 2839
rect 35357 2805 35391 2839
rect 35391 2805 35400 2839
rect 35624 2864 35676 2916
rect 35348 2796 35400 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 2964 2592 3016 2644
rect 14740 2567 14792 2576
rect 11704 2499 11756 2508
rect 11704 2465 11713 2499
rect 11713 2465 11747 2499
rect 11747 2465 11756 2499
rect 11704 2456 11756 2465
rect 11888 2499 11940 2508
rect 11888 2465 11897 2499
rect 11897 2465 11931 2499
rect 11931 2465 11940 2499
rect 11888 2456 11940 2465
rect 14740 2533 14749 2567
rect 14749 2533 14783 2567
rect 14783 2533 14792 2567
rect 14740 2524 14792 2533
rect 20444 2592 20496 2644
rect 22560 2592 22612 2644
rect 23572 2592 23624 2644
rect 26332 2592 26384 2644
rect 28080 2592 28132 2644
rect 19340 2524 19392 2576
rect 28908 2524 28960 2576
rect 30472 2592 30524 2644
rect 46388 2592 46440 2644
rect 34520 2524 34572 2576
rect 35440 2524 35492 2576
rect 38752 2567 38804 2576
rect 38752 2533 38761 2567
rect 38761 2533 38795 2567
rect 38795 2533 38804 2567
rect 38752 2524 38804 2533
rect 19432 2456 19484 2508
rect 20536 2456 20588 2508
rect 30380 2456 30432 2508
rect 41972 2456 42024 2508
rect 42616 2499 42668 2508
rect 42616 2465 42625 2499
rect 42625 2465 42659 2499
rect 42659 2465 42668 2499
rect 42616 2456 42668 2465
rect 42708 2456 42760 2508
rect 44640 2456 44692 2508
rect 45192 2499 45244 2508
rect 45192 2465 45201 2499
rect 45201 2465 45235 2499
rect 45235 2465 45244 2499
rect 45192 2456 45244 2465
rect 45376 2456 45428 2508
rect 1400 2431 1452 2440
rect 1400 2397 1409 2431
rect 1409 2397 1443 2431
rect 1443 2397 1452 2431
rect 1400 2388 1452 2397
rect 1952 2388 2004 2440
rect 7104 2388 7156 2440
rect 7472 2431 7524 2440
rect 7472 2397 7481 2431
rect 7481 2397 7515 2431
rect 7515 2397 7524 2431
rect 7472 2388 7524 2397
rect 7748 2388 7800 2440
rect 9680 2388 9732 2440
rect 4528 2320 4580 2372
rect 4988 2295 5040 2304
rect 4988 2261 4997 2295
rect 4997 2261 5031 2295
rect 5031 2261 5040 2295
rect 4988 2252 5040 2261
rect 10416 2295 10468 2304
rect 10416 2261 10425 2295
rect 10425 2261 10459 2295
rect 10459 2261 10468 2295
rect 10416 2252 10468 2261
rect 12256 2320 12308 2372
rect 14188 2320 14240 2372
rect 17408 2388 17460 2440
rect 17776 2431 17828 2440
rect 17776 2397 17785 2431
rect 17785 2397 17819 2431
rect 17819 2397 17828 2431
rect 17776 2388 17828 2397
rect 19984 2388 20036 2440
rect 22560 2320 22612 2372
rect 23204 2388 23256 2440
rect 24400 2388 24452 2440
rect 27068 2388 27120 2440
rect 32864 2388 32916 2440
rect 34152 2431 34204 2440
rect 34152 2397 34161 2431
rect 34161 2397 34195 2431
rect 34195 2397 34204 2431
rect 34152 2388 34204 2397
rect 34796 2388 34848 2440
rect 38660 2388 38712 2440
rect 24492 2363 24544 2372
rect 24492 2329 24501 2363
rect 24501 2329 24535 2363
rect 24535 2329 24544 2363
rect 24492 2320 24544 2329
rect 25136 2320 25188 2372
rect 20076 2252 20128 2304
rect 27712 2320 27764 2372
rect 36084 2320 36136 2372
rect 47768 2363 47820 2372
rect 47768 2329 47777 2363
rect 47777 2329 47811 2363
rect 47811 2329 47820 2363
rect 47768 2320 47820 2329
rect 28172 2252 28224 2304
rect 47860 2295 47912 2304
rect 47860 2261 47869 2295
rect 47869 2261 47903 2295
rect 47903 2261 47912 2295
rect 47860 2252 47912 2261
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 3424 1980 3476 2032
rect 39028 1980 39080 2032
rect 7472 1912 7524 1964
rect 22284 1912 22336 1964
rect 23940 1912 23992 1964
rect 47860 1912 47912 1964
rect 4988 1844 5040 1896
rect 28448 1844 28500 1896
rect 17776 1776 17828 1828
rect 35348 1776 35400 1828
<< metal2 >>
rect 18 51200 74 52000
rect 662 51200 718 52000
rect 1306 51200 1362 52000
rect 1950 51200 2006 52000
rect 2594 51200 2650 52000
rect 3238 51354 3294 52000
rect 3790 51776 3846 51785
rect 3790 51711 3846 51720
rect 3238 51326 3648 51354
rect 3238 51200 3294 51326
rect 32 48822 60 51200
rect 20 48816 72 48822
rect 20 48758 72 48764
rect 676 48754 704 51200
rect 1320 49298 1348 51200
rect 1308 49292 1360 49298
rect 1308 49234 1360 49240
rect 664 48748 716 48754
rect 664 48690 716 48696
rect 1492 48680 1544 48686
rect 1492 48622 1544 48628
rect 1400 48136 1452 48142
rect 1400 48078 1452 48084
rect 1412 47258 1440 48078
rect 1400 47252 1452 47258
rect 1400 47194 1452 47200
rect 1400 46368 1452 46374
rect 1400 46310 1452 46316
rect 1412 46034 1440 46310
rect 1400 46028 1452 46034
rect 1400 45970 1452 45976
rect 1398 45656 1454 45665
rect 1398 45591 1454 45600
rect 1412 45490 1440 45591
rect 1400 45484 1452 45490
rect 1400 45426 1452 45432
rect 1400 44872 1452 44878
rect 1400 44814 1452 44820
rect 1412 44305 1440 44814
rect 1398 44296 1454 44305
rect 1398 44231 1454 44240
rect 1400 43784 1452 43790
rect 1400 43726 1452 43732
rect 1412 43625 1440 43726
rect 1398 43616 1454 43625
rect 1398 43551 1454 43560
rect 1400 42016 1452 42022
rect 1400 41958 1452 41964
rect 1412 41682 1440 41958
rect 1400 41676 1452 41682
rect 1400 41618 1452 41624
rect 1400 41132 1452 41138
rect 1400 41074 1452 41080
rect 1412 40905 1440 41074
rect 1398 40896 1454 40905
rect 1398 40831 1454 40840
rect 1400 39840 1452 39846
rect 1400 39782 1452 39788
rect 1412 39506 1440 39782
rect 1400 39500 1452 39506
rect 1400 39442 1452 39448
rect 1400 38956 1452 38962
rect 1400 38898 1452 38904
rect 1412 37890 1440 38898
rect 1320 37862 1440 37890
rect 1320 37346 1348 37862
rect 1400 37800 1452 37806
rect 1400 37742 1452 37748
rect 1412 37505 1440 37742
rect 1398 37496 1454 37505
rect 1398 37431 1454 37440
rect 1320 37318 1440 37346
rect 1412 31754 1440 37318
rect 1504 35894 1532 48622
rect 1964 48278 1992 51200
rect 3422 51096 3478 51105
rect 3422 51031 3478 51040
rect 3436 49910 3464 51031
rect 3424 49904 3476 49910
rect 3424 49846 3476 49852
rect 3620 49230 3648 51326
rect 3608 49224 3660 49230
rect 3608 49166 3660 49172
rect 2596 49156 2648 49162
rect 2596 49098 2648 49104
rect 1952 48272 2004 48278
rect 1952 48214 2004 48220
rect 1584 48068 1636 48074
rect 1584 48010 1636 48016
rect 1596 47802 1624 48010
rect 1584 47796 1636 47802
rect 1584 47738 1636 47744
rect 2608 47734 2636 49098
rect 2778 49056 2834 49065
rect 2778 48991 2834 49000
rect 2792 48210 2820 48991
rect 3148 48680 3200 48686
rect 3148 48622 3200 48628
rect 3160 48346 3188 48622
rect 3148 48340 3200 48346
rect 3148 48282 3200 48288
rect 2780 48204 2832 48210
rect 2780 48146 2832 48152
rect 3804 48006 3832 51711
rect 3882 51200 3938 52000
rect 4526 51354 4582 52000
rect 5170 51354 5226 52000
rect 4526 51326 4936 51354
rect 4526 51200 4582 51326
rect 4066 50416 4122 50425
rect 4066 50351 4122 50360
rect 4080 49314 4108 50351
rect 4214 49532 4522 49552
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49456 4522 49476
rect 4080 49286 4200 49314
rect 3976 49088 4028 49094
rect 3976 49030 4028 49036
rect 3884 48816 3936 48822
rect 3884 48758 3936 48764
rect 3896 48385 3924 48758
rect 3882 48376 3938 48385
rect 3882 48311 3938 48320
rect 3792 48000 3844 48006
rect 3792 47942 3844 47948
rect 2596 47728 2648 47734
rect 1858 47696 1914 47705
rect 2596 47670 2648 47676
rect 2688 47728 2740 47734
rect 2688 47670 2740 47676
rect 1858 47631 1860 47640
rect 1912 47631 1914 47640
rect 2504 47660 2556 47666
rect 1860 47602 1912 47608
rect 2504 47602 2556 47608
rect 2412 47524 2464 47530
rect 2412 47466 2464 47472
rect 2228 47048 2280 47054
rect 2228 46990 2280 46996
rect 1584 46912 1636 46918
rect 1584 46854 1636 46860
rect 1596 46034 1624 46854
rect 1952 46504 2004 46510
rect 1952 46446 2004 46452
rect 1584 46028 1636 46034
rect 1584 45970 1636 45976
rect 1964 45082 1992 46446
rect 2240 45490 2268 46990
rect 2228 45484 2280 45490
rect 2228 45426 2280 45432
rect 2424 45422 2452 47466
rect 2412 45416 2464 45422
rect 2412 45358 2464 45364
rect 2412 45280 2464 45286
rect 2412 45222 2464 45228
rect 1952 45076 2004 45082
rect 1952 45018 2004 45024
rect 2228 44872 2280 44878
rect 2228 44814 2280 44820
rect 2044 44804 2096 44810
rect 2044 44746 2096 44752
rect 1676 44736 1728 44742
rect 1676 44678 1728 44684
rect 1584 41540 1636 41546
rect 1584 41482 1636 41488
rect 1596 41274 1624 41482
rect 1584 41268 1636 41274
rect 1584 41210 1636 41216
rect 1504 35866 1624 35894
rect 1412 31726 1532 31754
rect 1398 31376 1454 31385
rect 1398 31311 1400 31320
rect 1452 31311 1454 31320
rect 1400 31282 1452 31288
rect 1400 30048 1452 30054
rect 1400 29990 1452 29996
rect 1412 29714 1440 29990
rect 1400 29708 1452 29714
rect 1400 29650 1452 29656
rect 1398 25936 1454 25945
rect 1398 25871 1400 25880
rect 1452 25871 1454 25880
rect 1400 25842 1452 25848
rect 1400 24200 1452 24206
rect 1400 24142 1452 24148
rect 1412 23905 1440 24142
rect 1398 23896 1454 23905
rect 1398 23831 1454 23840
rect 1504 23662 1532 31726
rect 1492 23656 1544 23662
rect 1492 23598 1544 23604
rect 1492 23520 1544 23526
rect 1492 23462 1544 23468
rect 20 20256 72 20262
rect 20 20198 72 20204
rect 32 800 60 20198
rect 1400 19168 1452 19174
rect 1400 19110 1452 19116
rect 1412 18834 1440 19110
rect 1400 18828 1452 18834
rect 1400 18770 1452 18776
rect 1504 16114 1532 23462
rect 1596 21434 1624 35866
rect 1688 28014 1716 44678
rect 2056 44402 2084 44746
rect 2044 44396 2096 44402
rect 2044 44338 2096 44344
rect 1768 43716 1820 43722
rect 1768 43658 1820 43664
rect 1780 35222 1808 43658
rect 1860 41676 1912 41682
rect 1860 41618 1912 41624
rect 1872 41585 1900 41618
rect 1858 41576 1914 41585
rect 1858 41511 1914 41520
rect 1952 40928 2004 40934
rect 1952 40870 2004 40876
rect 1860 40452 1912 40458
rect 1860 40394 1912 40400
rect 1872 40225 1900 40394
rect 1858 40216 1914 40225
rect 1858 40151 1914 40160
rect 1860 37188 1912 37194
rect 1860 37130 1912 37136
rect 1872 36825 1900 37130
rect 1858 36816 1914 36825
rect 1858 36751 1914 36760
rect 1964 36666 1992 40870
rect 2136 39364 2188 39370
rect 2136 39306 2188 39312
rect 2148 39098 2176 39306
rect 2136 39092 2188 39098
rect 2136 39034 2188 39040
rect 2240 38978 2268 44814
rect 2320 41132 2372 41138
rect 2320 41074 2372 41080
rect 2148 38950 2268 38978
rect 2044 37188 2096 37194
rect 2044 37130 2096 37136
rect 2056 36854 2084 37130
rect 2044 36848 2096 36854
rect 2044 36790 2096 36796
rect 1964 36638 2084 36666
rect 1952 36576 2004 36582
rect 1952 36518 2004 36524
rect 1964 35698 1992 36518
rect 1952 35692 2004 35698
rect 1952 35634 2004 35640
rect 1768 35216 1820 35222
rect 1768 35158 1820 35164
rect 1768 35080 1820 35086
rect 1768 35022 1820 35028
rect 1780 34610 1808 35022
rect 1860 35012 1912 35018
rect 1860 34954 1912 34960
rect 1872 34785 1900 34954
rect 1858 34776 1914 34785
rect 1858 34711 1914 34720
rect 1768 34604 1820 34610
rect 1768 34546 1820 34552
rect 1768 33856 1820 33862
rect 1768 33798 1820 33804
rect 1780 33522 1808 33798
rect 1768 33516 1820 33522
rect 1768 33458 1820 33464
rect 1952 33448 2004 33454
rect 1952 33390 2004 33396
rect 1964 33114 1992 33390
rect 1952 33108 2004 33114
rect 1952 33050 2004 33056
rect 1952 32904 2004 32910
rect 1952 32846 2004 32852
rect 1964 32434 1992 32846
rect 1952 32428 2004 32434
rect 1952 32370 2004 32376
rect 1952 32292 2004 32298
rect 1952 32234 2004 32240
rect 1768 31340 1820 31346
rect 1768 31282 1820 31288
rect 1676 28008 1728 28014
rect 1676 27950 1728 27956
rect 1780 27554 1808 31282
rect 1860 30184 1912 30190
rect 1860 30126 1912 30132
rect 1688 27526 1808 27554
rect 1688 25922 1716 27526
rect 1768 27464 1820 27470
rect 1768 27406 1820 27412
rect 1780 26994 1808 27406
rect 1768 26988 1820 26994
rect 1768 26930 1820 26936
rect 1688 25894 1808 25922
rect 1676 25832 1728 25838
rect 1676 25774 1728 25780
rect 1688 25498 1716 25774
rect 1676 25492 1728 25498
rect 1676 25434 1728 25440
rect 1780 24290 1808 25894
rect 1872 24750 1900 30126
rect 1964 27418 1992 32234
rect 2056 31906 2084 36638
rect 2148 32910 2176 38950
rect 2332 38570 2360 41074
rect 2240 38542 2360 38570
rect 2136 32904 2188 32910
rect 2136 32846 2188 32852
rect 2136 32768 2188 32774
rect 2136 32710 2188 32716
rect 2148 32502 2176 32710
rect 2136 32496 2188 32502
rect 2136 32438 2188 32444
rect 2056 31878 2176 31906
rect 2044 31748 2096 31754
rect 2044 31690 2096 31696
rect 2056 30938 2084 31690
rect 2044 30932 2096 30938
rect 2044 30874 2096 30880
rect 2044 28960 2096 28966
rect 2044 28902 2096 28908
rect 2056 28626 2084 28902
rect 2044 28620 2096 28626
rect 2044 28562 2096 28568
rect 1964 27390 2084 27418
rect 1952 27328 2004 27334
rect 1952 27270 2004 27276
rect 1964 27062 1992 27270
rect 1952 27056 2004 27062
rect 1952 26998 2004 27004
rect 1860 24744 1912 24750
rect 1860 24686 1912 24692
rect 1952 24608 2004 24614
rect 1952 24550 2004 24556
rect 1780 24262 1900 24290
rect 1676 24200 1728 24206
rect 1676 24142 1728 24148
rect 1768 24200 1820 24206
rect 1768 24142 1820 24148
rect 1688 23594 1716 24142
rect 1780 23730 1808 24142
rect 1768 23724 1820 23730
rect 1768 23666 1820 23672
rect 1676 23588 1728 23594
rect 1676 23530 1728 23536
rect 1872 23526 1900 24262
rect 1964 23798 1992 24550
rect 1952 23792 2004 23798
rect 1952 23734 2004 23740
rect 1952 23656 2004 23662
rect 1952 23598 2004 23604
rect 1860 23520 1912 23526
rect 1860 23462 1912 23468
rect 1860 22636 1912 22642
rect 1860 22578 1912 22584
rect 1872 22545 1900 22578
rect 1858 22536 1914 22545
rect 1858 22471 1914 22480
rect 1596 21406 1716 21434
rect 1584 18080 1636 18086
rect 1584 18022 1636 18028
rect 1596 17746 1624 18022
rect 1584 17740 1636 17746
rect 1584 17682 1636 17688
rect 1584 16516 1636 16522
rect 1584 16458 1636 16464
rect 1596 16250 1624 16458
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 1492 16108 1544 16114
rect 1492 16050 1544 16056
rect 296 16040 348 16046
rect 296 15982 348 15988
rect 18 0 74 800
rect 308 762 336 15982
rect 1688 15162 1716 21406
rect 1964 18290 1992 23598
rect 2056 22710 2084 27390
rect 2148 27130 2176 31878
rect 2240 30190 2268 38542
rect 2424 34678 2452 45222
rect 2412 34672 2464 34678
rect 2412 34614 2464 34620
rect 2412 32904 2464 32910
rect 2412 32846 2464 32852
rect 2424 31754 2452 32846
rect 2332 31726 2452 31754
rect 2228 30184 2280 30190
rect 2228 30126 2280 30132
rect 2228 30048 2280 30054
rect 2228 29990 2280 29996
rect 2240 29714 2268 29990
rect 2228 29708 2280 29714
rect 2228 29650 2280 29656
rect 2332 28608 2360 31726
rect 2412 30252 2464 30258
rect 2412 30194 2464 30200
rect 2240 28580 2360 28608
rect 2136 27124 2188 27130
rect 2136 27066 2188 27072
rect 2136 25900 2188 25906
rect 2136 25842 2188 25848
rect 2148 24818 2176 25842
rect 2136 24812 2188 24818
rect 2136 24754 2188 24760
rect 2044 22704 2096 22710
rect 2044 22646 2096 22652
rect 2240 22094 2268 28580
rect 2320 28484 2372 28490
rect 2320 28426 2372 28432
rect 2332 28218 2360 28426
rect 2320 28212 2372 28218
rect 2320 28154 2372 28160
rect 2320 28008 2372 28014
rect 2320 27950 2372 27956
rect 2332 24410 2360 27950
rect 2320 24404 2372 24410
rect 2320 24346 2372 24352
rect 2148 22066 2268 22094
rect 2148 20398 2176 22066
rect 2424 20806 2452 30194
rect 2516 25770 2544 47602
rect 2700 47054 2728 47670
rect 3148 47660 3200 47666
rect 3148 47602 3200 47608
rect 2688 47048 2740 47054
rect 2872 47048 2924 47054
rect 2688 46990 2740 46996
rect 2778 47016 2834 47025
rect 2872 46990 2924 46996
rect 2778 46951 2834 46960
rect 2792 46510 2820 46951
rect 2884 46646 2912 46990
rect 2872 46640 2924 46646
rect 2872 46582 2924 46588
rect 2780 46504 2832 46510
rect 2780 46446 2832 46452
rect 2778 46336 2834 46345
rect 2778 46271 2834 46280
rect 2792 46034 2820 46271
rect 2780 46028 2832 46034
rect 2780 45970 2832 45976
rect 2596 45416 2648 45422
rect 2596 45358 2648 45364
rect 2608 36242 2636 45358
rect 3054 44976 3110 44985
rect 3054 44911 3110 44920
rect 3068 44334 3096 44911
rect 2964 44328 3016 44334
rect 2964 44270 3016 44276
rect 3056 44328 3108 44334
rect 3056 44270 3108 44276
rect 2976 43994 3004 44270
rect 2964 43988 3016 43994
rect 2964 43930 3016 43936
rect 2778 39536 2834 39545
rect 2778 39471 2780 39480
rect 2832 39471 2834 39480
rect 2780 39442 2832 39448
rect 2596 36236 2648 36242
rect 2596 36178 2648 36184
rect 2778 36136 2834 36145
rect 2778 36071 2834 36080
rect 2792 35630 2820 36071
rect 2872 36032 2924 36038
rect 2872 35974 2924 35980
rect 2884 35766 2912 35974
rect 2872 35760 2924 35766
rect 2872 35702 2924 35708
rect 2780 35624 2832 35630
rect 2780 35566 2832 35572
rect 2596 35216 2648 35222
rect 2596 35158 2648 35164
rect 2608 27538 2636 35158
rect 2780 34536 2832 34542
rect 2780 34478 2832 34484
rect 2792 34105 2820 34478
rect 2778 34096 2834 34105
rect 2778 34031 2834 34040
rect 2780 33448 2832 33454
rect 2778 33416 2780 33425
rect 2832 33416 2834 33425
rect 2778 33351 2834 33360
rect 2688 32904 2740 32910
rect 2688 32846 2740 32852
rect 2596 27532 2648 27538
rect 2596 27474 2648 27480
rect 2596 27396 2648 27402
rect 2596 27338 2648 27344
rect 2504 25764 2556 25770
rect 2504 25706 2556 25712
rect 2504 25424 2556 25430
rect 2504 25366 2556 25372
rect 2516 21554 2544 25366
rect 2504 21548 2556 21554
rect 2504 21490 2556 21496
rect 2412 20800 2464 20806
rect 2412 20742 2464 20748
rect 2608 20618 2636 27338
rect 2240 20590 2636 20618
rect 2136 20392 2188 20398
rect 2136 20334 2188 20340
rect 1952 18284 2004 18290
rect 1952 18226 2004 18232
rect 1860 17196 1912 17202
rect 1860 17138 1912 17144
rect 1872 17105 1900 17138
rect 1858 17096 1914 17105
rect 1858 17031 1914 17040
rect 1860 16720 1912 16726
rect 1860 16662 1912 16668
rect 1872 16425 1900 16662
rect 1964 16574 1992 18226
rect 2136 16992 2188 16998
rect 2136 16934 2188 16940
rect 2148 16658 2176 16934
rect 2136 16652 2188 16658
rect 2136 16594 2188 16600
rect 1964 16546 2084 16574
rect 1858 16416 1914 16425
rect 1858 16351 1914 16360
rect 1676 15156 1728 15162
rect 1676 15098 1728 15104
rect 1768 14408 1820 14414
rect 1768 14350 1820 14356
rect 1780 13938 1808 14350
rect 1768 13932 1820 13938
rect 1768 13874 1820 13880
rect 1952 13864 2004 13870
rect 1952 13806 2004 13812
rect 1964 13530 1992 13806
rect 1952 13524 2004 13530
rect 1952 13466 2004 13472
rect 1584 13388 1636 13394
rect 1584 13330 1636 13336
rect 1596 12986 1624 13330
rect 2056 13326 2084 16546
rect 2044 13320 2096 13326
rect 2044 13262 2096 13268
rect 2056 12986 2084 13262
rect 1584 12980 1636 12986
rect 1584 12922 1636 12928
rect 2044 12980 2096 12986
rect 2044 12922 2096 12928
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1412 12345 1440 12786
rect 1398 12336 1454 12345
rect 1398 12271 1454 12280
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 1596 11218 1624 11494
rect 1584 11212 1636 11218
rect 1584 11154 1636 11160
rect 1398 10976 1454 10985
rect 1398 10911 1454 10920
rect 1412 10674 1440 10911
rect 1400 10668 1452 10674
rect 1400 10610 1452 10616
rect 2240 10554 2268 20590
rect 2700 20482 2728 32846
rect 2778 32736 2834 32745
rect 2778 32671 2834 32680
rect 2792 32366 2820 32671
rect 2780 32360 2832 32366
rect 2780 32302 2832 32308
rect 2870 32056 2926 32065
rect 2870 31991 2926 32000
rect 2884 31890 2912 31991
rect 2780 31884 2832 31890
rect 2780 31826 2832 31832
rect 2872 31884 2924 31890
rect 2872 31826 2924 31832
rect 2792 31482 2820 31826
rect 2780 31476 2832 31482
rect 2780 31418 2832 31424
rect 2778 30016 2834 30025
rect 2778 29951 2834 29960
rect 2792 29714 2820 29951
rect 2780 29708 2832 29714
rect 2780 29650 2832 29656
rect 2778 28656 2834 28665
rect 2778 28591 2780 28600
rect 2832 28591 2834 28600
rect 2780 28562 2832 28568
rect 3160 28082 3188 47602
rect 3988 47258 4016 49030
rect 4172 48686 4200 49286
rect 4620 49156 4672 49162
rect 4620 49098 4672 49104
rect 4068 48680 4120 48686
rect 4068 48622 4120 48628
rect 4160 48680 4212 48686
rect 4160 48622 4212 48628
rect 4080 48328 4108 48622
rect 4214 48444 4522 48464
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48368 4522 48388
rect 4080 48300 4200 48328
rect 4172 47802 4200 48300
rect 4160 47796 4212 47802
rect 4160 47738 4212 47744
rect 4068 47660 4120 47666
rect 4068 47602 4120 47608
rect 3976 47252 4028 47258
rect 3976 47194 4028 47200
rect 3332 43784 3384 43790
rect 3332 43726 3384 43732
rect 2872 28076 2924 28082
rect 2872 28018 2924 28024
rect 3148 28076 3200 28082
rect 3148 28018 3200 28024
rect 2778 27296 2834 27305
rect 2778 27231 2834 27240
rect 2792 26926 2820 27231
rect 2780 26920 2832 26926
rect 2780 26862 2832 26868
rect 2778 26616 2834 26625
rect 2778 26551 2834 26560
rect 2792 26450 2820 26551
rect 2780 26444 2832 26450
rect 2780 26386 2832 26392
rect 2780 26308 2832 26314
rect 2780 26250 2832 26256
rect 2792 26042 2820 26250
rect 2780 26036 2832 26042
rect 2780 25978 2832 25984
rect 2884 25430 2912 28018
rect 2964 27532 3016 27538
rect 2964 27474 3016 27480
rect 2976 26586 3004 27474
rect 3056 27464 3108 27470
rect 3056 27406 3108 27412
rect 2964 26580 3016 26586
rect 2964 26522 3016 26528
rect 3068 26518 3096 27406
rect 3056 26512 3108 26518
rect 3056 26454 3108 26460
rect 2872 25424 2924 25430
rect 2872 25366 2924 25372
rect 2780 23656 2832 23662
rect 2780 23598 2832 23604
rect 2792 23225 2820 23598
rect 2778 23216 2834 23225
rect 2778 23151 2834 23160
rect 2872 22092 2924 22098
rect 2872 22034 2924 22040
rect 2884 21865 2912 22034
rect 2870 21856 2926 21865
rect 2870 21791 2926 21800
rect 2608 20454 2728 20482
rect 2412 19372 2464 19378
rect 2412 19314 2464 19320
rect 2320 19168 2372 19174
rect 2320 19110 2372 19116
rect 2332 18834 2360 19110
rect 2320 18828 2372 18834
rect 2320 18770 2372 18776
rect 2320 11076 2372 11082
rect 2320 11018 2372 11024
rect 2332 10674 2360 11018
rect 2320 10668 2372 10674
rect 2320 10610 2372 10616
rect 2240 10526 2360 10554
rect 1768 10056 1820 10062
rect 1768 9998 1820 10004
rect 1780 9586 1808 9998
rect 1768 9580 1820 9586
rect 1768 9522 1820 9528
rect 2228 9512 2280 9518
rect 2228 9454 2280 9460
rect 2240 9178 2268 9454
rect 2228 9172 2280 9178
rect 2228 9114 2280 9120
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 1872 8265 1900 8434
rect 1858 8256 1914 8265
rect 1858 8191 1914 8200
rect 1860 7812 1912 7818
rect 1860 7754 1912 7760
rect 1872 7585 1900 7754
rect 1858 7576 1914 7585
rect 1858 7511 1914 7520
rect 2044 7200 2096 7206
rect 2044 7142 2096 7148
rect 2056 6322 2084 7142
rect 2228 6656 2280 6662
rect 2228 6598 2280 6604
rect 2240 6390 2268 6598
rect 2228 6384 2280 6390
rect 2228 6326 2280 6332
rect 2044 6316 2096 6322
rect 2044 6258 2096 6264
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1596 5234 1624 6054
rect 2332 5778 2360 10526
rect 2424 6186 2452 19314
rect 2608 16522 2636 20454
rect 2780 20324 2832 20330
rect 2780 20266 2832 20272
rect 2792 19825 2820 20266
rect 2778 19816 2834 19825
rect 2778 19751 2834 19760
rect 2778 19136 2834 19145
rect 2778 19071 2834 19080
rect 2792 18834 2820 19071
rect 2780 18828 2832 18834
rect 2780 18770 2832 18776
rect 2872 18080 2924 18086
rect 2872 18022 2924 18028
rect 2884 17814 2912 18022
rect 2872 17808 2924 17814
rect 2778 17776 2834 17785
rect 2872 17750 2924 17756
rect 2778 17711 2780 17720
rect 2832 17711 2834 17720
rect 2780 17682 2832 17688
rect 3344 16658 3372 43726
rect 3700 40452 3752 40458
rect 3700 40394 3752 40400
rect 3514 38176 3570 38185
rect 3514 38111 3570 38120
rect 3424 36168 3476 36174
rect 3424 36110 3476 36116
rect 3436 30394 3464 36110
rect 3528 35894 3556 38111
rect 3528 35866 3648 35894
rect 3620 30546 3648 35866
rect 3712 31346 3740 40394
rect 3700 31340 3752 31346
rect 3700 31282 3752 31288
rect 3620 30518 3740 30546
rect 3424 30388 3476 30394
rect 3424 30330 3476 30336
rect 3436 29458 3464 30330
rect 3436 29430 3556 29458
rect 3422 29336 3478 29345
rect 3422 29271 3478 29280
rect 3436 29034 3464 29271
rect 3424 29028 3476 29034
rect 3424 28970 3476 28976
rect 3528 28914 3556 29430
rect 3436 28886 3556 28914
rect 3436 22642 3464 28886
rect 3712 28778 3740 30518
rect 3528 28750 3740 28778
rect 3528 23526 3556 28750
rect 3516 23520 3568 23526
rect 3516 23462 3568 23468
rect 3424 22636 3476 22642
rect 3424 22578 3476 22584
rect 3436 22030 3464 22578
rect 3516 22432 3568 22438
rect 3516 22374 3568 22380
rect 3424 22024 3476 22030
rect 3424 21966 3476 21972
rect 3528 21622 3556 22374
rect 3792 22024 3844 22030
rect 3792 21966 3844 21972
rect 3804 21690 3832 21966
rect 3792 21684 3844 21690
rect 3792 21626 3844 21632
rect 3516 21616 3568 21622
rect 3516 21558 3568 21564
rect 3422 21176 3478 21185
rect 3422 21111 3478 21120
rect 3436 21010 3464 21111
rect 3424 21004 3476 21010
rect 3424 20946 3476 20952
rect 3422 18456 3478 18465
rect 3422 18391 3478 18400
rect 3436 18154 3464 18391
rect 3424 18148 3476 18154
rect 3424 18090 3476 18096
rect 3332 16652 3384 16658
rect 3332 16594 3384 16600
rect 2596 16516 2648 16522
rect 2596 16458 2648 16464
rect 4080 14890 4108 47602
rect 4214 47356 4522 47376
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47280 4522 47300
rect 4214 46268 4522 46288
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46192 4522 46212
rect 4214 45180 4522 45200
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45104 4522 45124
rect 4214 44092 4522 44112
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44016 4522 44036
rect 4214 43004 4522 43024
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42928 4522 42948
rect 4214 41916 4522 41936
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41840 4522 41860
rect 4214 40828 4522 40848
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40752 4522 40772
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 4632 15706 4660 49098
rect 4908 48822 4936 51326
rect 5170 51326 5488 51354
rect 5170 51200 5226 51326
rect 5172 49156 5224 49162
rect 5172 49098 5224 49104
rect 4896 48816 4948 48822
rect 4896 48758 4948 48764
rect 5184 48278 5212 49098
rect 5264 49088 5316 49094
rect 5264 49030 5316 49036
rect 5172 48272 5224 48278
rect 5172 48214 5224 48220
rect 4804 47524 4856 47530
rect 4804 47466 4856 47472
rect 4816 47122 4844 47466
rect 4988 47456 5040 47462
rect 4988 47398 5040 47404
rect 5000 47122 5028 47398
rect 4804 47116 4856 47122
rect 4804 47058 4856 47064
rect 4988 47116 5040 47122
rect 4988 47058 5040 47064
rect 5276 25974 5304 49030
rect 5460 47802 5488 51326
rect 5814 51200 5870 52000
rect 6458 51354 6514 52000
rect 7102 51354 7158 52000
rect 7746 51354 7802 52000
rect 8390 51354 8446 52000
rect 6458 51326 6592 51354
rect 6458 51200 6514 51326
rect 5816 49292 5868 49298
rect 5816 49234 5868 49240
rect 5540 48680 5592 48686
rect 5540 48622 5592 48628
rect 5448 47796 5500 47802
rect 5448 47738 5500 47744
rect 5552 47122 5580 48622
rect 5632 48544 5684 48550
rect 5632 48486 5684 48492
rect 5540 47116 5592 47122
rect 5540 47058 5592 47064
rect 5540 38888 5592 38894
rect 5540 38830 5592 38836
rect 5264 25968 5316 25974
rect 5264 25910 5316 25916
rect 5172 21480 5224 21486
rect 5172 21422 5224 21428
rect 5184 20330 5212 21422
rect 5172 20324 5224 20330
rect 5172 20266 5224 20272
rect 5552 16574 5580 38830
rect 5644 38418 5672 48486
rect 5828 48210 5856 49234
rect 6564 49230 6592 51326
rect 7102 51326 7236 51354
rect 7102 51200 7158 51326
rect 6552 49224 6604 49230
rect 6552 49166 6604 49172
rect 6736 49088 6788 49094
rect 6736 49030 6788 49036
rect 5816 48204 5868 48210
rect 5816 48146 5868 48152
rect 6184 48068 6236 48074
rect 6184 48010 6236 48016
rect 6196 47462 6224 48010
rect 6644 48000 6696 48006
rect 6644 47942 6696 47948
rect 6656 47734 6684 47942
rect 6644 47728 6696 47734
rect 6644 47670 6696 47676
rect 6184 47456 6236 47462
rect 6184 47398 6236 47404
rect 6196 47054 6224 47398
rect 6184 47048 6236 47054
rect 6184 46990 6236 46996
rect 6644 39432 6696 39438
rect 6644 39374 6696 39380
rect 6656 38962 6684 39374
rect 6644 38956 6696 38962
rect 6644 38898 6696 38904
rect 5632 38412 5684 38418
rect 5632 38354 5684 38360
rect 6748 24682 6776 49030
rect 7208 48686 7236 51326
rect 7746 51326 7880 51354
rect 7746 51200 7802 51326
rect 7472 49224 7524 49230
rect 7472 49166 7524 49172
rect 7484 48822 7512 49166
rect 7472 48816 7524 48822
rect 7472 48758 7524 48764
rect 6920 48680 6972 48686
rect 6920 48622 6972 48628
rect 7196 48680 7248 48686
rect 7196 48622 7248 48628
rect 6932 48346 6960 48622
rect 6920 48340 6972 48346
rect 6920 48282 6972 48288
rect 7012 48136 7064 48142
rect 7012 48078 7064 48084
rect 7380 48136 7432 48142
rect 7380 48078 7432 48084
rect 6828 47592 6880 47598
rect 6828 47534 6880 47540
rect 6840 39386 6868 47534
rect 6840 39358 6960 39386
rect 6828 39296 6880 39302
rect 6828 39238 6880 39244
rect 6840 39030 6868 39238
rect 6828 39024 6880 39030
rect 6828 38966 6880 38972
rect 6932 38842 6960 39358
rect 6840 38814 6960 38842
rect 6840 25226 6868 38814
rect 7024 27606 7052 48078
rect 7392 47666 7420 48078
rect 7380 47660 7432 47666
rect 7380 47602 7432 47608
rect 7852 47598 7880 51326
rect 8312 51326 8446 51354
rect 8208 49904 8260 49910
rect 8208 49846 8260 49852
rect 8220 48822 8248 49846
rect 8208 48816 8260 48822
rect 8208 48758 8260 48764
rect 7840 47592 7892 47598
rect 7840 47534 7892 47540
rect 7472 45892 7524 45898
rect 7472 45834 7524 45840
rect 7484 39438 7512 45834
rect 7472 39432 7524 39438
rect 7472 39374 7524 39380
rect 7012 27600 7064 27606
rect 7012 27542 7064 27548
rect 8312 27334 8340 51326
rect 8390 51200 8446 51326
rect 9034 51200 9090 52000
rect 9678 51200 9734 52000
rect 10322 51200 10378 52000
rect 10966 51354 11022 52000
rect 10704 51326 11022 51354
rect 9128 48680 9180 48686
rect 9128 48622 9180 48628
rect 9140 48346 9168 48622
rect 9128 48340 9180 48346
rect 9128 48282 9180 48288
rect 9692 48278 9720 51200
rect 10336 49298 10364 51200
rect 10324 49292 10376 49298
rect 10324 49234 10376 49240
rect 10140 49088 10192 49094
rect 10140 49030 10192 49036
rect 9680 48272 9732 48278
rect 9680 48214 9732 48220
rect 10152 48210 10180 49030
rect 10232 48680 10284 48686
rect 10232 48622 10284 48628
rect 10140 48204 10192 48210
rect 10140 48146 10192 48152
rect 10244 47802 10272 48622
rect 10508 48000 10560 48006
rect 10508 47942 10560 47948
rect 10232 47796 10284 47802
rect 10232 47738 10284 47744
rect 10520 47598 10548 47942
rect 10508 47592 10560 47598
rect 10508 47534 10560 47540
rect 9956 47524 10008 47530
rect 9956 47466 10008 47472
rect 9968 46578 9996 47466
rect 10520 47054 10548 47534
rect 10508 47048 10560 47054
rect 10508 46990 10560 46996
rect 9956 46572 10008 46578
rect 9956 46514 10008 46520
rect 10704 46442 10732 51326
rect 10966 51200 11022 51326
rect 11610 51200 11666 52000
rect 12254 51354 12310 52000
rect 12898 51354 12954 52000
rect 13542 51354 13598 52000
rect 12254 51326 12388 51354
rect 12254 51200 12310 51326
rect 11624 48754 11652 51200
rect 12360 49586 12388 51326
rect 12898 51326 13124 51354
rect 12898 51200 12954 51326
rect 12360 49558 12664 49586
rect 12348 49292 12400 49298
rect 12348 49234 12400 49240
rect 11704 49156 11756 49162
rect 11704 49098 11756 49104
rect 11612 48748 11664 48754
rect 11612 48690 11664 48696
rect 11716 48278 11744 49098
rect 12360 48754 12388 49234
rect 12348 48748 12400 48754
rect 12348 48690 12400 48696
rect 12636 48686 12664 49558
rect 12532 48680 12584 48686
rect 12532 48622 12584 48628
rect 12624 48680 12676 48686
rect 12624 48622 12676 48628
rect 11796 48544 11848 48550
rect 11796 48486 11848 48492
rect 11704 48272 11756 48278
rect 11704 48214 11756 48220
rect 10876 48068 10928 48074
rect 10876 48010 10928 48016
rect 10888 47802 10916 48010
rect 10876 47796 10928 47802
rect 10876 47738 10928 47744
rect 10784 47660 10836 47666
rect 10784 47602 10836 47608
rect 10968 47660 11020 47666
rect 10968 47602 11020 47608
rect 10796 47122 10824 47602
rect 10784 47116 10836 47122
rect 10784 47058 10836 47064
rect 10692 46436 10744 46442
rect 10692 46378 10744 46384
rect 8852 29164 8904 29170
rect 8852 29106 8904 29112
rect 8300 27328 8352 27334
rect 8300 27270 8352 27276
rect 6828 25220 6880 25226
rect 6828 25162 6880 25168
rect 6736 24676 6788 24682
rect 6736 24618 6788 24624
rect 5552 16546 6132 16574
rect 4620 15700 4672 15706
rect 4620 15642 4672 15648
rect 4068 14884 4120 14890
rect 4068 14826 4120 14832
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 2792 13705 2820 13806
rect 3056 13796 3108 13802
rect 3056 13738 3108 13744
rect 2778 13696 2834 13705
rect 2778 13631 2834 13640
rect 3068 13025 3096 13738
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 3054 13016 3110 13025
rect 3054 12951 3110 12960
rect 3516 12776 3568 12782
rect 3516 12718 3568 12724
rect 2780 11212 2832 11218
rect 2780 11154 2832 11160
rect 2792 10305 2820 11154
rect 2778 10296 2834 10305
rect 2778 10231 2834 10240
rect 3148 9648 3200 9654
rect 2778 9616 2834 9625
rect 3148 9590 3200 9596
rect 2778 9551 2834 9560
rect 2792 9518 2820 9551
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 3160 8945 3188 9590
rect 3146 8936 3202 8945
rect 3146 8871 3202 8880
rect 2778 6896 2834 6905
rect 2778 6831 2834 6840
rect 3424 6860 3476 6866
rect 2792 6254 2820 6831
rect 3424 6802 3476 6808
rect 2780 6248 2832 6254
rect 3436 6225 3464 6802
rect 2780 6190 2832 6196
rect 3422 6216 3478 6225
rect 2412 6180 2464 6186
rect 2412 6122 2464 6128
rect 2688 6180 2740 6186
rect 3422 6151 3478 6160
rect 2688 6122 2740 6128
rect 2320 5772 2372 5778
rect 2320 5714 2372 5720
rect 2700 5710 2728 6122
rect 1768 5704 1820 5710
rect 1768 5646 1820 5652
rect 2688 5704 2740 5710
rect 2688 5646 2740 5652
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 1780 4690 1808 5646
rect 1952 5568 2004 5574
rect 2964 5568 3016 5574
rect 1952 5510 2004 5516
rect 2778 5536 2834 5545
rect 1964 5302 1992 5510
rect 2964 5510 3016 5516
rect 2778 5471 2834 5480
rect 1952 5296 2004 5302
rect 1952 5238 2004 5244
rect 2792 5166 2820 5471
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 2778 4856 2834 4865
rect 2778 4791 2834 4800
rect 2792 4690 2820 4791
rect 1768 4684 1820 4690
rect 1768 4626 1820 4632
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 2976 4554 3004 5510
rect 3424 5364 3476 5370
rect 3424 5306 3476 5312
rect 2964 4548 3016 4554
rect 2964 4490 3016 4496
rect 3436 4185 3464 5306
rect 3422 4176 3478 4185
rect 1584 4140 1636 4146
rect 1584 4082 1636 4088
rect 3056 4140 3108 4146
rect 3422 4111 3478 4120
rect 3056 4082 3108 4088
rect 1596 3398 1624 4082
rect 1952 3936 2004 3942
rect 1952 3878 2004 3884
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 1860 3596 1912 3602
rect 1860 3538 1912 3544
rect 1872 3505 1900 3538
rect 1858 3496 1914 3505
rect 1858 3431 1914 3440
rect 1584 3392 1636 3398
rect 1584 3334 1636 3340
rect 1964 3126 1992 3878
rect 2332 3670 2360 3878
rect 2320 3664 2372 3670
rect 2320 3606 2372 3612
rect 2596 3460 2648 3466
rect 2596 3402 2648 3408
rect 1952 3120 2004 3126
rect 1952 3062 2004 3068
rect 1308 2916 1360 2922
rect 1308 2858 1360 2864
rect 584 870 704 898
rect 584 762 612 870
rect 676 800 704 870
rect 1320 800 1348 2858
rect 1400 2440 1452 2446
rect 1400 2382 1452 2388
rect 1952 2440 2004 2446
rect 1952 2382 2004 2388
rect 308 734 612 762
rect 662 0 718 800
rect 1306 0 1362 800
rect 1412 785 1440 2382
rect 1964 800 1992 2382
rect 2608 800 2636 3402
rect 3068 3194 3096 4082
rect 3148 3936 3200 3942
rect 3148 3878 3200 3884
rect 3160 3602 3188 3878
rect 3240 3664 3292 3670
rect 3240 3606 3292 3612
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 3056 3188 3108 3194
rect 3056 3130 3108 3136
rect 2964 2984 3016 2990
rect 2964 2926 3016 2932
rect 2976 2650 3004 2926
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 3252 800 3280 3606
rect 3422 2136 3478 2145
rect 3422 2071 3478 2080
rect 3436 2038 3464 2071
rect 3424 2032 3476 2038
rect 3424 1974 3476 1980
rect 1398 776 1454 785
rect 1398 711 1454 720
rect 1950 0 2006 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3528 762 3556 12718
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 3884 3936 3936 3942
rect 3884 3878 3936 3884
rect 3896 3738 3924 3878
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 5816 3664 5868 3670
rect 5816 3606 5868 3612
rect 3792 3528 3844 3534
rect 3792 3470 3844 3476
rect 3804 3058 3832 3470
rect 3792 3052 3844 3058
rect 3792 2994 3844 3000
rect 5172 2916 5224 2922
rect 5172 2858 5224 2864
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 4528 2372 4580 2378
rect 4528 2314 4580 2320
rect 3804 870 3924 898
rect 3804 762 3832 870
rect 3896 800 3924 870
rect 4540 800 4568 2314
rect 4988 2304 5040 2310
rect 4988 2246 5040 2252
rect 5000 1902 5028 2246
rect 4988 1896 5040 1902
rect 4988 1838 5040 1844
rect 5184 800 5212 2858
rect 5828 800 5856 3606
rect 3528 734 3832 762
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6104 762 6132 16546
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 6196 3602 6224 4558
rect 6552 3936 6604 3942
rect 6552 3878 6604 3884
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 6184 3596 6236 3602
rect 6184 3538 6236 3544
rect 6564 3126 6592 3878
rect 7116 3602 7144 3878
rect 7104 3596 7156 3602
rect 7104 3538 7156 3544
rect 6552 3120 6604 3126
rect 6552 3062 6604 3068
rect 8392 3052 8444 3058
rect 8392 2994 8444 3000
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 6380 870 6500 898
rect 6380 762 6408 870
rect 6472 800 6500 870
rect 7116 800 7144 2382
rect 7484 1970 7512 2382
rect 7472 1964 7524 1970
rect 7472 1906 7524 1912
rect 7760 800 7788 2382
rect 8404 800 8432 2994
rect 8864 2922 8892 29106
rect 10796 19854 10824 47058
rect 10980 46986 11008 47602
rect 10968 46980 11020 46986
rect 10968 46922 11020 46928
rect 10980 46714 11008 46922
rect 10968 46708 11020 46714
rect 10968 46650 11020 46656
rect 10980 45966 11008 46650
rect 10968 45960 11020 45966
rect 10968 45902 11020 45908
rect 11808 35894 11836 48486
rect 12544 47802 12572 48622
rect 13096 48142 13124 51326
rect 13542 51326 13768 51354
rect 13542 51200 13598 51326
rect 13740 48906 13768 51326
rect 14186 51200 14242 52000
rect 14830 51354 14886 52000
rect 15474 51354 15530 52000
rect 14830 51326 14964 51354
rect 14830 51200 14886 51326
rect 14200 49230 14228 51200
rect 14188 49224 14240 49230
rect 14188 49166 14240 49172
rect 13740 48878 13860 48906
rect 13832 48822 13860 48878
rect 13820 48816 13872 48822
rect 13820 48758 13872 48764
rect 14832 48544 14884 48550
rect 14832 48486 14884 48492
rect 13084 48136 13136 48142
rect 13084 48078 13136 48084
rect 14464 48136 14516 48142
rect 14464 48078 14516 48084
rect 14372 48068 14424 48074
rect 14372 48010 14424 48016
rect 14384 47802 14412 48010
rect 12532 47796 12584 47802
rect 12532 47738 12584 47744
rect 14372 47796 14424 47802
rect 14372 47738 14424 47744
rect 13176 47728 13228 47734
rect 13176 47670 13228 47676
rect 12348 47592 12400 47598
rect 12348 47534 12400 47540
rect 12360 47190 12388 47534
rect 12348 47184 12400 47190
rect 12348 47126 12400 47132
rect 12256 46980 12308 46986
rect 12256 46922 12308 46928
rect 11808 35866 11928 35894
rect 11796 26920 11848 26926
rect 11796 26862 11848 26868
rect 11060 26852 11112 26858
rect 11060 26794 11112 26800
rect 10784 19848 10836 19854
rect 10784 19790 10836 19796
rect 11072 16574 11100 26794
rect 11808 26586 11836 26862
rect 11796 26580 11848 26586
rect 11796 26522 11848 26528
rect 11808 26042 11836 26522
rect 11796 26036 11848 26042
rect 11796 25978 11848 25984
rect 11900 25498 11928 35866
rect 12268 27402 12296 46922
rect 12256 27396 12308 27402
rect 12256 27338 12308 27344
rect 11888 25492 11940 25498
rect 11888 25434 11940 25440
rect 11888 20392 11940 20398
rect 11888 20334 11940 20340
rect 11900 20058 11928 20334
rect 11888 20052 11940 20058
rect 11888 19994 11940 20000
rect 12360 19378 12388 47126
rect 13188 46714 13216 47670
rect 14476 47666 14504 48078
rect 13268 47660 13320 47666
rect 13268 47602 13320 47608
rect 14464 47660 14516 47666
rect 14464 47602 14516 47608
rect 13176 46708 13228 46714
rect 13176 46650 13228 46656
rect 13188 45554 13216 46650
rect 13004 45526 13216 45554
rect 13004 45490 13032 45526
rect 12992 45484 13044 45490
rect 12992 45426 13044 45432
rect 12624 32428 12676 32434
rect 12624 32370 12676 32376
rect 12636 28082 12664 32370
rect 12624 28076 12676 28082
rect 12624 28018 12676 28024
rect 12716 27872 12768 27878
rect 12716 27814 12768 27820
rect 12728 27062 12756 27814
rect 12716 27056 12768 27062
rect 12716 26998 12768 27004
rect 13004 22094 13032 45426
rect 12912 22066 13032 22094
rect 12348 19372 12400 19378
rect 12348 19314 12400 19320
rect 11072 16546 11284 16574
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 8852 2916 8904 2922
rect 8852 2858 8904 2864
rect 9048 800 9076 3674
rect 10324 3664 10376 3670
rect 10324 3606 10376 3612
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 9692 800 9720 2382
rect 10336 800 10364 3606
rect 10968 2916 11020 2922
rect 10968 2858 11020 2864
rect 10414 2408 10470 2417
rect 10414 2343 10470 2352
rect 10428 2310 10456 2343
rect 10416 2304 10468 2310
rect 10416 2246 10468 2252
rect 10980 800 11008 2858
rect 6104 734 6408 762
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11256 762 11284 16546
rect 12912 12434 12940 22066
rect 12992 15904 13044 15910
rect 12992 15846 13044 15852
rect 12820 12406 12940 12434
rect 12256 4140 12308 4146
rect 12256 4082 12308 4088
rect 11612 4004 11664 4010
rect 11612 3946 11664 3952
rect 11980 4004 12032 4010
rect 11980 3946 12032 3952
rect 11624 3534 11652 3946
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 11612 3528 11664 3534
rect 11612 3470 11664 3476
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 11624 2854 11652 3334
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 11716 2514 11744 3878
rect 11888 3392 11940 3398
rect 11888 3334 11940 3340
rect 11900 2514 11928 3334
rect 11992 3058 12020 3946
rect 12268 3534 12296 4082
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 12636 3602 12664 3878
rect 12624 3596 12676 3602
rect 12624 3538 12676 3544
rect 12256 3528 12308 3534
rect 12820 3516 12848 12406
rect 12900 3664 12952 3670
rect 13004 3652 13032 15846
rect 13280 15502 13308 47602
rect 14844 30258 14872 48486
rect 14936 48210 14964 51326
rect 15212 51326 15530 51354
rect 15016 49088 15068 49094
rect 15016 49030 15068 49036
rect 14924 48204 14976 48210
rect 14924 48146 14976 48152
rect 14924 48000 14976 48006
rect 14924 47942 14976 47948
rect 14936 47802 14964 47942
rect 14924 47796 14976 47802
rect 14924 47738 14976 47744
rect 15028 31142 15056 49030
rect 15212 32978 15240 51326
rect 15474 51200 15530 51326
rect 16118 51354 16174 52000
rect 16118 51326 16528 51354
rect 16118 51200 16174 51326
rect 16500 49212 16528 51326
rect 16762 51200 16818 52000
rect 17406 51354 17462 52000
rect 17406 51326 17908 51354
rect 17406 51200 17462 51326
rect 16776 49722 16804 51200
rect 16776 49694 16988 49722
rect 16580 49224 16632 49230
rect 16500 49184 16580 49212
rect 16580 49166 16632 49172
rect 16960 48686 16988 49694
rect 17224 49088 17276 49094
rect 17224 49030 17276 49036
rect 16856 48680 16908 48686
rect 16856 48622 16908 48628
rect 16948 48680 17000 48686
rect 16948 48622 17000 48628
rect 16868 48346 16896 48622
rect 16856 48340 16908 48346
rect 16856 48282 16908 48288
rect 15844 47660 15896 47666
rect 15844 47602 15896 47608
rect 15200 32972 15252 32978
rect 15200 32914 15252 32920
rect 15568 32904 15620 32910
rect 15568 32846 15620 32852
rect 15580 32026 15608 32846
rect 15752 32836 15804 32842
rect 15752 32778 15804 32784
rect 15764 32570 15792 32778
rect 15752 32564 15804 32570
rect 15752 32506 15804 32512
rect 15660 32224 15712 32230
rect 15660 32166 15712 32172
rect 15568 32020 15620 32026
rect 15568 31962 15620 31968
rect 15672 31754 15700 32166
rect 15856 31754 15884 47602
rect 15936 46572 15988 46578
rect 15936 46514 15988 46520
rect 15948 41414 15976 46514
rect 16764 44872 16816 44878
rect 16764 44814 16816 44820
rect 15948 41386 16068 41414
rect 15660 31748 15712 31754
rect 15856 31726 15976 31754
rect 15660 31690 15712 31696
rect 15016 31136 15068 31142
rect 15016 31078 15068 31084
rect 14832 30252 14884 30258
rect 14832 30194 14884 30200
rect 15476 29028 15528 29034
rect 15476 28970 15528 28976
rect 13820 22568 13872 22574
rect 13820 22510 13872 22516
rect 13728 21684 13780 21690
rect 13728 21626 13780 21632
rect 13740 21418 13768 21626
rect 13832 21554 13860 22510
rect 15200 22500 15252 22506
rect 15200 22442 15252 22448
rect 13912 21956 13964 21962
rect 13912 21898 13964 21904
rect 13924 21690 13952 21898
rect 13912 21684 13964 21690
rect 13912 21626 13964 21632
rect 13820 21548 13872 21554
rect 13820 21490 13872 21496
rect 14924 21548 14976 21554
rect 14924 21490 14976 21496
rect 13728 21412 13780 21418
rect 13728 21354 13780 21360
rect 13832 20330 13860 21490
rect 14936 20942 14964 21490
rect 14924 20936 14976 20942
rect 14924 20878 14976 20884
rect 15212 20466 15240 22442
rect 15488 22098 15516 28970
rect 15752 27600 15804 27606
rect 15752 27542 15804 27548
rect 15764 26994 15792 27542
rect 15752 26988 15804 26994
rect 15752 26930 15804 26936
rect 15844 26784 15896 26790
rect 15844 26726 15896 26732
rect 15856 26450 15884 26726
rect 15844 26444 15896 26450
rect 15844 26386 15896 26392
rect 15660 25696 15712 25702
rect 15660 25638 15712 25644
rect 15672 24818 15700 25638
rect 15660 24812 15712 24818
rect 15660 24754 15712 24760
rect 15568 23860 15620 23866
rect 15568 23802 15620 23808
rect 15476 22092 15528 22098
rect 15476 22034 15528 22040
rect 15476 21480 15528 21486
rect 15476 21422 15528 21428
rect 15200 20460 15252 20466
rect 15200 20402 15252 20408
rect 13820 20324 13872 20330
rect 13820 20266 13872 20272
rect 13832 19854 13860 20266
rect 13820 19848 13872 19854
rect 13820 19790 13872 19796
rect 15212 16590 15240 20402
rect 15384 18352 15436 18358
rect 15384 18294 15436 18300
rect 15396 17882 15424 18294
rect 15384 17876 15436 17882
rect 15384 17818 15436 17824
rect 15200 16584 15252 16590
rect 15200 16526 15252 16532
rect 15384 16584 15436 16590
rect 15384 16526 15436 16532
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 13832 16182 13860 16390
rect 13820 16176 13872 16182
rect 13820 16118 13872 16124
rect 14188 16040 14240 16046
rect 14188 15982 14240 15988
rect 14200 15706 14228 15982
rect 14188 15700 14240 15706
rect 14188 15642 14240 15648
rect 15396 15502 15424 16526
rect 15488 16454 15516 21422
rect 15476 16448 15528 16454
rect 15476 16390 15528 16396
rect 15488 16182 15516 16390
rect 15476 16176 15528 16182
rect 15476 16118 15528 16124
rect 13268 15496 13320 15502
rect 13268 15438 13320 15444
rect 14096 15496 14148 15502
rect 14096 15438 14148 15444
rect 15384 15496 15436 15502
rect 15384 15438 15436 15444
rect 14108 13870 14136 15438
rect 15580 15314 15608 23802
rect 15672 23730 15700 24754
rect 15752 24200 15804 24206
rect 15752 24142 15804 24148
rect 15764 23730 15792 24142
rect 15948 23798 15976 31726
rect 16040 25906 16068 41386
rect 16580 31816 16632 31822
rect 16580 31758 16632 31764
rect 16592 30802 16620 31758
rect 16580 30796 16632 30802
rect 16580 30738 16632 30744
rect 16672 30660 16724 30666
rect 16672 30602 16724 30608
rect 16684 30326 16712 30602
rect 16672 30320 16724 30326
rect 16672 30262 16724 30268
rect 16672 29572 16724 29578
rect 16672 29514 16724 29520
rect 16684 29306 16712 29514
rect 16672 29300 16724 29306
rect 16672 29242 16724 29248
rect 16580 27328 16632 27334
rect 16580 27270 16632 27276
rect 16592 27062 16620 27270
rect 16580 27056 16632 27062
rect 16580 26998 16632 27004
rect 16120 26988 16172 26994
rect 16120 26930 16172 26936
rect 16028 25900 16080 25906
rect 16028 25842 16080 25848
rect 16028 25220 16080 25226
rect 16028 25162 16080 25168
rect 16040 23798 16068 25162
rect 15936 23792 15988 23798
rect 15936 23734 15988 23740
rect 16028 23792 16080 23798
rect 16028 23734 16080 23740
rect 15660 23724 15712 23730
rect 15660 23666 15712 23672
rect 15752 23724 15804 23730
rect 15752 23666 15804 23672
rect 15948 22094 15976 23734
rect 15856 22066 15976 22094
rect 15660 21072 15712 21078
rect 15660 21014 15712 21020
rect 15672 20874 15700 21014
rect 15660 20868 15712 20874
rect 15660 20810 15712 20816
rect 15304 15286 15608 15314
rect 14096 13864 14148 13870
rect 14096 13806 14148 13812
rect 14740 5296 14792 5302
rect 14740 5238 14792 5244
rect 13176 4616 13228 4622
rect 13176 4558 13228 4564
rect 13188 4146 13216 4558
rect 13176 4140 13228 4146
rect 13176 4082 13228 4088
rect 13084 4072 13136 4078
rect 13084 4014 13136 4020
rect 13544 4072 13596 4078
rect 13544 4014 13596 4020
rect 13096 3670 13124 4014
rect 12952 3624 13032 3652
rect 13084 3664 13136 3670
rect 12900 3606 12952 3612
rect 13084 3606 13136 3612
rect 13176 3664 13228 3670
rect 13176 3606 13228 3612
rect 12992 3528 13044 3534
rect 12820 3488 12992 3516
rect 12256 3470 12308 3476
rect 13188 3516 13216 3606
rect 13044 3488 13216 3516
rect 12992 3470 13044 3476
rect 12164 3392 12216 3398
rect 12164 3334 12216 3340
rect 12176 3126 12204 3334
rect 12164 3120 12216 3126
rect 12164 3062 12216 3068
rect 11980 3052 12032 3058
rect 11980 2994 12032 3000
rect 12900 2984 12952 2990
rect 12900 2926 12952 2932
rect 11704 2508 11756 2514
rect 11704 2450 11756 2456
rect 11888 2508 11940 2514
rect 11888 2450 11940 2456
rect 12256 2372 12308 2378
rect 12256 2314 12308 2320
rect 11532 870 11652 898
rect 11532 762 11560 870
rect 11624 800 11652 870
rect 12268 800 12296 2314
rect 12912 800 12940 2926
rect 13556 800 13584 4014
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 14292 3058 14320 3470
rect 14464 3392 14516 3398
rect 14464 3334 14516 3340
rect 14476 3126 14504 3334
rect 14464 3120 14516 3126
rect 14464 3062 14516 3068
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14752 2582 14780 5238
rect 15304 4010 15332 15286
rect 15292 4004 15344 4010
rect 15292 3946 15344 3952
rect 15672 3534 15700 20810
rect 15752 19848 15804 19854
rect 15752 19790 15804 19796
rect 15764 18766 15792 19790
rect 15752 18760 15804 18766
rect 15752 18702 15804 18708
rect 15764 18426 15792 18702
rect 15752 18420 15804 18426
rect 15752 18362 15804 18368
rect 15856 17678 15884 22066
rect 15936 20392 15988 20398
rect 15936 20334 15988 20340
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 15856 16522 15884 17614
rect 15948 17202 15976 20334
rect 16132 17882 16160 26930
rect 16580 26920 16632 26926
rect 16776 26874 16804 44814
rect 17236 44198 17264 49030
rect 17592 48204 17644 48210
rect 17592 48146 17644 48152
rect 17224 44192 17276 44198
rect 17224 44134 17276 44140
rect 17604 41414 17632 48146
rect 17604 41386 17724 41414
rect 16856 32224 16908 32230
rect 16856 32166 16908 32172
rect 16868 32026 16896 32166
rect 16856 32020 16908 32026
rect 16856 31962 16908 31968
rect 16856 31748 16908 31754
rect 16856 31690 16908 31696
rect 16868 31482 16896 31690
rect 16856 31476 16908 31482
rect 16856 31418 16908 31424
rect 17500 31340 17552 31346
rect 17500 31282 17552 31288
rect 17512 30938 17540 31282
rect 17592 31272 17644 31278
rect 17592 31214 17644 31220
rect 17500 30932 17552 30938
rect 17500 30874 17552 30880
rect 17132 30592 17184 30598
rect 17132 30534 17184 30540
rect 17144 30258 17172 30534
rect 17512 30258 17540 30874
rect 17604 30802 17632 31214
rect 17592 30796 17644 30802
rect 17592 30738 17644 30744
rect 17132 30252 17184 30258
rect 17132 30194 17184 30200
rect 17500 30252 17552 30258
rect 17500 30194 17552 30200
rect 17040 30116 17092 30122
rect 17040 30058 17092 30064
rect 16856 29640 16908 29646
rect 16856 29582 16908 29588
rect 16868 28014 16896 29582
rect 17052 29173 17080 30058
rect 17037 29167 17089 29173
rect 17512 29170 17540 30194
rect 17604 30122 17632 30738
rect 17592 30116 17644 30122
rect 17592 30058 17644 30064
rect 17037 29109 17089 29115
rect 17500 29164 17552 29170
rect 17500 29106 17552 29112
rect 17316 28484 17368 28490
rect 17316 28426 17368 28432
rect 16856 28008 16908 28014
rect 16856 27950 16908 27956
rect 16868 27402 16896 27950
rect 17328 27606 17356 28426
rect 17316 27600 17368 27606
rect 17316 27542 17368 27548
rect 16856 27396 16908 27402
rect 16856 27338 16908 27344
rect 16580 26862 16632 26868
rect 16592 25906 16620 26862
rect 16684 26846 16804 26874
rect 16212 25900 16264 25906
rect 16212 25842 16264 25848
rect 16580 25900 16632 25906
rect 16580 25842 16632 25848
rect 16224 25702 16252 25842
rect 16212 25696 16264 25702
rect 16212 25638 16264 25644
rect 16592 25294 16620 25842
rect 16580 25288 16632 25294
rect 16580 25230 16632 25236
rect 16592 24818 16620 25230
rect 16580 24812 16632 24818
rect 16580 24754 16632 24760
rect 16304 24064 16356 24070
rect 16304 24006 16356 24012
rect 16316 23050 16344 24006
rect 16488 23656 16540 23662
rect 16488 23598 16540 23604
rect 16304 23044 16356 23050
rect 16304 22986 16356 22992
rect 16212 20868 16264 20874
rect 16212 20810 16264 20816
rect 16224 20602 16252 20810
rect 16212 20596 16264 20602
rect 16212 20538 16264 20544
rect 16500 20346 16528 23598
rect 16580 22636 16632 22642
rect 16580 22578 16632 22584
rect 16592 21622 16620 22578
rect 16580 21616 16632 21622
rect 16580 21558 16632 21564
rect 16592 20602 16620 21558
rect 16580 20596 16632 20602
rect 16684 20584 16712 26846
rect 16868 23118 16896 27338
rect 17040 26920 17092 26926
rect 17040 26862 17092 26868
rect 17052 26450 17080 26862
rect 17328 26518 17356 27542
rect 17316 26512 17368 26518
rect 17316 26454 17368 26460
rect 17040 26444 17092 26450
rect 17040 26386 17092 26392
rect 17052 25838 17080 26386
rect 17592 26240 17644 26246
rect 17592 26182 17644 26188
rect 17040 25832 17092 25838
rect 17040 25774 17092 25780
rect 17224 25764 17276 25770
rect 17224 25706 17276 25712
rect 16948 24064 17000 24070
rect 16948 24006 17000 24012
rect 16856 23112 16908 23118
rect 16856 23054 16908 23060
rect 16764 23044 16816 23050
rect 16764 22986 16816 22992
rect 16776 20754 16804 22986
rect 16868 22030 16896 23054
rect 16856 22024 16908 22030
rect 16856 21966 16908 21972
rect 16776 20726 16896 20754
rect 16684 20556 16804 20584
rect 16580 20538 16632 20544
rect 16592 20466 16620 20538
rect 16580 20460 16632 20466
rect 16580 20402 16632 20408
rect 16672 20460 16724 20466
rect 16672 20402 16724 20408
rect 16684 20346 16712 20402
rect 16776 20398 16804 20556
rect 16500 20318 16712 20346
rect 16764 20392 16816 20398
rect 16764 20334 16816 20340
rect 16684 20040 16712 20318
rect 16592 20012 16712 20040
rect 16120 17876 16172 17882
rect 16120 17818 16172 17824
rect 15936 17196 15988 17202
rect 15936 17138 15988 17144
rect 15752 16516 15804 16522
rect 15752 16458 15804 16464
rect 15844 16516 15896 16522
rect 15844 16458 15896 16464
rect 15764 15706 15792 16458
rect 15752 15700 15804 15706
rect 15752 15642 15804 15648
rect 15856 15026 15884 16458
rect 15844 15020 15896 15026
rect 15844 14962 15896 14968
rect 15856 13938 15884 14962
rect 15844 13932 15896 13938
rect 15844 13874 15896 13880
rect 15948 11762 15976 17138
rect 15936 11756 15988 11762
rect 15936 11698 15988 11704
rect 16132 3602 16160 17818
rect 16592 17610 16620 20012
rect 16672 18624 16724 18630
rect 16672 18566 16724 18572
rect 16580 17604 16632 17610
rect 16580 17546 16632 17552
rect 16212 16176 16264 16182
rect 16212 16118 16264 16124
rect 16224 4078 16252 16118
rect 16592 15502 16620 17546
rect 16684 17202 16712 18566
rect 16672 17196 16724 17202
rect 16672 17138 16724 17144
rect 16672 16788 16724 16794
rect 16672 16730 16724 16736
rect 16580 15496 16632 15502
rect 16580 15438 16632 15444
rect 16580 15360 16632 15366
rect 16580 15302 16632 15308
rect 16592 14414 16620 15302
rect 16580 14408 16632 14414
rect 16580 14350 16632 14356
rect 16684 13410 16712 16730
rect 16868 15450 16896 20726
rect 16776 15422 16896 15450
rect 16776 14618 16804 15422
rect 16960 14958 16988 24006
rect 17132 23656 17184 23662
rect 17132 23598 17184 23604
rect 17144 22778 17172 23598
rect 17132 22772 17184 22778
rect 17132 22714 17184 22720
rect 17236 22094 17264 25706
rect 17604 25294 17632 26182
rect 17592 25288 17644 25294
rect 17592 25230 17644 25236
rect 17408 25152 17460 25158
rect 17408 25094 17460 25100
rect 17420 24970 17448 25094
rect 17604 24970 17632 25230
rect 17420 24942 17632 24970
rect 17316 24744 17368 24750
rect 17316 24686 17368 24692
rect 17328 23866 17356 24686
rect 17316 23860 17368 23866
rect 17316 23802 17368 23808
rect 17144 22066 17264 22094
rect 17040 16448 17092 16454
rect 17040 16390 17092 16396
rect 17052 16182 17080 16390
rect 17040 16176 17092 16182
rect 17040 16118 17092 16124
rect 16948 14952 17000 14958
rect 16948 14894 17000 14900
rect 16764 14612 16816 14618
rect 16764 14554 16816 14560
rect 16776 13530 16804 14554
rect 16856 13728 16908 13734
rect 16856 13670 16908 13676
rect 16764 13524 16816 13530
rect 16764 13466 16816 13472
rect 16684 13382 16804 13410
rect 16672 12776 16724 12782
rect 16672 12718 16724 12724
rect 16684 12442 16712 12718
rect 16672 12436 16724 12442
rect 16672 12378 16724 12384
rect 16776 4146 16804 13382
rect 16868 12918 16896 13670
rect 16856 12912 16908 12918
rect 16856 12854 16908 12860
rect 17040 9376 17092 9382
rect 17040 9318 17092 9324
rect 17052 9042 17080 9318
rect 17040 9036 17092 9042
rect 17040 8978 17092 8984
rect 16764 4140 16816 4146
rect 16764 4082 16816 4088
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 17144 3942 17172 22066
rect 17224 19984 17276 19990
rect 17224 19926 17276 19932
rect 17236 19446 17264 19926
rect 17224 19440 17276 19446
rect 17224 19382 17276 19388
rect 17328 12434 17356 23802
rect 17420 22094 17448 24942
rect 17500 24812 17552 24818
rect 17500 24754 17552 24760
rect 17512 23662 17540 24754
rect 17592 24268 17644 24274
rect 17592 24210 17644 24216
rect 17500 23656 17552 23662
rect 17500 23598 17552 23604
rect 17604 23322 17632 24210
rect 17592 23316 17644 23322
rect 17592 23258 17644 23264
rect 17420 22066 17540 22094
rect 17408 22024 17460 22030
rect 17408 21966 17460 21972
rect 17420 21554 17448 21966
rect 17408 21548 17460 21554
rect 17408 21490 17460 21496
rect 17408 20936 17460 20942
rect 17408 20878 17460 20884
rect 17420 20806 17448 20878
rect 17408 20800 17460 20806
rect 17408 20742 17460 20748
rect 17420 20058 17448 20742
rect 17408 20052 17460 20058
rect 17408 19994 17460 20000
rect 17408 19372 17460 19378
rect 17408 19314 17460 19320
rect 17420 18630 17448 19314
rect 17408 18624 17460 18630
rect 17408 18566 17460 18572
rect 17328 12406 17448 12434
rect 17420 9178 17448 12406
rect 17408 9172 17460 9178
rect 17408 9114 17460 9120
rect 17316 9036 17368 9042
rect 17316 8978 17368 8984
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 17236 4758 17264 6734
rect 17224 4752 17276 4758
rect 17224 4694 17276 4700
rect 17132 3936 17184 3942
rect 17132 3878 17184 3884
rect 16120 3596 16172 3602
rect 16120 3538 16172 3544
rect 15200 3528 15252 3534
rect 15200 3470 15252 3476
rect 15660 3528 15712 3534
rect 15660 3470 15712 3476
rect 15212 2854 15240 3470
rect 15476 2984 15528 2990
rect 15476 2926 15528 2932
rect 15200 2848 15252 2854
rect 15200 2790 15252 2796
rect 14740 2576 14792 2582
rect 14740 2518 14792 2524
rect 14188 2372 14240 2378
rect 14188 2314 14240 2320
rect 14200 800 14228 2314
rect 15488 800 15516 2926
rect 17328 2922 17356 8978
rect 17420 6610 17448 9114
rect 17512 6798 17540 22066
rect 17592 20256 17644 20262
rect 17592 20198 17644 20204
rect 17604 20058 17632 20198
rect 17592 20052 17644 20058
rect 17592 19994 17644 20000
rect 17696 15706 17724 41386
rect 17776 37732 17828 37738
rect 17776 37674 17828 37680
rect 17788 37262 17816 37674
rect 17776 37256 17828 37262
rect 17776 37198 17828 37204
rect 17776 30048 17828 30054
rect 17776 29990 17828 29996
rect 17788 29170 17816 29990
rect 17776 29164 17828 29170
rect 17776 29106 17828 29112
rect 17776 26308 17828 26314
rect 17776 26250 17828 26256
rect 17684 15700 17736 15706
rect 17684 15642 17736 15648
rect 17684 15088 17736 15094
rect 17684 15030 17736 15036
rect 17696 14414 17724 15030
rect 17684 14408 17736 14414
rect 17684 14350 17736 14356
rect 17696 13938 17724 14350
rect 17684 13932 17736 13938
rect 17684 13874 17736 13880
rect 17788 12434 17816 26250
rect 17880 24818 17908 51326
rect 18050 51200 18106 52000
rect 18694 51200 18750 52000
rect 19338 51200 19394 52000
rect 19982 51354 20038 52000
rect 19982 51326 20208 51354
rect 19982 51200 20038 51326
rect 18064 49298 18092 51200
rect 18052 49292 18104 49298
rect 18052 49234 18104 49240
rect 19352 49230 19380 51200
rect 20180 49230 20208 51326
rect 20626 51200 20682 52000
rect 21270 51200 21326 52000
rect 21914 51354 21970 52000
rect 21914 51326 22048 51354
rect 21914 51200 21970 51326
rect 19340 49224 19392 49230
rect 19340 49166 19392 49172
rect 20168 49224 20220 49230
rect 20168 49166 20220 49172
rect 20076 49088 20128 49094
rect 20076 49030 20128 49036
rect 20260 49088 20312 49094
rect 20260 49030 20312 49036
rect 19574 48988 19882 49008
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48912 19882 48932
rect 19432 48816 19484 48822
rect 19432 48758 19484 48764
rect 19444 48278 19472 48758
rect 19524 48680 19576 48686
rect 19524 48622 19576 48628
rect 19432 48272 19484 48278
rect 19432 48214 19484 48220
rect 19536 47988 19564 48622
rect 19984 48272 20036 48278
rect 19984 48214 20036 48220
rect 19444 47960 19564 47988
rect 19444 47802 19472 47960
rect 19574 47900 19882 47920
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47824 19882 47844
rect 18512 47796 18564 47802
rect 18512 47738 18564 47744
rect 19432 47796 19484 47802
rect 19432 47738 19484 47744
rect 18052 47660 18104 47666
rect 18052 47602 18104 47608
rect 18064 41414 18092 47602
rect 18524 47258 18552 47738
rect 19996 47734 20024 48214
rect 19984 47728 20036 47734
rect 19984 47670 20036 47676
rect 18512 47252 18564 47258
rect 18512 47194 18564 47200
rect 19574 46812 19882 46832
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46736 19882 46756
rect 19574 45724 19882 45744
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45648 19882 45668
rect 19432 45280 19484 45286
rect 19432 45222 19484 45228
rect 18064 41386 18276 41414
rect 18144 37120 18196 37126
rect 18144 37062 18196 37068
rect 18156 36786 18184 37062
rect 18144 36780 18196 36786
rect 18144 36722 18196 36728
rect 18052 36712 18104 36718
rect 18248 36666 18276 41386
rect 19340 37868 19392 37874
rect 19340 37810 19392 37816
rect 19352 37466 19380 37810
rect 19340 37460 19392 37466
rect 19340 37402 19392 37408
rect 19340 37120 19392 37126
rect 19340 37062 19392 37068
rect 18052 36654 18104 36660
rect 18064 35766 18092 36654
rect 18156 36638 18276 36666
rect 18052 35760 18104 35766
rect 18052 35702 18104 35708
rect 17960 32224 18012 32230
rect 17960 32166 18012 32172
rect 17972 31414 18000 32166
rect 18156 31754 18184 36638
rect 19352 36224 19380 37062
rect 19260 36196 19380 36224
rect 19260 36122 19288 36196
rect 19168 36106 19288 36122
rect 19156 36100 19288 36106
rect 19208 36094 19288 36100
rect 19340 36100 19392 36106
rect 19156 36042 19208 36048
rect 19340 36042 19392 36048
rect 18236 36032 18288 36038
rect 18236 35974 18288 35980
rect 18248 35698 18276 35974
rect 18236 35692 18288 35698
rect 18236 35634 18288 35640
rect 19168 35630 19196 36042
rect 19156 35624 19208 35630
rect 19156 35566 19208 35572
rect 19352 35290 19380 36042
rect 19340 35284 19392 35290
rect 19340 35226 19392 35232
rect 19444 34762 19472 45222
rect 19574 44636 19882 44656
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44560 19882 44580
rect 19574 43548 19882 43568
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43472 19882 43492
rect 19574 42460 19882 42480
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42384 19882 42404
rect 19574 41372 19882 41392
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41296 19882 41316
rect 19574 40284 19882 40304
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40208 19882 40228
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 19800 37800 19852 37806
rect 19800 37742 19852 37748
rect 19708 37664 19760 37670
rect 19708 37606 19760 37612
rect 19720 37194 19748 37606
rect 19812 37194 19840 37742
rect 20088 37466 20116 49030
rect 20272 45554 20300 49030
rect 20640 48686 20668 51200
rect 22020 49298 22048 51326
rect 22558 51200 22614 52000
rect 23202 51354 23258 52000
rect 23846 51354 23902 52000
rect 24490 51354 24546 52000
rect 23202 51326 23428 51354
rect 23202 51200 23258 51326
rect 22008 49292 22060 49298
rect 22008 49234 22060 49240
rect 22284 49224 22336 49230
rect 22284 49166 22336 49172
rect 20628 48680 20680 48686
rect 20628 48622 20680 48628
rect 22100 48204 22152 48210
rect 22100 48146 22152 48152
rect 22112 48074 22140 48146
rect 22008 48068 22060 48074
rect 22008 48010 22060 48016
rect 22100 48068 22152 48074
rect 22100 48010 22152 48016
rect 22020 47802 22048 48010
rect 22008 47796 22060 47802
rect 22008 47738 22060 47744
rect 22100 47456 22152 47462
rect 22100 47398 22152 47404
rect 22112 45898 22140 47398
rect 22100 45892 22152 45898
rect 22100 45834 22152 45840
rect 22100 45620 22152 45626
rect 22100 45562 22152 45568
rect 20180 45526 20300 45554
rect 20076 37460 20128 37466
rect 20076 37402 20128 37408
rect 20076 37324 20128 37330
rect 20076 37266 20128 37272
rect 19708 37188 19760 37194
rect 19708 37130 19760 37136
rect 19800 37188 19852 37194
rect 19800 37130 19852 37136
rect 19984 37120 20036 37126
rect 19984 37062 20036 37068
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 19996 36582 20024 37062
rect 19984 36576 20036 36582
rect 19984 36518 20036 36524
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19708 35760 19760 35766
rect 19708 35702 19760 35708
rect 19616 35624 19668 35630
rect 19616 35566 19668 35572
rect 19524 35488 19576 35494
rect 19524 35430 19576 35436
rect 19536 35018 19564 35430
rect 19628 35222 19656 35566
rect 19720 35494 19748 35702
rect 19708 35488 19760 35494
rect 19708 35430 19760 35436
rect 19616 35216 19668 35222
rect 19616 35158 19668 35164
rect 19720 35057 19748 35430
rect 19706 35048 19762 35057
rect 19524 35012 19576 35018
rect 19706 34983 19762 34992
rect 19524 34954 19576 34960
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 19260 34734 19472 34762
rect 18236 32428 18288 32434
rect 18236 32370 18288 32376
rect 18420 32428 18472 32434
rect 18420 32370 18472 32376
rect 18064 31726 18184 31754
rect 17960 31408 18012 31414
rect 17960 31350 18012 31356
rect 18064 30682 18092 31726
rect 18248 31482 18276 32370
rect 18432 32298 18460 32370
rect 18420 32292 18472 32298
rect 18420 32234 18472 32240
rect 19260 31770 19288 34734
rect 19338 34640 19394 34649
rect 19338 34575 19394 34584
rect 19432 34604 19484 34610
rect 19352 34406 19380 34575
rect 19432 34546 19484 34552
rect 19340 34400 19392 34406
rect 19340 34342 19392 34348
rect 19352 33590 19380 34342
rect 19340 33584 19392 33590
rect 19340 33526 19392 33532
rect 19352 31890 19380 33526
rect 19444 32570 19472 34546
rect 19800 34060 19852 34066
rect 19800 34002 19852 34008
rect 19812 33930 19840 34002
rect 19800 33924 19852 33930
rect 19800 33866 19852 33872
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 19892 33312 19944 33318
rect 19892 33254 19944 33260
rect 19904 32994 19932 33254
rect 19996 33114 20024 36518
rect 20088 35562 20116 37266
rect 20076 35556 20128 35562
rect 20076 35498 20128 35504
rect 20088 35154 20116 35498
rect 20076 35148 20128 35154
rect 20076 35090 20128 35096
rect 20076 34944 20128 34950
rect 20076 34886 20128 34892
rect 19984 33108 20036 33114
rect 19984 33050 20036 33056
rect 19904 32978 20024 32994
rect 19904 32972 20036 32978
rect 19904 32966 19984 32972
rect 19984 32914 20036 32920
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 19432 32564 19484 32570
rect 19432 32506 19484 32512
rect 19996 32230 20024 32914
rect 20088 32910 20116 34886
rect 20076 32904 20128 32910
rect 20076 32846 20128 32852
rect 19432 32224 19484 32230
rect 19432 32166 19484 32172
rect 19984 32224 20036 32230
rect 19984 32166 20036 32172
rect 20076 32224 20128 32230
rect 20076 32166 20128 32172
rect 19340 31884 19392 31890
rect 19340 31826 19392 31832
rect 19260 31742 19380 31770
rect 18512 31680 18564 31686
rect 18512 31622 18564 31628
rect 18236 31476 18288 31482
rect 18236 31418 18288 31424
rect 18524 31346 18552 31622
rect 18512 31340 18564 31346
rect 18512 31282 18564 31288
rect 19156 31272 19208 31278
rect 19156 31214 19208 31220
rect 18420 30864 18472 30870
rect 18420 30806 18472 30812
rect 17972 30654 18092 30682
rect 18144 30660 18196 30666
rect 17868 24812 17920 24818
rect 17868 24754 17920 24760
rect 17868 24268 17920 24274
rect 17868 24210 17920 24216
rect 17880 23526 17908 24210
rect 17868 23520 17920 23526
rect 17868 23462 17920 23468
rect 17972 23202 18000 30654
rect 18144 30602 18196 30608
rect 18156 30122 18184 30602
rect 18432 30258 18460 30806
rect 18420 30252 18472 30258
rect 18420 30194 18472 30200
rect 18144 30116 18196 30122
rect 18144 30058 18196 30064
rect 18328 28484 18380 28490
rect 18328 28426 18380 28432
rect 18340 28218 18368 28426
rect 18328 28212 18380 28218
rect 18328 28154 18380 28160
rect 18236 27872 18288 27878
rect 18236 27814 18288 27820
rect 18248 26994 18276 27814
rect 18236 26988 18288 26994
rect 18236 26930 18288 26936
rect 18248 26382 18276 26930
rect 18340 26382 18368 28154
rect 18432 27470 18460 30194
rect 19168 30122 19196 31214
rect 19352 30734 19380 31742
rect 19444 31482 19472 32166
rect 20088 31754 20116 32166
rect 20076 31748 20128 31754
rect 20076 31690 20128 31696
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 20180 31482 20208 45526
rect 20536 39024 20588 39030
rect 20536 38966 20588 38972
rect 20548 37874 20576 38966
rect 20904 38956 20956 38962
rect 20904 38898 20956 38904
rect 20812 38480 20864 38486
rect 20812 38422 20864 38428
rect 20536 37868 20588 37874
rect 20536 37810 20588 37816
rect 20352 37460 20404 37466
rect 20352 37402 20404 37408
rect 20260 35692 20312 35698
rect 20260 35634 20312 35640
rect 19432 31476 19484 31482
rect 19432 31418 19484 31424
rect 20168 31476 20220 31482
rect 20168 31418 20220 31424
rect 20168 31204 20220 31210
rect 20168 31146 20220 31152
rect 19340 30728 19392 30734
rect 19340 30670 19392 30676
rect 19984 30728 20036 30734
rect 19984 30670 20036 30676
rect 19432 30660 19484 30666
rect 19432 30602 19484 30608
rect 19444 30546 19472 30602
rect 19352 30518 19472 30546
rect 19156 30116 19208 30122
rect 19156 30058 19208 30064
rect 19352 30025 19380 30518
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19708 30252 19760 30258
rect 19708 30194 19760 30200
rect 19338 30016 19394 30025
rect 19338 29951 19394 29960
rect 19352 29170 19380 29951
rect 19720 29850 19748 30194
rect 19432 29844 19484 29850
rect 19432 29786 19484 29792
rect 19708 29844 19760 29850
rect 19708 29786 19760 29792
rect 19340 29164 19392 29170
rect 19340 29106 19392 29112
rect 18696 28416 18748 28422
rect 18696 28358 18748 28364
rect 19340 28416 19392 28422
rect 19340 28358 19392 28364
rect 18512 27600 18564 27606
rect 18512 27542 18564 27548
rect 18524 27470 18552 27542
rect 18708 27470 18736 28358
rect 18420 27464 18472 27470
rect 18420 27406 18472 27412
rect 18512 27464 18564 27470
rect 18512 27406 18564 27412
rect 18696 27464 18748 27470
rect 18696 27406 18748 27412
rect 18524 26382 18552 27406
rect 19248 27328 19300 27334
rect 19248 27270 19300 27276
rect 19260 26586 19288 27270
rect 19352 27062 19380 28358
rect 19444 28064 19472 29786
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19996 28422 20024 30670
rect 19984 28416 20036 28422
rect 19984 28358 20036 28364
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 19521 28076 19573 28082
rect 19444 28036 19521 28064
rect 19521 28018 19573 28024
rect 20076 28076 20128 28082
rect 20076 28018 20128 28024
rect 19800 27940 19852 27946
rect 19800 27882 19852 27888
rect 19616 27872 19668 27878
rect 19616 27814 19668 27820
rect 19432 27464 19484 27470
rect 19432 27406 19484 27412
rect 19340 27056 19392 27062
rect 19340 26998 19392 27004
rect 19444 26586 19472 27406
rect 19628 27316 19656 27814
rect 19812 27674 19840 27882
rect 19984 27872 20036 27878
rect 19984 27814 20036 27820
rect 19800 27668 19852 27674
rect 19800 27610 19852 27616
rect 19505 27288 19656 27316
rect 19505 27112 19533 27288
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 19505 27084 19564 27112
rect 19248 26580 19300 26586
rect 19248 26522 19300 26528
rect 19432 26580 19484 26586
rect 19432 26522 19484 26528
rect 19536 26382 19564 27084
rect 19892 26988 19944 26994
rect 19892 26930 19944 26936
rect 18236 26376 18288 26382
rect 18236 26318 18288 26324
rect 18328 26376 18380 26382
rect 18328 26318 18380 26324
rect 18512 26376 18564 26382
rect 18512 26318 18564 26324
rect 19248 26376 19300 26382
rect 19248 26318 19300 26324
rect 19524 26376 19576 26382
rect 19524 26318 19576 26324
rect 19708 26376 19760 26382
rect 19708 26318 19760 26324
rect 19260 26234 19288 26318
rect 19720 26234 19748 26318
rect 19260 26206 19748 26234
rect 19904 26228 19932 26930
rect 19996 26382 20024 27814
rect 20088 26518 20116 28018
rect 20076 26512 20128 26518
rect 20076 26454 20128 26460
rect 20180 26450 20208 31146
rect 20272 26874 20300 35634
rect 20364 35034 20392 37402
rect 20548 36786 20576 37810
rect 20824 37806 20852 38422
rect 20916 38010 20944 38898
rect 21088 38752 21140 38758
rect 21088 38694 21140 38700
rect 20904 38004 20956 38010
rect 20904 37946 20956 37952
rect 21100 37874 21128 38694
rect 21456 38412 21508 38418
rect 21456 38354 21508 38360
rect 21272 38344 21324 38350
rect 21272 38286 21324 38292
rect 21284 37874 21312 38286
rect 21088 37868 21140 37874
rect 21088 37810 21140 37816
rect 21272 37868 21324 37874
rect 21272 37810 21324 37816
rect 20812 37800 20864 37806
rect 20812 37742 20864 37748
rect 20996 37732 21048 37738
rect 20996 37674 21048 37680
rect 20904 37664 20956 37670
rect 20904 37606 20956 37612
rect 20916 37262 20944 37606
rect 20628 37256 20680 37262
rect 20628 37198 20680 37204
rect 20904 37256 20956 37262
rect 20904 37198 20956 37204
rect 20536 36780 20588 36786
rect 20536 36722 20588 36728
rect 20364 35006 20484 35034
rect 20352 34604 20404 34610
rect 20352 34546 20404 34552
rect 20364 34202 20392 34546
rect 20352 34196 20404 34202
rect 20352 34138 20404 34144
rect 20352 33924 20404 33930
rect 20352 33866 20404 33872
rect 20364 32978 20392 33866
rect 20456 33318 20484 35006
rect 20548 34610 20576 36722
rect 20640 36242 20668 37198
rect 21008 37194 21036 37674
rect 20996 37188 21048 37194
rect 20996 37130 21048 37136
rect 20812 36576 20864 36582
rect 20812 36518 20864 36524
rect 20628 36236 20680 36242
rect 20628 36178 20680 36184
rect 20640 35494 20668 36178
rect 20720 36100 20772 36106
rect 20720 36042 20772 36048
rect 20732 35834 20760 36042
rect 20720 35828 20772 35834
rect 20720 35770 20772 35776
rect 20824 35766 20852 36518
rect 21008 36106 21036 37130
rect 21468 36922 21496 38354
rect 21548 38344 21600 38350
rect 21548 38286 21600 38292
rect 21560 37466 21588 38286
rect 21548 37460 21600 37466
rect 21548 37402 21600 37408
rect 21456 36916 21508 36922
rect 21456 36858 21508 36864
rect 21824 36780 21876 36786
rect 21824 36722 21876 36728
rect 21916 36780 21968 36786
rect 21916 36722 21968 36728
rect 21272 36712 21324 36718
rect 21272 36654 21324 36660
rect 20996 36100 21048 36106
rect 20996 36042 21048 36048
rect 20812 35760 20864 35766
rect 20812 35702 20864 35708
rect 21008 35698 21036 36042
rect 21284 35834 21312 36654
rect 21836 36378 21864 36722
rect 21824 36372 21876 36378
rect 21824 36314 21876 36320
rect 21928 36038 21956 36722
rect 21456 36032 21508 36038
rect 21456 35974 21508 35980
rect 21916 36032 21968 36038
rect 21916 35974 21968 35980
rect 21272 35828 21324 35834
rect 21272 35770 21324 35776
rect 20996 35692 21048 35698
rect 20996 35634 21048 35640
rect 20628 35488 20680 35494
rect 20628 35430 20680 35436
rect 21008 35290 21036 35634
rect 20996 35284 21048 35290
rect 20996 35226 21048 35232
rect 20904 35012 20956 35018
rect 20904 34954 20956 34960
rect 20536 34604 20588 34610
rect 20536 34546 20588 34552
rect 20628 34536 20680 34542
rect 20628 34478 20680 34484
rect 20640 34066 20668 34478
rect 20628 34060 20680 34066
rect 20628 34002 20680 34008
rect 20536 33992 20588 33998
rect 20536 33934 20588 33940
rect 20640 33946 20668 34002
rect 20548 33658 20576 33934
rect 20640 33918 20852 33946
rect 20628 33856 20680 33862
rect 20628 33798 20680 33804
rect 20536 33652 20588 33658
rect 20536 33594 20588 33600
rect 20444 33312 20496 33318
rect 20444 33254 20496 33260
rect 20444 33108 20496 33114
rect 20444 33050 20496 33056
rect 20456 32994 20484 33050
rect 20352 32972 20404 32978
rect 20456 32966 20576 32994
rect 20352 32914 20404 32920
rect 20548 32910 20576 32966
rect 20536 32904 20588 32910
rect 20536 32846 20588 32852
rect 20350 32464 20406 32473
rect 20350 32399 20352 32408
rect 20404 32399 20406 32408
rect 20352 32370 20404 32376
rect 20444 30592 20496 30598
rect 20444 30534 20496 30540
rect 20456 29646 20484 30534
rect 20548 30326 20576 32846
rect 20640 32434 20668 33798
rect 20824 32910 20852 33918
rect 20812 32904 20864 32910
rect 20812 32846 20864 32852
rect 20916 32842 20944 34954
rect 21272 34944 21324 34950
rect 21272 34886 21324 34892
rect 21178 34096 21234 34105
rect 21178 34031 21180 34040
rect 21232 34031 21234 34040
rect 21180 34002 21232 34008
rect 21088 33516 21140 33522
rect 21088 33458 21140 33464
rect 20996 33040 21048 33046
rect 21100 32994 21128 33458
rect 21192 33454 21220 34002
rect 21180 33448 21232 33454
rect 21180 33390 21232 33396
rect 21048 32988 21220 32994
rect 20996 32982 21220 32988
rect 21008 32966 21220 32982
rect 20720 32836 20772 32842
rect 20720 32778 20772 32784
rect 20904 32836 20956 32842
rect 20904 32778 20956 32784
rect 20628 32428 20680 32434
rect 20628 32370 20680 32376
rect 20628 31476 20680 31482
rect 20628 31418 20680 31424
rect 20536 30320 20588 30326
rect 20536 30262 20588 30268
rect 20444 29640 20496 29646
rect 20444 29582 20496 29588
rect 20352 28416 20404 28422
rect 20352 28358 20404 28364
rect 20364 26994 20392 28358
rect 20352 26988 20404 26994
rect 20352 26930 20404 26936
rect 20272 26846 20484 26874
rect 20168 26444 20220 26450
rect 20168 26386 20220 26392
rect 19984 26376 20036 26382
rect 19984 26318 20036 26324
rect 18788 25356 18840 25362
rect 18788 25298 18840 25304
rect 18800 24818 18828 25298
rect 18788 24812 18840 24818
rect 18788 24754 18840 24760
rect 18052 24132 18104 24138
rect 18052 24074 18104 24080
rect 18064 23322 18092 24074
rect 18052 23316 18104 23322
rect 18052 23258 18104 23264
rect 17972 23174 18092 23202
rect 18064 21078 18092 23174
rect 18604 22976 18656 22982
rect 18604 22918 18656 22924
rect 18328 22636 18380 22642
rect 18328 22578 18380 22584
rect 18512 22636 18564 22642
rect 18512 22578 18564 22584
rect 18144 22568 18196 22574
rect 18144 22510 18196 22516
rect 18156 22098 18184 22510
rect 18236 22432 18288 22438
rect 18236 22374 18288 22380
rect 18144 22092 18196 22098
rect 18144 22034 18196 22040
rect 18248 22030 18276 22374
rect 18340 22166 18368 22578
rect 18524 22506 18552 22578
rect 18512 22500 18564 22506
rect 18512 22442 18564 22448
rect 18512 22228 18564 22234
rect 18512 22170 18564 22176
rect 18328 22160 18380 22166
rect 18328 22102 18380 22108
rect 18236 22024 18288 22030
rect 18236 21966 18288 21972
rect 18340 21842 18368 22102
rect 18420 22092 18472 22098
rect 18420 22034 18472 22040
rect 18248 21814 18368 21842
rect 18248 21298 18276 21814
rect 18328 21616 18380 21622
rect 18328 21558 18380 21564
rect 18340 21350 18368 21558
rect 18156 21270 18276 21298
rect 18328 21344 18380 21350
rect 18328 21286 18380 21292
rect 18052 21072 18104 21078
rect 18052 21014 18104 21020
rect 17960 20256 18012 20262
rect 17960 20198 18012 20204
rect 17972 19854 18000 20198
rect 17960 19848 18012 19854
rect 17960 19790 18012 19796
rect 18052 19712 18104 19718
rect 18052 19654 18104 19660
rect 17958 19408 18014 19417
rect 17958 19343 17960 19352
rect 18012 19343 18014 19352
rect 17960 19314 18012 19320
rect 17960 19168 18012 19174
rect 17960 19110 18012 19116
rect 17972 18698 18000 19110
rect 17960 18692 18012 18698
rect 17960 18634 18012 18640
rect 17868 18624 17920 18630
rect 17868 18566 17920 18572
rect 17880 18154 17908 18566
rect 18064 18358 18092 19654
rect 18052 18352 18104 18358
rect 18052 18294 18104 18300
rect 17868 18148 17920 18154
rect 17868 18090 17920 18096
rect 17880 15570 17908 18090
rect 17960 17604 18012 17610
rect 17960 17546 18012 17552
rect 17972 16658 18000 17546
rect 17960 16652 18012 16658
rect 17960 16594 18012 16600
rect 18156 15978 18184 21270
rect 18432 20890 18460 22034
rect 18524 21894 18552 22170
rect 18512 21888 18564 21894
rect 18512 21830 18564 21836
rect 18340 20874 18552 20890
rect 18328 20868 18552 20874
rect 18380 20862 18552 20868
rect 18328 20810 18380 20816
rect 18524 19990 18552 20862
rect 18236 19984 18288 19990
rect 18236 19926 18288 19932
rect 18512 19984 18564 19990
rect 18512 19926 18564 19932
rect 18248 18698 18276 19926
rect 18420 19848 18472 19854
rect 18420 19790 18472 19796
rect 18432 18970 18460 19790
rect 18616 19718 18644 22918
rect 18696 22772 18748 22778
rect 18696 22714 18748 22720
rect 18708 22642 18736 22714
rect 18972 22704 19024 22710
rect 18972 22646 19024 22652
rect 18696 22636 18748 22642
rect 18696 22578 18748 22584
rect 18880 22636 18932 22642
rect 18880 22578 18932 22584
rect 18696 21956 18748 21962
rect 18696 21898 18748 21904
rect 18708 21622 18736 21898
rect 18696 21616 18748 21622
rect 18696 21558 18748 21564
rect 18892 21078 18920 22578
rect 18880 21072 18932 21078
rect 18880 21014 18932 21020
rect 18984 20874 19012 22646
rect 19260 22642 19288 26206
rect 19904 26200 20024 26228
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19800 25288 19852 25294
rect 19798 25256 19800 25265
rect 19852 25256 19854 25265
rect 19340 25220 19392 25226
rect 19798 25191 19854 25200
rect 19340 25162 19392 25168
rect 19352 24342 19380 25162
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19996 24818 20024 26200
rect 20352 25900 20404 25906
rect 20352 25842 20404 25848
rect 20168 25492 20220 25498
rect 20168 25434 20220 25440
rect 20076 25356 20128 25362
rect 20076 25298 20128 25304
rect 20088 24886 20116 25298
rect 20076 24880 20128 24886
rect 20076 24822 20128 24828
rect 19984 24812 20036 24818
rect 19984 24754 20036 24760
rect 19706 24712 19762 24721
rect 19706 24647 19708 24656
rect 19760 24647 19762 24656
rect 19708 24618 19760 24624
rect 19340 24336 19392 24342
rect 19340 24278 19392 24284
rect 19800 24268 19852 24274
rect 19800 24210 19852 24216
rect 19892 24268 19944 24274
rect 19996 24256 20024 24754
rect 19944 24228 20024 24256
rect 19892 24210 19944 24216
rect 19340 24200 19392 24206
rect 19340 24142 19392 24148
rect 19352 23662 19380 24142
rect 19432 24132 19484 24138
rect 19432 24074 19484 24080
rect 19340 23656 19392 23662
rect 19340 23598 19392 23604
rect 19444 23594 19472 24074
rect 19812 24052 19840 24210
rect 20076 24200 20128 24206
rect 20076 24142 20128 24148
rect 19812 24024 20024 24052
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 19892 23724 19944 23730
rect 19892 23666 19944 23672
rect 19708 23656 19760 23662
rect 19904 23633 19932 23666
rect 19708 23598 19760 23604
rect 19890 23624 19946 23633
rect 19432 23588 19484 23594
rect 19432 23530 19484 23536
rect 19340 23180 19392 23186
rect 19444 23168 19472 23530
rect 19720 23322 19748 23598
rect 19890 23559 19946 23568
rect 19892 23520 19944 23526
rect 19890 23488 19892 23497
rect 19944 23488 19946 23497
rect 19890 23423 19946 23432
rect 19708 23316 19760 23322
rect 19708 23258 19760 23264
rect 19904 23254 19932 23423
rect 19892 23248 19944 23254
rect 19892 23190 19944 23196
rect 19444 23140 19564 23168
rect 19340 23122 19392 23128
rect 19248 22636 19300 22642
rect 19248 22578 19300 22584
rect 19352 22438 19380 23122
rect 19432 23044 19484 23050
rect 19432 22986 19484 22992
rect 19444 22574 19472 22986
rect 19536 22964 19564 23140
rect 19505 22936 19564 22964
rect 19505 22760 19533 22936
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19505 22732 19564 22760
rect 19536 22642 19564 22732
rect 19524 22636 19576 22642
rect 19524 22578 19576 22584
rect 19892 22636 19944 22642
rect 19996 22624 20024 24024
rect 20088 23526 20116 24142
rect 20076 23520 20128 23526
rect 20076 23462 20128 23468
rect 20180 23338 20208 25434
rect 20260 25152 20312 25158
rect 20260 25094 20312 25100
rect 20272 24886 20300 25094
rect 20260 24880 20312 24886
rect 20260 24822 20312 24828
rect 20260 24608 20312 24614
rect 20260 24550 20312 24556
rect 20272 24290 20300 24550
rect 20364 24410 20392 25842
rect 20352 24404 20404 24410
rect 20352 24346 20404 24352
rect 20272 24262 20392 24290
rect 20364 23798 20392 24262
rect 20352 23792 20404 23798
rect 20352 23734 20404 23740
rect 20260 23724 20312 23730
rect 20260 23666 20312 23672
rect 20088 23322 20208 23338
rect 20272 23322 20300 23666
rect 20076 23316 20208 23322
rect 20128 23310 20208 23316
rect 20260 23316 20312 23322
rect 20076 23258 20128 23264
rect 20260 23258 20312 23264
rect 19944 22596 20024 22624
rect 19892 22578 19944 22584
rect 19432 22568 19484 22574
rect 19904 22545 19932 22578
rect 19432 22510 19484 22516
rect 19890 22536 19946 22545
rect 19340 22432 19392 22438
rect 19340 22374 19392 22380
rect 19352 21706 19380 22374
rect 19076 21678 19380 21706
rect 18972 20868 19024 20874
rect 18972 20810 19024 20816
rect 18696 20800 18748 20806
rect 18696 20742 18748 20748
rect 18708 20398 18736 20742
rect 18984 20602 19012 20810
rect 18788 20596 18840 20602
rect 18788 20538 18840 20544
rect 18972 20596 19024 20602
rect 18972 20538 19024 20544
rect 18696 20392 18748 20398
rect 18696 20334 18748 20340
rect 18800 19922 18828 20538
rect 18880 20460 18932 20466
rect 18880 20402 18932 20408
rect 18788 19916 18840 19922
rect 18708 19876 18788 19904
rect 18604 19712 18656 19718
rect 18604 19654 18656 19660
rect 18708 19514 18736 19876
rect 18788 19858 18840 19864
rect 18892 19854 18920 20402
rect 18972 20392 19024 20398
rect 18972 20334 19024 20340
rect 18880 19848 18932 19854
rect 18880 19790 18932 19796
rect 18696 19508 18748 19514
rect 18696 19450 18748 19456
rect 18788 19440 18840 19446
rect 18786 19408 18788 19417
rect 18840 19408 18842 19417
rect 18892 19378 18920 19790
rect 18984 19718 19012 20334
rect 18972 19712 19024 19718
rect 18972 19654 19024 19660
rect 18786 19343 18842 19352
rect 18880 19372 18932 19378
rect 18880 19314 18932 19320
rect 18420 18964 18472 18970
rect 18420 18906 18472 18912
rect 18236 18692 18288 18698
rect 18236 18634 18288 18640
rect 18880 18080 18932 18086
rect 18880 18022 18932 18028
rect 18328 17128 18380 17134
rect 18328 17070 18380 17076
rect 18144 15972 18196 15978
rect 18144 15914 18196 15920
rect 17868 15564 17920 15570
rect 17868 15506 17920 15512
rect 18144 15564 18196 15570
rect 18144 15506 18196 15512
rect 18052 14884 18104 14890
rect 18052 14826 18104 14832
rect 17960 14476 18012 14482
rect 17960 14418 18012 14424
rect 17696 12406 17816 12434
rect 17592 11688 17644 11694
rect 17592 11630 17644 11636
rect 17604 10062 17632 11630
rect 17592 10056 17644 10062
rect 17592 9998 17644 10004
rect 17604 9042 17632 9998
rect 17592 9036 17644 9042
rect 17592 8978 17644 8984
rect 17604 8498 17632 8978
rect 17592 8492 17644 8498
rect 17592 8434 17644 8440
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 17420 6582 17540 6610
rect 17408 3936 17460 3942
rect 17408 3878 17460 3884
rect 17420 2922 17448 3878
rect 17316 2916 17368 2922
rect 17316 2858 17368 2864
rect 17408 2916 17460 2922
rect 17408 2858 17460 2864
rect 17512 2854 17540 6582
rect 17696 3534 17724 12406
rect 17972 12238 18000 14418
rect 18064 13870 18092 14826
rect 18052 13864 18104 13870
rect 18052 13806 18104 13812
rect 18156 13802 18184 15506
rect 18236 14952 18288 14958
rect 18236 14894 18288 14900
rect 18144 13796 18196 13802
rect 18144 13738 18196 13744
rect 18144 13524 18196 13530
rect 18144 13466 18196 13472
rect 18052 13184 18104 13190
rect 18052 13126 18104 13132
rect 17960 12232 18012 12238
rect 17960 12174 18012 12180
rect 18064 12170 18092 13126
rect 18156 12918 18184 13466
rect 18144 12912 18196 12918
rect 18144 12854 18196 12860
rect 18052 12164 18104 12170
rect 18052 12106 18104 12112
rect 18156 10146 18184 12854
rect 17972 10118 18184 10146
rect 17972 9602 18000 10118
rect 18248 10010 18276 14894
rect 18156 9982 18276 10010
rect 18156 9654 18184 9982
rect 18236 9920 18288 9926
rect 18236 9862 18288 9868
rect 17880 9586 18000 9602
rect 18144 9648 18196 9654
rect 18144 9590 18196 9596
rect 18248 9586 18276 9862
rect 17868 9580 18000 9586
rect 17920 9574 18000 9580
rect 17868 9522 17920 9528
rect 17972 7410 18000 9574
rect 18052 9580 18104 9586
rect 18052 9522 18104 9528
rect 18236 9580 18288 9586
rect 18236 9522 18288 9528
rect 18064 7886 18092 9522
rect 18248 9110 18276 9522
rect 18236 9104 18288 9110
rect 18236 9046 18288 9052
rect 18340 8106 18368 17070
rect 18892 14482 18920 18022
rect 18880 14476 18932 14482
rect 18880 14418 18932 14424
rect 18604 14340 18656 14346
rect 18604 14282 18656 14288
rect 18420 13864 18472 13870
rect 18420 13806 18472 13812
rect 18156 8078 18368 8106
rect 18052 7880 18104 7886
rect 18052 7822 18104 7828
rect 17960 7404 18012 7410
rect 17960 7346 18012 7352
rect 18156 5370 18184 8078
rect 18432 7970 18460 13806
rect 18512 13320 18564 13326
rect 18512 13262 18564 13268
rect 18524 12442 18552 13262
rect 18616 12986 18644 14282
rect 18604 12980 18656 12986
rect 18604 12922 18656 12928
rect 18512 12436 18564 12442
rect 18512 12378 18564 12384
rect 18512 10464 18564 10470
rect 18512 10406 18564 10412
rect 18524 9994 18552 10406
rect 18512 9988 18564 9994
rect 18512 9930 18564 9936
rect 18616 8004 18644 12922
rect 18984 12782 19012 19654
rect 19076 17338 19104 21678
rect 19340 21616 19392 21622
rect 19340 21558 19392 21564
rect 19352 21146 19380 21558
rect 19340 21140 19392 21146
rect 19340 21082 19392 21088
rect 19340 19916 19392 19922
rect 19340 19858 19392 19864
rect 19156 19848 19208 19854
rect 19156 19790 19208 19796
rect 19064 17332 19116 17338
rect 19064 17274 19116 17280
rect 19168 16810 19196 19790
rect 19352 18766 19380 19858
rect 19340 18760 19392 18766
rect 19340 18702 19392 18708
rect 19352 16998 19380 18702
rect 19340 16992 19392 16998
rect 19340 16934 19392 16940
rect 19168 16782 19380 16810
rect 19248 16584 19300 16590
rect 19248 16526 19300 16532
rect 19064 16516 19116 16522
rect 19064 16458 19116 16464
rect 18972 12776 19024 12782
rect 18972 12718 19024 12724
rect 18788 11008 18840 11014
rect 18788 10950 18840 10956
rect 18800 10674 18828 10950
rect 18788 10668 18840 10674
rect 18788 10610 18840 10616
rect 18972 10668 19024 10674
rect 18972 10610 19024 10616
rect 18984 9722 19012 10610
rect 18972 9716 19024 9722
rect 18972 9658 19024 9664
rect 18972 8288 19024 8294
rect 18972 8230 19024 8236
rect 18248 7942 18460 7970
rect 18524 7976 18644 8004
rect 18788 8016 18840 8022
rect 18144 5364 18196 5370
rect 18144 5306 18196 5312
rect 17684 3528 17736 3534
rect 17684 3470 17736 3476
rect 17776 3528 17828 3534
rect 17776 3470 17828 3476
rect 17788 3058 17816 3470
rect 18248 3398 18276 7942
rect 18420 7404 18472 7410
rect 18420 7346 18472 7352
rect 18432 6798 18460 7346
rect 18420 6792 18472 6798
rect 18420 6734 18472 6740
rect 18524 3670 18552 7976
rect 18788 7958 18840 7964
rect 18604 7812 18656 7818
rect 18604 7754 18656 7760
rect 18616 7546 18644 7754
rect 18696 7744 18748 7750
rect 18696 7686 18748 7692
rect 18604 7540 18656 7546
rect 18604 7482 18656 7488
rect 18708 7478 18736 7686
rect 18696 7472 18748 7478
rect 18696 7414 18748 7420
rect 18512 3664 18564 3670
rect 18512 3606 18564 3612
rect 17960 3392 18012 3398
rect 17960 3334 18012 3340
rect 18236 3392 18288 3398
rect 18236 3334 18288 3340
rect 17972 3126 18000 3334
rect 17960 3120 18012 3126
rect 17960 3062 18012 3068
rect 17776 3052 17828 3058
rect 17776 2994 17828 3000
rect 18052 2984 18104 2990
rect 18052 2926 18104 2932
rect 17500 2848 17552 2854
rect 17500 2790 17552 2796
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 17776 2440 17828 2446
rect 17776 2382 17828 2388
rect 17420 800 17448 2382
rect 17788 1834 17816 2382
rect 17776 1828 17828 1834
rect 17776 1770 17828 1776
rect 18064 800 18092 2926
rect 18800 2774 18828 7958
rect 18984 7954 19012 8230
rect 18972 7948 19024 7954
rect 18972 7890 19024 7896
rect 19076 7274 19104 16458
rect 19260 16114 19288 16526
rect 19248 16108 19300 16114
rect 19248 16050 19300 16056
rect 19260 15502 19288 16050
rect 19248 15496 19300 15502
rect 19248 15438 19300 15444
rect 19352 13394 19380 16782
rect 19444 14521 19472 22510
rect 19890 22471 19946 22480
rect 20088 22438 20116 23258
rect 20168 23112 20220 23118
rect 20168 23054 20220 23060
rect 20076 22432 20128 22438
rect 20076 22374 20128 22380
rect 20074 21992 20130 22001
rect 20074 21927 20130 21936
rect 19984 21888 20036 21894
rect 19984 21830 20036 21836
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19996 21010 20024 21830
rect 19984 21004 20036 21010
rect 19984 20946 20036 20952
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19890 19408 19946 19417
rect 19890 19343 19946 19352
rect 19984 19372 20036 19378
rect 19616 19168 19668 19174
rect 19616 19110 19668 19116
rect 19628 18766 19656 19110
rect 19616 18760 19668 18766
rect 19616 18702 19668 18708
rect 19904 18698 19932 19343
rect 19984 19314 20036 19320
rect 19892 18692 19944 18698
rect 19892 18634 19944 18640
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19996 18426 20024 19314
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19984 17264 20036 17270
rect 19984 17206 20036 17212
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19892 16040 19944 16046
rect 19890 16008 19892 16017
rect 19944 16008 19946 16017
rect 19890 15943 19946 15952
rect 19904 15706 19932 15943
rect 19892 15700 19944 15706
rect 19892 15642 19944 15648
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19430 14512 19486 14521
rect 19430 14447 19486 14456
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19156 13388 19208 13394
rect 19156 13330 19208 13336
rect 19340 13388 19392 13394
rect 19340 13330 19392 13336
rect 19168 12850 19196 13330
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19340 13252 19392 13258
rect 19340 13194 19392 13200
rect 19156 12844 19208 12850
rect 19156 12786 19208 12792
rect 19352 12594 19380 13194
rect 19444 12646 19472 13262
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 19260 12566 19380 12594
rect 19432 12640 19484 12646
rect 19432 12582 19484 12588
rect 19708 12640 19760 12646
rect 19708 12582 19760 12588
rect 19260 12374 19288 12566
rect 19248 12368 19300 12374
rect 19248 12310 19300 12316
rect 19156 12232 19208 12238
rect 19156 12174 19208 12180
rect 19168 11898 19196 12174
rect 19720 12170 19748 12582
rect 19708 12164 19760 12170
rect 19708 12106 19760 12112
rect 19340 12096 19392 12102
rect 19340 12038 19392 12044
rect 19156 11892 19208 11898
rect 19156 11834 19208 11840
rect 19168 11150 19196 11834
rect 19156 11144 19208 11150
rect 19156 11086 19208 11092
rect 19352 11082 19380 12038
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19432 11756 19484 11762
rect 19432 11698 19484 11704
rect 19340 11076 19392 11082
rect 19340 11018 19392 11024
rect 19352 10062 19380 11018
rect 19444 10674 19472 11698
rect 19996 11098 20024 17206
rect 20088 15094 20116 21927
rect 20076 15088 20128 15094
rect 20076 15030 20128 15036
rect 20076 14816 20128 14822
rect 20074 14784 20076 14793
rect 20128 14784 20130 14793
rect 20074 14719 20130 14728
rect 20076 14340 20128 14346
rect 20076 14282 20128 14288
rect 20088 14074 20116 14282
rect 20076 14068 20128 14074
rect 20076 14010 20128 14016
rect 20076 11756 20128 11762
rect 20076 11698 20128 11704
rect 20088 11354 20116 11698
rect 20076 11348 20128 11354
rect 20076 11290 20128 11296
rect 19996 11070 20116 11098
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19432 10668 19484 10674
rect 19432 10610 19484 10616
rect 19444 10130 19472 10610
rect 19524 10600 19576 10606
rect 19524 10542 19576 10548
rect 19432 10124 19484 10130
rect 19432 10066 19484 10072
rect 19340 10056 19392 10062
rect 19536 10033 19564 10542
rect 19708 10056 19760 10062
rect 19340 9998 19392 10004
rect 19522 10024 19578 10033
rect 19352 9586 19380 9998
rect 19432 9988 19484 9994
rect 19522 9959 19578 9968
rect 19706 10024 19708 10033
rect 19760 10024 19762 10033
rect 19706 9959 19762 9968
rect 19432 9930 19484 9936
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 19444 9466 19472 9930
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19616 9686 19668 9692
rect 19616 9628 19668 9634
rect 19798 9688 19854 9697
rect 19982 9688 20038 9697
rect 19854 9646 19932 9674
rect 19352 9438 19472 9466
rect 19352 8838 19380 9438
rect 19524 9376 19576 9382
rect 19524 9318 19576 9324
rect 19536 8974 19564 9318
rect 19524 8968 19576 8974
rect 19524 8910 19576 8916
rect 19340 8832 19392 8838
rect 19628 8820 19656 9628
rect 19798 9623 19854 9632
rect 19904 9432 19932 9646
rect 19982 9623 20038 9632
rect 19996 9586 20024 9623
rect 19984 9580 20036 9586
rect 19984 9522 20036 9528
rect 19984 9444 20036 9450
rect 19904 9404 19984 9432
rect 19984 9386 20036 9392
rect 19340 8774 19392 8780
rect 19444 8792 19656 8820
rect 19248 8492 19300 8498
rect 19248 8434 19300 8440
rect 19260 7546 19288 8434
rect 19352 8430 19380 8774
rect 19340 8424 19392 8430
rect 19340 8366 19392 8372
rect 19340 8288 19392 8294
rect 19340 8230 19392 8236
rect 19248 7540 19300 7546
rect 19248 7482 19300 7488
rect 19064 7268 19116 7274
rect 19064 7210 19116 7216
rect 19352 7002 19380 8230
rect 19340 6996 19392 7002
rect 19340 6938 19392 6944
rect 19444 6746 19472 8792
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19996 7546 20024 9386
rect 19984 7540 20036 7546
rect 19984 7482 20036 7488
rect 19616 7404 19668 7410
rect 19616 7346 19668 7352
rect 19628 6798 19656 7346
rect 19982 7304 20038 7313
rect 19982 7239 20038 7248
rect 19352 6718 19472 6746
rect 19616 6792 19668 6798
rect 19616 6734 19668 6740
rect 19352 5658 19380 6718
rect 19432 6656 19484 6662
rect 19432 6598 19484 6604
rect 19260 5630 19380 5658
rect 19260 5302 19288 5630
rect 19248 5296 19300 5302
rect 19248 5238 19300 5244
rect 19340 5228 19392 5234
rect 19340 5170 19392 5176
rect 18708 2746 18828 2774
rect 18708 800 18736 2746
rect 19352 2582 19380 5170
rect 19340 2576 19392 2582
rect 19340 2518 19392 2524
rect 19444 2514 19472 6598
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 19996 3194 20024 7239
rect 19984 3188 20036 3194
rect 19984 3130 20036 3136
rect 19432 2508 19484 2514
rect 19432 2450 19484 2456
rect 19984 2440 20036 2446
rect 19984 2382 20036 2388
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 19996 800 20024 2382
rect 20088 2310 20116 11070
rect 20180 6662 20208 23054
rect 20272 17270 20300 23258
rect 20364 17678 20392 23734
rect 20352 17672 20404 17678
rect 20352 17614 20404 17620
rect 20352 17536 20404 17542
rect 20352 17478 20404 17484
rect 20260 17264 20312 17270
rect 20260 17206 20312 17212
rect 20364 16998 20392 17478
rect 20260 16992 20312 16998
rect 20260 16934 20312 16940
rect 20352 16992 20404 16998
rect 20352 16934 20404 16940
rect 20272 16658 20300 16934
rect 20260 16652 20312 16658
rect 20260 16594 20312 16600
rect 20272 15706 20300 16594
rect 20260 15700 20312 15706
rect 20260 15642 20312 15648
rect 20260 15360 20312 15366
rect 20260 15302 20312 15308
rect 20352 15360 20404 15366
rect 20352 15302 20404 15308
rect 20272 13938 20300 15302
rect 20364 14550 20392 15302
rect 20352 14544 20404 14550
rect 20352 14486 20404 14492
rect 20260 13932 20312 13938
rect 20260 13874 20312 13880
rect 20260 12776 20312 12782
rect 20260 12718 20312 12724
rect 20272 11676 20300 12718
rect 20352 12368 20404 12374
rect 20352 12310 20404 12316
rect 20364 12170 20392 12310
rect 20352 12164 20404 12170
rect 20352 12106 20404 12112
rect 20364 11830 20392 12106
rect 20352 11824 20404 11830
rect 20352 11766 20404 11772
rect 20352 11688 20404 11694
rect 20272 11648 20352 11676
rect 20272 10606 20300 11648
rect 20352 11630 20404 11636
rect 20350 11520 20406 11529
rect 20350 11455 20406 11464
rect 20260 10600 20312 10606
rect 20260 10542 20312 10548
rect 20260 10124 20312 10130
rect 20260 10066 20312 10072
rect 20272 9586 20300 10066
rect 20260 9580 20312 9586
rect 20260 9522 20312 9528
rect 20258 9480 20314 9489
rect 20258 9415 20314 9424
rect 20168 6656 20220 6662
rect 20168 6598 20220 6604
rect 20168 3936 20220 3942
rect 20168 3878 20220 3884
rect 20180 3602 20208 3878
rect 20168 3596 20220 3602
rect 20168 3538 20220 3544
rect 20272 3126 20300 9415
rect 20364 7562 20392 11455
rect 20456 7721 20484 26846
rect 20536 25900 20588 25906
rect 20536 25842 20588 25848
rect 20548 24954 20576 25842
rect 20640 25362 20668 31418
rect 20732 31278 20760 32778
rect 20812 32768 20864 32774
rect 20812 32710 20864 32716
rect 20824 32434 20852 32710
rect 20812 32428 20864 32434
rect 20812 32370 20864 32376
rect 21192 31958 21220 32966
rect 21180 31952 21232 31958
rect 21180 31894 21232 31900
rect 20812 31884 20864 31890
rect 20812 31826 20864 31832
rect 20720 31272 20772 31278
rect 20720 31214 20772 31220
rect 20720 31136 20772 31142
rect 20720 31078 20772 31084
rect 20732 25498 20760 31078
rect 20824 30326 20852 31826
rect 21088 31136 21140 31142
rect 21088 31078 21140 31084
rect 20996 30932 21048 30938
rect 21100 30920 21128 31078
rect 21048 30892 21128 30920
rect 20996 30874 21048 30880
rect 21100 30734 21128 30892
rect 21088 30728 21140 30734
rect 21088 30670 21140 30676
rect 21192 30326 21220 31894
rect 20812 30320 20864 30326
rect 20812 30262 20864 30268
rect 21180 30320 21232 30326
rect 21180 30262 21232 30268
rect 20904 30252 20956 30258
rect 20904 30194 20956 30200
rect 20916 29510 20944 30194
rect 20904 29504 20956 29510
rect 20904 29446 20956 29452
rect 21180 28484 21232 28490
rect 21180 28426 21232 28432
rect 20812 28212 20864 28218
rect 20812 28154 20864 28160
rect 20824 27606 20852 28154
rect 21088 28076 21140 28082
rect 21088 28018 21140 28024
rect 21100 27946 21128 28018
rect 21088 27940 21140 27946
rect 21088 27882 21140 27888
rect 20812 27600 20864 27606
rect 20812 27542 20864 27548
rect 21100 27062 21128 27882
rect 21192 27470 21220 28426
rect 21284 28014 21312 34886
rect 21364 33312 21416 33318
rect 21364 33254 21416 33260
rect 21272 28008 21324 28014
rect 21272 27950 21324 27956
rect 21180 27464 21232 27470
rect 21180 27406 21232 27412
rect 21272 27396 21324 27402
rect 21272 27338 21324 27344
rect 21284 27062 21312 27338
rect 21088 27056 21140 27062
rect 21088 26998 21140 27004
rect 21272 27056 21324 27062
rect 21272 26998 21324 27004
rect 21088 25764 21140 25770
rect 21088 25706 21140 25712
rect 20824 25622 21036 25650
rect 20720 25492 20772 25498
rect 20720 25434 20772 25440
rect 20824 25362 20852 25622
rect 20904 25492 20956 25498
rect 20904 25434 20956 25440
rect 20628 25356 20680 25362
rect 20628 25298 20680 25304
rect 20812 25356 20864 25362
rect 20812 25298 20864 25304
rect 20732 25226 20852 25242
rect 20720 25220 20852 25226
rect 20772 25214 20852 25220
rect 20720 25162 20772 25168
rect 20824 24970 20852 25214
rect 20732 24954 20852 24970
rect 20536 24948 20588 24954
rect 20536 24890 20588 24896
rect 20720 24948 20852 24954
rect 20772 24942 20852 24948
rect 20720 24890 20772 24896
rect 20812 24880 20864 24886
rect 20812 24822 20864 24828
rect 20628 24812 20680 24818
rect 20628 24754 20680 24760
rect 20720 24812 20772 24818
rect 20720 24754 20772 24760
rect 20640 24290 20668 24754
rect 20732 24721 20760 24754
rect 20718 24712 20774 24721
rect 20718 24647 20774 24656
rect 20548 24262 20668 24290
rect 20720 24336 20772 24342
rect 20720 24278 20772 24284
rect 20548 22778 20576 24262
rect 20628 24132 20680 24138
rect 20628 24074 20680 24080
rect 20640 23322 20668 24074
rect 20732 23730 20760 24278
rect 20824 24274 20852 24822
rect 20812 24268 20864 24274
rect 20812 24210 20864 24216
rect 20916 24206 20944 25434
rect 21008 24410 21036 25622
rect 21100 25430 21128 25706
rect 21088 25424 21140 25430
rect 21088 25366 21140 25372
rect 21088 24744 21140 24750
rect 21088 24686 21140 24692
rect 20996 24404 21048 24410
rect 20996 24346 21048 24352
rect 20904 24200 20956 24206
rect 20904 24142 20956 24148
rect 20902 23896 20958 23905
rect 21100 23866 21128 24686
rect 21376 24410 21404 33254
rect 21468 32230 21496 35974
rect 21640 33516 21692 33522
rect 21640 33458 21692 33464
rect 21548 32496 21600 32502
rect 21548 32438 21600 32444
rect 21456 32224 21508 32230
rect 21456 32166 21508 32172
rect 21468 30802 21496 32166
rect 21456 30796 21508 30802
rect 21456 30738 21508 30744
rect 21560 30122 21588 32438
rect 21652 32434 21680 33458
rect 21916 33448 21968 33454
rect 21916 33390 21968 33396
rect 21640 32428 21692 32434
rect 21640 32370 21692 32376
rect 21824 31816 21876 31822
rect 21824 31758 21876 31764
rect 21732 31680 21784 31686
rect 21732 31622 21784 31628
rect 21640 30932 21692 30938
rect 21640 30874 21692 30880
rect 21548 30116 21600 30122
rect 21548 30058 21600 30064
rect 21652 28994 21680 30874
rect 21744 30870 21772 31622
rect 21732 30864 21784 30870
rect 21732 30806 21784 30812
rect 21732 30728 21784 30734
rect 21732 30670 21784 30676
rect 21744 30190 21772 30670
rect 21732 30184 21784 30190
rect 21732 30126 21784 30132
rect 21836 29714 21864 31758
rect 21928 31414 21956 33390
rect 22008 32972 22060 32978
rect 22008 32914 22060 32920
rect 22020 32434 22048 32914
rect 22008 32428 22060 32434
rect 22008 32370 22060 32376
rect 21916 31408 21968 31414
rect 21916 31350 21968 31356
rect 22020 30870 22048 32370
rect 22008 30864 22060 30870
rect 22008 30806 22060 30812
rect 21916 30660 21968 30666
rect 21916 30602 21968 30608
rect 21928 30258 21956 30602
rect 21916 30252 21968 30258
rect 21916 30194 21968 30200
rect 22008 30116 22060 30122
rect 22008 30058 22060 30064
rect 21824 29708 21876 29714
rect 21824 29650 21876 29656
rect 21732 29504 21784 29510
rect 21732 29446 21784 29452
rect 21560 28966 21680 28994
rect 21456 28076 21508 28082
rect 21456 28018 21508 28024
rect 21468 27470 21496 28018
rect 21456 27464 21508 27470
rect 21456 27406 21508 27412
rect 21456 24608 21508 24614
rect 21456 24550 21508 24556
rect 21180 24404 21232 24410
rect 21180 24346 21232 24352
rect 21364 24404 21416 24410
rect 21364 24346 21416 24352
rect 20902 23831 20904 23840
rect 20956 23831 20958 23840
rect 21088 23860 21140 23866
rect 20904 23802 20956 23808
rect 21088 23802 21140 23808
rect 20720 23724 20772 23730
rect 20720 23666 20772 23672
rect 20996 23724 21048 23730
rect 20996 23666 21048 23672
rect 20628 23316 20680 23322
rect 20628 23258 20680 23264
rect 20628 23180 20680 23186
rect 20628 23122 20680 23128
rect 20536 22772 20588 22778
rect 20536 22714 20588 22720
rect 20536 22432 20588 22438
rect 20536 22374 20588 22380
rect 20548 22103 20576 22374
rect 20534 22094 20590 22103
rect 20534 22029 20590 22038
rect 20536 21956 20588 21962
rect 20536 21898 20588 21904
rect 20548 21418 20576 21898
rect 20536 21412 20588 21418
rect 20536 21354 20588 21360
rect 20536 20936 20588 20942
rect 20536 20878 20588 20884
rect 20548 20330 20576 20878
rect 20536 20324 20588 20330
rect 20536 20266 20588 20272
rect 20640 19334 20668 23122
rect 21008 23118 21036 23666
rect 20996 23112 21048 23118
rect 20996 23054 21048 23060
rect 20720 21956 20772 21962
rect 20720 21898 20772 21904
rect 20732 19854 20760 21898
rect 20720 19848 20772 19854
rect 20720 19790 20772 19796
rect 20548 19306 20668 19334
rect 20548 13734 20576 19306
rect 21088 18692 21140 18698
rect 21088 18634 21140 18640
rect 20628 18624 20680 18630
rect 20628 18566 20680 18572
rect 20640 18290 20668 18566
rect 20628 18284 20680 18290
rect 20628 18226 20680 18232
rect 20996 18216 21048 18222
rect 20996 18158 21048 18164
rect 20812 17808 20864 17814
rect 20812 17750 20864 17756
rect 20628 17604 20680 17610
rect 20628 17546 20680 17552
rect 20640 17320 20668 17546
rect 20640 17292 20760 17320
rect 20628 17196 20680 17202
rect 20628 17138 20680 17144
rect 20640 16250 20668 17138
rect 20628 16244 20680 16250
rect 20628 16186 20680 16192
rect 20732 15994 20760 17292
rect 20824 16114 20852 17750
rect 21008 17746 21036 18158
rect 20996 17740 21048 17746
rect 20996 17682 21048 17688
rect 20904 16992 20956 16998
rect 20904 16934 20956 16940
rect 20916 16794 20944 16934
rect 20904 16788 20956 16794
rect 20904 16730 20956 16736
rect 20812 16108 20864 16114
rect 20812 16050 20864 16056
rect 20732 15966 20852 15994
rect 20628 15088 20680 15094
rect 20628 15030 20680 15036
rect 20536 13728 20588 13734
rect 20536 13670 20588 13676
rect 20640 12714 20668 15030
rect 20628 12708 20680 12714
rect 20628 12650 20680 12656
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20732 12442 20760 12582
rect 20720 12436 20772 12442
rect 20720 12378 20772 12384
rect 20824 12186 20852 15966
rect 21008 15570 21036 17682
rect 20996 15564 21048 15570
rect 20996 15506 21048 15512
rect 20904 12708 20956 12714
rect 20904 12650 20956 12656
rect 20548 12158 20852 12186
rect 20548 7750 20576 12158
rect 20916 12084 20944 12650
rect 20640 12056 20944 12084
rect 20640 9450 20668 12056
rect 21100 11914 21128 18634
rect 21192 16028 21220 24346
rect 21468 23594 21496 24550
rect 21456 23588 21508 23594
rect 21456 23530 21508 23536
rect 21192 16000 21312 16028
rect 21180 15020 21232 15026
rect 21180 14962 21232 14968
rect 21192 14074 21220 14962
rect 21180 14068 21232 14074
rect 21180 14010 21232 14016
rect 21180 13728 21232 13734
rect 21180 13670 21232 13676
rect 20916 11886 21128 11914
rect 20916 9674 20944 11886
rect 21192 9722 21220 13670
rect 20732 9646 20944 9674
rect 21180 9716 21232 9722
rect 21180 9658 21232 9664
rect 20996 9648 21048 9654
rect 20628 9444 20680 9450
rect 20628 9386 20680 9392
rect 20732 9330 20760 9646
rect 20996 9590 21048 9596
rect 20640 9302 20760 9330
rect 20536 7744 20588 7750
rect 20442 7712 20498 7721
rect 20536 7686 20588 7692
rect 20442 7647 20498 7656
rect 20364 7534 20576 7562
rect 20442 7304 20498 7313
rect 20352 7268 20404 7274
rect 20442 7239 20498 7248
rect 20352 7210 20404 7216
rect 20364 4010 20392 7210
rect 20352 4004 20404 4010
rect 20352 3946 20404 3952
rect 20352 3596 20404 3602
rect 20352 3538 20404 3544
rect 20364 3194 20392 3538
rect 20352 3188 20404 3194
rect 20352 3130 20404 3136
rect 20260 3120 20312 3126
rect 20260 3062 20312 3068
rect 20456 2650 20484 7239
rect 20444 2644 20496 2650
rect 20444 2586 20496 2592
rect 20548 2514 20576 7534
rect 20640 3754 20668 9302
rect 20904 6724 20956 6730
rect 20904 6666 20956 6672
rect 20916 6458 20944 6666
rect 20904 6452 20956 6458
rect 20904 6394 20956 6400
rect 21008 6390 21036 9590
rect 21284 8514 21312 16000
rect 21456 15428 21508 15434
rect 21456 15370 21508 15376
rect 21468 15094 21496 15370
rect 21456 15088 21508 15094
rect 21456 15030 21508 15036
rect 21454 14920 21510 14929
rect 21454 14855 21456 14864
rect 21508 14855 21510 14864
rect 21456 14826 21508 14832
rect 21364 14612 21416 14618
rect 21364 14554 21416 14560
rect 21376 14346 21404 14554
rect 21456 14544 21508 14550
rect 21456 14486 21508 14492
rect 21364 14340 21416 14346
rect 21364 14282 21416 14288
rect 21376 13734 21404 14282
rect 21468 13870 21496 14486
rect 21456 13864 21508 13870
rect 21456 13806 21508 13812
rect 21364 13728 21416 13734
rect 21364 13670 21416 13676
rect 21560 12434 21588 28966
rect 21744 27606 21772 29446
rect 22020 28558 22048 30058
rect 22008 28552 22060 28558
rect 22008 28494 22060 28500
rect 21732 27600 21784 27606
rect 21732 27542 21784 27548
rect 21916 27328 21968 27334
rect 21916 27270 21968 27276
rect 21928 26994 21956 27270
rect 21916 26988 21968 26994
rect 21916 26930 21968 26936
rect 21916 26308 21968 26314
rect 21916 26250 21968 26256
rect 21824 24812 21876 24818
rect 21824 24754 21876 24760
rect 21836 24206 21864 24754
rect 21928 24274 21956 26250
rect 21916 24268 21968 24274
rect 21916 24210 21968 24216
rect 21824 24200 21876 24206
rect 21824 24142 21876 24148
rect 21928 23730 21956 24210
rect 21916 23724 21968 23730
rect 21744 23684 21916 23712
rect 21638 21856 21694 21865
rect 21638 21791 21694 21800
rect 21652 21554 21680 21791
rect 21744 21554 21772 23684
rect 21916 23666 21968 23672
rect 22112 22098 22140 45562
rect 22192 34468 22244 34474
rect 22192 34410 22244 34416
rect 22204 33504 22232 34410
rect 22296 33862 22324 49166
rect 22572 48210 22600 51200
rect 23400 48770 23428 51326
rect 23846 51326 24256 51354
rect 23846 51200 23902 51326
rect 24228 49298 24256 51326
rect 24490 51326 24624 51354
rect 24490 51200 24546 51326
rect 24216 49292 24268 49298
rect 24216 49234 24268 49240
rect 23848 49224 23900 49230
rect 23848 49166 23900 49172
rect 23400 48742 23520 48770
rect 23492 48686 23520 48742
rect 22744 48680 22796 48686
rect 22744 48622 22796 48628
rect 23480 48680 23532 48686
rect 23480 48622 23532 48628
rect 22560 48204 22612 48210
rect 22560 48146 22612 48152
rect 22756 47802 22784 48622
rect 23860 48210 23888 49166
rect 24492 49156 24544 49162
rect 24492 49098 24544 49104
rect 23848 48204 23900 48210
rect 23848 48146 23900 48152
rect 24308 48136 24360 48142
rect 24308 48078 24360 48084
rect 24216 48068 24268 48074
rect 24216 48010 24268 48016
rect 24228 47802 24256 48010
rect 24320 47802 24348 48078
rect 22744 47796 22796 47802
rect 22744 47738 22796 47744
rect 24216 47796 24268 47802
rect 24216 47738 24268 47744
rect 24308 47796 24360 47802
rect 24308 47738 24360 47744
rect 22836 47660 22888 47666
rect 22836 47602 22888 47608
rect 23664 47660 23716 47666
rect 23664 47602 23716 47608
rect 22848 46646 22876 47602
rect 23112 47592 23164 47598
rect 23112 47534 23164 47540
rect 22836 46640 22888 46646
rect 22836 46582 22888 46588
rect 22848 45626 22876 46582
rect 22836 45620 22888 45626
rect 22836 45562 22888 45568
rect 22744 38208 22796 38214
rect 22744 38150 22796 38156
rect 22376 37868 22428 37874
rect 22376 37810 22428 37816
rect 22388 37126 22416 37810
rect 22468 37800 22520 37806
rect 22468 37742 22520 37748
rect 22376 37120 22428 37126
rect 22376 37062 22428 37068
rect 22480 36242 22508 37742
rect 22468 36236 22520 36242
rect 22468 36178 22520 36184
rect 22652 36236 22704 36242
rect 22652 36178 22704 36184
rect 22468 36032 22520 36038
rect 22468 35974 22520 35980
rect 22480 35698 22508 35974
rect 22468 35692 22520 35698
rect 22468 35634 22520 35640
rect 22664 35630 22692 36178
rect 22756 36038 22784 38150
rect 22744 36032 22796 36038
rect 22744 35974 22796 35980
rect 22652 35624 22704 35630
rect 22652 35566 22704 35572
rect 22652 35012 22704 35018
rect 22652 34954 22704 34960
rect 22468 34604 22520 34610
rect 22468 34546 22520 34552
rect 22480 34202 22508 34546
rect 22468 34196 22520 34202
rect 22468 34138 22520 34144
rect 22284 33856 22336 33862
rect 22284 33798 22336 33804
rect 22376 33856 22428 33862
rect 22376 33798 22428 33804
rect 22560 33856 22612 33862
rect 22560 33798 22612 33804
rect 22284 33516 22336 33522
rect 22204 33476 22284 33504
rect 22284 33458 22336 33464
rect 22388 33454 22416 33798
rect 22572 33590 22600 33798
rect 22560 33584 22612 33590
rect 22560 33526 22612 33532
rect 22376 33448 22428 33454
rect 22376 33390 22428 33396
rect 22560 33448 22612 33454
rect 22560 33390 22612 33396
rect 22192 32360 22244 32366
rect 22192 32302 22244 32308
rect 22204 32026 22232 32302
rect 22388 32298 22416 33390
rect 22572 32502 22600 33390
rect 22560 32496 22612 32502
rect 22560 32438 22612 32444
rect 22376 32292 22428 32298
rect 22376 32234 22428 32240
rect 22192 32020 22244 32026
rect 22192 31962 22244 31968
rect 22388 31958 22416 32234
rect 22572 32230 22600 32438
rect 22560 32224 22612 32230
rect 22560 32166 22612 32172
rect 22376 31952 22428 31958
rect 22376 31894 22428 31900
rect 22284 31816 22336 31822
rect 22282 31784 22284 31793
rect 22664 31793 22692 34954
rect 22336 31784 22338 31793
rect 22282 31719 22338 31728
rect 22650 31784 22706 31793
rect 22650 31719 22706 31728
rect 22756 31754 22784 35974
rect 22836 35692 22888 35698
rect 22836 35634 22888 35640
rect 22848 32230 22876 35634
rect 22928 33516 22980 33522
rect 22928 33458 22980 33464
rect 22940 33114 22968 33458
rect 22928 33108 22980 33114
rect 22928 33050 22980 33056
rect 22926 32600 22982 32609
rect 22926 32535 22982 32544
rect 22940 32502 22968 32535
rect 22928 32496 22980 32502
rect 22928 32438 22980 32444
rect 22836 32224 22888 32230
rect 22836 32166 22888 32172
rect 23020 32020 23072 32026
rect 23020 31962 23072 31968
rect 23032 31754 23060 31962
rect 22756 31726 22876 31754
rect 22192 31680 22244 31686
rect 22192 31622 22244 31628
rect 22204 29238 22232 31622
rect 22376 31408 22428 31414
rect 22376 31350 22428 31356
rect 22284 30592 22336 30598
rect 22284 30534 22336 30540
rect 22296 30326 22324 30534
rect 22284 30320 22336 30326
rect 22284 30262 22336 30268
rect 22284 29572 22336 29578
rect 22284 29514 22336 29520
rect 22296 29306 22324 29514
rect 22284 29300 22336 29306
rect 22284 29242 22336 29248
rect 22192 29232 22244 29238
rect 22192 29174 22244 29180
rect 22284 28416 22336 28422
rect 22284 28358 22336 28364
rect 22296 26450 22324 28358
rect 22284 26444 22336 26450
rect 22284 26386 22336 26392
rect 21824 22092 21876 22098
rect 21824 22034 21876 22040
rect 22100 22092 22152 22098
rect 22388 22094 22416 31350
rect 22560 31136 22612 31142
rect 22560 31078 22612 31084
rect 22468 30592 22520 30598
rect 22468 30534 22520 30540
rect 22480 29170 22508 30534
rect 22572 29238 22600 31078
rect 22744 30796 22796 30802
rect 22744 30738 22796 30744
rect 22652 30592 22704 30598
rect 22652 30534 22704 30540
rect 22664 30054 22692 30534
rect 22756 30054 22784 30738
rect 22652 30048 22704 30054
rect 22652 29990 22704 29996
rect 22744 30048 22796 30054
rect 22744 29990 22796 29996
rect 22560 29232 22612 29238
rect 22560 29174 22612 29180
rect 22468 29164 22520 29170
rect 22468 29106 22520 29112
rect 22652 29028 22704 29034
rect 22652 28970 22704 28976
rect 22560 28076 22612 28082
rect 22560 28018 22612 28024
rect 22572 27538 22600 28018
rect 22560 27532 22612 27538
rect 22560 27474 22612 27480
rect 22468 26988 22520 26994
rect 22468 26930 22520 26936
rect 22480 26382 22508 26930
rect 22468 26376 22520 26382
rect 22468 26318 22520 26324
rect 22664 24614 22692 28970
rect 22848 28626 22876 31726
rect 23020 31748 23072 31754
rect 23020 31690 23072 31696
rect 22836 28620 22888 28626
rect 22836 28562 22888 28568
rect 22744 27872 22796 27878
rect 22744 27814 22796 27820
rect 22756 26314 22784 27814
rect 22834 26616 22890 26625
rect 22834 26551 22836 26560
rect 22888 26551 22890 26560
rect 22836 26522 22888 26528
rect 22744 26308 22796 26314
rect 22744 26250 22796 26256
rect 22836 26308 22888 26314
rect 22836 26250 22888 26256
rect 22560 24608 22612 24614
rect 22560 24550 22612 24556
rect 22652 24608 22704 24614
rect 22652 24550 22704 24556
rect 22572 24206 22600 24550
rect 22560 24200 22612 24206
rect 22560 24142 22612 24148
rect 22652 23316 22704 23322
rect 22652 23258 22704 23264
rect 22388 22066 22508 22094
rect 22100 22034 22152 22040
rect 21640 21548 21692 21554
rect 21640 21490 21692 21496
rect 21732 21548 21784 21554
rect 21732 21490 21784 21496
rect 21732 19984 21784 19990
rect 21732 19926 21784 19932
rect 21744 19718 21772 19926
rect 21836 19825 21864 22034
rect 21916 21548 21968 21554
rect 21916 21490 21968 21496
rect 21928 21146 21956 21490
rect 21916 21140 21968 21146
rect 21916 21082 21968 21088
rect 22100 20936 22152 20942
rect 22100 20878 22152 20884
rect 22284 20936 22336 20942
rect 22284 20878 22336 20884
rect 22112 20602 22140 20878
rect 22100 20596 22152 20602
rect 22100 20538 22152 20544
rect 21916 20324 21968 20330
rect 21916 20266 21968 20272
rect 21928 20233 21956 20266
rect 22100 20256 22152 20262
rect 21914 20224 21970 20233
rect 22100 20198 22152 20204
rect 21914 20159 21970 20168
rect 21914 20088 21970 20097
rect 21914 20023 21916 20032
rect 21968 20023 21970 20032
rect 21916 19994 21968 20000
rect 22112 19854 22140 20198
rect 22192 19984 22244 19990
rect 22192 19926 22244 19932
rect 22100 19848 22152 19854
rect 21822 19816 21878 19825
rect 22204 19825 22232 19926
rect 22100 19790 22152 19796
rect 22190 19816 22246 19825
rect 21822 19751 21878 19760
rect 21916 19780 21968 19786
rect 21916 19722 21968 19728
rect 21732 19712 21784 19718
rect 21732 19654 21784 19660
rect 21928 18426 21956 19722
rect 22112 19334 22140 19790
rect 22190 19751 22246 19760
rect 22112 19306 22232 19334
rect 22100 19236 22152 19242
rect 22100 19178 22152 19184
rect 22112 18766 22140 19178
rect 22204 19174 22232 19306
rect 22192 19168 22244 19174
rect 22192 19110 22244 19116
rect 22204 18902 22232 19110
rect 22192 18896 22244 18902
rect 22192 18838 22244 18844
rect 22100 18760 22152 18766
rect 22100 18702 22152 18708
rect 22192 18624 22244 18630
rect 22192 18566 22244 18572
rect 21916 18420 21968 18426
rect 21916 18362 21968 18368
rect 22204 18290 22232 18566
rect 22192 18284 22244 18290
rect 22192 18226 22244 18232
rect 22296 17338 22324 20878
rect 22376 19780 22428 19786
rect 22376 19722 22428 19728
rect 22388 19310 22416 19722
rect 22376 19304 22428 19310
rect 22376 19246 22428 19252
rect 22388 18834 22416 19246
rect 22376 18828 22428 18834
rect 22376 18770 22428 18776
rect 21732 17332 21784 17338
rect 21732 17274 21784 17280
rect 22284 17332 22336 17338
rect 22284 17274 22336 17280
rect 21640 16448 21692 16454
rect 21640 16390 21692 16396
rect 21652 16182 21680 16390
rect 21640 16176 21692 16182
rect 21640 16118 21692 16124
rect 21652 15570 21680 16118
rect 21744 16046 21772 17274
rect 22376 17264 22428 17270
rect 22376 17206 22428 17212
rect 22192 16584 22244 16590
rect 22192 16526 22244 16532
rect 21824 16448 21876 16454
rect 21824 16390 21876 16396
rect 21836 16114 21864 16390
rect 21824 16108 21876 16114
rect 21824 16050 21876 16056
rect 21732 16040 21784 16046
rect 21732 15982 21784 15988
rect 21640 15564 21692 15570
rect 21640 15506 21692 15512
rect 21640 14816 21692 14822
rect 21640 14758 21692 14764
rect 21652 14550 21680 14758
rect 21640 14544 21692 14550
rect 21640 14486 21692 14492
rect 21652 13938 21680 14486
rect 21640 13932 21692 13938
rect 21640 13874 21692 13880
rect 21652 13394 21680 13874
rect 21640 13388 21692 13394
rect 21640 13330 21692 13336
rect 21652 12986 21680 13330
rect 21640 12980 21692 12986
rect 21640 12922 21692 12928
rect 21640 12844 21692 12850
rect 21640 12786 21692 12792
rect 21652 12442 21680 12786
rect 21468 12406 21588 12434
rect 21640 12436 21692 12442
rect 21364 11552 21416 11558
rect 21364 11494 21416 11500
rect 21376 11082 21404 11494
rect 21364 11076 21416 11082
rect 21364 11018 21416 11024
rect 21284 8486 21404 8514
rect 21272 8424 21324 8430
rect 21272 8366 21324 8372
rect 21284 8090 21312 8366
rect 21272 8084 21324 8090
rect 21272 8026 21324 8032
rect 21376 7834 21404 8486
rect 21468 8022 21496 12406
rect 21640 12378 21692 12384
rect 21744 11744 21772 15982
rect 21824 15428 21876 15434
rect 21824 15370 21876 15376
rect 21836 14414 21864 15370
rect 22204 15366 22232 16526
rect 22388 15978 22416 17206
rect 22376 15972 22428 15978
rect 22376 15914 22428 15920
rect 22284 15564 22336 15570
rect 22284 15506 22336 15512
rect 22192 15360 22244 15366
rect 22192 15302 22244 15308
rect 21916 14952 21968 14958
rect 21916 14894 21968 14900
rect 21824 14408 21876 14414
rect 21824 14350 21876 14356
rect 21836 14074 21864 14350
rect 21824 14068 21876 14074
rect 21824 14010 21876 14016
rect 21928 13938 21956 14894
rect 22008 14884 22060 14890
rect 22008 14826 22060 14832
rect 21916 13932 21968 13938
rect 21916 13874 21968 13880
rect 21824 13524 21876 13530
rect 21824 13466 21876 13472
rect 21836 12782 21864 13466
rect 21824 12776 21876 12782
rect 21824 12718 21876 12724
rect 21928 12730 21956 13874
rect 22020 13802 22048 14826
rect 22204 14822 22232 15302
rect 22192 14816 22244 14822
rect 22192 14758 22244 14764
rect 22296 14498 22324 15506
rect 22112 14482 22324 14498
rect 22112 14476 22336 14482
rect 22112 14470 22284 14476
rect 22008 13796 22060 13802
rect 22008 13738 22060 13744
rect 22020 13530 22048 13738
rect 22008 13524 22060 13530
rect 22008 13466 22060 13472
rect 22112 13326 22140 14470
rect 22284 14418 22336 14424
rect 22192 14408 22244 14414
rect 22192 14350 22244 14356
rect 22008 13320 22060 13326
rect 22008 13262 22060 13268
rect 22100 13320 22152 13326
rect 22100 13262 22152 13268
rect 22020 12850 22048 13262
rect 22204 13258 22232 14350
rect 22284 13864 22336 13870
rect 22284 13806 22336 13812
rect 22296 13394 22324 13806
rect 22284 13388 22336 13394
rect 22284 13330 22336 13336
rect 22376 13320 22428 13326
rect 22376 13262 22428 13268
rect 22192 13252 22244 13258
rect 22192 13194 22244 13200
rect 22008 12844 22060 12850
rect 22008 12786 22060 12792
rect 21928 12702 22048 12730
rect 21916 11756 21968 11762
rect 21744 11716 21916 11744
rect 21916 11698 21968 11704
rect 21824 11144 21876 11150
rect 21824 11086 21876 11092
rect 21836 9926 21864 11086
rect 21824 9920 21876 9926
rect 21824 9862 21876 9868
rect 21548 9376 21600 9382
rect 21548 9318 21600 9324
rect 21560 9042 21588 9318
rect 21548 9036 21600 9042
rect 21548 8978 21600 8984
rect 21836 8906 21864 9862
rect 21928 9042 21956 11698
rect 22020 9654 22048 12702
rect 22388 12238 22416 13262
rect 22480 12434 22508 22066
rect 22560 20528 22612 20534
rect 22558 20496 22560 20505
rect 22612 20496 22614 20505
rect 22558 20431 22614 20440
rect 22558 20360 22614 20369
rect 22558 20295 22614 20304
rect 22572 20058 22600 20295
rect 22560 20052 22612 20058
rect 22560 19994 22612 20000
rect 22558 19952 22614 19961
rect 22558 19887 22614 19896
rect 22572 19378 22600 19887
rect 22560 19372 22612 19378
rect 22560 19314 22612 19320
rect 22560 18964 22612 18970
rect 22560 18906 22612 18912
rect 22572 18290 22600 18906
rect 22560 18284 22612 18290
rect 22560 18226 22612 18232
rect 22560 17740 22612 17746
rect 22560 17682 22612 17688
rect 22572 17610 22600 17682
rect 22560 17604 22612 17610
rect 22560 17546 22612 17552
rect 22572 16998 22600 17546
rect 22560 16992 22612 16998
rect 22560 16934 22612 16940
rect 22560 16516 22612 16522
rect 22560 16458 22612 16464
rect 22572 16046 22600 16458
rect 22560 16040 22612 16046
rect 22560 15982 22612 15988
rect 22560 15496 22612 15502
rect 22560 15438 22612 15444
rect 22572 13734 22600 15438
rect 22664 14278 22692 23258
rect 22848 22386 22876 26250
rect 23032 24970 23060 31690
rect 22940 24942 23060 24970
rect 22940 23118 22968 24942
rect 23020 24812 23072 24818
rect 23020 24754 23072 24760
rect 23032 24070 23060 24754
rect 23020 24064 23072 24070
rect 23020 24006 23072 24012
rect 23124 23322 23152 47534
rect 23296 37120 23348 37126
rect 23296 37062 23348 37068
rect 23308 33318 23336 37062
rect 23572 36032 23624 36038
rect 23572 35974 23624 35980
rect 23584 34746 23612 35974
rect 23572 34740 23624 34746
rect 23572 34682 23624 34688
rect 23480 34400 23532 34406
rect 23480 34342 23532 34348
rect 23492 33590 23520 34342
rect 23480 33584 23532 33590
rect 23480 33526 23532 33532
rect 23296 33312 23348 33318
rect 23296 33254 23348 33260
rect 23572 33312 23624 33318
rect 23572 33254 23624 33260
rect 23204 32768 23256 32774
rect 23204 32710 23256 32716
rect 23216 32570 23244 32710
rect 23204 32564 23256 32570
rect 23204 32506 23256 32512
rect 23204 32224 23256 32230
rect 23204 32166 23256 32172
rect 23216 29170 23244 32166
rect 23308 31890 23336 33254
rect 23584 32910 23612 33254
rect 23572 32904 23624 32910
rect 23572 32846 23624 32852
rect 23480 32836 23532 32842
rect 23480 32778 23532 32784
rect 23492 32570 23520 32778
rect 23388 32564 23440 32570
rect 23388 32506 23440 32512
rect 23480 32564 23532 32570
rect 23480 32506 23532 32512
rect 23296 31884 23348 31890
rect 23296 31826 23348 31832
rect 23400 31278 23428 32506
rect 23572 32412 23624 32418
rect 23572 32354 23624 32360
rect 23480 32224 23532 32230
rect 23480 32166 23532 32172
rect 23492 31822 23520 32166
rect 23584 31958 23612 32354
rect 23572 31952 23624 31958
rect 23572 31894 23624 31900
rect 23480 31816 23532 31822
rect 23480 31758 23532 31764
rect 23492 31414 23520 31758
rect 23676 31754 23704 47602
rect 24308 47252 24360 47258
rect 24308 47194 24360 47200
rect 24032 38956 24084 38962
rect 24032 38898 24084 38904
rect 23940 38888 23992 38894
rect 23940 38830 23992 38836
rect 23952 38350 23980 38830
rect 23940 38344 23992 38350
rect 23940 38286 23992 38292
rect 24044 38010 24072 38898
rect 24032 38004 24084 38010
rect 24032 37946 24084 37952
rect 24320 37874 24348 47194
rect 24400 39500 24452 39506
rect 24400 39442 24452 39448
rect 24412 38010 24440 39442
rect 24504 39438 24532 49098
rect 24596 48210 24624 51326
rect 25134 51200 25190 52000
rect 25778 51354 25834 52000
rect 26422 51354 26478 52000
rect 25608 51326 25834 51354
rect 24676 49224 24728 49230
rect 24676 49166 24728 49172
rect 24688 48890 24716 49166
rect 24676 48884 24728 48890
rect 24676 48826 24728 48832
rect 25412 48748 25464 48754
rect 25412 48690 25464 48696
rect 24584 48204 24636 48210
rect 24584 48146 24636 48152
rect 24676 48068 24728 48074
rect 24676 48010 24728 48016
rect 24688 47666 24716 48010
rect 24676 47660 24728 47666
rect 24676 47602 24728 47608
rect 24952 47660 25004 47666
rect 24952 47602 25004 47608
rect 24964 47054 24992 47602
rect 25424 47258 25452 48690
rect 25412 47252 25464 47258
rect 25412 47194 25464 47200
rect 25608 47054 25636 51326
rect 25778 51200 25834 51326
rect 26252 51326 26478 51354
rect 26148 47796 26200 47802
rect 26148 47738 26200 47744
rect 26056 47660 26108 47666
rect 26056 47602 26108 47608
rect 25872 47592 25924 47598
rect 25872 47534 25924 47540
rect 25964 47592 26016 47598
rect 25964 47534 26016 47540
rect 24952 47048 25004 47054
rect 24952 46990 25004 46996
rect 25596 47048 25648 47054
rect 25596 46990 25648 46996
rect 24492 39432 24544 39438
rect 24492 39374 24544 39380
rect 24952 39432 25004 39438
rect 24952 39374 25004 39380
rect 24492 39296 24544 39302
rect 24492 39238 24544 39244
rect 24504 38350 24532 39238
rect 24492 38344 24544 38350
rect 24492 38286 24544 38292
rect 24768 38208 24820 38214
rect 24768 38150 24820 38156
rect 24400 38004 24452 38010
rect 24400 37946 24452 37952
rect 24308 37868 24360 37874
rect 24308 37810 24360 37816
rect 24124 37732 24176 37738
rect 24124 37674 24176 37680
rect 24136 37398 24164 37674
rect 24124 37392 24176 37398
rect 24124 37334 24176 37340
rect 24136 35018 24164 37334
rect 24412 36174 24440 37946
rect 24584 36848 24636 36854
rect 24584 36790 24636 36796
rect 24596 36378 24624 36790
rect 24584 36372 24636 36378
rect 24584 36314 24636 36320
rect 24780 36242 24808 38150
rect 24964 37874 24992 39374
rect 25044 38752 25096 38758
rect 25044 38694 25096 38700
rect 24952 37868 25004 37874
rect 24952 37810 25004 37816
rect 24964 36582 24992 37810
rect 25056 36854 25084 38694
rect 25780 38208 25832 38214
rect 25780 38150 25832 38156
rect 25136 37868 25188 37874
rect 25136 37810 25188 37816
rect 25148 36922 25176 37810
rect 25504 37324 25556 37330
rect 25504 37266 25556 37272
rect 25136 36916 25188 36922
rect 25136 36858 25188 36864
rect 25228 36916 25280 36922
rect 25228 36858 25280 36864
rect 25044 36848 25096 36854
rect 25044 36790 25096 36796
rect 24952 36576 25004 36582
rect 24952 36518 25004 36524
rect 24768 36236 24820 36242
rect 24768 36178 24820 36184
rect 24400 36168 24452 36174
rect 24400 36110 24452 36116
rect 24216 35692 24268 35698
rect 24216 35634 24268 35640
rect 24308 35692 24360 35698
rect 24308 35634 24360 35640
rect 24228 35222 24256 35634
rect 24216 35216 24268 35222
rect 24216 35158 24268 35164
rect 24124 35012 24176 35018
rect 24124 34954 24176 34960
rect 24032 34400 24084 34406
rect 24032 34342 24084 34348
rect 24044 33998 24072 34342
rect 24032 33992 24084 33998
rect 24032 33934 24084 33940
rect 24124 33992 24176 33998
rect 24124 33934 24176 33940
rect 23756 33856 23808 33862
rect 23756 33798 23808 33804
rect 23768 32910 23796 33798
rect 24136 33658 24164 33934
rect 24228 33930 24256 35158
rect 24320 35086 24348 35634
rect 24412 35630 24440 36110
rect 24400 35624 24452 35630
rect 24400 35566 24452 35572
rect 24492 35148 24544 35154
rect 24492 35090 24544 35096
rect 24308 35080 24360 35086
rect 24308 35022 24360 35028
rect 24504 34746 24532 35090
rect 24676 35080 24728 35086
rect 24676 35022 24728 35028
rect 24492 34740 24544 34746
rect 24492 34682 24544 34688
rect 24584 34536 24636 34542
rect 24584 34478 24636 34484
rect 24596 34202 24624 34478
rect 24584 34196 24636 34202
rect 24584 34138 24636 34144
rect 24596 34105 24624 34138
rect 24582 34096 24638 34105
rect 24582 34031 24638 34040
rect 24216 33924 24268 33930
rect 24216 33866 24268 33872
rect 24492 33924 24544 33930
rect 24492 33866 24544 33872
rect 24124 33652 24176 33658
rect 24124 33594 24176 33600
rect 23940 33516 23992 33522
rect 23940 33458 23992 33464
rect 24216 33516 24268 33522
rect 24216 33458 24268 33464
rect 23848 33108 23900 33114
rect 23848 33050 23900 33056
rect 23756 32904 23808 32910
rect 23756 32846 23808 32852
rect 23756 32360 23808 32366
rect 23860 32348 23888 33050
rect 23952 32434 23980 33458
rect 24228 33046 24256 33458
rect 24400 33312 24452 33318
rect 24400 33254 24452 33260
rect 24216 33040 24268 33046
rect 24216 32982 24268 32988
rect 24308 32972 24360 32978
rect 24308 32914 24360 32920
rect 24032 32496 24084 32502
rect 24030 32464 24032 32473
rect 24084 32464 24086 32473
rect 23940 32428 23992 32434
rect 24030 32399 24086 32408
rect 23940 32370 23992 32376
rect 23808 32320 23888 32348
rect 23756 32302 23808 32308
rect 23952 32026 23980 32370
rect 23940 32020 23992 32026
rect 23940 31962 23992 31968
rect 24124 31816 24176 31822
rect 24124 31758 24176 31764
rect 23584 31726 23704 31754
rect 23480 31408 23532 31414
rect 23480 31350 23532 31356
rect 23388 31272 23440 31278
rect 23388 31214 23440 31220
rect 23388 31136 23440 31142
rect 23388 31078 23440 31084
rect 23296 30660 23348 30666
rect 23296 30602 23348 30608
rect 23308 30190 23336 30602
rect 23400 30598 23428 31078
rect 23388 30592 23440 30598
rect 23388 30534 23440 30540
rect 23400 30190 23428 30534
rect 23296 30184 23348 30190
rect 23296 30126 23348 30132
rect 23388 30184 23440 30190
rect 23388 30126 23440 30132
rect 23204 29164 23256 29170
rect 23204 29106 23256 29112
rect 23388 29096 23440 29102
rect 23388 29038 23440 29044
rect 23400 28490 23428 29038
rect 23388 28484 23440 28490
rect 23388 28426 23440 28432
rect 23480 28076 23532 28082
rect 23480 28018 23532 28024
rect 23204 26580 23256 26586
rect 23204 26522 23256 26528
rect 23216 24018 23244 26522
rect 23492 25974 23520 28018
rect 23584 26625 23612 31726
rect 23940 30252 23992 30258
rect 23940 30194 23992 30200
rect 23952 29782 23980 30194
rect 23940 29776 23992 29782
rect 23940 29718 23992 29724
rect 23664 28416 23716 28422
rect 23664 28358 23716 28364
rect 23676 27946 23704 28358
rect 23952 28150 23980 29718
rect 23940 28144 23992 28150
rect 23940 28086 23992 28092
rect 24032 28076 24084 28082
rect 24032 28018 24084 28024
rect 23664 27940 23716 27946
rect 23664 27882 23716 27888
rect 23570 26616 23626 26625
rect 23570 26551 23626 26560
rect 23572 26512 23624 26518
rect 23572 26454 23624 26460
rect 23296 25968 23348 25974
rect 23296 25910 23348 25916
rect 23480 25968 23532 25974
rect 23480 25910 23532 25916
rect 23308 25294 23336 25910
rect 23388 25900 23440 25906
rect 23388 25842 23440 25848
rect 23400 25786 23428 25842
rect 23584 25786 23612 26454
rect 23400 25758 23612 25786
rect 23296 25288 23348 25294
rect 23296 25230 23348 25236
rect 23480 24812 23532 24818
rect 23480 24754 23532 24760
rect 23388 24608 23440 24614
rect 23388 24550 23440 24556
rect 23400 24342 23428 24550
rect 23388 24336 23440 24342
rect 23388 24278 23440 24284
rect 23216 23990 23336 24018
rect 23204 23724 23256 23730
rect 23204 23666 23256 23672
rect 23112 23316 23164 23322
rect 23112 23258 23164 23264
rect 22928 23112 22980 23118
rect 22928 23054 22980 23060
rect 23216 22506 23244 23666
rect 23308 23050 23336 23990
rect 23492 23662 23520 24754
rect 23572 24744 23624 24750
rect 23572 24686 23624 24692
rect 23584 24614 23612 24686
rect 23572 24608 23624 24614
rect 23572 24550 23624 24556
rect 23480 23656 23532 23662
rect 23480 23598 23532 23604
rect 23296 23044 23348 23050
rect 23296 22986 23348 22992
rect 23204 22500 23256 22506
rect 23204 22442 23256 22448
rect 22848 22358 23244 22386
rect 23020 20868 23072 20874
rect 23020 20810 23072 20816
rect 22928 20392 22980 20398
rect 22928 20334 22980 20340
rect 22744 20052 22796 20058
rect 22744 19994 22796 20000
rect 22756 19242 22784 19994
rect 22836 19848 22888 19854
rect 22834 19816 22836 19825
rect 22888 19816 22890 19825
rect 22834 19751 22890 19760
rect 22836 19712 22888 19718
rect 22836 19654 22888 19660
rect 22848 19310 22876 19654
rect 22940 19514 22968 20334
rect 22928 19508 22980 19514
rect 22928 19450 22980 19456
rect 22926 19408 22982 19417
rect 22926 19343 22982 19352
rect 22836 19304 22888 19310
rect 22836 19246 22888 19252
rect 22744 19236 22796 19242
rect 22744 19178 22796 19184
rect 22744 18760 22796 18766
rect 22744 18702 22796 18708
rect 22756 17592 22784 18702
rect 22848 18426 22876 19246
rect 22836 18420 22888 18426
rect 22836 18362 22888 18368
rect 22836 17604 22888 17610
rect 22756 17564 22836 17592
rect 22836 17546 22888 17552
rect 22848 17354 22876 17546
rect 22940 17542 22968 19343
rect 23032 18426 23060 20810
rect 23112 20800 23164 20806
rect 23112 20742 23164 20748
rect 23124 20398 23152 20742
rect 23112 20392 23164 20398
rect 23112 20334 23164 20340
rect 23124 19802 23152 20334
rect 23216 19938 23244 22358
rect 23308 22094 23336 22986
rect 23492 22794 23520 23598
rect 23676 22930 23704 27882
rect 23940 27872 23992 27878
rect 23940 27814 23992 27820
rect 23952 26994 23980 27814
rect 24044 27674 24072 28018
rect 24032 27668 24084 27674
rect 24032 27610 24084 27616
rect 23940 26988 23992 26994
rect 23940 26930 23992 26936
rect 24136 26874 24164 31758
rect 24216 31272 24268 31278
rect 24216 31214 24268 31220
rect 23952 26846 24164 26874
rect 23756 23520 23808 23526
rect 23756 23462 23808 23468
rect 23768 23118 23796 23462
rect 23756 23112 23808 23118
rect 23756 23054 23808 23060
rect 23676 22902 23796 22930
rect 23492 22766 23612 22794
rect 23584 22710 23612 22766
rect 23572 22704 23624 22710
rect 23572 22646 23624 22652
rect 23664 22636 23716 22642
rect 23664 22578 23716 22584
rect 23572 22568 23624 22574
rect 23572 22510 23624 22516
rect 23308 22066 23428 22094
rect 23296 21344 23348 21350
rect 23296 21286 23348 21292
rect 23308 20874 23336 21286
rect 23400 21010 23428 22066
rect 23584 21962 23612 22510
rect 23572 21956 23624 21962
rect 23572 21898 23624 21904
rect 23572 21548 23624 21554
rect 23572 21490 23624 21496
rect 23480 21344 23532 21350
rect 23480 21286 23532 21292
rect 23388 21004 23440 21010
rect 23388 20946 23440 20952
rect 23296 20868 23348 20874
rect 23296 20810 23348 20816
rect 23296 20392 23348 20398
rect 23296 20334 23348 20340
rect 23308 20058 23336 20334
rect 23400 20058 23428 20946
rect 23492 20466 23520 21286
rect 23584 21010 23612 21490
rect 23572 21004 23624 21010
rect 23572 20946 23624 20952
rect 23572 20800 23624 20806
rect 23572 20742 23624 20748
rect 23584 20466 23612 20742
rect 23480 20460 23532 20466
rect 23480 20402 23532 20408
rect 23572 20460 23624 20466
rect 23572 20402 23624 20408
rect 23296 20052 23348 20058
rect 23296 19994 23348 20000
rect 23388 20052 23440 20058
rect 23388 19994 23440 20000
rect 23216 19910 23336 19938
rect 23124 19774 23244 19802
rect 23216 19718 23244 19774
rect 23112 19712 23164 19718
rect 23112 19654 23164 19660
rect 23204 19712 23256 19718
rect 23204 19654 23256 19660
rect 23124 18834 23152 19654
rect 23112 18828 23164 18834
rect 23112 18770 23164 18776
rect 23020 18420 23072 18426
rect 23020 18362 23072 18368
rect 23204 18284 23256 18290
rect 23032 18244 23204 18272
rect 23032 18154 23060 18244
rect 23204 18226 23256 18232
rect 23308 18170 23336 19910
rect 23400 19310 23428 19994
rect 23584 19961 23612 20402
rect 23570 19952 23626 19961
rect 23570 19887 23626 19896
rect 23480 19372 23532 19378
rect 23480 19314 23532 19320
rect 23388 19304 23440 19310
rect 23388 19246 23440 19252
rect 23400 18290 23428 19246
rect 23492 18766 23520 19314
rect 23480 18760 23532 18766
rect 23480 18702 23532 18708
rect 23388 18284 23440 18290
rect 23388 18226 23440 18232
rect 23020 18148 23072 18154
rect 23020 18090 23072 18096
rect 23124 18142 23336 18170
rect 22928 17536 22980 17542
rect 22928 17478 22980 17484
rect 22848 17326 22968 17354
rect 22940 17202 22968 17326
rect 22928 17196 22980 17202
rect 22928 17138 22980 17144
rect 22940 16522 22968 17138
rect 23020 16584 23072 16590
rect 23020 16526 23072 16532
rect 22928 16516 22980 16522
rect 22928 16458 22980 16464
rect 22744 16448 22796 16454
rect 22744 16390 22796 16396
rect 22756 15502 22784 16390
rect 22744 15496 22796 15502
rect 22744 15438 22796 15444
rect 22652 14272 22704 14278
rect 22652 14214 22704 14220
rect 22744 14272 22796 14278
rect 22744 14214 22796 14220
rect 22560 13728 22612 13734
rect 22560 13670 22612 13676
rect 22652 13184 22704 13190
rect 22652 13126 22704 13132
rect 22664 12850 22692 13126
rect 22652 12844 22704 12850
rect 22652 12786 22704 12792
rect 22480 12406 22600 12434
rect 22100 12232 22152 12238
rect 22100 12174 22152 12180
rect 22376 12232 22428 12238
rect 22376 12174 22428 12180
rect 22112 11762 22140 12174
rect 22376 12096 22428 12102
rect 22376 12038 22428 12044
rect 22192 11892 22244 11898
rect 22192 11834 22244 11840
rect 22100 11756 22152 11762
rect 22100 11698 22152 11704
rect 22112 11354 22140 11698
rect 22204 11694 22232 11834
rect 22388 11762 22416 12038
rect 22376 11756 22428 11762
rect 22376 11698 22428 11704
rect 22192 11688 22244 11694
rect 22192 11630 22244 11636
rect 22100 11348 22152 11354
rect 22100 11290 22152 11296
rect 22468 9716 22520 9722
rect 22468 9658 22520 9664
rect 22008 9648 22060 9654
rect 22008 9590 22060 9596
rect 22480 9178 22508 9658
rect 22468 9172 22520 9178
rect 22468 9114 22520 9120
rect 22100 9104 22152 9110
rect 22100 9046 22152 9052
rect 21916 9036 21968 9042
rect 21916 8978 21968 8984
rect 21824 8900 21876 8906
rect 21824 8842 21876 8848
rect 21836 8430 21864 8842
rect 21824 8424 21876 8430
rect 21824 8366 21876 8372
rect 21456 8016 21508 8022
rect 21456 7958 21508 7964
rect 21376 7806 21496 7834
rect 21088 6656 21140 6662
rect 21088 6598 21140 6604
rect 20996 6384 21048 6390
rect 20996 6326 21048 6332
rect 21100 5234 21128 6598
rect 21088 5228 21140 5234
rect 21088 5170 21140 5176
rect 20812 4072 20864 4078
rect 20812 4014 20864 4020
rect 21180 4072 21232 4078
rect 21180 4014 21232 4020
rect 20640 3726 20760 3754
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 20536 2508 20588 2514
rect 20536 2450 20588 2456
rect 20076 2304 20128 2310
rect 20076 2246 20128 2252
rect 20640 800 20668 3538
rect 20732 3194 20760 3726
rect 20824 3602 20852 4014
rect 20812 3596 20864 3602
rect 20812 3538 20864 3544
rect 20720 3188 20772 3194
rect 20720 3130 20772 3136
rect 21192 3058 21220 4014
rect 21272 4004 21324 4010
rect 21272 3946 21324 3952
rect 21180 3052 21232 3058
rect 21180 2994 21232 3000
rect 21178 2952 21234 2961
rect 21178 2887 21180 2896
rect 21232 2887 21234 2896
rect 21180 2858 21232 2864
rect 21284 800 21312 3946
rect 21468 2922 21496 7806
rect 21640 5772 21692 5778
rect 21640 5714 21692 5720
rect 21652 5098 21680 5714
rect 21836 5710 21864 8366
rect 22112 8022 22140 9046
rect 22192 8968 22244 8974
rect 22190 8936 22192 8945
rect 22376 8968 22428 8974
rect 22244 8936 22246 8945
rect 22376 8910 22428 8916
rect 22468 8968 22520 8974
rect 22468 8910 22520 8916
rect 22190 8871 22246 8880
rect 22388 8838 22416 8910
rect 22376 8832 22428 8838
rect 22376 8774 22428 8780
rect 22100 8016 22152 8022
rect 22100 7958 22152 7964
rect 22480 7750 22508 8910
rect 22468 7744 22520 7750
rect 22468 7686 22520 7692
rect 22480 6798 22508 7686
rect 22468 6792 22520 6798
rect 22468 6734 22520 6740
rect 22008 6384 22060 6390
rect 22008 6326 22060 6332
rect 22020 5846 22048 6326
rect 22008 5840 22060 5846
rect 22008 5782 22060 5788
rect 21824 5704 21876 5710
rect 21824 5646 21876 5652
rect 22284 5704 22336 5710
rect 22284 5646 22336 5652
rect 21836 5234 21864 5646
rect 21824 5228 21876 5234
rect 21824 5170 21876 5176
rect 21640 5092 21692 5098
rect 21640 5034 21692 5040
rect 22008 4004 22060 4010
rect 21928 3964 22008 3992
rect 21928 3602 21956 3964
rect 22008 3946 22060 3952
rect 21916 3596 21968 3602
rect 21916 3538 21968 3544
rect 21456 2916 21508 2922
rect 21456 2858 21508 2864
rect 22296 1970 22324 5646
rect 22480 5370 22508 6734
rect 22468 5364 22520 5370
rect 22468 5306 22520 5312
rect 22376 4072 22428 4078
rect 22376 4014 22428 4020
rect 22388 2990 22416 4014
rect 22468 3188 22520 3194
rect 22468 3130 22520 3136
rect 22376 2984 22428 2990
rect 22376 2926 22428 2932
rect 22480 2854 22508 3130
rect 22468 2848 22520 2854
rect 22468 2790 22520 2796
rect 22572 2650 22600 12406
rect 22756 10538 22784 14214
rect 22836 12776 22888 12782
rect 22836 12718 22888 12724
rect 22848 12238 22876 12718
rect 22940 12594 22968 16458
rect 23032 16250 23060 16526
rect 23020 16244 23072 16250
rect 23020 16186 23072 16192
rect 23124 16114 23152 18142
rect 23204 18080 23256 18086
rect 23204 18022 23256 18028
rect 23216 17678 23244 18022
rect 23676 17882 23704 22578
rect 23664 17876 23716 17882
rect 23664 17818 23716 17824
rect 23572 17808 23624 17814
rect 23572 17750 23624 17756
rect 23204 17672 23256 17678
rect 23204 17614 23256 17620
rect 23296 17672 23348 17678
rect 23348 17620 23428 17626
rect 23296 17614 23428 17620
rect 23216 16794 23244 17614
rect 23308 17598 23428 17614
rect 23296 17536 23348 17542
rect 23296 17478 23348 17484
rect 23400 17490 23428 17598
rect 23308 16810 23336 17478
rect 23400 17462 23520 17490
rect 23308 16794 23428 16810
rect 23204 16788 23256 16794
rect 23204 16730 23256 16736
rect 23308 16788 23440 16794
rect 23308 16782 23388 16788
rect 23112 16108 23164 16114
rect 23112 16050 23164 16056
rect 23124 14414 23152 16050
rect 23204 15360 23256 15366
rect 23204 15302 23256 15308
rect 23216 15026 23244 15302
rect 23204 15020 23256 15026
rect 23204 14962 23256 14968
rect 23308 14822 23336 16782
rect 23388 16730 23440 16736
rect 23492 16674 23520 17462
rect 23584 16726 23612 17750
rect 23664 16992 23716 16998
rect 23664 16934 23716 16940
rect 23400 16658 23520 16674
rect 23572 16720 23624 16726
rect 23572 16662 23624 16668
rect 23388 16652 23520 16658
rect 23440 16646 23520 16652
rect 23388 16594 23440 16600
rect 23388 14952 23440 14958
rect 23388 14894 23440 14900
rect 23296 14816 23348 14822
rect 23296 14758 23348 14764
rect 23112 14408 23164 14414
rect 23112 14350 23164 14356
rect 23400 14278 23428 14894
rect 23492 14550 23520 16646
rect 23480 14544 23532 14550
rect 23480 14486 23532 14492
rect 23388 14272 23440 14278
rect 23388 14214 23440 14220
rect 23480 13796 23532 13802
rect 23480 13738 23532 13744
rect 23296 13524 23348 13530
rect 23296 13466 23348 13472
rect 23308 13394 23336 13466
rect 23296 13388 23348 13394
rect 23296 13330 23348 13336
rect 23204 12708 23256 12714
rect 23256 12668 23336 12696
rect 23204 12650 23256 12656
rect 22940 12566 23244 12594
rect 22928 12436 22980 12442
rect 22928 12378 22980 12384
rect 22836 12232 22888 12238
rect 22836 12174 22888 12180
rect 22836 11552 22888 11558
rect 22836 11494 22888 11500
rect 22848 10674 22876 11494
rect 22836 10668 22888 10674
rect 22836 10610 22888 10616
rect 22940 10538 22968 12378
rect 23216 11762 23244 12566
rect 23308 12238 23336 12668
rect 23492 12434 23520 13738
rect 23584 13530 23612 16662
rect 23676 15978 23704 16934
rect 23768 16658 23796 22902
rect 23848 21412 23900 21418
rect 23848 21354 23900 21360
rect 23860 20874 23888 21354
rect 23848 20868 23900 20874
rect 23848 20810 23900 20816
rect 23848 18692 23900 18698
rect 23848 18634 23900 18640
rect 23860 17202 23888 18634
rect 23848 17196 23900 17202
rect 23848 17138 23900 17144
rect 23756 16652 23808 16658
rect 23756 16594 23808 16600
rect 23664 15972 23716 15978
rect 23664 15914 23716 15920
rect 23756 15904 23808 15910
rect 23756 15846 23808 15852
rect 23664 15632 23716 15638
rect 23664 15574 23716 15580
rect 23572 13524 23624 13530
rect 23572 13466 23624 13472
rect 23492 12406 23612 12434
rect 23584 12306 23612 12406
rect 23572 12300 23624 12306
rect 23572 12242 23624 12248
rect 23296 12232 23348 12238
rect 23296 12174 23348 12180
rect 23388 12096 23440 12102
rect 23388 12038 23440 12044
rect 23400 11830 23428 12038
rect 23388 11824 23440 11830
rect 23388 11766 23440 11772
rect 23204 11756 23256 11762
rect 23204 11698 23256 11704
rect 23480 11756 23532 11762
rect 23480 11698 23532 11704
rect 23216 11150 23244 11698
rect 23308 11218 23428 11234
rect 23308 11212 23440 11218
rect 23308 11206 23388 11212
rect 23204 11144 23256 11150
rect 23204 11086 23256 11092
rect 23020 10668 23072 10674
rect 23020 10610 23072 10616
rect 22744 10532 22796 10538
rect 22744 10474 22796 10480
rect 22928 10532 22980 10538
rect 22928 10474 22980 10480
rect 22652 9580 22704 9586
rect 22652 9522 22704 9528
rect 22664 9110 22692 9522
rect 22940 9518 22968 10474
rect 23032 10266 23060 10610
rect 23020 10260 23072 10266
rect 23020 10202 23072 10208
rect 23308 10062 23336 11206
rect 23388 11154 23440 11160
rect 23388 11076 23440 11082
rect 23388 11018 23440 11024
rect 23400 10810 23428 11018
rect 23492 11014 23520 11698
rect 23480 11008 23532 11014
rect 23480 10950 23532 10956
rect 23388 10804 23440 10810
rect 23388 10746 23440 10752
rect 23480 10464 23532 10470
rect 23480 10406 23532 10412
rect 23584 10418 23612 12242
rect 23676 10606 23704 15574
rect 23768 12238 23796 15846
rect 23848 15360 23900 15366
rect 23848 15302 23900 15308
rect 23860 15094 23888 15302
rect 23848 15088 23900 15094
rect 23848 15030 23900 15036
rect 23860 14482 23888 15030
rect 23848 14476 23900 14482
rect 23848 14418 23900 14424
rect 23848 13388 23900 13394
rect 23848 13330 23900 13336
rect 23756 12232 23808 12238
rect 23756 12174 23808 12180
rect 23756 11824 23808 11830
rect 23756 11766 23808 11772
rect 23768 11558 23796 11766
rect 23756 11552 23808 11558
rect 23756 11494 23808 11500
rect 23860 11354 23888 13330
rect 23848 11348 23900 11354
rect 23848 11290 23900 11296
rect 23860 10810 23888 11290
rect 23848 10804 23900 10810
rect 23848 10746 23900 10752
rect 23664 10600 23716 10606
rect 23664 10542 23716 10548
rect 23492 10130 23520 10406
rect 23584 10390 23704 10418
rect 23480 10124 23532 10130
rect 23480 10066 23532 10072
rect 23296 10056 23348 10062
rect 23296 9998 23348 10004
rect 23308 9722 23336 9998
rect 23480 9920 23532 9926
rect 23480 9862 23532 9868
rect 23296 9716 23348 9722
rect 23296 9658 23348 9664
rect 22928 9512 22980 9518
rect 22928 9454 22980 9460
rect 22652 9104 22704 9110
rect 22652 9046 22704 9052
rect 22744 9104 22796 9110
rect 22744 9046 22796 9052
rect 22650 8936 22706 8945
rect 22650 8871 22652 8880
rect 22704 8871 22706 8880
rect 22652 8842 22704 8848
rect 22756 8566 22784 9046
rect 23204 9036 23256 9042
rect 23204 8978 23256 8984
rect 22744 8560 22796 8566
rect 22744 8502 22796 8508
rect 23216 8294 23244 8978
rect 23204 8288 23256 8294
rect 23204 8230 23256 8236
rect 23216 7886 23244 8230
rect 23492 7886 23520 9862
rect 23572 8968 23624 8974
rect 23572 8910 23624 8916
rect 23584 8634 23612 8910
rect 23572 8628 23624 8634
rect 23572 8570 23624 8576
rect 23676 7954 23704 10390
rect 23848 9580 23900 9586
rect 23848 9522 23900 9528
rect 23756 9376 23808 9382
rect 23756 9318 23808 9324
rect 23768 8945 23796 9318
rect 23860 8974 23888 9522
rect 23848 8968 23900 8974
rect 23754 8936 23810 8945
rect 23848 8910 23900 8916
rect 23754 8871 23810 8880
rect 23664 7948 23716 7954
rect 23664 7890 23716 7896
rect 23204 7880 23256 7886
rect 23204 7822 23256 7828
rect 23480 7880 23532 7886
rect 23480 7822 23532 7828
rect 23492 7410 23520 7822
rect 23480 7404 23532 7410
rect 23480 7346 23532 7352
rect 23572 6316 23624 6322
rect 23572 6258 23624 6264
rect 23848 6316 23900 6322
rect 23848 6258 23900 6264
rect 22928 6112 22980 6118
rect 22928 6054 22980 6060
rect 23388 6112 23440 6118
rect 23388 6054 23440 6060
rect 22940 5710 22968 6054
rect 23400 5710 23428 6054
rect 22928 5704 22980 5710
rect 22928 5646 22980 5652
rect 23112 5704 23164 5710
rect 23112 5646 23164 5652
rect 23388 5704 23440 5710
rect 23388 5646 23440 5652
rect 23124 5234 23152 5646
rect 23112 5228 23164 5234
rect 23112 5170 23164 5176
rect 22744 3528 22796 3534
rect 22744 3470 22796 3476
rect 22652 3188 22704 3194
rect 22652 3130 22704 3136
rect 22664 2961 22692 3130
rect 22756 3058 22784 3470
rect 22744 3052 22796 3058
rect 22744 2994 22796 3000
rect 22650 2952 22706 2961
rect 22650 2887 22706 2896
rect 23584 2650 23612 6258
rect 23860 5370 23888 6258
rect 23848 5364 23900 5370
rect 23848 5306 23900 5312
rect 23664 3392 23716 3398
rect 23664 3334 23716 3340
rect 23756 3392 23808 3398
rect 23756 3334 23808 3340
rect 23676 3126 23704 3334
rect 23664 3120 23716 3126
rect 23664 3062 23716 3068
rect 23768 2990 23796 3334
rect 23756 2984 23808 2990
rect 23756 2926 23808 2932
rect 23848 2984 23900 2990
rect 23848 2926 23900 2932
rect 22560 2644 22612 2650
rect 22560 2586 22612 2592
rect 23572 2644 23624 2650
rect 23572 2586 23624 2592
rect 23204 2440 23256 2446
rect 23204 2382 23256 2388
rect 22560 2372 22612 2378
rect 22560 2314 22612 2320
rect 22284 1964 22336 1970
rect 22284 1906 22336 1912
rect 22572 800 22600 2314
rect 23216 800 23244 2382
rect 23860 800 23888 2926
rect 23952 1970 23980 26846
rect 24124 26444 24176 26450
rect 24124 26386 24176 26392
rect 24136 21554 24164 26386
rect 24228 22094 24256 31214
rect 24320 30802 24348 32914
rect 24412 32609 24440 33254
rect 24398 32600 24454 32609
rect 24398 32535 24454 32544
rect 24412 31754 24440 32535
rect 24504 32434 24532 33866
rect 24596 33454 24624 34031
rect 24584 33448 24636 33454
rect 24584 33390 24636 33396
rect 24492 32428 24544 32434
rect 24492 32370 24544 32376
rect 24504 32230 24532 32370
rect 24596 32366 24624 33390
rect 24688 32570 24716 35022
rect 24780 34678 24808 36178
rect 24860 36100 24912 36106
rect 24860 36042 24912 36048
rect 24872 35834 24900 36042
rect 25056 35834 25084 36790
rect 25240 36582 25268 36858
rect 25516 36718 25544 37266
rect 25792 37194 25820 38150
rect 25780 37188 25832 37194
rect 25780 37130 25832 37136
rect 25504 36712 25556 36718
rect 25504 36654 25556 36660
rect 25228 36576 25280 36582
rect 25228 36518 25280 36524
rect 24860 35828 24912 35834
rect 24860 35770 24912 35776
rect 25044 35828 25096 35834
rect 25044 35770 25096 35776
rect 25056 35290 25084 35770
rect 25240 35698 25268 36518
rect 25320 36032 25372 36038
rect 25320 35974 25372 35980
rect 25228 35692 25280 35698
rect 25228 35634 25280 35640
rect 25044 35284 25096 35290
rect 25044 35226 25096 35232
rect 24860 34944 24912 34950
rect 24860 34886 24912 34892
rect 24768 34672 24820 34678
rect 24768 34614 24820 34620
rect 24780 33658 24808 34614
rect 24872 34066 24900 34886
rect 25228 34536 25280 34542
rect 25228 34478 25280 34484
rect 25240 34134 25268 34478
rect 25332 34406 25360 35974
rect 25516 35562 25544 36654
rect 25504 35556 25556 35562
rect 25504 35498 25556 35504
rect 25516 35290 25544 35498
rect 25504 35284 25556 35290
rect 25504 35226 25556 35232
rect 25596 34944 25648 34950
rect 25596 34886 25648 34892
rect 25412 34604 25464 34610
rect 25412 34546 25464 34552
rect 25320 34400 25372 34406
rect 25320 34342 25372 34348
rect 25228 34128 25280 34134
rect 25228 34070 25280 34076
rect 24860 34060 24912 34066
rect 24860 34002 24912 34008
rect 24768 33652 24820 33658
rect 24768 33594 24820 33600
rect 24780 33114 24808 33594
rect 25332 33386 25360 34342
rect 25424 34134 25452 34546
rect 25412 34128 25464 34134
rect 25412 34070 25464 34076
rect 25424 33522 25452 34070
rect 25504 33992 25556 33998
rect 25608 33980 25636 34886
rect 25792 34610 25820 37130
rect 25780 34604 25832 34610
rect 25780 34546 25832 34552
rect 25556 33952 25636 33980
rect 25504 33934 25556 33940
rect 25412 33516 25464 33522
rect 25412 33458 25464 33464
rect 25320 33380 25372 33386
rect 25320 33322 25372 33328
rect 24768 33108 24820 33114
rect 24768 33050 24820 33056
rect 25780 32836 25832 32842
rect 25780 32778 25832 32784
rect 24860 32768 24912 32774
rect 24860 32710 24912 32716
rect 24676 32564 24728 32570
rect 24676 32506 24728 32512
rect 24584 32360 24636 32366
rect 24584 32302 24636 32308
rect 24492 32224 24544 32230
rect 24492 32166 24544 32172
rect 24688 32042 24716 32506
rect 24688 32014 24808 32042
rect 24412 31726 24716 31754
rect 24492 31680 24544 31686
rect 24492 31622 24544 31628
rect 24308 30796 24360 30802
rect 24308 30738 24360 30744
rect 24504 30734 24532 31622
rect 24584 31136 24636 31142
rect 24584 31078 24636 31084
rect 24492 30728 24544 30734
rect 24492 30670 24544 30676
rect 24596 30258 24624 31078
rect 24584 30252 24636 30258
rect 24584 30194 24636 30200
rect 24308 29572 24360 29578
rect 24308 29514 24360 29520
rect 24320 29306 24348 29514
rect 24308 29300 24360 29306
rect 24308 29242 24360 29248
rect 24596 28490 24624 30194
rect 24688 28694 24716 31726
rect 24780 30666 24808 32014
rect 24872 31822 24900 32710
rect 25792 32230 25820 32778
rect 25780 32224 25832 32230
rect 25780 32166 25832 32172
rect 24860 31816 24912 31822
rect 25228 31816 25280 31822
rect 24860 31758 24912 31764
rect 25226 31784 25228 31793
rect 25280 31784 25282 31793
rect 25226 31719 25282 31728
rect 25792 31346 25820 32166
rect 25044 31340 25096 31346
rect 25044 31282 25096 31288
rect 25780 31340 25832 31346
rect 25780 31282 25832 31288
rect 25056 31226 25084 31282
rect 25056 31198 25176 31226
rect 24768 30660 24820 30666
rect 24768 30602 24820 30608
rect 24860 30252 24912 30258
rect 24860 30194 24912 30200
rect 24872 29850 24900 30194
rect 24952 30048 25004 30054
rect 24952 29990 25004 29996
rect 24860 29844 24912 29850
rect 24860 29786 24912 29792
rect 24964 29170 24992 29990
rect 25044 29640 25096 29646
rect 25044 29582 25096 29588
rect 24768 29164 24820 29170
rect 24768 29106 24820 29112
rect 24952 29164 25004 29170
rect 24952 29106 25004 29112
rect 24676 28688 24728 28694
rect 24676 28630 24728 28636
rect 24688 28558 24716 28630
rect 24676 28552 24728 28558
rect 24676 28494 24728 28500
rect 24780 28540 24808 29106
rect 24860 28552 24912 28558
rect 24780 28512 24860 28540
rect 24584 28484 24636 28490
rect 24584 28426 24636 28432
rect 24400 28416 24452 28422
rect 24400 28358 24452 28364
rect 24412 28150 24440 28358
rect 24400 28144 24452 28150
rect 24400 28086 24452 28092
rect 24596 27402 24624 28426
rect 24688 27470 24716 28494
rect 24780 28014 24808 28512
rect 24860 28494 24912 28500
rect 25056 28082 25084 29582
rect 25044 28076 25096 28082
rect 25044 28018 25096 28024
rect 24768 28008 24820 28014
rect 24768 27950 24820 27956
rect 24676 27464 24728 27470
rect 24676 27406 24728 27412
rect 24584 27396 24636 27402
rect 24584 27338 24636 27344
rect 24596 25906 24624 27338
rect 24688 26994 24716 27406
rect 24676 26988 24728 26994
rect 24676 26930 24728 26936
rect 24584 25900 24636 25906
rect 24584 25842 24636 25848
rect 24492 25356 24544 25362
rect 24492 25298 24544 25304
rect 24504 24206 24532 25298
rect 24676 24608 24728 24614
rect 24676 24550 24728 24556
rect 24688 24206 24716 24550
rect 24492 24200 24544 24206
rect 24492 24142 24544 24148
rect 24676 24200 24728 24206
rect 24676 24142 24728 24148
rect 24308 24064 24360 24070
rect 24308 24006 24360 24012
rect 24320 23730 24348 24006
rect 24308 23724 24360 23730
rect 24308 23666 24360 23672
rect 24400 23520 24452 23526
rect 24400 23462 24452 23468
rect 24412 22778 24440 23462
rect 24400 22772 24452 22778
rect 24400 22714 24452 22720
rect 24504 22710 24532 24142
rect 24674 23760 24730 23769
rect 24674 23695 24676 23704
rect 24728 23695 24730 23704
rect 24676 23666 24728 23672
rect 24584 23044 24636 23050
rect 24584 22986 24636 22992
rect 24492 22704 24544 22710
rect 24492 22646 24544 22652
rect 24228 22066 24440 22094
rect 24124 21548 24176 21554
rect 24044 21508 24124 21536
rect 24044 14822 24072 21508
rect 24124 21490 24176 21496
rect 24124 21004 24176 21010
rect 24124 20946 24176 20952
rect 24136 18970 24164 20946
rect 24306 20496 24362 20505
rect 24306 20431 24362 20440
rect 24320 20262 24348 20431
rect 24308 20256 24360 20262
rect 24308 20198 24360 20204
rect 24124 18964 24176 18970
rect 24124 18906 24176 18912
rect 24136 16538 24164 18906
rect 24216 18080 24268 18086
rect 24216 18022 24268 18028
rect 24228 17678 24256 18022
rect 24216 17672 24268 17678
rect 24216 17614 24268 17620
rect 24308 17196 24360 17202
rect 24308 17138 24360 17144
rect 24136 16510 24256 16538
rect 24124 16244 24176 16250
rect 24124 16186 24176 16192
rect 24136 16114 24164 16186
rect 24124 16108 24176 16114
rect 24124 16050 24176 16056
rect 24228 15638 24256 16510
rect 24216 15632 24268 15638
rect 24216 15574 24268 15580
rect 24320 15450 24348 17138
rect 24412 16454 24440 22066
rect 24492 20324 24544 20330
rect 24492 20266 24544 20272
rect 24504 20233 24532 20266
rect 24490 20224 24546 20233
rect 24490 20159 24546 20168
rect 24492 17332 24544 17338
rect 24492 17274 24544 17280
rect 24400 16448 24452 16454
rect 24400 16390 24452 16396
rect 24400 16108 24452 16114
rect 24400 16050 24452 16056
rect 24412 15502 24440 16050
rect 24136 15422 24348 15450
rect 24400 15496 24452 15502
rect 24400 15438 24452 15444
rect 24032 14816 24084 14822
rect 24032 14758 24084 14764
rect 24044 11642 24072 14758
rect 24136 11830 24164 15422
rect 24412 15026 24440 15438
rect 24400 15020 24452 15026
rect 24400 14962 24452 14968
rect 24400 14272 24452 14278
rect 24400 14214 24452 14220
rect 24412 13938 24440 14214
rect 24308 13932 24360 13938
rect 24308 13874 24360 13880
rect 24400 13932 24452 13938
rect 24400 13874 24452 13880
rect 24216 13524 24268 13530
rect 24216 13466 24268 13472
rect 24228 13258 24256 13466
rect 24216 13252 24268 13258
rect 24216 13194 24268 13200
rect 24320 12986 24348 13874
rect 24504 13190 24532 17274
rect 24596 16250 24624 22986
rect 24780 22094 24808 27950
rect 25056 27062 25084 28018
rect 25044 27056 25096 27062
rect 25044 26998 25096 27004
rect 24860 26920 24912 26926
rect 24860 26862 24912 26868
rect 24872 26586 24900 26862
rect 25056 26586 25084 26998
rect 24860 26580 24912 26586
rect 24860 26522 24912 26528
rect 25044 26580 25096 26586
rect 25044 26522 25096 26528
rect 24952 25900 25004 25906
rect 24952 25842 25004 25848
rect 24860 25696 24912 25702
rect 24860 25638 24912 25644
rect 24872 24449 24900 25638
rect 24858 24440 24914 24449
rect 24858 24375 24914 24384
rect 24964 22982 24992 25842
rect 25056 24818 25084 26522
rect 25148 26314 25176 31198
rect 25596 30252 25648 30258
rect 25596 30194 25648 30200
rect 25608 29102 25636 30194
rect 25596 29096 25648 29102
rect 25596 29038 25648 29044
rect 25780 28620 25832 28626
rect 25780 28562 25832 28568
rect 25228 28552 25280 28558
rect 25228 28494 25280 28500
rect 25240 28422 25268 28494
rect 25228 28416 25280 28422
rect 25228 28358 25280 28364
rect 25792 28218 25820 28562
rect 25780 28212 25832 28218
rect 25780 28154 25832 28160
rect 25228 27328 25280 27334
rect 25228 27270 25280 27276
rect 25240 26858 25268 27270
rect 25228 26852 25280 26858
rect 25228 26794 25280 26800
rect 25136 26308 25188 26314
rect 25136 26250 25188 26256
rect 25780 26240 25832 26246
rect 25780 26182 25832 26188
rect 25596 25696 25648 25702
rect 25596 25638 25648 25644
rect 25608 25498 25636 25638
rect 25792 25498 25820 26182
rect 25596 25492 25648 25498
rect 25596 25434 25648 25440
rect 25780 25492 25832 25498
rect 25780 25434 25832 25440
rect 25688 25288 25740 25294
rect 25688 25230 25740 25236
rect 25596 25152 25648 25158
rect 25596 25094 25648 25100
rect 25044 24812 25096 24818
rect 25044 24754 25096 24760
rect 25228 24812 25280 24818
rect 25228 24754 25280 24760
rect 25056 24206 25084 24754
rect 25044 24200 25096 24206
rect 25044 24142 25096 24148
rect 24952 22976 25004 22982
rect 24952 22918 25004 22924
rect 24860 22636 24912 22642
rect 24860 22578 24912 22584
rect 24872 22409 24900 22578
rect 24952 22432 25004 22438
rect 24858 22400 24914 22409
rect 24952 22374 25004 22380
rect 24858 22335 24914 22344
rect 24688 22066 24808 22094
rect 24688 17270 24716 22066
rect 24964 21962 24992 22374
rect 25056 22234 25084 24142
rect 25136 24064 25188 24070
rect 25136 24006 25188 24012
rect 25148 23798 25176 24006
rect 25240 23866 25268 24754
rect 25320 24336 25372 24342
rect 25320 24278 25372 24284
rect 25332 24070 25360 24278
rect 25608 24138 25636 25094
rect 25596 24132 25648 24138
rect 25596 24074 25648 24080
rect 25320 24064 25372 24070
rect 25320 24006 25372 24012
rect 25228 23860 25280 23866
rect 25228 23802 25280 23808
rect 25136 23792 25188 23798
rect 25136 23734 25188 23740
rect 25228 23724 25280 23730
rect 25228 23666 25280 23672
rect 25136 22636 25188 22642
rect 25136 22578 25188 22584
rect 25044 22228 25096 22234
rect 25044 22170 25096 22176
rect 24952 21956 25004 21962
rect 24952 21898 25004 21904
rect 24952 21684 25004 21690
rect 24952 21626 25004 21632
rect 24860 20936 24912 20942
rect 24860 20878 24912 20884
rect 24768 18760 24820 18766
rect 24768 18702 24820 18708
rect 24780 18426 24808 18702
rect 24768 18420 24820 18426
rect 24768 18362 24820 18368
rect 24676 17264 24728 17270
rect 24676 17206 24728 17212
rect 24584 16244 24636 16250
rect 24584 16186 24636 16192
rect 24596 15502 24624 16186
rect 24584 15496 24636 15502
rect 24584 15438 24636 15444
rect 24584 15360 24636 15366
rect 24584 15302 24636 15308
rect 24596 13802 24624 15302
rect 24872 15178 24900 20878
rect 24964 20806 24992 21626
rect 25056 21554 25084 22170
rect 25044 21548 25096 21554
rect 25044 21490 25096 21496
rect 24952 20800 25004 20806
rect 24952 20742 25004 20748
rect 25148 20602 25176 22578
rect 25136 20596 25188 20602
rect 25136 20538 25188 20544
rect 24952 20460 25004 20466
rect 24952 20402 25004 20408
rect 25136 20460 25188 20466
rect 25136 20402 25188 20408
rect 24964 18766 24992 20402
rect 25148 19378 25176 20402
rect 25136 19372 25188 19378
rect 25136 19314 25188 19320
rect 25044 18896 25096 18902
rect 25044 18838 25096 18844
rect 24952 18760 25004 18766
rect 24952 18702 25004 18708
rect 25056 18086 25084 18838
rect 25136 18216 25188 18222
rect 25136 18158 25188 18164
rect 25044 18080 25096 18086
rect 25044 18022 25096 18028
rect 25148 17882 25176 18158
rect 25136 17876 25188 17882
rect 25136 17818 25188 17824
rect 24952 16652 25004 16658
rect 24952 16594 25004 16600
rect 24964 16114 24992 16594
rect 25136 16448 25188 16454
rect 25136 16390 25188 16396
rect 24952 16108 25004 16114
rect 24952 16050 25004 16056
rect 24964 15570 24992 16050
rect 24952 15564 25004 15570
rect 24952 15506 25004 15512
rect 24688 15150 24900 15178
rect 25148 15162 25176 16390
rect 25136 15156 25188 15162
rect 24584 13796 24636 13802
rect 24584 13738 24636 13744
rect 24596 13258 24624 13738
rect 24584 13252 24636 13258
rect 24584 13194 24636 13200
rect 24400 13184 24452 13190
rect 24400 13126 24452 13132
rect 24492 13184 24544 13190
rect 24492 13126 24544 13132
rect 24308 12980 24360 12986
rect 24308 12922 24360 12928
rect 24124 11824 24176 11830
rect 24124 11766 24176 11772
rect 24044 11614 24256 11642
rect 24032 11552 24084 11558
rect 24032 11494 24084 11500
rect 24044 11354 24072 11494
rect 24032 11348 24084 11354
rect 24032 11290 24084 11296
rect 24228 10742 24256 11614
rect 24216 10736 24268 10742
rect 24216 10678 24268 10684
rect 24214 10296 24270 10305
rect 24214 10231 24270 10240
rect 24032 9920 24084 9926
rect 24032 9862 24084 9868
rect 24044 9654 24072 9862
rect 24032 9648 24084 9654
rect 24032 9590 24084 9596
rect 24044 9042 24072 9590
rect 24032 9036 24084 9042
rect 24032 8978 24084 8984
rect 24228 8566 24256 10231
rect 24320 10062 24348 12922
rect 24412 12646 24440 13126
rect 24400 12640 24452 12646
rect 24400 12582 24452 12588
rect 24504 11762 24532 13126
rect 24584 12640 24636 12646
rect 24584 12582 24636 12588
rect 24596 12442 24624 12582
rect 24584 12436 24636 12442
rect 24584 12378 24636 12384
rect 24492 11756 24544 11762
rect 24492 11698 24544 11704
rect 24400 11688 24452 11694
rect 24400 11630 24452 11636
rect 24308 10056 24360 10062
rect 24308 9998 24360 10004
rect 24412 9058 24440 11630
rect 24596 11082 24624 12378
rect 24584 11076 24636 11082
rect 24584 11018 24636 11024
rect 24492 10736 24544 10742
rect 24492 10678 24544 10684
rect 24504 10146 24532 10678
rect 24596 10674 24624 11018
rect 24584 10668 24636 10674
rect 24584 10610 24636 10616
rect 24596 10266 24624 10610
rect 24584 10260 24636 10266
rect 24584 10202 24636 10208
rect 24504 10118 24624 10146
rect 24596 9489 24624 10118
rect 24582 9480 24638 9489
rect 24582 9415 24638 9424
rect 24492 9376 24544 9382
rect 24492 9318 24544 9324
rect 24584 9376 24636 9382
rect 24584 9318 24636 9324
rect 24504 9178 24532 9318
rect 24492 9172 24544 9178
rect 24492 9114 24544 9120
rect 24308 9036 24360 9042
rect 24412 9030 24532 9058
rect 24308 8978 24360 8984
rect 24320 8838 24348 8978
rect 24400 8968 24452 8974
rect 24400 8910 24452 8916
rect 24412 8838 24440 8910
rect 24308 8832 24360 8838
rect 24308 8774 24360 8780
rect 24400 8832 24452 8838
rect 24400 8774 24452 8780
rect 24400 8628 24452 8634
rect 24400 8570 24452 8576
rect 24216 8560 24268 8566
rect 24412 8537 24440 8570
rect 24216 8502 24268 8508
rect 24398 8528 24454 8537
rect 24398 8463 24454 8472
rect 24400 7880 24452 7886
rect 24400 7822 24452 7828
rect 24124 6384 24176 6390
rect 24124 6326 24176 6332
rect 24032 6316 24084 6322
rect 24032 6258 24084 6264
rect 24044 5778 24072 6258
rect 24032 5772 24084 5778
rect 24032 5714 24084 5720
rect 24044 5098 24072 5714
rect 24136 5302 24164 6326
rect 24216 6248 24268 6254
rect 24216 6190 24268 6196
rect 24228 5846 24256 6190
rect 24216 5840 24268 5846
rect 24216 5782 24268 5788
rect 24228 5302 24256 5782
rect 24412 5778 24440 7822
rect 24504 6322 24532 9030
rect 24596 8838 24624 9318
rect 24584 8832 24636 8838
rect 24584 8774 24636 8780
rect 24584 8424 24636 8430
rect 24584 8366 24636 8372
rect 24596 7954 24624 8366
rect 24584 7948 24636 7954
rect 24584 7890 24636 7896
rect 24492 6316 24544 6322
rect 24492 6258 24544 6264
rect 24400 5772 24452 5778
rect 24400 5714 24452 5720
rect 24412 5642 24440 5714
rect 24400 5636 24452 5642
rect 24400 5578 24452 5584
rect 24124 5296 24176 5302
rect 24124 5238 24176 5244
rect 24216 5296 24268 5302
rect 24216 5238 24268 5244
rect 24032 5092 24084 5098
rect 24032 5034 24084 5040
rect 24688 2774 24716 15150
rect 25136 15098 25188 15104
rect 25240 14958 25268 23666
rect 25412 22704 25464 22710
rect 25412 22646 25464 22652
rect 25424 22234 25452 22646
rect 25700 22642 25728 25230
rect 25780 23792 25832 23798
rect 25780 23734 25832 23740
rect 25792 23633 25820 23734
rect 25778 23624 25834 23633
rect 25778 23559 25834 23568
rect 25688 22636 25740 22642
rect 25608 22596 25688 22624
rect 25412 22228 25464 22234
rect 25412 22170 25464 22176
rect 25320 21548 25372 21554
rect 25320 21490 25372 21496
rect 25332 21078 25360 21490
rect 25320 21072 25372 21078
rect 25320 21014 25372 21020
rect 25424 20942 25452 22170
rect 25608 22080 25636 22596
rect 25688 22578 25740 22584
rect 25688 22092 25740 22098
rect 25608 22052 25688 22080
rect 25608 20942 25636 22052
rect 25688 22034 25740 22040
rect 25688 21888 25740 21894
rect 25688 21830 25740 21836
rect 25412 20936 25464 20942
rect 25412 20878 25464 20884
rect 25596 20936 25648 20942
rect 25596 20878 25648 20884
rect 25320 20596 25372 20602
rect 25320 20538 25372 20544
rect 25332 20369 25360 20538
rect 25700 20466 25728 21830
rect 25688 20460 25740 20466
rect 25688 20402 25740 20408
rect 25318 20360 25374 20369
rect 25318 20295 25374 20304
rect 25884 19938 25912 47534
rect 25976 47462 26004 47534
rect 25964 47456 26016 47462
rect 25964 47398 26016 47404
rect 26068 47258 26096 47602
rect 26160 47462 26188 47738
rect 26148 47456 26200 47462
rect 26148 47398 26200 47404
rect 26056 47252 26108 47258
rect 26056 47194 26108 47200
rect 26252 47054 26280 51326
rect 26422 51200 26478 51326
rect 27066 51354 27122 52000
rect 27710 51354 27766 52000
rect 27066 51326 27568 51354
rect 27066 51200 27122 51326
rect 27540 49586 27568 51326
rect 27710 51326 27936 51354
rect 27710 51200 27766 51326
rect 27540 49558 27660 49586
rect 27632 49298 27660 49558
rect 27620 49292 27672 49298
rect 27620 49234 27672 49240
rect 26424 49224 26476 49230
rect 26424 49166 26476 49172
rect 26976 49224 27028 49230
rect 26976 49166 27028 49172
rect 26436 48754 26464 49166
rect 26424 48748 26476 48754
rect 26424 48690 26476 48696
rect 26516 48680 26568 48686
rect 26516 48622 26568 48628
rect 26528 48142 26556 48622
rect 26516 48136 26568 48142
rect 26516 48078 26568 48084
rect 26988 47258 27016 49166
rect 27160 49156 27212 49162
rect 27160 49098 27212 49104
rect 27172 47802 27200 49098
rect 27908 48686 27936 51326
rect 28354 51200 28410 52000
rect 28998 51200 29054 52000
rect 29642 51354 29698 52000
rect 29642 51326 29960 51354
rect 29642 51200 29698 51326
rect 27620 48680 27672 48686
rect 27620 48622 27672 48628
rect 27896 48680 27948 48686
rect 27896 48622 27948 48628
rect 27528 48544 27580 48550
rect 27528 48486 27580 48492
rect 27160 47796 27212 47802
rect 27160 47738 27212 47744
rect 27252 47660 27304 47666
rect 27252 47602 27304 47608
rect 27264 47462 27292 47602
rect 27252 47456 27304 47462
rect 27252 47398 27304 47404
rect 26976 47252 27028 47258
rect 26976 47194 27028 47200
rect 26240 47048 26292 47054
rect 26240 46990 26292 46996
rect 26148 44192 26200 44198
rect 26148 44134 26200 44140
rect 25964 37868 26016 37874
rect 25964 37810 26016 37816
rect 25976 37466 26004 37810
rect 26056 37800 26108 37806
rect 26056 37742 26108 37748
rect 25964 37460 26016 37466
rect 25964 37402 26016 37408
rect 25964 34400 26016 34406
rect 25964 34342 26016 34348
rect 25976 33998 26004 34342
rect 25964 33992 26016 33998
rect 25964 33934 26016 33940
rect 26068 33930 26096 37742
rect 26056 33924 26108 33930
rect 26056 33866 26108 33872
rect 25964 33856 26016 33862
rect 25964 33798 26016 33804
rect 25976 27606 26004 33798
rect 26068 33658 26096 33866
rect 26056 33652 26108 33658
rect 26056 33594 26108 33600
rect 26160 32910 26188 44134
rect 26332 39364 26384 39370
rect 26332 39306 26384 39312
rect 26344 38010 26372 39306
rect 26700 38276 26752 38282
rect 26700 38218 26752 38224
rect 26332 38004 26384 38010
rect 26332 37946 26384 37952
rect 26712 37466 26740 38218
rect 26700 37460 26752 37466
rect 26700 37402 26752 37408
rect 27252 37324 27304 37330
rect 27252 37266 27304 37272
rect 26516 37256 26568 37262
rect 26516 37198 26568 37204
rect 26240 36780 26292 36786
rect 26240 36722 26292 36728
rect 26252 35698 26280 36722
rect 26240 35692 26292 35698
rect 26240 35634 26292 35640
rect 26252 33930 26280 35634
rect 26240 33924 26292 33930
rect 26240 33866 26292 33872
rect 26148 32904 26200 32910
rect 26148 32846 26200 32852
rect 26252 32298 26280 33866
rect 26424 33516 26476 33522
rect 26424 33458 26476 33464
rect 26436 32434 26464 33458
rect 26424 32428 26476 32434
rect 26424 32370 26476 32376
rect 26240 32292 26292 32298
rect 26240 32234 26292 32240
rect 26436 30258 26464 32370
rect 26424 30252 26476 30258
rect 26424 30194 26476 30200
rect 26424 28756 26476 28762
rect 26424 28698 26476 28704
rect 26436 28626 26464 28698
rect 26424 28620 26476 28626
rect 26424 28562 26476 28568
rect 26332 28552 26384 28558
rect 26332 28494 26384 28500
rect 25964 27600 26016 27606
rect 25964 27542 26016 27548
rect 26056 27600 26108 27606
rect 26056 27542 26108 27548
rect 25976 26994 26004 27542
rect 25964 26988 26016 26994
rect 25964 26930 26016 26936
rect 26068 26586 26096 27542
rect 26148 27464 26200 27470
rect 26148 27406 26200 27412
rect 26160 27130 26188 27406
rect 26148 27124 26200 27130
rect 26148 27066 26200 27072
rect 26240 26920 26292 26926
rect 26240 26862 26292 26868
rect 26252 26790 26280 26862
rect 26240 26784 26292 26790
rect 26240 26726 26292 26732
rect 26056 26580 26108 26586
rect 26056 26522 26108 26528
rect 26068 25294 26096 26522
rect 26148 26512 26200 26518
rect 26200 26460 26280 26466
rect 26148 26454 26280 26460
rect 26160 26438 26280 26454
rect 26252 26314 26280 26438
rect 26148 26308 26200 26314
rect 26148 26250 26200 26256
rect 26240 26308 26292 26314
rect 26240 26250 26292 26256
rect 26056 25288 26108 25294
rect 26056 25230 26108 25236
rect 26056 23724 26108 23730
rect 26056 23666 26108 23672
rect 26068 23633 26096 23666
rect 26054 23624 26110 23633
rect 26054 23559 26110 23568
rect 26160 21128 26188 26250
rect 26240 25152 26292 25158
rect 26240 25094 26292 25100
rect 26252 23866 26280 25094
rect 26240 23860 26292 23866
rect 26240 23802 26292 23808
rect 26240 21344 26292 21350
rect 26240 21286 26292 21292
rect 26068 21100 26188 21128
rect 25884 19910 26004 19938
rect 25780 19780 25832 19786
rect 25780 19722 25832 19728
rect 25792 19553 25820 19722
rect 25778 19544 25834 19553
rect 25778 19479 25834 19488
rect 25596 19304 25648 19310
rect 25596 19246 25648 19252
rect 25320 18760 25372 18766
rect 25320 18702 25372 18708
rect 25332 18290 25360 18702
rect 25412 18624 25464 18630
rect 25412 18566 25464 18572
rect 25320 18284 25372 18290
rect 25320 18226 25372 18232
rect 25332 17490 25360 18226
rect 25424 17678 25452 18566
rect 25608 18358 25636 19246
rect 25688 19168 25740 19174
rect 25688 19110 25740 19116
rect 25700 18766 25728 19110
rect 25792 18970 25820 19479
rect 25780 18964 25832 18970
rect 25780 18906 25832 18912
rect 25688 18760 25740 18766
rect 25688 18702 25740 18708
rect 25596 18352 25648 18358
rect 25596 18294 25648 18300
rect 25780 18216 25832 18222
rect 25780 18158 25832 18164
rect 25504 18080 25556 18086
rect 25504 18022 25556 18028
rect 25516 17678 25544 18022
rect 25412 17672 25464 17678
rect 25412 17614 25464 17620
rect 25504 17672 25556 17678
rect 25504 17614 25556 17620
rect 25688 17604 25740 17610
rect 25688 17546 25740 17552
rect 25332 17462 25452 17490
rect 25424 17202 25452 17462
rect 25412 17196 25464 17202
rect 25412 17138 25464 17144
rect 25228 14952 25280 14958
rect 25228 14894 25280 14900
rect 25320 13932 25372 13938
rect 25320 13874 25372 13880
rect 24952 13728 25004 13734
rect 24952 13670 25004 13676
rect 24768 13320 24820 13326
rect 24768 13262 24820 13268
rect 24780 8634 24808 13262
rect 24860 12776 24912 12782
rect 24860 12718 24912 12724
rect 24872 11082 24900 12718
rect 24964 12714 24992 13670
rect 24952 12708 25004 12714
rect 24952 12650 25004 12656
rect 24952 12232 25004 12238
rect 24952 12174 25004 12180
rect 24964 11898 24992 12174
rect 25332 12170 25360 13874
rect 25424 12646 25452 17138
rect 25596 16992 25648 16998
rect 25596 16934 25648 16940
rect 25608 16658 25636 16934
rect 25596 16652 25648 16658
rect 25596 16594 25648 16600
rect 25700 16590 25728 17546
rect 25792 17542 25820 18158
rect 25976 17678 26004 19910
rect 26068 17814 26096 21100
rect 26148 20936 26200 20942
rect 26148 20878 26200 20884
rect 26160 20534 26188 20878
rect 26252 20874 26280 21286
rect 26240 20868 26292 20874
rect 26240 20810 26292 20816
rect 26148 20528 26200 20534
rect 26148 20470 26200 20476
rect 26148 19848 26200 19854
rect 26148 19790 26200 19796
rect 26160 19310 26188 19790
rect 26252 19378 26280 20810
rect 26240 19372 26292 19378
rect 26240 19314 26292 19320
rect 26148 19304 26200 19310
rect 26148 19246 26200 19252
rect 26160 18204 26188 19246
rect 26240 18216 26292 18222
rect 26160 18176 26240 18204
rect 26056 17808 26108 17814
rect 26056 17750 26108 17756
rect 25964 17672 26016 17678
rect 25964 17614 26016 17620
rect 25780 17536 25832 17542
rect 25780 17478 25832 17484
rect 25792 17202 25820 17478
rect 25780 17196 25832 17202
rect 25780 17138 25832 17144
rect 25976 16726 26004 17614
rect 25964 16720 26016 16726
rect 25964 16662 26016 16668
rect 25688 16584 25740 16590
rect 25688 16526 25740 16532
rect 25872 16584 25924 16590
rect 25872 16526 25924 16532
rect 25780 15564 25832 15570
rect 25780 15506 25832 15512
rect 25792 15366 25820 15506
rect 25780 15360 25832 15366
rect 25780 15302 25832 15308
rect 25780 15020 25832 15026
rect 25780 14962 25832 14968
rect 25792 14414 25820 14962
rect 25884 14618 25912 16526
rect 26160 15570 26188 18176
rect 26240 18158 26292 18164
rect 26240 17876 26292 17882
rect 26240 17818 26292 17824
rect 26252 17270 26280 17818
rect 26240 17264 26292 17270
rect 26240 17206 26292 17212
rect 26252 16794 26280 17206
rect 26240 16788 26292 16794
rect 26240 16730 26292 16736
rect 26240 16584 26292 16590
rect 26240 16526 26292 16532
rect 26148 15564 26200 15570
rect 26148 15506 26200 15512
rect 26252 15502 26280 16526
rect 26240 15496 26292 15502
rect 26240 15438 26292 15444
rect 25964 15360 26016 15366
rect 25964 15302 26016 15308
rect 25872 14612 25924 14618
rect 25872 14554 25924 14560
rect 25976 14414 26004 15302
rect 26240 14952 26292 14958
rect 26240 14894 26292 14900
rect 26148 14816 26200 14822
rect 26148 14758 26200 14764
rect 26160 14482 26188 14758
rect 26148 14476 26200 14482
rect 26148 14418 26200 14424
rect 25780 14408 25832 14414
rect 25780 14350 25832 14356
rect 25964 14408 26016 14414
rect 25964 14350 26016 14356
rect 25792 13938 25820 14350
rect 25976 14006 26004 14350
rect 25964 14000 26016 14006
rect 25964 13942 26016 13948
rect 25780 13932 25832 13938
rect 25780 13874 25832 13880
rect 26160 13734 26188 14418
rect 26252 14346 26280 14894
rect 26240 14340 26292 14346
rect 26240 14282 26292 14288
rect 26252 13870 26280 14282
rect 26240 13864 26292 13870
rect 26240 13806 26292 13812
rect 25504 13728 25556 13734
rect 25504 13670 25556 13676
rect 26148 13728 26200 13734
rect 26148 13670 26200 13676
rect 25516 12918 25544 13670
rect 26160 13394 26188 13670
rect 26148 13388 26200 13394
rect 26148 13330 26200 13336
rect 26252 13326 26280 13806
rect 26240 13320 26292 13326
rect 26240 13262 26292 13268
rect 25504 12912 25556 12918
rect 25504 12854 25556 12860
rect 26252 12850 26280 13262
rect 26240 12844 26292 12850
rect 26240 12786 26292 12792
rect 25688 12776 25740 12782
rect 25688 12718 25740 12724
rect 25412 12640 25464 12646
rect 25412 12582 25464 12588
rect 25700 12434 25728 12718
rect 26252 12442 26280 12786
rect 25516 12406 25728 12434
rect 26240 12436 26292 12442
rect 25516 12238 25544 12406
rect 26240 12378 26292 12384
rect 25504 12232 25556 12238
rect 25504 12174 25556 12180
rect 25780 12232 25832 12238
rect 25780 12174 25832 12180
rect 25320 12164 25372 12170
rect 25320 12106 25372 12112
rect 24952 11892 25004 11898
rect 24952 11834 25004 11840
rect 24860 11076 24912 11082
rect 24860 11018 24912 11024
rect 24872 10810 24900 11018
rect 24860 10804 24912 10810
rect 24860 10746 24912 10752
rect 24964 10554 24992 11834
rect 25516 11558 25544 12174
rect 25688 12096 25740 12102
rect 25688 12038 25740 12044
rect 25700 11762 25728 12038
rect 25688 11756 25740 11762
rect 25688 11698 25740 11704
rect 25504 11552 25556 11558
rect 25504 11494 25556 11500
rect 25044 11008 25096 11014
rect 25044 10950 25096 10956
rect 25056 10674 25084 10950
rect 25688 10804 25740 10810
rect 25792 10792 25820 12174
rect 25964 11688 26016 11694
rect 25964 11630 26016 11636
rect 25872 11552 25924 11558
rect 25872 11494 25924 11500
rect 25740 10764 25820 10792
rect 25688 10746 25740 10752
rect 25044 10668 25096 10674
rect 25044 10610 25096 10616
rect 25136 10668 25188 10674
rect 25136 10610 25188 10616
rect 25412 10668 25464 10674
rect 25412 10610 25464 10616
rect 24964 10526 25084 10554
rect 24952 10260 25004 10266
rect 24952 10202 25004 10208
rect 24860 8900 24912 8906
rect 24860 8842 24912 8848
rect 24768 8628 24820 8634
rect 24768 8570 24820 8576
rect 24872 8566 24900 8842
rect 24860 8560 24912 8566
rect 24860 8502 24912 8508
rect 24872 7546 24900 8502
rect 24964 8362 24992 10202
rect 25056 9625 25084 10526
rect 25042 9616 25098 9625
rect 25042 9551 25098 9560
rect 25056 9110 25084 9551
rect 25148 9178 25176 10610
rect 25424 10130 25452 10610
rect 25504 10464 25556 10470
rect 25504 10406 25556 10412
rect 25412 10124 25464 10130
rect 25412 10066 25464 10072
rect 25228 9988 25280 9994
rect 25228 9930 25280 9936
rect 25240 9722 25268 9930
rect 25228 9716 25280 9722
rect 25228 9658 25280 9664
rect 25226 9480 25282 9489
rect 25226 9415 25282 9424
rect 25136 9172 25188 9178
rect 25136 9114 25188 9120
rect 25240 9110 25268 9415
rect 25044 9104 25096 9110
rect 25044 9046 25096 9052
rect 25228 9104 25280 9110
rect 25228 9046 25280 9052
rect 25044 8832 25096 8838
rect 25044 8774 25096 8780
rect 25228 8832 25280 8838
rect 25228 8774 25280 8780
rect 25056 8537 25084 8774
rect 25042 8528 25098 8537
rect 25042 8463 25098 8472
rect 25136 8492 25188 8498
rect 25136 8434 25188 8440
rect 25148 8401 25176 8434
rect 25134 8392 25190 8401
rect 24952 8356 25004 8362
rect 25134 8327 25190 8336
rect 24952 8298 25004 8304
rect 24860 7540 24912 7546
rect 24860 7482 24912 7488
rect 25240 7410 25268 8774
rect 25320 8424 25372 8430
rect 25372 8384 25452 8412
rect 25320 8366 25372 8372
rect 25424 8294 25452 8384
rect 25412 8288 25464 8294
rect 25412 8230 25464 8236
rect 25516 7818 25544 10406
rect 25596 10260 25648 10266
rect 25596 10202 25648 10208
rect 25608 9994 25636 10202
rect 25700 10062 25728 10746
rect 25688 10056 25740 10062
rect 25688 9998 25740 10004
rect 25596 9988 25648 9994
rect 25596 9930 25648 9936
rect 25884 9926 25912 11494
rect 25976 11082 26004 11630
rect 26056 11144 26108 11150
rect 26056 11086 26108 11092
rect 25964 11076 26016 11082
rect 25964 11018 26016 11024
rect 25964 10736 26016 10742
rect 25964 10678 26016 10684
rect 25872 9920 25924 9926
rect 25872 9862 25924 9868
rect 25780 9716 25832 9722
rect 25780 9658 25832 9664
rect 25792 8974 25820 9658
rect 25884 9586 25912 9862
rect 25976 9722 26004 10678
rect 25964 9716 26016 9722
rect 25964 9658 26016 9664
rect 25872 9580 25924 9586
rect 25872 9522 25924 9528
rect 25872 9172 25924 9178
rect 25872 9114 25924 9120
rect 25884 8974 25912 9114
rect 25780 8968 25832 8974
rect 25686 8936 25742 8945
rect 25780 8910 25832 8916
rect 25872 8968 25924 8974
rect 25872 8910 25924 8916
rect 25686 8871 25688 8880
rect 25740 8871 25742 8880
rect 25688 8842 25740 8848
rect 25778 8528 25834 8537
rect 25778 8463 25834 8472
rect 25504 7812 25556 7818
rect 25504 7754 25556 7760
rect 25228 7404 25280 7410
rect 25228 7346 25280 7352
rect 25792 5846 25820 8463
rect 25976 8294 26004 9658
rect 26068 9586 26096 11086
rect 26344 10826 26372 28494
rect 26422 26616 26478 26625
rect 26422 26551 26478 26560
rect 26436 26518 26464 26551
rect 26424 26512 26476 26518
rect 26424 26454 26476 26460
rect 26424 25356 26476 25362
rect 26424 25298 26476 25304
rect 26436 23866 26464 25298
rect 26424 23860 26476 23866
rect 26424 23802 26476 23808
rect 26422 23624 26478 23633
rect 26422 23559 26478 23568
rect 26436 20942 26464 23559
rect 26424 20936 26476 20942
rect 26424 20878 26476 20884
rect 26424 20052 26476 20058
rect 26424 19994 26476 20000
rect 26436 19718 26464 19994
rect 26424 19712 26476 19718
rect 26424 19654 26476 19660
rect 26424 19372 26476 19378
rect 26424 19314 26476 19320
rect 26436 18358 26464 19314
rect 26424 18352 26476 18358
rect 26424 18294 26476 18300
rect 26436 17610 26464 18294
rect 26424 17604 26476 17610
rect 26424 17546 26476 17552
rect 26424 17128 26476 17134
rect 26424 17070 26476 17076
rect 26436 15366 26464 17070
rect 26424 15360 26476 15366
rect 26422 15328 26424 15337
rect 26476 15328 26478 15337
rect 26422 15263 26478 15272
rect 26424 14816 26476 14822
rect 26424 14758 26476 14764
rect 26436 14414 26464 14758
rect 26424 14408 26476 14414
rect 26424 14350 26476 14356
rect 26528 12434 26556 37198
rect 26700 37120 26752 37126
rect 26700 37062 26752 37068
rect 26792 37120 26844 37126
rect 26792 37062 26844 37068
rect 26608 36168 26660 36174
rect 26608 36110 26660 36116
rect 26620 31754 26648 36110
rect 26712 35816 26740 37062
rect 26804 36854 26832 37062
rect 26792 36848 26844 36854
rect 26792 36790 26844 36796
rect 27264 36242 27292 37266
rect 27344 37256 27396 37262
rect 27344 37198 27396 37204
rect 27356 36922 27384 37198
rect 27344 36916 27396 36922
rect 27344 36858 27396 36864
rect 27252 36236 27304 36242
rect 27252 36178 27304 36184
rect 27344 36032 27396 36038
rect 27344 35974 27396 35980
rect 27068 35828 27120 35834
rect 26712 35788 27068 35816
rect 27068 35770 27120 35776
rect 27356 35698 27384 35974
rect 27344 35692 27396 35698
rect 27344 35634 27396 35640
rect 27252 33856 27304 33862
rect 27252 33798 27304 33804
rect 26976 33516 27028 33522
rect 26976 33458 27028 33464
rect 27068 33516 27120 33522
rect 27068 33458 27120 33464
rect 26988 32434 27016 33458
rect 27080 33114 27108 33458
rect 27068 33108 27120 33114
rect 27068 33050 27120 33056
rect 27264 32910 27292 33798
rect 27344 32972 27396 32978
rect 27344 32914 27396 32920
rect 27252 32904 27304 32910
rect 27252 32846 27304 32852
rect 26976 32428 27028 32434
rect 26976 32370 27028 32376
rect 27356 31958 27384 32914
rect 27436 32428 27488 32434
rect 27436 32370 27488 32376
rect 27448 32026 27476 32370
rect 27436 32020 27488 32026
rect 27436 31962 27488 31968
rect 27344 31952 27396 31958
rect 27344 31894 27396 31900
rect 27344 31816 27396 31822
rect 27344 31758 27396 31764
rect 26608 31748 26660 31754
rect 26608 31690 26660 31696
rect 27252 31748 27304 31754
rect 27252 31690 27304 31696
rect 26620 28762 26648 31690
rect 26976 31408 27028 31414
rect 26976 31350 27028 31356
rect 26988 31210 27016 31350
rect 26976 31204 27028 31210
rect 26976 31146 27028 31152
rect 27160 30728 27212 30734
rect 27160 30670 27212 30676
rect 26608 28756 26660 28762
rect 26608 28698 26660 28704
rect 27172 28626 27200 30670
rect 27160 28620 27212 28626
rect 27160 28562 27212 28568
rect 27172 26994 27200 28562
rect 27160 26988 27212 26994
rect 27160 26930 27212 26936
rect 26700 26784 26752 26790
rect 26700 26726 26752 26732
rect 26608 24608 26660 24614
rect 26608 24550 26660 24556
rect 26620 23769 26648 24550
rect 26606 23760 26662 23769
rect 26606 23695 26662 23704
rect 26608 19916 26660 19922
rect 26608 19858 26660 19864
rect 26620 19514 26648 19858
rect 26608 19508 26660 19514
rect 26608 19450 26660 19456
rect 26608 18284 26660 18290
rect 26608 18226 26660 18232
rect 26620 18086 26648 18226
rect 26608 18080 26660 18086
rect 26608 18022 26660 18028
rect 26712 17252 26740 26726
rect 27264 24614 27292 31690
rect 27356 30938 27384 31758
rect 27344 30932 27396 30938
rect 27344 30874 27396 30880
rect 27436 30252 27488 30258
rect 27436 30194 27488 30200
rect 27344 30048 27396 30054
rect 27342 30016 27344 30025
rect 27396 30016 27398 30025
rect 27342 29951 27398 29960
rect 27448 29850 27476 30194
rect 27436 29844 27488 29850
rect 27436 29786 27488 29792
rect 27436 28484 27488 28490
rect 27436 28426 27488 28432
rect 27448 27878 27476 28426
rect 27436 27872 27488 27878
rect 27436 27814 27488 27820
rect 27252 24608 27304 24614
rect 27252 24550 27304 24556
rect 27434 24440 27490 24449
rect 27434 24375 27490 24384
rect 27448 24342 27476 24375
rect 27436 24336 27488 24342
rect 27436 24278 27488 24284
rect 27540 24274 27568 48486
rect 27632 47802 27660 48622
rect 28368 48210 28396 51200
rect 29012 49230 29040 51200
rect 29000 49224 29052 49230
rect 29000 49166 29052 49172
rect 29736 49156 29788 49162
rect 29736 49098 29788 49104
rect 29276 49088 29328 49094
rect 29276 49030 29328 49036
rect 28080 48204 28132 48210
rect 28080 48146 28132 48152
rect 28356 48204 28408 48210
rect 28356 48146 28408 48152
rect 27896 48068 27948 48074
rect 27896 48010 27948 48016
rect 27620 47796 27672 47802
rect 27620 47738 27672 47744
rect 27908 47258 27936 48010
rect 28092 47802 28120 48146
rect 28172 48068 28224 48074
rect 28172 48010 28224 48016
rect 28080 47796 28132 47802
rect 28080 47738 28132 47744
rect 28184 47666 28212 48010
rect 28172 47660 28224 47666
rect 28172 47602 28224 47608
rect 27988 47592 28040 47598
rect 27988 47534 28040 47540
rect 28540 47592 28592 47598
rect 28540 47534 28592 47540
rect 28000 47258 28028 47534
rect 27896 47252 27948 47258
rect 27896 47194 27948 47200
rect 27988 47252 28040 47258
rect 27988 47194 28040 47200
rect 28552 47122 28580 47534
rect 28540 47116 28592 47122
rect 28540 47058 28592 47064
rect 28448 42084 28500 42090
rect 28448 42026 28500 42032
rect 27988 38208 28040 38214
rect 27988 38150 28040 38156
rect 27804 37868 27856 37874
rect 27804 37810 27856 37816
rect 27712 37256 27764 37262
rect 27712 37198 27764 37204
rect 27620 36644 27672 36650
rect 27620 36586 27672 36592
rect 27632 35766 27660 36586
rect 27724 35766 27752 37198
rect 27816 36378 27844 37810
rect 28000 37398 28028 38150
rect 28172 37664 28224 37670
rect 28092 37624 28172 37652
rect 27988 37392 28040 37398
rect 27988 37334 28040 37340
rect 28000 36786 28028 37334
rect 28092 37126 28120 37624
rect 28172 37606 28224 37612
rect 28356 37324 28408 37330
rect 28356 37266 28408 37272
rect 28080 37120 28132 37126
rect 28080 37062 28132 37068
rect 27988 36780 28040 36786
rect 27988 36722 28040 36728
rect 27896 36712 27948 36718
rect 27896 36654 27948 36660
rect 27804 36372 27856 36378
rect 27804 36314 27856 36320
rect 27908 36258 27936 36654
rect 27908 36230 28028 36258
rect 27896 36168 27948 36174
rect 27896 36110 27948 36116
rect 27620 35760 27672 35766
rect 27620 35702 27672 35708
rect 27712 35760 27764 35766
rect 27712 35702 27764 35708
rect 27804 34672 27856 34678
rect 27804 34614 27856 34620
rect 27712 32904 27764 32910
rect 27712 32846 27764 32852
rect 27724 32026 27752 32846
rect 27712 32020 27764 32026
rect 27712 31962 27764 31968
rect 27724 31822 27752 31962
rect 27712 31816 27764 31822
rect 27712 31758 27764 31764
rect 27712 27396 27764 27402
rect 27712 27338 27764 27344
rect 27724 26586 27752 27338
rect 27816 26586 27844 34614
rect 27712 26580 27764 26586
rect 27712 26522 27764 26528
rect 27804 26580 27856 26586
rect 27804 26522 27856 26528
rect 27620 25220 27672 25226
rect 27620 25162 27672 25168
rect 27528 24268 27580 24274
rect 27528 24210 27580 24216
rect 27528 24132 27580 24138
rect 27528 24074 27580 24080
rect 26884 24064 26936 24070
rect 26884 24006 26936 24012
rect 26896 23730 26924 24006
rect 27540 23769 27568 24074
rect 27526 23760 27582 23769
rect 26884 23724 26936 23730
rect 27526 23695 27582 23704
rect 26884 23666 26936 23672
rect 26792 19780 26844 19786
rect 26792 19722 26844 19728
rect 26804 19310 26832 19722
rect 26792 19304 26844 19310
rect 26792 19246 26844 19252
rect 26804 18698 26832 19246
rect 26792 18692 26844 18698
rect 26792 18634 26844 18640
rect 26804 18426 26832 18634
rect 26792 18420 26844 18426
rect 26792 18362 26844 18368
rect 26896 18086 26924 23666
rect 27160 23656 27212 23662
rect 27160 23598 27212 23604
rect 27172 23497 27200 23598
rect 27158 23488 27214 23497
rect 27158 23423 27214 23432
rect 27344 22976 27396 22982
rect 27344 22918 27396 22924
rect 27356 22234 27384 22918
rect 27344 22228 27396 22234
rect 27344 22170 27396 22176
rect 27356 22030 27384 22170
rect 27344 22024 27396 22030
rect 27344 21966 27396 21972
rect 27528 22024 27580 22030
rect 27528 21966 27580 21972
rect 27436 21888 27488 21894
rect 27436 21830 27488 21836
rect 27448 21554 27476 21830
rect 27436 21548 27488 21554
rect 27436 21490 27488 21496
rect 27160 21344 27212 21350
rect 27160 21286 27212 21292
rect 27172 21078 27200 21286
rect 27540 21078 27568 21966
rect 27160 21072 27212 21078
rect 27160 21014 27212 21020
rect 27528 21072 27580 21078
rect 27528 21014 27580 21020
rect 27344 20256 27396 20262
rect 27344 20198 27396 20204
rect 27356 19718 27384 20198
rect 27160 19712 27212 19718
rect 27160 19654 27212 19660
rect 27344 19712 27396 19718
rect 27344 19654 27396 19660
rect 27066 19544 27122 19553
rect 27066 19479 27122 19488
rect 26974 19408 27030 19417
rect 27080 19378 27108 19479
rect 26974 19343 26976 19352
rect 27028 19343 27030 19352
rect 27068 19372 27120 19378
rect 26976 19314 27028 19320
rect 27068 19314 27120 19320
rect 27172 18290 27200 19654
rect 27436 18624 27488 18630
rect 27436 18566 27488 18572
rect 27160 18284 27212 18290
rect 27160 18226 27212 18232
rect 27344 18284 27396 18290
rect 27344 18226 27396 18232
rect 26884 18080 26936 18086
rect 26884 18022 26936 18028
rect 26252 10798 26372 10826
rect 26436 12406 26556 12434
rect 26620 17224 26740 17252
rect 26792 17264 26844 17270
rect 26252 10305 26280 10798
rect 26332 10668 26384 10674
rect 26332 10610 26384 10616
rect 26238 10296 26294 10305
rect 26238 10231 26294 10240
rect 26344 9722 26372 10610
rect 26332 9716 26384 9722
rect 26332 9658 26384 9664
rect 26056 9580 26108 9586
rect 26056 9522 26108 9528
rect 26068 8838 26096 9522
rect 26240 9512 26292 9518
rect 26240 9454 26292 9460
rect 26252 9382 26280 9454
rect 26240 9376 26292 9382
rect 26240 9318 26292 9324
rect 26344 8906 26372 9658
rect 26332 8900 26384 8906
rect 26332 8842 26384 8848
rect 26056 8832 26108 8838
rect 26056 8774 26108 8780
rect 26054 8528 26110 8537
rect 26054 8463 26110 8472
rect 26068 8362 26096 8463
rect 26056 8356 26108 8362
rect 26056 8298 26108 8304
rect 25964 8288 26016 8294
rect 25964 8230 26016 8236
rect 26240 8288 26292 8294
rect 26240 8230 26292 8236
rect 26252 8022 26280 8230
rect 26240 8016 26292 8022
rect 26240 7958 26292 7964
rect 26436 7562 26464 12406
rect 26516 10804 26568 10810
rect 26516 10746 26568 10752
rect 26528 10470 26556 10746
rect 26516 10464 26568 10470
rect 26516 10406 26568 10412
rect 26528 10266 26556 10406
rect 26516 10260 26568 10266
rect 26516 10202 26568 10208
rect 26344 7534 26464 7562
rect 25780 5840 25832 5846
rect 25780 5782 25832 5788
rect 25792 5234 25820 5782
rect 25780 5228 25832 5234
rect 25780 5170 25832 5176
rect 26240 4140 26292 4146
rect 26240 4082 26292 4088
rect 26252 3602 26280 4082
rect 26240 3596 26292 3602
rect 26240 3538 26292 3544
rect 25872 3528 25924 3534
rect 25872 3470 25924 3476
rect 25884 3058 25912 3470
rect 25872 3052 25924 3058
rect 25872 2994 25924 3000
rect 24412 2746 24716 2774
rect 24412 2446 24440 2746
rect 26344 2650 26372 7534
rect 26620 4146 26648 17224
rect 26792 17206 26844 17212
rect 26804 15910 26832 17206
rect 26884 17060 26936 17066
rect 26884 17002 26936 17008
rect 26896 16794 26924 17002
rect 26884 16788 26936 16794
rect 26884 16730 26936 16736
rect 27356 16726 27384 18226
rect 27448 18222 27476 18566
rect 27632 18290 27660 25162
rect 27802 24712 27858 24721
rect 27802 24647 27858 24656
rect 27712 24064 27764 24070
rect 27712 24006 27764 24012
rect 27724 22982 27752 24006
rect 27816 23905 27844 24647
rect 27802 23896 27858 23905
rect 27802 23831 27858 23840
rect 27804 23044 27856 23050
rect 27804 22986 27856 22992
rect 27712 22976 27764 22982
rect 27712 22918 27764 22924
rect 27724 22642 27752 22918
rect 27816 22778 27844 22986
rect 27804 22772 27856 22778
rect 27804 22714 27856 22720
rect 27712 22636 27764 22642
rect 27712 22578 27764 22584
rect 27908 22094 27936 36110
rect 28000 34406 28028 36230
rect 28092 34474 28120 37062
rect 28264 36780 28316 36786
rect 28264 36722 28316 36728
rect 28276 36038 28304 36722
rect 28368 36718 28396 37266
rect 28356 36712 28408 36718
rect 28356 36654 28408 36660
rect 28356 36576 28408 36582
rect 28356 36518 28408 36524
rect 28368 36174 28396 36518
rect 28356 36168 28408 36174
rect 28356 36110 28408 36116
rect 28264 36032 28316 36038
rect 28264 35974 28316 35980
rect 28172 35692 28224 35698
rect 28172 35634 28224 35640
rect 28080 34468 28132 34474
rect 28080 34410 28132 34416
rect 27988 34400 28040 34406
rect 27988 34342 28040 34348
rect 28000 32434 28028 34342
rect 28080 34060 28132 34066
rect 28080 34002 28132 34008
rect 28092 32842 28120 34002
rect 28184 33266 28212 35634
rect 28276 34610 28304 35974
rect 28264 34604 28316 34610
rect 28264 34546 28316 34552
rect 28356 33992 28408 33998
rect 28356 33934 28408 33940
rect 28368 33658 28396 33934
rect 28356 33652 28408 33658
rect 28356 33594 28408 33600
rect 28184 33238 28304 33266
rect 28080 32836 28132 32842
rect 28080 32778 28132 32784
rect 28172 32768 28224 32774
rect 28172 32710 28224 32716
rect 27988 32428 28040 32434
rect 27988 32370 28040 32376
rect 28184 31822 28212 32710
rect 28276 32314 28304 33238
rect 28356 32360 28408 32366
rect 28276 32308 28356 32314
rect 28276 32302 28408 32308
rect 28276 32286 28396 32302
rect 28172 31816 28224 31822
rect 28172 31758 28224 31764
rect 27988 31408 28040 31414
rect 27988 31350 28040 31356
rect 28000 30054 28028 31350
rect 27988 30048 28040 30054
rect 27988 29990 28040 29996
rect 27988 29572 28040 29578
rect 27988 29514 28040 29520
rect 28000 28762 28028 29514
rect 27988 28756 28040 28762
rect 27988 28698 28040 28704
rect 28172 27328 28224 27334
rect 28172 27270 28224 27276
rect 28184 27130 28212 27270
rect 28172 27124 28224 27130
rect 28172 27066 28224 27072
rect 28080 26988 28132 26994
rect 28080 26930 28132 26936
rect 28092 26790 28120 26930
rect 28080 26784 28132 26790
rect 28080 26726 28132 26732
rect 27988 24948 28040 24954
rect 27988 24890 28040 24896
rect 28000 24818 28028 24890
rect 27988 24812 28040 24818
rect 27988 24754 28040 24760
rect 28000 24410 28028 24754
rect 27988 24404 28040 24410
rect 27988 24346 28040 24352
rect 28276 24290 28304 32286
rect 28356 32224 28408 32230
rect 28356 32166 28408 32172
rect 28368 31822 28396 32166
rect 28356 31816 28408 31822
rect 28356 31758 28408 31764
rect 28460 31482 28488 42026
rect 29184 37188 29236 37194
rect 29184 37130 29236 37136
rect 29196 36922 29224 37130
rect 29184 36916 29236 36922
rect 29184 36858 29236 36864
rect 28540 36168 28592 36174
rect 28540 36110 28592 36116
rect 28552 35766 28580 36110
rect 28540 35760 28592 35766
rect 28540 35702 28592 35708
rect 29000 35692 29052 35698
rect 29000 35634 29052 35640
rect 28724 35080 28776 35086
rect 28724 35022 28776 35028
rect 28736 34746 28764 35022
rect 28724 34740 28776 34746
rect 28724 34682 28776 34688
rect 28632 34604 28684 34610
rect 28632 34546 28684 34552
rect 28644 32774 28672 34546
rect 29012 33862 29040 35634
rect 29000 33856 29052 33862
rect 29000 33798 29052 33804
rect 28816 32972 28868 32978
rect 28816 32914 28868 32920
rect 28632 32768 28684 32774
rect 28632 32710 28684 32716
rect 28644 32570 28672 32710
rect 28632 32564 28684 32570
rect 28632 32506 28684 32512
rect 28828 32298 28856 32914
rect 28908 32564 28960 32570
rect 28908 32506 28960 32512
rect 28920 32366 28948 32506
rect 28908 32360 28960 32366
rect 28908 32302 28960 32308
rect 28816 32292 28868 32298
rect 28816 32234 28868 32240
rect 28448 31476 28500 31482
rect 28448 31418 28500 31424
rect 28908 31136 28960 31142
rect 28908 31078 28960 31084
rect 28920 30870 28948 31078
rect 29012 30938 29040 33798
rect 29184 31136 29236 31142
rect 29184 31078 29236 31084
rect 29000 30932 29052 30938
rect 29000 30874 29052 30880
rect 28908 30864 28960 30870
rect 28908 30806 28960 30812
rect 28632 30660 28684 30666
rect 28632 30602 28684 30608
rect 28644 30190 28672 30602
rect 28908 30252 28960 30258
rect 29012 30240 29040 30874
rect 29092 30864 29144 30870
rect 29092 30806 29144 30812
rect 28960 30212 29040 30240
rect 28908 30194 28960 30200
rect 28632 30184 28684 30190
rect 28632 30126 28684 30132
rect 29000 30048 29052 30054
rect 29000 29990 29052 29996
rect 29012 29714 29040 29990
rect 29000 29708 29052 29714
rect 29000 29650 29052 29656
rect 28724 29504 28776 29510
rect 28724 29446 28776 29452
rect 28736 29170 28764 29446
rect 29012 29306 29040 29650
rect 29000 29300 29052 29306
rect 29000 29242 29052 29248
rect 28448 29164 28500 29170
rect 28448 29106 28500 29112
rect 28724 29164 28776 29170
rect 28724 29106 28776 29112
rect 28460 27402 28488 29106
rect 29000 29028 29052 29034
rect 29000 28970 29052 28976
rect 29012 28694 29040 28970
rect 29104 28966 29132 30806
rect 29196 30258 29224 31078
rect 29184 30252 29236 30258
rect 29184 30194 29236 30200
rect 29184 29300 29236 29306
rect 29184 29242 29236 29248
rect 29092 28960 29144 28966
rect 29092 28902 29144 28908
rect 29000 28688 29052 28694
rect 29000 28630 29052 28636
rect 28540 28484 28592 28490
rect 28540 28426 28592 28432
rect 28552 28082 28580 28426
rect 28540 28076 28592 28082
rect 28540 28018 28592 28024
rect 28448 27396 28500 27402
rect 28448 27338 28500 27344
rect 28724 27396 28776 27402
rect 28724 27338 28776 27344
rect 28448 26988 28500 26994
rect 28448 26930 28500 26936
rect 28460 24886 28488 26930
rect 28736 26790 28764 27338
rect 28908 27328 28960 27334
rect 28908 27270 28960 27276
rect 28920 26926 28948 27270
rect 28908 26920 28960 26926
rect 28908 26862 28960 26868
rect 28724 26784 28776 26790
rect 28724 26726 28776 26732
rect 28632 26580 28684 26586
rect 28632 26522 28684 26528
rect 28448 24880 28500 24886
rect 28448 24822 28500 24828
rect 28540 24744 28592 24750
rect 28540 24686 28592 24692
rect 28356 24608 28408 24614
rect 28356 24550 28408 24556
rect 27816 22066 27936 22094
rect 28000 24262 28304 24290
rect 28368 24274 28396 24550
rect 28552 24410 28580 24686
rect 28540 24404 28592 24410
rect 28540 24346 28592 24352
rect 28356 24268 28408 24274
rect 27710 19408 27766 19417
rect 27710 19343 27766 19352
rect 27620 18284 27672 18290
rect 27620 18226 27672 18232
rect 27436 18216 27488 18222
rect 27436 18158 27488 18164
rect 27632 16726 27660 18226
rect 27344 16720 27396 16726
rect 27344 16662 27396 16668
rect 27620 16720 27672 16726
rect 27620 16662 27672 16668
rect 26884 15972 26936 15978
rect 26884 15914 26936 15920
rect 26792 15904 26844 15910
rect 26792 15846 26844 15852
rect 26700 15632 26752 15638
rect 26700 15574 26752 15580
rect 26712 14618 26740 15574
rect 26896 15434 26924 15914
rect 26884 15428 26936 15434
rect 26884 15370 26936 15376
rect 27068 15156 27120 15162
rect 27068 15098 27120 15104
rect 26700 14612 26752 14618
rect 26700 14554 26752 14560
rect 26712 14498 26740 14554
rect 27080 14550 27108 15098
rect 27252 15088 27304 15094
rect 27252 15030 27304 15036
rect 27264 14958 27292 15030
rect 27252 14952 27304 14958
rect 27252 14894 27304 14900
rect 27068 14544 27120 14550
rect 26712 14470 26832 14498
rect 27068 14486 27120 14492
rect 26700 14408 26752 14414
rect 26700 14350 26752 14356
rect 26712 13802 26740 14350
rect 26700 13796 26752 13802
rect 26700 13738 26752 13744
rect 26700 12776 26752 12782
rect 26700 12718 26752 12724
rect 26712 11898 26740 12718
rect 26804 12646 26832 14470
rect 27264 14056 27292 14894
rect 27356 14482 27384 16662
rect 27528 15156 27580 15162
rect 27528 15098 27580 15104
rect 27540 14929 27568 15098
rect 27526 14920 27582 14929
rect 27526 14855 27582 14864
rect 27344 14476 27396 14482
rect 27344 14418 27396 14424
rect 27724 14362 27752 19343
rect 27632 14334 27752 14362
rect 27264 14028 27384 14056
rect 26792 12640 26844 12646
rect 26792 12582 26844 12588
rect 27252 12640 27304 12646
rect 27252 12582 27304 12588
rect 26804 12434 26832 12582
rect 26804 12406 27016 12434
rect 26700 11892 26752 11898
rect 26700 11834 26752 11840
rect 26700 10736 26752 10742
rect 26700 10678 26752 10684
rect 26712 9926 26740 10678
rect 26988 9994 27016 12406
rect 27264 11150 27292 12582
rect 27356 12306 27384 14028
rect 27436 13524 27488 13530
rect 27436 13466 27488 13472
rect 27448 13326 27476 13466
rect 27436 13320 27488 13326
rect 27436 13262 27488 13268
rect 27632 13190 27660 14334
rect 27712 14272 27764 14278
rect 27712 14214 27764 14220
rect 27620 13184 27672 13190
rect 27620 13126 27672 13132
rect 27632 12646 27660 13126
rect 27620 12640 27672 12646
rect 27620 12582 27672 12588
rect 27344 12300 27396 12306
rect 27344 12242 27396 12248
rect 27252 11144 27304 11150
rect 27252 11086 27304 11092
rect 27068 10668 27120 10674
rect 27068 10610 27120 10616
rect 26976 9988 27028 9994
rect 26976 9930 27028 9936
rect 26700 9920 26752 9926
rect 26700 9862 26752 9868
rect 26712 9654 26740 9862
rect 26700 9648 26752 9654
rect 26700 9590 26752 9596
rect 26712 8906 26740 9590
rect 26884 9444 26936 9450
rect 26884 9386 26936 9392
rect 26896 9178 26924 9386
rect 26988 9382 27016 9930
rect 26976 9376 27028 9382
rect 26976 9318 27028 9324
rect 26884 9172 26936 9178
rect 26884 9114 26936 9120
rect 27080 9110 27108 10610
rect 27160 10464 27212 10470
rect 27160 10406 27212 10412
rect 27068 9104 27120 9110
rect 27068 9046 27120 9052
rect 26700 8900 26752 8906
rect 26700 8842 26752 8848
rect 27172 8498 27200 10406
rect 27356 9586 27384 12242
rect 27620 12232 27672 12238
rect 27620 12174 27672 12180
rect 27436 11688 27488 11694
rect 27436 11630 27488 11636
rect 27344 9580 27396 9586
rect 27344 9522 27396 9528
rect 27252 9512 27304 9518
rect 27252 9454 27304 9460
rect 27264 8838 27292 9454
rect 27448 9042 27476 11630
rect 27632 11286 27660 12174
rect 27620 11280 27672 11286
rect 27620 11222 27672 11228
rect 27620 11144 27672 11150
rect 27540 11104 27620 11132
rect 27540 9625 27568 11104
rect 27620 11086 27672 11092
rect 27724 11082 27752 14214
rect 27712 11076 27764 11082
rect 27712 11018 27764 11024
rect 27620 10056 27672 10062
rect 27620 9998 27672 10004
rect 27632 9654 27660 9998
rect 27620 9648 27672 9654
rect 27526 9616 27582 9625
rect 27620 9590 27672 9596
rect 27526 9551 27582 9560
rect 27436 9036 27488 9042
rect 27436 8978 27488 8984
rect 27252 8832 27304 8838
rect 27252 8774 27304 8780
rect 27160 8492 27212 8498
rect 27160 8434 27212 8440
rect 27264 8430 27292 8774
rect 27252 8424 27304 8430
rect 27250 8392 27252 8401
rect 27304 8392 27306 8401
rect 27250 8327 27306 8336
rect 27448 7886 27476 8978
rect 27540 8430 27568 9551
rect 27632 8634 27660 9590
rect 27620 8628 27672 8634
rect 27620 8570 27672 8576
rect 27620 8492 27672 8498
rect 27724 8480 27752 11018
rect 27672 8452 27752 8480
rect 27620 8434 27672 8440
rect 27528 8424 27580 8430
rect 27528 8366 27580 8372
rect 27436 7880 27488 7886
rect 27436 7822 27488 7828
rect 27448 7342 27476 7822
rect 27816 7546 27844 22066
rect 27896 18692 27948 18698
rect 27896 18634 27948 18640
rect 27908 18426 27936 18634
rect 27896 18420 27948 18426
rect 27896 18362 27948 18368
rect 27896 17672 27948 17678
rect 27896 17614 27948 17620
rect 27908 17202 27936 17614
rect 27896 17196 27948 17202
rect 27896 17138 27948 17144
rect 27908 16810 27936 17138
rect 28000 16998 28028 24262
rect 28356 24210 28408 24216
rect 28264 24200 28316 24206
rect 28264 24142 28316 24148
rect 28080 24132 28132 24138
rect 28080 24074 28132 24080
rect 28092 23866 28120 24074
rect 28080 23860 28132 23866
rect 28080 23802 28132 23808
rect 28092 23662 28120 23802
rect 28172 23724 28224 23730
rect 28172 23666 28224 23672
rect 28080 23656 28132 23662
rect 28080 23598 28132 23604
rect 28184 23361 28212 23666
rect 28170 23352 28226 23361
rect 28170 23287 28226 23296
rect 28276 23254 28304 24142
rect 28264 23248 28316 23254
rect 28264 23190 28316 23196
rect 28368 23100 28396 24210
rect 28448 24200 28500 24206
rect 28552 24177 28580 24346
rect 28448 24142 28500 24148
rect 28538 24168 28594 24177
rect 28460 23526 28488 24142
rect 28538 24103 28594 24112
rect 28538 24032 28594 24041
rect 28538 23967 28594 23976
rect 28552 23730 28580 23967
rect 28540 23724 28592 23730
rect 28540 23666 28592 23672
rect 28448 23520 28500 23526
rect 28644 23474 28672 26522
rect 28448 23462 28500 23468
rect 28276 23072 28396 23100
rect 28080 22704 28132 22710
rect 28080 22646 28132 22652
rect 28092 22438 28120 22646
rect 28080 22432 28132 22438
rect 28080 22374 28132 22380
rect 28276 22094 28304 23072
rect 28356 22432 28408 22438
rect 28356 22374 28408 22380
rect 28092 22066 28304 22094
rect 27988 16992 28040 16998
rect 27988 16934 28040 16940
rect 27908 16782 28028 16810
rect 27896 16720 27948 16726
rect 27896 16662 27948 16668
rect 27908 14414 27936 16662
rect 28000 16658 28028 16782
rect 27988 16652 28040 16658
rect 27988 16594 28040 16600
rect 27988 14544 28040 14550
rect 27988 14486 28040 14492
rect 27896 14408 27948 14414
rect 27896 14350 27948 14356
rect 27908 11150 27936 14350
rect 28000 14074 28028 14486
rect 27988 14068 28040 14074
rect 27988 14010 28040 14016
rect 27988 13796 28040 13802
rect 27988 13738 28040 13744
rect 28000 13326 28028 13738
rect 27988 13320 28040 13326
rect 27988 13262 28040 13268
rect 28000 12986 28028 13262
rect 27988 12980 28040 12986
rect 27988 12922 28040 12928
rect 28092 12434 28120 22066
rect 28172 22024 28224 22030
rect 28172 21966 28224 21972
rect 28264 22024 28316 22030
rect 28264 21966 28316 21972
rect 28184 21894 28212 21966
rect 28172 21888 28224 21894
rect 28276 21865 28304 21966
rect 28172 21830 28224 21836
rect 28262 21856 28318 21865
rect 28262 21791 28318 21800
rect 28262 21720 28318 21729
rect 28262 21655 28318 21664
rect 28276 19786 28304 21655
rect 28368 20942 28396 22374
rect 28356 20936 28408 20942
rect 28356 20878 28408 20884
rect 28264 19780 28316 19786
rect 28264 19722 28316 19728
rect 28276 18426 28304 19722
rect 28356 18692 28408 18698
rect 28356 18634 28408 18640
rect 28264 18420 28316 18426
rect 28264 18362 28316 18368
rect 28276 17882 28304 18362
rect 28368 18290 28396 18634
rect 28356 18284 28408 18290
rect 28356 18226 28408 18232
rect 28264 17876 28316 17882
rect 28264 17818 28316 17824
rect 28368 17678 28396 18226
rect 28356 17672 28408 17678
rect 28356 17614 28408 17620
rect 28264 15428 28316 15434
rect 28264 15370 28316 15376
rect 28172 15020 28224 15026
rect 28172 14962 28224 14968
rect 28184 14550 28212 14962
rect 28172 14544 28224 14550
rect 28172 14486 28224 14492
rect 28184 14414 28212 14486
rect 28276 14414 28304 15370
rect 28356 14952 28408 14958
rect 28356 14894 28408 14900
rect 28172 14408 28224 14414
rect 28172 14350 28224 14356
rect 28264 14408 28316 14414
rect 28264 14350 28316 14356
rect 28172 14272 28224 14278
rect 28172 14214 28224 14220
rect 28184 13394 28212 14214
rect 28368 13870 28396 14894
rect 28356 13864 28408 13870
rect 28356 13806 28408 13812
rect 28172 13388 28224 13394
rect 28172 13330 28224 13336
rect 28172 13184 28224 13190
rect 28172 13126 28224 13132
rect 28184 12850 28212 13126
rect 28172 12844 28224 12850
rect 28172 12786 28224 12792
rect 28264 12640 28316 12646
rect 28264 12582 28316 12588
rect 28000 12406 28120 12434
rect 28276 12434 28304 12582
rect 28276 12406 28396 12434
rect 27896 11144 27948 11150
rect 27896 11086 27948 11092
rect 27896 8900 27948 8906
rect 27896 8842 27948 8848
rect 27908 8634 27936 8842
rect 27896 8628 27948 8634
rect 27896 8570 27948 8576
rect 27804 7540 27856 7546
rect 27804 7482 27856 7488
rect 27436 7336 27488 7342
rect 27436 7278 27488 7284
rect 27804 6316 27856 6322
rect 27804 6258 27856 6264
rect 27816 5914 27844 6258
rect 27804 5908 27856 5914
rect 27804 5850 27856 5856
rect 27160 5772 27212 5778
rect 27160 5714 27212 5720
rect 27172 5642 27200 5714
rect 27160 5636 27212 5642
rect 27160 5578 27212 5584
rect 27712 5636 27764 5642
rect 27712 5578 27764 5584
rect 27724 5370 27752 5578
rect 27712 5364 27764 5370
rect 27712 5306 27764 5312
rect 26608 4140 26660 4146
rect 26608 4082 26660 4088
rect 26424 3596 26476 3602
rect 26424 3538 26476 3544
rect 26332 2644 26384 2650
rect 26332 2586 26384 2592
rect 24400 2440 24452 2446
rect 24400 2382 24452 2388
rect 24492 2372 24544 2378
rect 24492 2314 24544 2320
rect 25136 2372 25188 2378
rect 25136 2314 25188 2320
rect 23940 1964 23992 1970
rect 23940 1906 23992 1912
rect 24504 800 24532 2314
rect 25148 800 25176 2314
rect 26436 800 26464 3538
rect 28000 2530 28028 12406
rect 28264 12164 28316 12170
rect 28264 12106 28316 12112
rect 28172 12096 28224 12102
rect 28172 12038 28224 12044
rect 28184 11830 28212 12038
rect 28172 11824 28224 11830
rect 28172 11766 28224 11772
rect 28080 11756 28132 11762
rect 28080 11698 28132 11704
rect 28092 11354 28120 11698
rect 28080 11348 28132 11354
rect 28080 11290 28132 11296
rect 28184 11218 28212 11766
rect 28276 11354 28304 12106
rect 28264 11348 28316 11354
rect 28264 11290 28316 11296
rect 28172 11212 28224 11218
rect 28172 11154 28224 11160
rect 28368 10266 28396 12406
rect 28356 10260 28408 10266
rect 28356 10202 28408 10208
rect 28080 7540 28132 7546
rect 28080 7482 28132 7488
rect 28092 2650 28120 7482
rect 28172 6112 28224 6118
rect 28172 6054 28224 6060
rect 28184 5234 28212 6054
rect 28172 5228 28224 5234
rect 28172 5170 28224 5176
rect 28080 2644 28132 2650
rect 28080 2586 28132 2592
rect 28000 2502 28212 2530
rect 27068 2440 27120 2446
rect 27068 2382 27120 2388
rect 27080 800 27108 2382
rect 27712 2372 27764 2378
rect 27712 2314 27764 2320
rect 27724 800 27752 2314
rect 28184 2310 28212 2502
rect 28172 2304 28224 2310
rect 28172 2246 28224 2252
rect 28460 1902 28488 23462
rect 28552 23446 28672 23474
rect 28552 21729 28580 23446
rect 28736 23338 28764 26726
rect 29000 25764 29052 25770
rect 29000 25706 29052 25712
rect 29012 25362 29040 25706
rect 29000 25356 29052 25362
rect 29000 25298 29052 25304
rect 29092 24948 29144 24954
rect 29092 24890 29144 24896
rect 29000 24744 29052 24750
rect 29000 24686 29052 24692
rect 29012 24585 29040 24686
rect 28998 24576 29054 24585
rect 28998 24511 29054 24520
rect 29104 24410 29132 24890
rect 29092 24404 29144 24410
rect 29092 24346 29144 24352
rect 28998 24304 29054 24313
rect 28828 24248 28998 24256
rect 28828 24239 29054 24248
rect 28828 24228 29040 24239
rect 28828 23633 28856 24228
rect 28906 24168 28962 24177
rect 28906 24103 28962 24112
rect 29092 24132 29144 24138
rect 28814 23624 28870 23633
rect 28814 23559 28870 23568
rect 28644 23310 28764 23338
rect 28644 22506 28672 23310
rect 28724 23248 28776 23254
rect 28722 23216 28724 23225
rect 28776 23216 28778 23225
rect 28722 23151 28778 23160
rect 28724 22976 28776 22982
rect 28724 22918 28776 22924
rect 28736 22642 28764 22918
rect 28724 22636 28776 22642
rect 28724 22578 28776 22584
rect 28632 22500 28684 22506
rect 28632 22442 28684 22448
rect 28538 21720 28594 21729
rect 28538 21655 28594 21664
rect 28540 21548 28592 21554
rect 28540 21490 28592 21496
rect 28552 20942 28580 21490
rect 28540 20936 28592 20942
rect 28540 20878 28592 20884
rect 28644 17066 28672 22442
rect 28736 21554 28764 22578
rect 28828 22098 28856 23559
rect 28816 22092 28868 22098
rect 28816 22034 28868 22040
rect 28724 21548 28776 21554
rect 28724 21490 28776 21496
rect 28722 20088 28778 20097
rect 28722 20023 28778 20032
rect 28736 19786 28764 20023
rect 28724 19780 28776 19786
rect 28724 19722 28776 19728
rect 28540 17060 28592 17066
rect 28540 17002 28592 17008
rect 28632 17060 28684 17066
rect 28632 17002 28684 17008
rect 28552 13258 28580 17002
rect 28722 15328 28778 15337
rect 28722 15263 28778 15272
rect 28736 14958 28764 15263
rect 28816 15020 28868 15026
rect 28816 14962 28868 14968
rect 28724 14952 28776 14958
rect 28724 14894 28776 14900
rect 28724 14816 28776 14822
rect 28724 14758 28776 14764
rect 28736 13818 28764 14758
rect 28644 13790 28764 13818
rect 28540 13252 28592 13258
rect 28540 13194 28592 13200
rect 28644 12238 28672 13790
rect 28724 13728 28776 13734
rect 28724 13670 28776 13676
rect 28736 13258 28764 13670
rect 28724 13252 28776 13258
rect 28724 13194 28776 13200
rect 28828 12986 28856 14962
rect 28816 12980 28868 12986
rect 28816 12922 28868 12928
rect 28632 12232 28684 12238
rect 28632 12174 28684 12180
rect 28644 11898 28672 12174
rect 28632 11892 28684 11898
rect 28632 11834 28684 11840
rect 28724 11076 28776 11082
rect 28724 11018 28776 11024
rect 28736 10810 28764 11018
rect 28724 10804 28776 10810
rect 28724 10746 28776 10752
rect 28632 10600 28684 10606
rect 28632 10542 28684 10548
rect 28644 9994 28672 10542
rect 28632 9988 28684 9994
rect 28632 9930 28684 9936
rect 28644 6390 28672 9930
rect 28632 6384 28684 6390
rect 28632 6326 28684 6332
rect 28736 5234 28764 10746
rect 28724 5228 28776 5234
rect 28724 5170 28776 5176
rect 28736 5098 28764 5170
rect 28724 5092 28776 5098
rect 28724 5034 28776 5040
rect 28920 2582 28948 24103
rect 29092 24074 29144 24080
rect 28998 23896 29054 23905
rect 28998 23831 29000 23840
rect 29052 23831 29054 23840
rect 29000 23802 29052 23808
rect 29104 23746 29132 24074
rect 29196 24041 29224 29242
rect 29288 24274 29316 49030
rect 29748 48754 29776 49098
rect 29736 48748 29788 48754
rect 29736 48690 29788 48696
rect 29932 48210 29960 51326
rect 30930 51200 30986 52000
rect 31574 51200 31630 52000
rect 32218 51354 32274 52000
rect 31956 51326 32274 51354
rect 30012 48884 30064 48890
rect 30012 48826 30064 48832
rect 29828 48204 29880 48210
rect 29828 48146 29880 48152
rect 29920 48204 29972 48210
rect 29920 48146 29972 48152
rect 29840 48074 29868 48146
rect 29736 48068 29788 48074
rect 29736 48010 29788 48016
rect 29828 48068 29880 48074
rect 29828 48010 29880 48016
rect 29748 47258 29776 48010
rect 29736 47252 29788 47258
rect 29736 47194 29788 47200
rect 30024 45554 30052 48826
rect 30564 48680 30616 48686
rect 30564 48622 30616 48628
rect 30576 47802 30604 48622
rect 30748 48612 30800 48618
rect 30748 48554 30800 48560
rect 30380 47796 30432 47802
rect 30380 47738 30432 47744
rect 30564 47796 30616 47802
rect 30564 47738 30616 47744
rect 30392 47682 30420 47738
rect 30392 47654 30604 47682
rect 30576 47530 30604 47654
rect 30564 47524 30616 47530
rect 30564 47466 30616 47472
rect 29932 45526 30052 45554
rect 29932 37942 29960 45526
rect 29552 37936 29604 37942
rect 29552 37878 29604 37884
rect 29920 37936 29972 37942
rect 29920 37878 29972 37884
rect 29564 37262 29592 37878
rect 30104 37664 30156 37670
rect 30104 37606 30156 37612
rect 30288 37664 30340 37670
rect 30288 37606 30340 37612
rect 30116 37482 30144 37606
rect 30116 37466 30236 37482
rect 30116 37460 30248 37466
rect 30116 37454 30196 37460
rect 30196 37402 30248 37408
rect 29552 37256 29604 37262
rect 29552 37198 29604 37204
rect 29564 36786 29592 37198
rect 29828 37188 29880 37194
rect 29828 37130 29880 37136
rect 29552 36780 29604 36786
rect 29552 36722 29604 36728
rect 29368 35692 29420 35698
rect 29368 35634 29420 35640
rect 29380 35222 29408 35634
rect 29460 35488 29512 35494
rect 29460 35430 29512 35436
rect 29472 35290 29500 35430
rect 29460 35284 29512 35290
rect 29460 35226 29512 35232
rect 29368 35216 29420 35222
rect 29368 35158 29420 35164
rect 29564 34066 29592 36722
rect 29840 36378 29868 37130
rect 30104 37120 30156 37126
rect 30104 37062 30156 37068
rect 30012 36780 30064 36786
rect 30012 36722 30064 36728
rect 29828 36372 29880 36378
rect 29828 36314 29880 36320
rect 29920 36168 29972 36174
rect 29920 36110 29972 36116
rect 29932 35766 29960 36110
rect 30024 35834 30052 36722
rect 30116 36242 30144 37062
rect 30208 36378 30236 37402
rect 30196 36372 30248 36378
rect 30196 36314 30248 36320
rect 30104 36236 30156 36242
rect 30104 36178 30156 36184
rect 30012 35828 30064 35834
rect 30012 35770 30064 35776
rect 29920 35760 29972 35766
rect 29920 35702 29972 35708
rect 30116 35630 30144 36178
rect 30104 35624 30156 35630
rect 30104 35566 30156 35572
rect 30208 35578 30236 36314
rect 30300 36242 30328 37606
rect 30380 36576 30432 36582
rect 30380 36518 30432 36524
rect 30288 36236 30340 36242
rect 30288 36178 30340 36184
rect 30392 35698 30420 36518
rect 30564 36168 30616 36174
rect 30564 36110 30616 36116
rect 30380 35692 30432 35698
rect 30380 35634 30432 35640
rect 30208 35550 30328 35578
rect 30576 35562 30604 36110
rect 30300 35290 30328 35550
rect 30564 35556 30616 35562
rect 30564 35498 30616 35504
rect 30288 35284 30340 35290
rect 30288 35226 30340 35232
rect 30300 34610 30328 35226
rect 30472 35080 30524 35086
rect 30472 35022 30524 35028
rect 30288 34604 30340 34610
rect 30288 34546 30340 34552
rect 29644 34536 29696 34542
rect 29644 34478 29696 34484
rect 29552 34060 29604 34066
rect 29552 34002 29604 34008
rect 29564 33658 29592 34002
rect 29552 33652 29604 33658
rect 29552 33594 29604 33600
rect 29564 30734 29592 33594
rect 29656 31754 29684 34478
rect 30300 34474 30328 34546
rect 30288 34468 30340 34474
rect 30288 34410 30340 34416
rect 30380 34400 30432 34406
rect 30380 34342 30432 34348
rect 30392 33998 30420 34342
rect 30380 33992 30432 33998
rect 30380 33934 30432 33940
rect 30484 33114 30512 35022
rect 30576 34610 30604 35498
rect 30760 35086 30788 48554
rect 30944 48210 30972 51200
rect 31956 48822 31984 51326
rect 32218 51200 32274 51326
rect 32862 51200 32918 52000
rect 33506 51200 33562 52000
rect 34150 51354 34206 52000
rect 34794 51354 34850 52000
rect 34150 51326 34376 51354
rect 34150 51200 34206 51326
rect 32128 49088 32180 49094
rect 32128 49030 32180 49036
rect 31944 48816 31996 48822
rect 31944 48758 31996 48764
rect 32140 48754 32168 49030
rect 32128 48748 32180 48754
rect 32128 48690 32180 48696
rect 32876 48686 32904 51200
rect 33520 49314 33548 51200
rect 33520 49286 33732 49314
rect 33508 49224 33560 49230
rect 33508 49166 33560 49172
rect 32312 48680 32364 48686
rect 32312 48622 32364 48628
rect 32864 48680 32916 48686
rect 32864 48622 32916 48628
rect 30932 48204 30984 48210
rect 30932 48146 30984 48152
rect 31852 48136 31904 48142
rect 31852 48078 31904 48084
rect 31760 48068 31812 48074
rect 31760 48010 31812 48016
rect 31116 47660 31168 47666
rect 31116 47602 31168 47608
rect 31128 41414 31156 47602
rect 31772 47598 31800 48010
rect 31760 47592 31812 47598
rect 31760 47534 31812 47540
rect 31864 47258 31892 48078
rect 32036 48068 32088 48074
rect 32036 48010 32088 48016
rect 32048 47802 32076 48010
rect 32324 47802 32352 48622
rect 32036 47796 32088 47802
rect 32036 47738 32088 47744
rect 32312 47796 32364 47802
rect 32312 47738 32364 47744
rect 33520 47666 33548 49166
rect 32128 47660 32180 47666
rect 32128 47602 32180 47608
rect 33508 47660 33560 47666
rect 33508 47602 33560 47608
rect 31852 47252 31904 47258
rect 31852 47194 31904 47200
rect 32140 46986 32168 47602
rect 32496 47592 32548 47598
rect 32496 47534 32548 47540
rect 32128 46980 32180 46986
rect 32128 46922 32180 46928
rect 32128 44940 32180 44946
rect 32128 44882 32180 44888
rect 31036 41386 31156 41414
rect 32140 41414 32168 44882
rect 32140 41386 32352 41414
rect 30840 36304 30892 36310
rect 30840 36246 30892 36252
rect 30852 36038 30880 36246
rect 30840 36032 30892 36038
rect 30840 35974 30892 35980
rect 30748 35080 30800 35086
rect 30748 35022 30800 35028
rect 30840 35012 30892 35018
rect 30840 34954 30892 34960
rect 30852 34610 30880 34954
rect 30564 34604 30616 34610
rect 30564 34546 30616 34552
rect 30840 34604 30892 34610
rect 30840 34546 30892 34552
rect 30576 33522 30604 34546
rect 30748 34536 30800 34542
rect 31036 34490 31064 41386
rect 32220 39364 32272 39370
rect 32220 39306 32272 39312
rect 31116 37936 31168 37942
rect 31116 37878 31168 37884
rect 31128 37194 31156 37878
rect 32232 37194 32260 39306
rect 31116 37188 31168 37194
rect 31116 37130 31168 37136
rect 32220 37188 32272 37194
rect 32220 37130 32272 37136
rect 31128 36106 31156 37130
rect 31944 36780 31996 36786
rect 31944 36722 31996 36728
rect 31956 36378 31984 36722
rect 32128 36712 32180 36718
rect 32128 36654 32180 36660
rect 31944 36372 31996 36378
rect 31944 36314 31996 36320
rect 31668 36236 31720 36242
rect 31668 36178 31720 36184
rect 31116 36100 31168 36106
rect 31116 36042 31168 36048
rect 31128 35154 31156 36042
rect 31392 36032 31444 36038
rect 31392 35974 31444 35980
rect 31404 35698 31432 35974
rect 31392 35692 31444 35698
rect 31392 35634 31444 35640
rect 31116 35148 31168 35154
rect 31116 35090 31168 35096
rect 31128 34746 31156 35090
rect 31576 35080 31628 35086
rect 31576 35022 31628 35028
rect 31208 34944 31260 34950
rect 31208 34886 31260 34892
rect 31116 34740 31168 34746
rect 31116 34682 31168 34688
rect 31220 34610 31248 34886
rect 31484 34672 31536 34678
rect 31484 34614 31536 34620
rect 31208 34604 31260 34610
rect 31208 34546 31260 34552
rect 30748 34478 30800 34484
rect 30760 33946 30788 34478
rect 30944 34462 31064 34490
rect 30760 33918 30880 33946
rect 30852 33862 30880 33918
rect 30840 33856 30892 33862
rect 30840 33798 30892 33804
rect 30564 33516 30616 33522
rect 30564 33458 30616 33464
rect 30472 33108 30524 33114
rect 30472 33050 30524 33056
rect 30564 33108 30616 33114
rect 30564 33050 30616 33056
rect 30576 32502 30604 33050
rect 30852 32978 30880 33798
rect 30840 32972 30892 32978
rect 30840 32914 30892 32920
rect 30564 32496 30616 32502
rect 30564 32438 30616 32444
rect 29656 31726 29868 31754
rect 29736 31476 29788 31482
rect 29736 31418 29788 31424
rect 29552 30728 29604 30734
rect 29552 30670 29604 30676
rect 29368 30184 29420 30190
rect 29368 30126 29420 30132
rect 29380 29646 29408 30126
rect 29368 29640 29420 29646
rect 29368 29582 29420 29588
rect 29380 29034 29408 29582
rect 29748 29322 29776 31418
rect 29840 31278 29868 31726
rect 29828 31272 29880 31278
rect 29828 31214 29880 31220
rect 30012 31272 30064 31278
rect 30064 31220 30144 31226
rect 30012 31214 30144 31220
rect 29840 29714 29868 31214
rect 30024 31198 30144 31214
rect 30012 31136 30064 31142
rect 30012 31078 30064 31084
rect 30024 30734 30052 31078
rect 29920 30728 29972 30734
rect 29920 30670 29972 30676
rect 30012 30728 30064 30734
rect 30012 30670 30064 30676
rect 29932 30258 29960 30670
rect 29920 30252 29972 30258
rect 29920 30194 29972 30200
rect 30012 30252 30064 30258
rect 30012 30194 30064 30200
rect 30024 29850 30052 30194
rect 30012 29844 30064 29850
rect 30012 29786 30064 29792
rect 29828 29708 29880 29714
rect 29828 29650 29880 29656
rect 30012 29708 30064 29714
rect 30012 29650 30064 29656
rect 30024 29578 30052 29650
rect 30116 29628 30144 31198
rect 30196 29640 30248 29646
rect 30116 29600 30196 29628
rect 30196 29582 30248 29588
rect 30288 29640 30340 29646
rect 30288 29582 30340 29588
rect 30012 29572 30064 29578
rect 30012 29514 30064 29520
rect 29748 29306 29868 29322
rect 30300 29306 30328 29582
rect 30944 29492 30972 34462
rect 31024 33516 31076 33522
rect 31024 33458 31076 33464
rect 31036 31793 31064 33458
rect 31300 33040 31352 33046
rect 31300 32982 31352 32988
rect 31208 32836 31260 32842
rect 31208 32778 31260 32784
rect 31116 32768 31168 32774
rect 31116 32710 31168 32716
rect 31128 31822 31156 32710
rect 31116 31816 31168 31822
rect 31022 31784 31078 31793
rect 31116 31758 31168 31764
rect 31022 31719 31078 31728
rect 31036 31482 31064 31719
rect 31024 31476 31076 31482
rect 31024 31418 31076 31424
rect 31220 30122 31248 32778
rect 31312 32366 31340 32982
rect 31496 32910 31524 34614
rect 31484 32904 31536 32910
rect 31484 32846 31536 32852
rect 31300 32360 31352 32366
rect 31300 32302 31352 32308
rect 31312 31346 31340 32302
rect 31300 31340 31352 31346
rect 31300 31282 31352 31288
rect 31392 31340 31444 31346
rect 31392 31282 31444 31288
rect 31312 30938 31340 31282
rect 31300 30932 31352 30938
rect 31300 30874 31352 30880
rect 31208 30116 31260 30122
rect 31208 30058 31260 30064
rect 31220 29714 31248 30058
rect 31208 29708 31260 29714
rect 31208 29650 31260 29656
rect 30944 29464 31064 29492
rect 29748 29300 29880 29306
rect 29748 29294 29828 29300
rect 29828 29242 29880 29248
rect 30288 29300 30340 29306
rect 30288 29242 30340 29248
rect 30380 29164 30432 29170
rect 30380 29106 30432 29112
rect 29368 29028 29420 29034
rect 29368 28970 29420 28976
rect 29828 28960 29880 28966
rect 29828 28902 29880 28908
rect 29552 28076 29604 28082
rect 29552 28018 29604 28024
rect 29460 28008 29512 28014
rect 29366 27976 29422 27985
rect 29460 27950 29512 27956
rect 29366 27911 29422 27920
rect 29380 26994 29408 27911
rect 29472 27538 29500 27950
rect 29564 27674 29592 28018
rect 29644 27872 29696 27878
rect 29644 27814 29696 27820
rect 29552 27668 29604 27674
rect 29552 27610 29604 27616
rect 29460 27532 29512 27538
rect 29460 27474 29512 27480
rect 29368 26988 29420 26994
rect 29368 26930 29420 26936
rect 29472 26586 29500 27474
rect 29656 27470 29684 27814
rect 29644 27464 29696 27470
rect 29644 27406 29696 27412
rect 29736 26784 29788 26790
rect 29736 26726 29788 26732
rect 29460 26580 29512 26586
rect 29460 26522 29512 26528
rect 29748 26382 29776 26726
rect 29736 26376 29788 26382
rect 29736 26318 29788 26324
rect 29736 26240 29788 26246
rect 29736 26182 29788 26188
rect 29644 25968 29696 25974
rect 29644 25910 29696 25916
rect 29656 24818 29684 25910
rect 29748 25906 29776 26182
rect 29736 25900 29788 25906
rect 29736 25842 29788 25848
rect 29736 25696 29788 25702
rect 29736 25638 29788 25644
rect 29644 24812 29696 24818
rect 29644 24754 29696 24760
rect 29644 24676 29696 24682
rect 29644 24618 29696 24624
rect 29368 24608 29420 24614
rect 29368 24550 29420 24556
rect 29276 24268 29328 24274
rect 29276 24210 29328 24216
rect 29288 24177 29316 24210
rect 29274 24168 29330 24177
rect 29274 24103 29330 24112
rect 29276 24064 29328 24070
rect 29182 24032 29238 24041
rect 29276 24006 29328 24012
rect 29182 23967 29238 23976
rect 29104 23718 29224 23746
rect 29000 23656 29052 23662
rect 29092 23656 29144 23662
rect 29052 23616 29092 23644
rect 29000 23598 29052 23604
rect 29092 23598 29144 23604
rect 29196 23508 29224 23718
rect 29012 23480 29224 23508
rect 29012 23361 29040 23480
rect 28998 23352 29054 23361
rect 28998 23287 29054 23296
rect 29182 23352 29238 23361
rect 29182 23287 29238 23296
rect 29000 21888 29052 21894
rect 29000 21830 29052 21836
rect 29012 20806 29040 21830
rect 29000 20800 29052 20806
rect 29000 20742 29052 20748
rect 29012 18698 29040 20742
rect 29092 20052 29144 20058
rect 29092 19994 29144 20000
rect 29104 19378 29132 19994
rect 29092 19372 29144 19378
rect 29092 19314 29144 19320
rect 29000 18692 29052 18698
rect 29000 18634 29052 18640
rect 29196 16726 29224 23287
rect 29288 23225 29316 24006
rect 29380 23730 29408 24550
rect 29552 24132 29604 24138
rect 29552 24074 29604 24080
rect 29564 24041 29592 24074
rect 29550 24032 29606 24041
rect 29550 23967 29606 23976
rect 29368 23724 29420 23730
rect 29368 23666 29420 23672
rect 29552 23724 29604 23730
rect 29552 23666 29604 23672
rect 29564 23304 29592 23666
rect 29472 23276 29592 23304
rect 29274 23216 29330 23225
rect 29274 23151 29330 23160
rect 29472 23118 29500 23276
rect 29552 23180 29604 23186
rect 29552 23122 29604 23128
rect 29460 23112 29512 23118
rect 29460 23054 29512 23060
rect 29564 22642 29592 23122
rect 29552 22636 29604 22642
rect 29552 22578 29604 22584
rect 29564 21554 29592 22578
rect 29552 21548 29604 21554
rect 29552 21490 29604 21496
rect 29552 21344 29604 21350
rect 29552 21286 29604 21292
rect 29460 20528 29512 20534
rect 29460 20470 29512 20476
rect 29276 20324 29328 20330
rect 29276 20266 29328 20272
rect 29288 19514 29316 20266
rect 29472 19514 29500 20470
rect 29564 20466 29592 21286
rect 29552 20460 29604 20466
rect 29552 20402 29604 20408
rect 29276 19508 29328 19514
rect 29276 19450 29328 19456
rect 29460 19508 29512 19514
rect 29460 19450 29512 19456
rect 29368 18216 29420 18222
rect 29368 18158 29420 18164
rect 29276 18080 29328 18086
rect 29276 18022 29328 18028
rect 29288 17882 29316 18022
rect 29276 17876 29328 17882
rect 29276 17818 29328 17824
rect 29288 17270 29316 17818
rect 29380 17542 29408 18158
rect 29552 17876 29604 17882
rect 29552 17818 29604 17824
rect 29460 17808 29512 17814
rect 29460 17750 29512 17756
rect 29368 17536 29420 17542
rect 29368 17478 29420 17484
rect 29380 17338 29408 17478
rect 29368 17332 29420 17338
rect 29368 17274 29420 17280
rect 29276 17264 29328 17270
rect 29276 17206 29328 17212
rect 29184 16720 29236 16726
rect 29184 16662 29236 16668
rect 29472 16114 29500 17750
rect 29564 17678 29592 17818
rect 29552 17672 29604 17678
rect 29552 17614 29604 17620
rect 29460 16108 29512 16114
rect 29460 16050 29512 16056
rect 29564 15502 29592 17614
rect 29552 15496 29604 15502
rect 29552 15438 29604 15444
rect 29000 15360 29052 15366
rect 29000 15302 29052 15308
rect 29012 15094 29040 15302
rect 29000 15088 29052 15094
rect 29000 15030 29052 15036
rect 29012 14482 29040 15030
rect 29092 14816 29144 14822
rect 29092 14758 29144 14764
rect 29104 14618 29132 14758
rect 29092 14612 29144 14618
rect 29092 14554 29144 14560
rect 29000 14476 29052 14482
rect 29000 14418 29052 14424
rect 29092 14408 29144 14414
rect 29092 14350 29144 14356
rect 29104 13870 29132 14350
rect 29092 13864 29144 13870
rect 29092 13806 29144 13812
rect 29104 12918 29132 13806
rect 29092 12912 29144 12918
rect 29092 12854 29144 12860
rect 29276 12368 29328 12374
rect 29276 12310 29328 12316
rect 29288 11898 29316 12310
rect 29276 11892 29328 11898
rect 29276 11834 29328 11840
rect 29000 11008 29052 11014
rect 29000 10950 29052 10956
rect 29012 5302 29040 10950
rect 29460 9104 29512 9110
rect 29460 9046 29512 9052
rect 29472 8634 29500 9046
rect 29656 8786 29684 24618
rect 29748 23594 29776 25638
rect 29736 23588 29788 23594
rect 29736 23530 29788 23536
rect 29736 20596 29788 20602
rect 29736 20538 29788 20544
rect 29748 20262 29776 20538
rect 29736 20256 29788 20262
rect 29736 20198 29788 20204
rect 29736 18760 29788 18766
rect 29736 18702 29788 18708
rect 29748 17218 29776 18702
rect 29840 18086 29868 28902
rect 30196 27464 30248 27470
rect 30196 27406 30248 27412
rect 30010 26752 30066 26761
rect 30010 26687 30066 26696
rect 30024 26450 30052 26687
rect 30104 26512 30156 26518
rect 30102 26480 30104 26489
rect 30156 26480 30158 26489
rect 30012 26444 30064 26450
rect 30208 26450 30236 27406
rect 30288 26988 30340 26994
rect 30288 26930 30340 26936
rect 30102 26415 30158 26424
rect 30196 26444 30248 26450
rect 30012 26386 30064 26392
rect 30196 26386 30248 26392
rect 30104 25832 30156 25838
rect 30102 25800 30104 25809
rect 30156 25800 30158 25809
rect 30102 25735 30158 25744
rect 30012 25356 30064 25362
rect 30012 25298 30064 25304
rect 30024 25158 30052 25298
rect 30012 25152 30064 25158
rect 30012 25094 30064 25100
rect 30024 24886 30052 25094
rect 30012 24880 30064 24886
rect 30012 24822 30064 24828
rect 30208 24750 30236 26386
rect 30300 25974 30328 26930
rect 30288 25968 30340 25974
rect 30288 25910 30340 25916
rect 30288 25832 30340 25838
rect 30288 25774 30340 25780
rect 30104 24744 30156 24750
rect 30104 24686 30156 24692
rect 30196 24744 30248 24750
rect 30196 24686 30248 24692
rect 30116 24342 30144 24686
rect 30104 24336 30156 24342
rect 30104 24278 30156 24284
rect 30012 23792 30064 23798
rect 30012 23734 30064 23740
rect 30024 23594 30052 23734
rect 30012 23588 30064 23594
rect 30012 23530 30064 23536
rect 30104 23520 30156 23526
rect 30102 23488 30104 23497
rect 30156 23488 30158 23497
rect 30102 23423 30158 23432
rect 30012 23248 30064 23254
rect 30012 23190 30064 23196
rect 29920 20868 29972 20874
rect 29920 20810 29972 20816
rect 29932 20602 29960 20810
rect 29920 20596 29972 20602
rect 29920 20538 29972 20544
rect 30024 18290 30052 23190
rect 30208 21622 30236 24686
rect 30300 23730 30328 25774
rect 30288 23724 30340 23730
rect 30288 23666 30340 23672
rect 30300 23254 30328 23666
rect 30288 23248 30340 23254
rect 30288 23190 30340 23196
rect 30392 22166 30420 29106
rect 30472 26988 30524 26994
rect 30472 26930 30524 26936
rect 30484 26790 30512 26930
rect 30748 26920 30800 26926
rect 30748 26862 30800 26868
rect 30472 26784 30524 26790
rect 30472 26726 30524 26732
rect 30484 25770 30512 26726
rect 30760 26353 30788 26862
rect 30746 26344 30802 26353
rect 30746 26279 30802 26288
rect 30760 25974 30788 26279
rect 30748 25968 30800 25974
rect 30748 25910 30800 25916
rect 30472 25764 30524 25770
rect 30472 25706 30524 25712
rect 30472 25288 30524 25294
rect 30524 25248 30604 25276
rect 30472 25230 30524 25236
rect 30472 25152 30524 25158
rect 30472 25094 30524 25100
rect 30484 24818 30512 25094
rect 30472 24812 30524 24818
rect 30472 24754 30524 24760
rect 30576 24274 30604 25248
rect 30840 25220 30892 25226
rect 30840 25162 30892 25168
rect 30852 24818 30880 25162
rect 30840 24812 30892 24818
rect 30840 24754 30892 24760
rect 30564 24268 30616 24274
rect 30564 24210 30616 24216
rect 30472 24064 30524 24070
rect 30472 24006 30524 24012
rect 30484 23322 30512 24006
rect 30576 23526 30604 24210
rect 30852 24138 30880 24754
rect 30840 24132 30892 24138
rect 30840 24074 30892 24080
rect 30932 24132 30984 24138
rect 30932 24074 30984 24080
rect 30564 23520 30616 23526
rect 30564 23462 30616 23468
rect 30472 23316 30524 23322
rect 30472 23258 30524 23264
rect 30656 22228 30708 22234
rect 30656 22170 30708 22176
rect 30380 22160 30432 22166
rect 30380 22102 30432 22108
rect 30472 21956 30524 21962
rect 30472 21898 30524 21904
rect 30196 21616 30248 21622
rect 30196 21558 30248 21564
rect 30380 20868 30432 20874
rect 30380 20810 30432 20816
rect 30392 20618 30420 20810
rect 30208 20590 30420 20618
rect 30208 20466 30236 20590
rect 30196 20460 30248 20466
rect 30196 20402 30248 20408
rect 30380 20460 30432 20466
rect 30380 20402 30432 20408
rect 30392 20058 30420 20402
rect 30380 20052 30432 20058
rect 30380 19994 30432 20000
rect 30012 18284 30064 18290
rect 30012 18226 30064 18232
rect 29828 18080 29880 18086
rect 29828 18022 29880 18028
rect 29828 17604 29880 17610
rect 29828 17546 29880 17552
rect 29840 17338 29868 17546
rect 29828 17332 29880 17338
rect 29828 17274 29880 17280
rect 29748 17190 29868 17218
rect 29736 16992 29788 16998
rect 29736 16934 29788 16940
rect 29748 11762 29776 16934
rect 29840 13870 29868 17190
rect 29920 17128 29972 17134
rect 29920 17070 29972 17076
rect 29828 13864 29880 13870
rect 29828 13806 29880 13812
rect 29736 11756 29788 11762
rect 29736 11698 29788 11704
rect 29840 10674 29868 13806
rect 29828 10668 29880 10674
rect 29828 10610 29880 10616
rect 29828 10464 29880 10470
rect 29828 10406 29880 10412
rect 29840 9994 29868 10406
rect 29828 9988 29880 9994
rect 29828 9930 29880 9936
rect 29656 8758 29868 8786
rect 29460 8628 29512 8634
rect 29460 8570 29512 8576
rect 29736 8492 29788 8498
rect 29736 8434 29788 8440
rect 29552 8356 29604 8362
rect 29552 8298 29604 8304
rect 29092 8288 29144 8294
rect 29092 8230 29144 8236
rect 29184 8288 29236 8294
rect 29184 8230 29236 8236
rect 29104 7478 29132 8230
rect 29196 8090 29224 8230
rect 29564 8090 29592 8298
rect 29184 8084 29236 8090
rect 29184 8026 29236 8032
rect 29552 8084 29604 8090
rect 29552 8026 29604 8032
rect 29644 7744 29696 7750
rect 29644 7686 29696 7692
rect 29092 7472 29144 7478
rect 29092 7414 29144 7420
rect 29000 5296 29052 5302
rect 29000 5238 29052 5244
rect 29552 4140 29604 4146
rect 29552 4082 29604 4088
rect 29564 3942 29592 4082
rect 29552 3936 29604 3942
rect 29552 3878 29604 3884
rect 29000 3528 29052 3534
rect 29000 3470 29052 3476
rect 29458 3496 29514 3505
rect 29012 3058 29040 3470
rect 29458 3431 29460 3440
rect 29512 3431 29514 3440
rect 29460 3402 29512 3408
rect 29000 3052 29052 3058
rect 29000 2994 29052 3000
rect 28908 2576 28960 2582
rect 28908 2518 28960 2524
rect 28448 1896 28500 1902
rect 28448 1838 28500 1844
rect 29656 800 29684 7686
rect 29748 7546 29776 8434
rect 29736 7540 29788 7546
rect 29736 7482 29788 7488
rect 29736 7200 29788 7206
rect 29736 7142 29788 7148
rect 29748 6866 29776 7142
rect 29736 6860 29788 6866
rect 29736 6802 29788 6808
rect 29840 5098 29868 8758
rect 29932 6322 29960 17070
rect 30024 13326 30052 18226
rect 30288 18080 30340 18086
rect 30288 18022 30340 18028
rect 30300 17202 30328 18022
rect 30288 17196 30340 17202
rect 30288 17138 30340 17144
rect 30380 16516 30432 16522
rect 30380 16458 30432 16464
rect 30392 16182 30420 16458
rect 30380 16176 30432 16182
rect 30380 16118 30432 16124
rect 30104 15428 30156 15434
rect 30104 15370 30156 15376
rect 30116 15094 30144 15370
rect 30104 15088 30156 15094
rect 30104 15030 30156 15036
rect 30380 14952 30432 14958
rect 30380 14894 30432 14900
rect 30392 14346 30420 14894
rect 30380 14340 30432 14346
rect 30380 14282 30432 14288
rect 30392 13870 30420 14282
rect 30380 13864 30432 13870
rect 30380 13806 30432 13812
rect 30012 13320 30064 13326
rect 30012 13262 30064 13268
rect 30024 11150 30052 13262
rect 30288 11756 30340 11762
rect 30288 11698 30340 11704
rect 30012 11144 30064 11150
rect 30012 11086 30064 11092
rect 30300 11082 30328 11698
rect 30288 11076 30340 11082
rect 30288 11018 30340 11024
rect 30196 11008 30248 11014
rect 30196 10950 30248 10956
rect 30208 10674 30236 10950
rect 30196 10668 30248 10674
rect 30196 10610 30248 10616
rect 30380 10668 30432 10674
rect 30380 10610 30432 10616
rect 30288 10260 30340 10266
rect 30392 10248 30420 10610
rect 30340 10220 30420 10248
rect 30288 10202 30340 10208
rect 30196 10056 30248 10062
rect 30196 9998 30248 10004
rect 30208 8498 30236 9998
rect 30196 8492 30248 8498
rect 30196 8434 30248 8440
rect 30104 8084 30156 8090
rect 30104 8026 30156 8032
rect 30116 7886 30144 8026
rect 30104 7880 30156 7886
rect 30104 7822 30156 7828
rect 30288 7812 30340 7818
rect 30288 7754 30340 7760
rect 30300 7206 30328 7754
rect 30288 7200 30340 7206
rect 30288 7142 30340 7148
rect 30300 6934 30328 7142
rect 30288 6928 30340 6934
rect 30288 6870 30340 6876
rect 29920 6316 29972 6322
rect 29920 6258 29972 6264
rect 29828 5092 29880 5098
rect 29828 5034 29880 5040
rect 30380 4480 30432 4486
rect 30380 4422 30432 4428
rect 29736 4140 29788 4146
rect 29736 4082 29788 4088
rect 29748 3534 29776 4082
rect 30286 4040 30342 4049
rect 30286 3975 30342 3984
rect 30300 3670 30328 3975
rect 30288 3664 30340 3670
rect 30288 3606 30340 3612
rect 29736 3528 29788 3534
rect 29736 3470 29788 3476
rect 29920 3392 29972 3398
rect 29920 3334 29972 3340
rect 30012 3392 30064 3398
rect 30012 3334 30064 3340
rect 29932 3126 29960 3334
rect 30024 3194 30052 3334
rect 30012 3188 30064 3194
rect 30012 3130 30064 3136
rect 29920 3120 29972 3126
rect 29920 3062 29972 3068
rect 30288 2984 30340 2990
rect 30288 2926 30340 2932
rect 30300 800 30328 2926
rect 30392 2514 30420 4422
rect 30484 2650 30512 21898
rect 30668 21690 30696 22170
rect 30656 21684 30708 21690
rect 30656 21626 30708 21632
rect 30748 21684 30800 21690
rect 30748 21626 30800 21632
rect 30760 20806 30788 21626
rect 30748 20800 30800 20806
rect 30748 20742 30800 20748
rect 30564 20460 30616 20466
rect 30564 20402 30616 20408
rect 30576 20330 30604 20402
rect 30564 20324 30616 20330
rect 30564 20266 30616 20272
rect 30852 18766 30880 24074
rect 30944 23254 30972 24074
rect 30932 23248 30984 23254
rect 30932 23190 30984 23196
rect 30944 22642 30972 23190
rect 30932 22636 30984 22642
rect 30932 22578 30984 22584
rect 30932 22432 30984 22438
rect 30932 22374 30984 22380
rect 30944 21622 30972 22374
rect 31036 22030 31064 29464
rect 31404 29306 31432 31282
rect 31588 29850 31616 35022
rect 31680 35018 31708 36178
rect 32036 36168 32088 36174
rect 32036 36110 32088 36116
rect 32048 35766 32076 36110
rect 32036 35760 32088 35766
rect 32036 35702 32088 35708
rect 32048 35086 32076 35702
rect 32140 35630 32168 36654
rect 32220 35692 32272 35698
rect 32220 35634 32272 35640
rect 32128 35624 32180 35630
rect 32128 35566 32180 35572
rect 32036 35080 32088 35086
rect 32036 35022 32088 35028
rect 31668 35012 31720 35018
rect 31668 34954 31720 34960
rect 32036 34740 32088 34746
rect 32036 34682 32088 34688
rect 32048 34066 32076 34682
rect 32036 34060 32088 34066
rect 32036 34002 32088 34008
rect 31760 33992 31812 33998
rect 31760 33934 31812 33940
rect 31772 33590 31800 33934
rect 31760 33584 31812 33590
rect 31760 33526 31812 33532
rect 31668 32972 31720 32978
rect 31668 32914 31720 32920
rect 31680 32366 31708 32914
rect 31668 32360 31720 32366
rect 31668 32302 31720 32308
rect 31772 31822 31800 33526
rect 31944 33516 31996 33522
rect 31944 33458 31996 33464
rect 31956 32570 31984 33458
rect 32140 32978 32168 35566
rect 32232 35290 32260 35634
rect 32220 35284 32272 35290
rect 32220 35226 32272 35232
rect 32324 35170 32352 41386
rect 32232 35142 32352 35170
rect 32128 32972 32180 32978
rect 32128 32914 32180 32920
rect 31944 32564 31996 32570
rect 31944 32506 31996 32512
rect 32128 32564 32180 32570
rect 32128 32506 32180 32512
rect 32036 32224 32088 32230
rect 32036 32166 32088 32172
rect 32140 32178 32168 32506
rect 32232 32348 32260 35142
rect 32312 32904 32364 32910
rect 32312 32846 32364 32852
rect 32324 32502 32352 32846
rect 32404 32836 32456 32842
rect 32404 32778 32456 32784
rect 32312 32496 32364 32502
rect 32312 32438 32364 32444
rect 32232 32320 32352 32348
rect 32048 32042 32076 32166
rect 32140 32150 32260 32178
rect 32048 32014 32168 32042
rect 32036 31952 32088 31958
rect 32036 31894 32088 31900
rect 31760 31816 31812 31822
rect 31812 31764 31892 31770
rect 31760 31758 31892 31764
rect 31772 31726 31892 31758
rect 31576 29844 31628 29850
rect 31576 29786 31628 29792
rect 31772 29578 31800 31726
rect 32048 31278 32076 31894
rect 32140 31754 32168 32014
rect 32128 31748 32180 31754
rect 32128 31690 32180 31696
rect 32036 31272 32088 31278
rect 32036 31214 32088 31220
rect 31760 29572 31812 29578
rect 31760 29514 31812 29520
rect 31392 29300 31444 29306
rect 31392 29242 31444 29248
rect 31772 28694 31800 29514
rect 32232 28762 32260 32150
rect 32324 31754 32352 32320
rect 32416 31958 32444 32778
rect 32508 32570 32536 47534
rect 32588 37120 32640 37126
rect 32588 37062 32640 37068
rect 32600 36242 32628 37062
rect 33508 36576 33560 36582
rect 33508 36518 33560 36524
rect 32588 36236 32640 36242
rect 32588 36178 32640 36184
rect 33520 36174 33548 36518
rect 33508 36168 33560 36174
rect 33508 36110 33560 36116
rect 33508 35488 33560 35494
rect 33508 35430 33560 35436
rect 33520 35154 33548 35430
rect 33508 35148 33560 35154
rect 33508 35090 33560 35096
rect 32680 35080 32732 35086
rect 32680 35022 32732 35028
rect 32692 34746 32720 35022
rect 32680 34740 32732 34746
rect 32680 34682 32732 34688
rect 32864 33312 32916 33318
rect 32864 33254 32916 33260
rect 32588 32972 32640 32978
rect 32588 32914 32640 32920
rect 32600 32570 32628 32914
rect 32496 32564 32548 32570
rect 32496 32506 32548 32512
rect 32588 32564 32640 32570
rect 32588 32506 32640 32512
rect 32600 32434 32628 32506
rect 32588 32428 32640 32434
rect 32588 32370 32640 32376
rect 32496 32360 32548 32366
rect 32496 32302 32548 32308
rect 32404 31952 32456 31958
rect 32404 31894 32456 31900
rect 32324 31726 32444 31754
rect 32220 28756 32272 28762
rect 32220 28698 32272 28704
rect 31760 28688 31812 28694
rect 31760 28630 31812 28636
rect 31852 28484 31904 28490
rect 31852 28426 31904 28432
rect 31576 28416 31628 28422
rect 31576 28358 31628 28364
rect 31588 28082 31616 28358
rect 31576 28076 31628 28082
rect 31576 28018 31628 28024
rect 31864 27946 31892 28426
rect 31852 27940 31904 27946
rect 31852 27882 31904 27888
rect 31944 27940 31996 27946
rect 31944 27882 31996 27888
rect 31956 27402 31984 27882
rect 32128 27872 32180 27878
rect 32128 27814 32180 27820
rect 32140 27470 32168 27814
rect 32232 27606 32260 28698
rect 32312 28076 32364 28082
rect 32312 28018 32364 28024
rect 32324 27674 32352 28018
rect 32312 27668 32364 27674
rect 32312 27610 32364 27616
rect 32220 27600 32272 27606
rect 32220 27542 32272 27548
rect 32128 27464 32180 27470
rect 32128 27406 32180 27412
rect 31944 27396 31996 27402
rect 31944 27338 31996 27344
rect 32416 26874 32444 31726
rect 32508 31482 32536 32302
rect 32496 31476 32548 31482
rect 32496 31418 32548 31424
rect 32876 31346 32904 33254
rect 33232 31884 33284 31890
rect 33232 31826 33284 31832
rect 32956 31816 33008 31822
rect 32956 31758 33008 31764
rect 32968 31686 32996 31758
rect 32956 31680 33008 31686
rect 32956 31622 33008 31628
rect 33048 31680 33100 31686
rect 33048 31622 33100 31628
rect 32588 31340 32640 31346
rect 32588 31282 32640 31288
rect 32864 31340 32916 31346
rect 32864 31282 32916 31288
rect 32600 31249 32628 31282
rect 32586 31240 32642 31249
rect 32586 31175 32642 31184
rect 32956 29844 33008 29850
rect 32956 29786 33008 29792
rect 32588 29300 32640 29306
rect 32588 29242 32640 29248
rect 32600 27402 32628 29242
rect 32968 28558 32996 29786
rect 32956 28552 33008 28558
rect 32956 28494 33008 28500
rect 32680 28484 32732 28490
rect 32680 28426 32732 28432
rect 32692 27470 32720 28426
rect 33060 27614 33088 31622
rect 33244 31346 33272 31826
rect 33600 31816 33652 31822
rect 33598 31784 33600 31793
rect 33652 31784 33654 31793
rect 33598 31719 33654 31728
rect 33232 31340 33284 31346
rect 33232 31282 33284 31288
rect 33600 28416 33652 28422
rect 33600 28358 33652 28364
rect 33232 27872 33284 27878
rect 33232 27814 33284 27820
rect 33244 27674 33272 27814
rect 32772 27600 32824 27606
rect 32772 27542 32824 27548
rect 32876 27586 33088 27614
rect 33232 27668 33284 27674
rect 33232 27610 33284 27616
rect 32680 27464 32732 27470
rect 32680 27406 32732 27412
rect 32588 27396 32640 27402
rect 32588 27338 32640 27344
rect 32324 26846 32444 26874
rect 31300 26240 31352 26246
rect 31300 26182 31352 26188
rect 31208 24608 31260 24614
rect 31208 24550 31260 24556
rect 31116 23044 31168 23050
rect 31116 22986 31168 22992
rect 31024 22024 31076 22030
rect 31024 21966 31076 21972
rect 31128 21690 31156 22986
rect 31116 21684 31168 21690
rect 31116 21626 31168 21632
rect 30932 21616 30984 21622
rect 30932 21558 30984 21564
rect 31220 20874 31248 24550
rect 31312 22094 31340 26182
rect 31392 25220 31444 25226
rect 31392 25162 31444 25168
rect 32128 25220 32180 25226
rect 32128 25162 32180 25168
rect 31404 24614 31432 25162
rect 31392 24608 31444 24614
rect 31392 24550 31444 24556
rect 32140 24342 32168 25162
rect 32220 24880 32272 24886
rect 32220 24822 32272 24828
rect 32128 24336 32180 24342
rect 32128 24278 32180 24284
rect 32232 24206 32260 24822
rect 32220 24200 32272 24206
rect 32220 24142 32272 24148
rect 31668 24132 31720 24138
rect 31668 24074 31720 24080
rect 31852 24132 31904 24138
rect 31852 24074 31904 24080
rect 31680 23798 31708 24074
rect 31668 23792 31720 23798
rect 31668 23734 31720 23740
rect 31392 22976 31444 22982
rect 31392 22918 31444 22924
rect 31404 22642 31432 22918
rect 31484 22704 31536 22710
rect 31668 22704 31720 22710
rect 31536 22664 31668 22692
rect 31484 22646 31536 22652
rect 31668 22646 31720 22652
rect 31392 22636 31444 22642
rect 31392 22578 31444 22584
rect 31576 22160 31628 22166
rect 31576 22102 31628 22108
rect 31312 22066 31524 22094
rect 31300 20936 31352 20942
rect 31300 20878 31352 20884
rect 31208 20868 31260 20874
rect 31208 20810 31260 20816
rect 30932 20800 30984 20806
rect 30932 20742 30984 20748
rect 30944 19786 30972 20742
rect 31312 20262 31340 20878
rect 31496 20330 31524 22066
rect 31484 20324 31536 20330
rect 31484 20266 31536 20272
rect 31300 20256 31352 20262
rect 31300 20198 31352 20204
rect 30932 19780 30984 19786
rect 30932 19722 30984 19728
rect 31024 19780 31076 19786
rect 31024 19722 31076 19728
rect 31036 19378 31064 19722
rect 31024 19372 31076 19378
rect 31024 19314 31076 19320
rect 30840 18760 30892 18766
rect 30840 18702 30892 18708
rect 30852 17270 30880 18702
rect 30932 18692 30984 18698
rect 30932 18634 30984 18640
rect 30944 18426 30972 18634
rect 30932 18420 30984 18426
rect 30932 18362 30984 18368
rect 30840 17264 30892 17270
rect 30840 17206 30892 17212
rect 31312 17202 31340 20198
rect 31484 17604 31536 17610
rect 31484 17546 31536 17552
rect 31300 17196 31352 17202
rect 31300 17138 31352 17144
rect 30840 17128 30892 17134
rect 30840 17070 30892 17076
rect 30564 16108 30616 16114
rect 30564 16050 30616 16056
rect 30748 16108 30800 16114
rect 30748 16050 30800 16056
rect 30576 15706 30604 16050
rect 30656 15904 30708 15910
rect 30656 15846 30708 15852
rect 30564 15700 30616 15706
rect 30564 15642 30616 15648
rect 30668 15502 30696 15846
rect 30564 15496 30616 15502
rect 30564 15438 30616 15444
rect 30656 15496 30708 15502
rect 30656 15438 30708 15444
rect 30576 13530 30604 15438
rect 30656 15360 30708 15366
rect 30656 15302 30708 15308
rect 30564 13524 30616 13530
rect 30564 13466 30616 13472
rect 30564 10804 30616 10810
rect 30564 10746 30616 10752
rect 30576 10674 30604 10746
rect 30564 10668 30616 10674
rect 30564 10610 30616 10616
rect 30668 8974 30696 15302
rect 30760 15162 30788 16050
rect 30748 15156 30800 15162
rect 30748 15098 30800 15104
rect 30852 12238 30880 17070
rect 30932 16720 30984 16726
rect 30932 16662 30984 16668
rect 30840 12232 30892 12238
rect 30840 12174 30892 12180
rect 30944 10470 30972 16662
rect 31496 16590 31524 17546
rect 31484 16584 31536 16590
rect 31484 16526 31536 16532
rect 31024 16176 31076 16182
rect 31024 16118 31076 16124
rect 31036 15094 31064 16118
rect 31484 16040 31536 16046
rect 31484 15982 31536 15988
rect 31496 15094 31524 15982
rect 31024 15088 31076 15094
rect 31484 15088 31536 15094
rect 31076 15048 31156 15076
rect 31024 15030 31076 15036
rect 31128 14482 31156 15048
rect 31484 15030 31536 15036
rect 31392 15020 31444 15026
rect 31392 14962 31444 14968
rect 31208 14816 31260 14822
rect 31208 14758 31260 14764
rect 31220 14550 31248 14758
rect 31404 14618 31432 14962
rect 31392 14612 31444 14618
rect 31392 14554 31444 14560
rect 31208 14544 31260 14550
rect 31208 14486 31260 14492
rect 31116 14476 31168 14482
rect 31116 14418 31168 14424
rect 31024 13796 31076 13802
rect 31024 13738 31076 13744
rect 31036 11830 31064 13738
rect 31128 13394 31156 14418
rect 31220 14346 31248 14486
rect 31208 14340 31260 14346
rect 31208 14282 31260 14288
rect 31588 14006 31616 22102
rect 31680 20942 31708 22646
rect 31760 21004 31812 21010
rect 31760 20946 31812 20952
rect 31668 20936 31720 20942
rect 31668 20878 31720 20884
rect 31680 20602 31708 20878
rect 31668 20596 31720 20602
rect 31668 20538 31720 20544
rect 31668 19168 31720 19174
rect 31668 19110 31720 19116
rect 31680 18698 31708 19110
rect 31772 18766 31800 20946
rect 31760 18760 31812 18766
rect 31760 18702 31812 18708
rect 31668 18692 31720 18698
rect 31668 18634 31720 18640
rect 31680 18290 31708 18634
rect 31772 18290 31800 18702
rect 31864 18306 31892 24074
rect 31944 23112 31996 23118
rect 31944 23054 31996 23060
rect 31956 21350 31984 23054
rect 32036 23044 32088 23050
rect 32036 22986 32088 22992
rect 32048 22234 32076 22986
rect 32128 22500 32180 22506
rect 32128 22442 32180 22448
rect 32036 22228 32088 22234
rect 32036 22170 32088 22176
rect 32140 21554 32168 22442
rect 32220 22432 32272 22438
rect 32220 22374 32272 22380
rect 32232 21962 32260 22374
rect 32220 21956 32272 21962
rect 32220 21898 32272 21904
rect 32128 21548 32180 21554
rect 32128 21490 32180 21496
rect 32140 21434 32168 21490
rect 32048 21406 32168 21434
rect 31944 21344 31996 21350
rect 31944 21286 31996 21292
rect 31956 19854 31984 21286
rect 31944 19848 31996 19854
rect 31944 19790 31996 19796
rect 31668 18284 31720 18290
rect 31668 18226 31720 18232
rect 31760 18284 31812 18290
rect 31864 18278 31984 18306
rect 31760 18226 31812 18232
rect 31772 17882 31800 18226
rect 31852 18216 31904 18222
rect 31852 18158 31904 18164
rect 31760 17876 31812 17882
rect 31760 17818 31812 17824
rect 31864 17270 31892 18158
rect 31852 17264 31904 17270
rect 31852 17206 31904 17212
rect 31668 16584 31720 16590
rect 31668 16526 31720 16532
rect 31680 15910 31708 16526
rect 31956 16266 31984 18278
rect 32048 17746 32076 21406
rect 32324 18970 32352 26846
rect 32680 26580 32732 26586
rect 32680 26522 32732 26528
rect 32404 24812 32456 24818
rect 32404 24754 32456 24760
rect 32416 23730 32444 24754
rect 32692 24750 32720 26522
rect 32784 26450 32812 27542
rect 32772 26444 32824 26450
rect 32772 26386 32824 26392
rect 32772 25832 32824 25838
rect 32772 25774 32824 25780
rect 32784 24954 32812 25774
rect 32876 25106 32904 27586
rect 33230 27024 33286 27033
rect 33230 26959 33286 26968
rect 33244 26858 33272 26959
rect 33232 26852 33284 26858
rect 33232 26794 33284 26800
rect 32956 26444 33008 26450
rect 32956 26386 33008 26392
rect 32968 25906 32996 26386
rect 32956 25900 33008 25906
rect 32956 25842 33008 25848
rect 33140 25900 33192 25906
rect 33140 25842 33192 25848
rect 33321 25900 33373 25906
rect 33321 25842 33373 25848
rect 33152 25265 33180 25842
rect 33138 25256 33194 25265
rect 33336 25226 33364 25842
rect 33508 25696 33560 25702
rect 33508 25638 33560 25644
rect 33138 25191 33194 25200
rect 33324 25220 33376 25226
rect 33324 25162 33376 25168
rect 32876 25078 32996 25106
rect 32772 24948 32824 24954
rect 32772 24890 32824 24896
rect 32680 24744 32732 24750
rect 32680 24686 32732 24692
rect 32692 24274 32720 24686
rect 32680 24268 32732 24274
rect 32680 24210 32732 24216
rect 32864 24132 32916 24138
rect 32864 24074 32916 24080
rect 32876 23798 32904 24074
rect 32864 23792 32916 23798
rect 32864 23734 32916 23740
rect 32404 23724 32456 23730
rect 32404 23666 32456 23672
rect 32496 23316 32548 23322
rect 32496 23258 32548 23264
rect 32508 22642 32536 23258
rect 32680 22976 32732 22982
rect 32680 22918 32732 22924
rect 32692 22642 32720 22918
rect 32864 22772 32916 22778
rect 32864 22714 32916 22720
rect 32876 22642 32904 22714
rect 32496 22636 32548 22642
rect 32496 22578 32548 22584
rect 32680 22636 32732 22642
rect 32680 22578 32732 22584
rect 32864 22636 32916 22642
rect 32864 22578 32916 22584
rect 32404 22568 32456 22574
rect 32404 22510 32456 22516
rect 32416 20058 32444 22510
rect 32508 22506 32536 22578
rect 32496 22500 32548 22506
rect 32496 22442 32548 22448
rect 32588 22024 32640 22030
rect 32586 21992 32588 22001
rect 32640 21992 32642 22001
rect 32586 21927 32642 21936
rect 32772 21480 32824 21486
rect 32772 21422 32824 21428
rect 32784 21010 32812 21422
rect 32772 21004 32824 21010
rect 32772 20946 32824 20952
rect 32404 20052 32456 20058
rect 32404 19994 32456 20000
rect 32312 18964 32364 18970
rect 32312 18906 32364 18912
rect 32324 18290 32352 18906
rect 32128 18284 32180 18290
rect 32128 18226 32180 18232
rect 32312 18284 32364 18290
rect 32312 18226 32364 18232
rect 32036 17740 32088 17746
rect 32036 17682 32088 17688
rect 31864 16238 31984 16266
rect 31668 15904 31720 15910
rect 31668 15846 31720 15852
rect 31680 15026 31708 15846
rect 31668 15020 31720 15026
rect 31668 14962 31720 14968
rect 31576 14000 31628 14006
rect 31576 13942 31628 13948
rect 31668 13524 31720 13530
rect 31668 13466 31720 13472
rect 31116 13388 31168 13394
rect 31116 13330 31168 13336
rect 31576 13252 31628 13258
rect 31576 13194 31628 13200
rect 31588 12238 31616 13194
rect 31680 12850 31708 13466
rect 31864 13394 31892 16238
rect 31944 16108 31996 16114
rect 31944 16050 31996 16056
rect 31956 15706 31984 16050
rect 31944 15700 31996 15706
rect 31944 15642 31996 15648
rect 31852 13388 31904 13394
rect 31852 13330 31904 13336
rect 32048 12918 32076 17682
rect 32140 17610 32168 18226
rect 32864 18216 32916 18222
rect 32864 18158 32916 18164
rect 32876 17882 32904 18158
rect 32864 17876 32916 17882
rect 32864 17818 32916 17824
rect 32128 17604 32180 17610
rect 32128 17546 32180 17552
rect 32128 16516 32180 16522
rect 32128 16458 32180 16464
rect 32140 16250 32168 16458
rect 32588 16448 32640 16454
rect 32588 16390 32640 16396
rect 32128 16244 32180 16250
rect 32128 16186 32180 16192
rect 32600 16114 32628 16390
rect 32588 16108 32640 16114
rect 32588 16050 32640 16056
rect 32220 13864 32272 13870
rect 32220 13806 32272 13812
rect 32232 13326 32260 13806
rect 32496 13728 32548 13734
rect 32496 13670 32548 13676
rect 32508 13394 32536 13670
rect 32312 13388 32364 13394
rect 32312 13330 32364 13336
rect 32496 13388 32548 13394
rect 32496 13330 32548 13336
rect 32220 13320 32272 13326
rect 32220 13262 32272 13268
rect 32036 12912 32088 12918
rect 32036 12854 32088 12860
rect 31668 12844 31720 12850
rect 31668 12786 31720 12792
rect 32220 12844 32272 12850
rect 32220 12786 32272 12792
rect 31576 12232 31628 12238
rect 31576 12174 31628 12180
rect 31300 12164 31352 12170
rect 31300 12106 31352 12112
rect 31024 11824 31076 11830
rect 31024 11766 31076 11772
rect 31312 11762 31340 12106
rect 31300 11756 31352 11762
rect 31300 11698 31352 11704
rect 30932 10464 30984 10470
rect 30932 10406 30984 10412
rect 31024 9988 31076 9994
rect 31024 9930 31076 9936
rect 30932 9920 30984 9926
rect 30932 9862 30984 9868
rect 30944 9586 30972 9862
rect 31036 9722 31064 9930
rect 31312 9722 31340 11698
rect 31484 11620 31536 11626
rect 31484 11562 31536 11568
rect 31496 9722 31524 11562
rect 31576 11144 31628 11150
rect 31680 11132 31708 12786
rect 32128 12708 32180 12714
rect 32128 12650 32180 12656
rect 32140 12170 32168 12650
rect 32232 12442 32260 12786
rect 32324 12646 32352 13330
rect 32312 12640 32364 12646
rect 32312 12582 32364 12588
rect 32220 12436 32272 12442
rect 32220 12378 32272 12384
rect 32324 12238 32352 12582
rect 32968 12434 32996 25078
rect 33520 24886 33548 25638
rect 33612 25401 33640 28358
rect 33598 25392 33654 25401
rect 33598 25327 33654 25336
rect 33600 25288 33652 25294
rect 33600 25230 33652 25236
rect 33508 24880 33560 24886
rect 33508 24822 33560 24828
rect 33324 24812 33376 24818
rect 33324 24754 33376 24760
rect 33048 23724 33100 23730
rect 33048 23666 33100 23672
rect 33060 23322 33088 23666
rect 33336 23322 33364 24754
rect 33612 23866 33640 25230
rect 33600 23860 33652 23866
rect 33600 23802 33652 23808
rect 33048 23316 33100 23322
rect 33048 23258 33100 23264
rect 33324 23316 33376 23322
rect 33324 23258 33376 23264
rect 33140 22704 33192 22710
rect 33140 22646 33192 22652
rect 33048 21684 33100 21690
rect 33048 21626 33100 21632
rect 33060 21146 33088 21626
rect 33152 21554 33180 22646
rect 33336 22642 33364 23258
rect 33416 22772 33468 22778
rect 33416 22714 33468 22720
rect 33324 22636 33376 22642
rect 33324 22578 33376 22584
rect 33324 22432 33376 22438
rect 33324 22374 33376 22380
rect 33140 21548 33192 21554
rect 33140 21490 33192 21496
rect 33232 21548 33284 21554
rect 33232 21490 33284 21496
rect 33244 21162 33272 21490
rect 33152 21146 33272 21162
rect 33048 21140 33100 21146
rect 33048 21082 33100 21088
rect 33140 21140 33272 21146
rect 33192 21134 33272 21140
rect 33140 21082 33192 21088
rect 33336 20942 33364 22374
rect 33428 21554 33456 22714
rect 33416 21548 33468 21554
rect 33416 21490 33468 21496
rect 33324 20936 33376 20942
rect 33324 20878 33376 20884
rect 33140 20800 33192 20806
rect 33140 20742 33192 20748
rect 33152 20398 33180 20742
rect 33140 20392 33192 20398
rect 33140 20334 33192 20340
rect 33152 19854 33180 20334
rect 33140 19848 33192 19854
rect 33140 19790 33192 19796
rect 33428 19786 33456 21490
rect 33416 19780 33468 19786
rect 33416 19722 33468 19728
rect 33416 19508 33468 19514
rect 33416 19450 33468 19456
rect 33428 19378 33456 19450
rect 33416 19372 33468 19378
rect 33416 19314 33468 19320
rect 33600 19372 33652 19378
rect 33600 19314 33652 19320
rect 33508 19236 33560 19242
rect 33508 19178 33560 19184
rect 33140 19168 33192 19174
rect 33140 19110 33192 19116
rect 33048 18828 33100 18834
rect 33048 18770 33100 18776
rect 33060 17270 33088 18770
rect 33152 18358 33180 19110
rect 33520 18902 33548 19178
rect 33508 18896 33560 18902
rect 33508 18838 33560 18844
rect 33508 18760 33560 18766
rect 33508 18702 33560 18708
rect 33140 18352 33192 18358
rect 33140 18294 33192 18300
rect 33520 18154 33548 18702
rect 33508 18148 33560 18154
rect 33508 18090 33560 18096
rect 33612 17882 33640 19314
rect 33600 17876 33652 17882
rect 33600 17818 33652 17824
rect 33048 17264 33100 17270
rect 33048 17206 33100 17212
rect 33060 16658 33088 17206
rect 33232 16720 33284 16726
rect 33232 16662 33284 16668
rect 33048 16652 33100 16658
rect 33048 16594 33100 16600
rect 33060 16182 33088 16594
rect 33048 16176 33100 16182
rect 33048 16118 33100 16124
rect 33244 16114 33272 16662
rect 33416 16584 33468 16590
rect 33416 16526 33468 16532
rect 33232 16108 33284 16114
rect 33232 16050 33284 16056
rect 33140 14544 33192 14550
rect 33140 14486 33192 14492
rect 33048 14340 33100 14346
rect 33048 14282 33100 14288
rect 33060 13870 33088 14282
rect 33152 14006 33180 14486
rect 33140 14000 33192 14006
rect 33140 13942 33192 13948
rect 33048 13864 33100 13870
rect 33048 13806 33100 13812
rect 33244 12434 33272 16050
rect 33428 14822 33456 16526
rect 33600 16516 33652 16522
rect 33600 16458 33652 16464
rect 33508 16108 33560 16114
rect 33508 16050 33560 16056
rect 33416 14816 33468 14822
rect 33416 14758 33468 14764
rect 33520 14550 33548 16050
rect 33612 16046 33640 16458
rect 33600 16040 33652 16046
rect 33600 15982 33652 15988
rect 33508 14544 33560 14550
rect 33508 14486 33560 14492
rect 33508 14272 33560 14278
rect 33508 14214 33560 14220
rect 33520 14006 33548 14214
rect 33508 14000 33560 14006
rect 33508 13942 33560 13948
rect 33324 13932 33376 13938
rect 33324 13874 33376 13880
rect 32968 12406 33088 12434
rect 32312 12232 32364 12238
rect 32680 12232 32732 12238
rect 32312 12174 32364 12180
rect 32600 12192 32680 12220
rect 32128 12164 32180 12170
rect 32128 12106 32180 12112
rect 32140 11762 32168 12106
rect 32128 11756 32180 11762
rect 32128 11698 32180 11704
rect 31760 11552 31812 11558
rect 31760 11494 31812 11500
rect 31772 11150 31800 11494
rect 31628 11104 31708 11132
rect 31760 11144 31812 11150
rect 31576 11086 31628 11092
rect 31760 11086 31812 11092
rect 31588 10130 31616 11086
rect 31576 10124 31628 10130
rect 31576 10066 31628 10072
rect 31024 9716 31076 9722
rect 31024 9658 31076 9664
rect 31300 9716 31352 9722
rect 31300 9658 31352 9664
rect 31484 9716 31536 9722
rect 31484 9658 31536 9664
rect 30932 9580 30984 9586
rect 30932 9522 30984 9528
rect 31312 9110 31340 9658
rect 31300 9104 31352 9110
rect 31300 9046 31352 9052
rect 31496 8974 31524 9658
rect 32140 9586 32168 11698
rect 32600 10674 32628 12192
rect 32680 12174 32732 12180
rect 32864 11756 32916 11762
rect 32864 11698 32916 11704
rect 32876 11286 32904 11698
rect 32864 11280 32916 11286
rect 32864 11222 32916 11228
rect 32588 10668 32640 10674
rect 32588 10610 32640 10616
rect 32128 9580 32180 9586
rect 32128 9522 32180 9528
rect 30656 8968 30708 8974
rect 30656 8910 30708 8916
rect 31484 8968 31536 8974
rect 31484 8910 31536 8916
rect 30656 8832 30708 8838
rect 30656 8774 30708 8780
rect 30668 8566 30696 8774
rect 30656 8560 30708 8566
rect 30656 8502 30708 8508
rect 31496 8498 31524 8910
rect 31576 8628 31628 8634
rect 31576 8570 31628 8576
rect 31484 8492 31536 8498
rect 31484 8434 31536 8440
rect 31588 8430 31616 8570
rect 32140 8498 32168 9522
rect 32496 9036 32548 9042
rect 32496 8978 32548 8984
rect 32508 8634 32536 8978
rect 32496 8628 32548 8634
rect 32496 8570 32548 8576
rect 32128 8492 32180 8498
rect 32128 8434 32180 8440
rect 31576 8424 31628 8430
rect 31576 8366 31628 8372
rect 31588 7954 31616 8366
rect 32140 8090 32168 8434
rect 32128 8084 32180 8090
rect 32128 8026 32180 8032
rect 31576 7948 31628 7954
rect 31576 7890 31628 7896
rect 30932 7812 30984 7818
rect 30932 7754 30984 7760
rect 30944 7546 30972 7754
rect 30932 7540 30984 7546
rect 30932 7482 30984 7488
rect 32600 7410 32628 10610
rect 32956 10600 33008 10606
rect 32956 10542 33008 10548
rect 32968 10266 32996 10542
rect 32956 10260 33008 10266
rect 32956 10202 33008 10208
rect 32968 9654 32996 10202
rect 32956 9648 33008 9654
rect 32956 9590 33008 9596
rect 33060 8362 33088 12406
rect 33152 12406 33272 12434
rect 33152 12102 33180 12406
rect 33336 12238 33364 13874
rect 33704 13394 33732 49286
rect 34060 32768 34112 32774
rect 34060 32710 34112 32716
rect 33784 32564 33836 32570
rect 33784 32506 33836 32512
rect 33796 31754 33824 32506
rect 34072 31890 34100 32710
rect 34060 31884 34112 31890
rect 34060 31826 34112 31832
rect 33784 31748 33836 31754
rect 33784 31690 33836 31696
rect 33796 29714 33824 31690
rect 33784 29708 33836 29714
rect 33784 29650 33836 29656
rect 33876 29504 33928 29510
rect 33876 29446 33928 29452
rect 33888 28558 33916 29446
rect 34244 28960 34296 28966
rect 34164 28908 34244 28914
rect 34164 28902 34296 28908
rect 34164 28886 34284 28902
rect 34164 28558 34192 28886
rect 33876 28552 33928 28558
rect 33876 28494 33928 28500
rect 34152 28552 34204 28558
rect 34152 28494 34204 28500
rect 33888 28082 33916 28494
rect 33876 28076 33928 28082
rect 33876 28018 33928 28024
rect 34164 27962 34192 28494
rect 33796 27934 34192 27962
rect 33796 27130 33824 27934
rect 34060 27396 34112 27402
rect 34060 27338 34112 27344
rect 33784 27124 33836 27130
rect 33784 27066 33836 27072
rect 33874 26752 33930 26761
rect 33874 26687 33930 26696
rect 33888 26382 33916 26687
rect 33876 26376 33928 26382
rect 33876 26318 33928 26324
rect 33784 26308 33836 26314
rect 33784 26250 33836 26256
rect 33796 26194 33824 26250
rect 34072 26194 34100 27338
rect 33796 26166 34100 26194
rect 34072 25974 34100 26166
rect 34060 25968 34112 25974
rect 34060 25910 34112 25916
rect 33784 25900 33836 25906
rect 33784 25842 33836 25848
rect 33796 25294 33824 25842
rect 33784 25288 33836 25294
rect 33784 25230 33836 25236
rect 33796 24954 33824 25230
rect 33784 24948 33836 24954
rect 33784 24890 33836 24896
rect 33968 20392 34020 20398
rect 33968 20334 34020 20340
rect 33876 19304 33928 19310
rect 33876 19246 33928 19252
rect 33784 19168 33836 19174
rect 33784 19110 33836 19116
rect 33796 18766 33824 19110
rect 33784 18760 33836 18766
rect 33784 18702 33836 18708
rect 33888 17610 33916 19246
rect 33876 17604 33928 17610
rect 33876 17546 33928 17552
rect 33888 17270 33916 17546
rect 33876 17264 33928 17270
rect 33876 17206 33928 17212
rect 33876 16992 33928 16998
rect 33876 16934 33928 16940
rect 33888 16590 33916 16934
rect 33876 16584 33928 16590
rect 33876 16526 33928 16532
rect 33692 13388 33744 13394
rect 33692 13330 33744 13336
rect 33324 12232 33376 12238
rect 33324 12174 33376 12180
rect 33140 12096 33192 12102
rect 33140 12038 33192 12044
rect 33324 12096 33376 12102
rect 33324 12038 33376 12044
rect 33336 11830 33364 12038
rect 33324 11824 33376 11830
rect 33324 11766 33376 11772
rect 33048 8356 33100 8362
rect 33048 8298 33100 8304
rect 32588 7404 32640 7410
rect 32588 7346 32640 7352
rect 30932 4684 30984 4690
rect 30932 4626 30984 4632
rect 30656 4548 30708 4554
rect 30656 4490 30708 4496
rect 30668 3942 30696 4490
rect 30564 3936 30616 3942
rect 30564 3878 30616 3884
rect 30656 3936 30708 3942
rect 30656 3878 30708 3884
rect 30576 3466 30604 3878
rect 30564 3460 30616 3466
rect 30564 3402 30616 3408
rect 30472 2644 30524 2650
rect 30472 2586 30524 2592
rect 30380 2508 30432 2514
rect 30380 2450 30432 2456
rect 30944 800 30972 4626
rect 31392 3936 31444 3942
rect 31392 3878 31444 3884
rect 32772 3936 32824 3942
rect 32772 3878 32824 3884
rect 31404 3670 31432 3878
rect 32220 3732 32272 3738
rect 32220 3674 32272 3680
rect 31392 3664 31444 3670
rect 31392 3606 31444 3612
rect 31576 3596 31628 3602
rect 31576 3538 31628 3544
rect 31588 800 31616 3538
rect 32232 800 32260 3674
rect 32312 3664 32364 3670
rect 32312 3606 32364 3612
rect 32324 3505 32352 3606
rect 32310 3496 32366 3505
rect 32310 3431 32366 3440
rect 32784 3058 32812 3878
rect 33980 3738 34008 20334
rect 34152 20256 34204 20262
rect 34152 20198 34204 20204
rect 34060 19780 34112 19786
rect 34060 19722 34112 19728
rect 34072 19378 34100 19722
rect 34164 19446 34192 20198
rect 34152 19440 34204 19446
rect 34152 19382 34204 19388
rect 34060 19372 34112 19378
rect 34060 19314 34112 19320
rect 34060 18760 34112 18766
rect 34060 18702 34112 18708
rect 34072 16726 34100 18702
rect 34152 17672 34204 17678
rect 34152 17614 34204 17620
rect 34164 17202 34192 17614
rect 34152 17196 34204 17202
rect 34152 17138 34204 17144
rect 34060 16720 34112 16726
rect 34060 16662 34112 16668
rect 34164 16182 34192 17138
rect 34244 16448 34296 16454
rect 34244 16390 34296 16396
rect 34152 16176 34204 16182
rect 34152 16118 34204 16124
rect 34256 16114 34284 16390
rect 34244 16108 34296 16114
rect 34244 16050 34296 16056
rect 34152 15904 34204 15910
rect 34152 15846 34204 15852
rect 34164 15026 34192 15846
rect 34152 15020 34204 15026
rect 34152 14962 34204 14968
rect 34164 14550 34192 14962
rect 34152 14544 34204 14550
rect 34152 14486 34204 14492
rect 34164 13394 34192 14486
rect 34152 13388 34204 13394
rect 34152 13330 34204 13336
rect 34164 12850 34192 13330
rect 34152 12844 34204 12850
rect 34152 12786 34204 12792
rect 34348 11694 34376 51326
rect 34716 51326 34850 51354
rect 34716 47598 34744 51326
rect 34794 51200 34850 51326
rect 35438 51200 35494 52000
rect 36082 51200 36138 52000
rect 36726 51200 36782 52000
rect 37370 51354 37426 52000
rect 38014 51354 38070 52000
rect 38658 51354 38714 52000
rect 37370 51326 37688 51354
rect 37370 51200 37426 51326
rect 34934 49532 35242 49552
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49456 35242 49476
rect 34888 49224 34940 49230
rect 34888 49166 34940 49172
rect 34900 48754 34928 49166
rect 34888 48748 34940 48754
rect 34888 48690 34940 48696
rect 36096 48686 36124 51200
rect 36268 49224 36320 49230
rect 36268 49166 36320 49172
rect 36084 48680 36136 48686
rect 36084 48622 36136 48628
rect 35992 48544 36044 48550
rect 35992 48486 36044 48492
rect 34934 48444 35242 48464
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48368 35242 48388
rect 35808 48136 35860 48142
rect 35808 48078 35860 48084
rect 35820 47818 35848 48078
rect 35900 48000 35952 48006
rect 35900 47942 35952 47948
rect 35912 47818 35940 47942
rect 35820 47790 35940 47818
rect 36004 47802 36032 48486
rect 36280 48210 36308 49166
rect 36740 48210 36768 51200
rect 37660 48550 37688 51326
rect 38014 51326 38148 51354
rect 38014 51200 38070 51326
rect 38120 49230 38148 51326
rect 38658 51326 39160 51354
rect 38658 51200 38714 51326
rect 38108 49224 38160 49230
rect 38108 49166 38160 49172
rect 38292 49088 38344 49094
rect 38292 49030 38344 49036
rect 37648 48544 37700 48550
rect 37648 48486 37700 48492
rect 37280 48272 37332 48278
rect 37280 48214 37332 48220
rect 36268 48204 36320 48210
rect 36268 48146 36320 48152
rect 36728 48204 36780 48210
rect 36728 48146 36780 48152
rect 36544 48068 36596 48074
rect 36544 48010 36596 48016
rect 36452 48000 36504 48006
rect 36452 47942 36504 47948
rect 35992 47796 36044 47802
rect 35992 47738 36044 47744
rect 36464 47666 36492 47942
rect 36556 47802 36584 48010
rect 36544 47796 36596 47802
rect 36544 47738 36596 47744
rect 35808 47660 35860 47666
rect 35808 47602 35860 47608
rect 36452 47660 36504 47666
rect 36452 47602 36504 47608
rect 34704 47592 34756 47598
rect 34704 47534 34756 47540
rect 34934 47356 35242 47376
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47280 35242 47300
rect 35820 47190 35848 47602
rect 35808 47184 35860 47190
rect 35808 47126 35860 47132
rect 34934 46268 35242 46288
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46192 35242 46212
rect 34934 45180 35242 45200
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45104 35242 45124
rect 34934 44092 35242 44112
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44016 35242 44036
rect 36084 43784 36136 43790
rect 36084 43726 36136 43732
rect 34934 43004 35242 43024
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42928 35242 42948
rect 34934 41916 35242 41936
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41840 35242 41860
rect 36096 41414 36124 43726
rect 36464 43314 36492 47602
rect 37292 44946 37320 48214
rect 37280 44940 37332 44946
rect 37280 44882 37332 44888
rect 36544 43716 36596 43722
rect 36544 43658 36596 43664
rect 36556 43450 36584 43658
rect 36544 43444 36596 43450
rect 36544 43386 36596 43392
rect 36452 43308 36504 43314
rect 36452 43250 36504 43256
rect 36096 41386 36216 41414
rect 34934 40828 35242 40848
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40752 35242 40772
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 34612 37324 34664 37330
rect 34612 37266 34664 37272
rect 34520 29232 34572 29238
rect 34520 29174 34572 29180
rect 34532 27062 34560 29174
rect 34520 27056 34572 27062
rect 34520 26998 34572 27004
rect 34520 26920 34572 26926
rect 34520 26862 34572 26868
rect 34428 26784 34480 26790
rect 34426 26752 34428 26761
rect 34480 26752 34482 26761
rect 34426 26687 34482 26696
rect 34532 26450 34560 26862
rect 34520 26444 34572 26450
rect 34520 26386 34572 26392
rect 34532 25838 34560 26386
rect 34520 25832 34572 25838
rect 34520 25774 34572 25780
rect 34520 25696 34572 25702
rect 34520 25638 34572 25644
rect 34532 25430 34560 25638
rect 34520 25424 34572 25430
rect 34520 25366 34572 25372
rect 34520 24812 34572 24818
rect 34520 24754 34572 24760
rect 34532 23905 34560 24754
rect 34518 23896 34574 23905
rect 34518 23831 34574 23840
rect 34624 22094 34652 37266
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 35900 33108 35952 33114
rect 35900 33050 35952 33056
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 35912 31822 35940 33050
rect 35900 31816 35952 31822
rect 35952 31764 36032 31770
rect 35900 31758 36032 31764
rect 35912 31742 36032 31758
rect 35808 31680 35860 31686
rect 35808 31622 35860 31628
rect 35820 31278 35848 31622
rect 36004 31346 36032 31742
rect 35992 31340 36044 31346
rect 35992 31282 36044 31288
rect 35348 31272 35400 31278
rect 35808 31272 35860 31278
rect 35348 31214 35400 31220
rect 35622 31240 35678 31249
rect 35360 31142 35388 31214
rect 35808 31214 35860 31220
rect 35622 31175 35678 31184
rect 35636 31142 35664 31175
rect 35348 31136 35400 31142
rect 35348 31078 35400 31084
rect 35624 31136 35676 31142
rect 35624 31078 35676 31084
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 34796 29844 34848 29850
rect 34796 29786 34848 29792
rect 34704 29640 34756 29646
rect 34704 29582 34756 29588
rect 34716 29102 34744 29582
rect 34808 29238 34836 29786
rect 34888 29640 34940 29646
rect 34888 29582 34940 29588
rect 34796 29232 34848 29238
rect 34796 29174 34848 29180
rect 34704 29096 34756 29102
rect 34704 29038 34756 29044
rect 34716 28150 34744 29038
rect 34808 28966 34836 29174
rect 34900 29034 34928 29582
rect 34888 29028 34940 29034
rect 34888 28970 34940 28976
rect 34796 28960 34848 28966
rect 34796 28902 34848 28908
rect 34808 28490 34836 28902
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 34796 28484 34848 28490
rect 34796 28426 34848 28432
rect 35360 28370 35388 31078
rect 36004 30666 36032 31282
rect 35992 30660 36044 30666
rect 35992 30602 36044 30608
rect 35532 29164 35584 29170
rect 35532 29106 35584 29112
rect 34808 28342 35388 28370
rect 34704 28144 34756 28150
rect 34704 28086 34756 28092
rect 34704 26988 34756 26994
rect 34704 26930 34756 26936
rect 34716 26450 34744 26930
rect 34704 26444 34756 26450
rect 34704 26386 34756 26392
rect 34704 26240 34756 26246
rect 34702 26208 34704 26217
rect 34756 26208 34758 26217
rect 34702 26143 34758 26152
rect 34808 25702 34836 28342
rect 35544 28150 35572 29106
rect 35532 28144 35584 28150
rect 35532 28086 35584 28092
rect 35544 27985 35572 28086
rect 36004 28082 36032 30602
rect 35992 28076 36044 28082
rect 35992 28018 36044 28024
rect 35530 27976 35586 27985
rect 35530 27911 35586 27920
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 35808 27464 35860 27470
rect 35808 27406 35860 27412
rect 35164 27396 35216 27402
rect 35164 27338 35216 27344
rect 35624 27396 35676 27402
rect 35624 27338 35676 27344
rect 35176 26926 35204 27338
rect 35532 27328 35584 27334
rect 35532 27270 35584 27276
rect 35544 27169 35572 27270
rect 35530 27160 35586 27169
rect 35636 27130 35664 27338
rect 35530 27095 35586 27104
rect 35624 27124 35676 27130
rect 35624 27066 35676 27072
rect 35532 26988 35584 26994
rect 35532 26930 35584 26936
rect 35164 26920 35216 26926
rect 35164 26862 35216 26868
rect 35348 26852 35400 26858
rect 35348 26794 35400 26800
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 35360 26518 35388 26794
rect 35544 26586 35572 26930
rect 35532 26580 35584 26586
rect 35532 26522 35584 26528
rect 35072 26512 35124 26518
rect 35072 26454 35124 26460
rect 35348 26512 35400 26518
rect 35348 26454 35400 26460
rect 35084 26353 35112 26454
rect 35164 26376 35216 26382
rect 35070 26344 35126 26353
rect 35164 26318 35216 26324
rect 35070 26279 35126 26288
rect 35176 26217 35204 26318
rect 35532 26240 35584 26246
rect 35162 26208 35218 26217
rect 35532 26182 35584 26188
rect 35162 26143 35218 26152
rect 35440 25832 35492 25838
rect 35440 25774 35492 25780
rect 34796 25696 34848 25702
rect 34796 25638 34848 25644
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 35452 25226 35480 25774
rect 35544 25498 35572 26182
rect 35532 25492 35584 25498
rect 35532 25434 35584 25440
rect 35440 25220 35492 25226
rect 35440 25162 35492 25168
rect 34796 25152 34848 25158
rect 34796 25094 34848 25100
rect 34704 24744 34756 24750
rect 34704 24686 34756 24692
rect 34716 24274 34744 24686
rect 34704 24268 34756 24274
rect 34704 24210 34756 24216
rect 34532 22066 34652 22094
rect 34532 14498 34560 22066
rect 34716 22030 34744 24210
rect 34808 24206 34836 25094
rect 35532 24880 35584 24886
rect 35532 24822 35584 24828
rect 35348 24608 35400 24614
rect 35348 24550 35400 24556
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 34796 24200 34848 24206
rect 34796 24142 34848 24148
rect 34796 24064 34848 24070
rect 34796 24006 34848 24012
rect 34808 23118 34836 24006
rect 35360 23769 35388 24550
rect 35440 24200 35492 24206
rect 35440 24142 35492 24148
rect 35346 23760 35402 23769
rect 35346 23695 35402 23704
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 35452 23186 35480 24142
rect 35440 23180 35492 23186
rect 35440 23122 35492 23128
rect 34796 23112 34848 23118
rect 34796 23054 34848 23060
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 34704 22024 34756 22030
rect 34704 21966 34756 21972
rect 35348 21412 35400 21418
rect 35348 21354 35400 21360
rect 34796 21344 34848 21350
rect 34796 21286 34848 21292
rect 34808 20942 34836 21286
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 35360 20942 35388 21354
rect 34796 20936 34848 20942
rect 34796 20878 34848 20884
rect 35348 20936 35400 20942
rect 35348 20878 35400 20884
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 35348 18080 35400 18086
rect 35348 18022 35400 18028
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 35360 17610 35388 18022
rect 35348 17604 35400 17610
rect 35348 17546 35400 17552
rect 35544 17270 35572 24822
rect 35636 20602 35664 27066
rect 35820 27062 35848 27406
rect 35808 27056 35860 27062
rect 35808 26998 35860 27004
rect 36084 27056 36136 27062
rect 36084 26998 36136 27004
rect 35820 26382 35848 26998
rect 35808 26376 35860 26382
rect 36096 26353 36124 26998
rect 35808 26318 35860 26324
rect 36082 26344 36138 26353
rect 35820 25974 35848 26318
rect 36082 26279 36138 26288
rect 36096 25974 36124 26279
rect 35808 25968 35860 25974
rect 35808 25910 35860 25916
rect 36084 25968 36136 25974
rect 36084 25910 36136 25916
rect 35806 25528 35862 25537
rect 35806 25463 35808 25472
rect 35860 25463 35862 25472
rect 35808 25434 35860 25440
rect 35898 25256 35954 25265
rect 35808 25220 35860 25226
rect 35898 25191 35954 25200
rect 35808 25162 35860 25168
rect 35714 24712 35770 24721
rect 35714 24647 35770 24656
rect 35728 24342 35756 24647
rect 35716 24336 35768 24342
rect 35716 24278 35768 24284
rect 35820 23866 35848 25162
rect 35912 24954 35940 25191
rect 35900 24948 35952 24954
rect 35900 24890 35952 24896
rect 36188 24154 36216 41386
rect 36464 32570 36492 43250
rect 36452 32564 36504 32570
rect 36452 32506 36504 32512
rect 36360 32428 36412 32434
rect 36360 32370 36412 32376
rect 36372 31822 36400 32370
rect 37464 32360 37516 32366
rect 37464 32302 37516 32308
rect 37476 32026 37504 32302
rect 37464 32020 37516 32026
rect 37464 31962 37516 31968
rect 36360 31816 36412 31822
rect 36280 31764 36360 31770
rect 36280 31758 36412 31764
rect 36636 31816 36688 31822
rect 36636 31758 36688 31764
rect 37188 31816 37240 31822
rect 37188 31758 37240 31764
rect 36280 31742 36400 31758
rect 36280 31278 36308 31742
rect 36268 31272 36320 31278
rect 36268 31214 36320 31220
rect 36544 31272 36596 31278
rect 36544 31214 36596 31220
rect 36556 30734 36584 31214
rect 36648 30734 36676 31758
rect 36544 30728 36596 30734
rect 36544 30670 36596 30676
rect 36636 30728 36688 30734
rect 36636 30670 36688 30676
rect 36556 30258 36584 30670
rect 36648 30598 36676 30670
rect 36912 30660 36964 30666
rect 36912 30602 36964 30608
rect 36636 30592 36688 30598
rect 36636 30534 36688 30540
rect 36924 30394 36952 30602
rect 36912 30388 36964 30394
rect 36912 30330 36964 30336
rect 36544 30252 36596 30258
rect 36544 30194 36596 30200
rect 36636 28484 36688 28490
rect 36636 28426 36688 28432
rect 36648 28218 36676 28426
rect 36636 28212 36688 28218
rect 36636 28154 36688 28160
rect 37096 27464 37148 27470
rect 37016 27412 37096 27418
rect 37016 27406 37148 27412
rect 37016 27390 37136 27406
rect 37016 27130 37044 27390
rect 37004 27124 37056 27130
rect 37004 27066 37056 27072
rect 36820 27056 36872 27062
rect 36740 27004 36820 27010
rect 36740 26998 36872 27004
rect 36268 26988 36320 26994
rect 36740 26982 36860 26998
rect 36740 26976 36768 26982
rect 36320 26948 36768 26976
rect 36268 26930 36320 26936
rect 36820 26920 36872 26926
rect 37004 26920 37056 26926
rect 36820 26862 36872 26868
rect 37002 26888 37004 26897
rect 37056 26888 37058 26897
rect 36452 26784 36504 26790
rect 36452 26726 36504 26732
rect 36464 26382 36492 26726
rect 36268 26376 36320 26382
rect 36268 26318 36320 26324
rect 36452 26376 36504 26382
rect 36452 26318 36504 26324
rect 36280 25294 36308 26318
rect 36636 25968 36688 25974
rect 36636 25910 36688 25916
rect 36544 25900 36596 25906
rect 36544 25842 36596 25848
rect 36360 25696 36412 25702
rect 36360 25638 36412 25644
rect 36372 25294 36400 25638
rect 36556 25537 36584 25842
rect 36648 25838 36676 25910
rect 36832 25906 36860 26862
rect 37002 26823 37058 26832
rect 37096 26580 37148 26586
rect 37096 26522 37148 26528
rect 37004 26376 37056 26382
rect 37002 26344 37004 26353
rect 37056 26344 37058 26353
rect 37002 26279 37058 26288
rect 36820 25900 36872 25906
rect 36820 25842 36872 25848
rect 37004 25900 37056 25906
rect 37004 25842 37056 25848
rect 36636 25832 36688 25838
rect 36636 25774 36688 25780
rect 36912 25832 36964 25838
rect 37016 25809 37044 25842
rect 36912 25774 36964 25780
rect 37002 25800 37058 25809
rect 36542 25528 36598 25537
rect 36542 25463 36598 25472
rect 36268 25288 36320 25294
rect 36268 25230 36320 25236
rect 36360 25288 36412 25294
rect 36360 25230 36412 25236
rect 36280 24750 36308 25230
rect 36924 24886 36952 25774
rect 37002 25735 37058 25744
rect 36912 24880 36964 24886
rect 36912 24822 36964 24828
rect 36268 24744 36320 24750
rect 36268 24686 36320 24692
rect 36636 24404 36688 24410
rect 35912 24126 36216 24154
rect 36464 24364 36636 24392
rect 35808 23860 35860 23866
rect 35808 23802 35860 23808
rect 35716 23792 35768 23798
rect 35716 23734 35768 23740
rect 35728 22982 35756 23734
rect 35808 23112 35860 23118
rect 35808 23054 35860 23060
rect 35716 22976 35768 22982
rect 35716 22918 35768 22924
rect 35820 22642 35848 23054
rect 35808 22636 35860 22642
rect 35808 22578 35860 22584
rect 35624 20596 35676 20602
rect 35624 20538 35676 20544
rect 35636 19718 35664 20538
rect 35624 19712 35676 19718
rect 35624 19654 35676 19660
rect 35912 19446 35940 24126
rect 36084 24064 36136 24070
rect 36084 24006 36136 24012
rect 36096 23798 36124 24006
rect 36084 23792 36136 23798
rect 36084 23734 36136 23740
rect 35992 23724 36044 23730
rect 35992 23666 36044 23672
rect 36004 23610 36032 23666
rect 36004 23582 36124 23610
rect 35992 23316 36044 23322
rect 35992 23258 36044 23264
rect 36004 22642 36032 23258
rect 36096 23202 36124 23582
rect 36464 23526 36492 24364
rect 36636 24346 36688 24352
rect 36544 23656 36596 23662
rect 36544 23598 36596 23604
rect 36452 23520 36504 23526
rect 36452 23462 36504 23468
rect 36176 23248 36228 23254
rect 36096 23196 36176 23202
rect 36096 23190 36228 23196
rect 36096 23174 36216 23190
rect 36464 23186 36492 23462
rect 36556 23322 36584 23598
rect 36544 23316 36596 23322
rect 36544 23258 36596 23264
rect 36452 23180 36504 23186
rect 35992 22636 36044 22642
rect 35992 22578 36044 22584
rect 36096 22506 36124 23174
rect 36452 23122 36504 23128
rect 36268 23112 36320 23118
rect 36268 23054 36320 23060
rect 36176 22976 36228 22982
rect 36176 22918 36228 22924
rect 36188 22642 36216 22918
rect 36176 22636 36228 22642
rect 36176 22578 36228 22584
rect 36084 22500 36136 22506
rect 36084 22442 36136 22448
rect 36176 22432 36228 22438
rect 36176 22374 36228 22380
rect 36188 22030 36216 22374
rect 36280 22030 36308 23054
rect 36820 22636 36872 22642
rect 36820 22578 36872 22584
rect 36832 22098 36860 22578
rect 37108 22574 37136 26522
rect 37096 22568 37148 22574
rect 37096 22510 37148 22516
rect 36820 22092 36872 22098
rect 36820 22034 36872 22040
rect 36176 22024 36228 22030
rect 36176 21966 36228 21972
rect 36268 22024 36320 22030
rect 36268 21966 36320 21972
rect 36176 21684 36228 21690
rect 36176 21626 36228 21632
rect 36188 21078 36216 21626
rect 36176 21072 36228 21078
rect 36176 21014 36228 21020
rect 36188 20398 36216 21014
rect 36280 21010 36308 21966
rect 36360 21888 36412 21894
rect 36360 21830 36412 21836
rect 36372 21690 36400 21830
rect 36360 21684 36412 21690
rect 36360 21626 36412 21632
rect 36268 21004 36320 21010
rect 36268 20946 36320 20952
rect 36544 20460 36596 20466
rect 36544 20402 36596 20408
rect 36176 20392 36228 20398
rect 36176 20334 36228 20340
rect 36188 19854 36216 20334
rect 36556 20330 36584 20402
rect 36544 20324 36596 20330
rect 36544 20266 36596 20272
rect 36176 19848 36228 19854
rect 36176 19790 36228 19796
rect 35900 19440 35952 19446
rect 35900 19382 35952 19388
rect 35912 18970 35940 19382
rect 35900 18964 35952 18970
rect 35900 18906 35952 18912
rect 35992 18760 36044 18766
rect 35992 18702 36044 18708
rect 36004 17338 36032 18702
rect 36556 18290 36584 20266
rect 37108 20262 37136 22510
rect 37200 22098 37228 31758
rect 37372 31748 37424 31754
rect 37372 31690 37424 31696
rect 37384 31482 37412 31690
rect 37372 31476 37424 31482
rect 37372 31418 37424 31424
rect 38108 31272 38160 31278
rect 38108 31214 38160 31220
rect 38016 31204 38068 31210
rect 38016 31146 38068 31152
rect 37464 30048 37516 30054
rect 37464 29990 37516 29996
rect 37280 29572 37332 29578
rect 37280 29514 37332 29520
rect 37292 29170 37320 29514
rect 37280 29164 37332 29170
rect 37280 29106 37332 29112
rect 37476 29102 37504 29990
rect 37556 29572 37608 29578
rect 37556 29514 37608 29520
rect 37464 29096 37516 29102
rect 37464 29038 37516 29044
rect 37464 28688 37516 28694
rect 37464 28630 37516 28636
rect 37372 28416 37424 28422
rect 37372 28358 37424 28364
rect 37384 27962 37412 28358
rect 37476 28082 37504 28630
rect 37568 28218 37596 29514
rect 37556 28212 37608 28218
rect 37556 28154 37608 28160
rect 37464 28076 37516 28082
rect 37464 28018 37516 28024
rect 37384 27934 37596 27962
rect 37280 27396 37332 27402
rect 37280 27338 37332 27344
rect 37292 27130 37320 27338
rect 37464 27328 37516 27334
rect 37464 27270 37516 27276
rect 37476 27130 37504 27270
rect 37280 27124 37332 27130
rect 37280 27066 37332 27072
rect 37464 27124 37516 27130
rect 37464 27066 37516 27072
rect 37464 26920 37516 26926
rect 37464 26862 37516 26868
rect 37476 26382 37504 26862
rect 37464 26376 37516 26382
rect 37464 26318 37516 26324
rect 37280 25152 37332 25158
rect 37280 25094 37332 25100
rect 37292 24070 37320 25094
rect 37372 24200 37424 24206
rect 37372 24142 37424 24148
rect 37280 24064 37332 24070
rect 37280 24006 37332 24012
rect 37280 23792 37332 23798
rect 37280 23734 37332 23740
rect 37292 22778 37320 23734
rect 37280 22772 37332 22778
rect 37280 22714 37332 22720
rect 37384 22438 37412 24142
rect 37464 23520 37516 23526
rect 37464 23462 37516 23468
rect 37476 22506 37504 23462
rect 37568 23118 37596 27934
rect 37738 27024 37794 27033
rect 37738 26959 37794 26968
rect 37924 26988 37976 26994
rect 37752 26858 37780 26959
rect 37924 26930 37976 26936
rect 37936 26897 37964 26930
rect 37922 26888 37978 26897
rect 37740 26852 37792 26858
rect 37922 26823 37978 26832
rect 37740 26794 37792 26800
rect 37648 25152 37700 25158
rect 37648 25094 37700 25100
rect 37660 24206 37688 25094
rect 37648 24200 37700 24206
rect 37648 24142 37700 24148
rect 37924 24064 37976 24070
rect 37924 24006 37976 24012
rect 37648 23520 37700 23526
rect 37648 23462 37700 23468
rect 37660 23186 37688 23462
rect 37648 23180 37700 23186
rect 37648 23122 37700 23128
rect 37556 23112 37608 23118
rect 37556 23054 37608 23060
rect 37556 22976 37608 22982
rect 37556 22918 37608 22924
rect 37464 22500 37516 22506
rect 37464 22442 37516 22448
rect 37372 22432 37424 22438
rect 37372 22374 37424 22380
rect 37188 22092 37240 22098
rect 37188 22034 37240 22040
rect 37280 21344 37332 21350
rect 37280 21286 37332 21292
rect 37292 20398 37320 21286
rect 37568 21146 37596 22918
rect 37648 22432 37700 22438
rect 37648 22374 37700 22380
rect 37556 21140 37608 21146
rect 37556 21082 37608 21088
rect 37372 20800 37424 20806
rect 37372 20742 37424 20748
rect 37280 20392 37332 20398
rect 37280 20334 37332 20340
rect 37096 20256 37148 20262
rect 37096 20198 37148 20204
rect 37292 19922 37320 20334
rect 37280 19916 37332 19922
rect 37280 19858 37332 19864
rect 37004 19848 37056 19854
rect 37004 19790 37056 19796
rect 37016 19378 37044 19790
rect 37004 19372 37056 19378
rect 37004 19314 37056 19320
rect 37292 19242 37320 19858
rect 37280 19236 37332 19242
rect 37280 19178 37332 19184
rect 37384 18970 37412 20742
rect 37464 20256 37516 20262
rect 37464 20198 37516 20204
rect 37476 19310 37504 20198
rect 37660 20058 37688 22374
rect 37832 22024 37884 22030
rect 37832 21966 37884 21972
rect 37844 21554 37872 21966
rect 37832 21548 37884 21554
rect 37832 21490 37884 21496
rect 37740 21412 37792 21418
rect 37740 21354 37792 21360
rect 37752 21146 37780 21354
rect 37844 21350 37872 21490
rect 37832 21344 37884 21350
rect 37832 21286 37884 21292
rect 37740 21140 37792 21146
rect 37740 21082 37792 21088
rect 37936 21078 37964 24006
rect 38028 21486 38056 31146
rect 38120 30938 38148 31214
rect 38108 30932 38160 30938
rect 38108 30874 38160 30880
rect 38106 27160 38162 27169
rect 38106 27095 38162 27104
rect 38120 26926 38148 27095
rect 38108 26920 38160 26926
rect 38108 26862 38160 26868
rect 38106 25392 38162 25401
rect 38106 25327 38162 25336
rect 38120 24206 38148 25327
rect 38304 24682 38332 49030
rect 38568 48544 38620 48550
rect 38568 48486 38620 48492
rect 38476 46504 38528 46510
rect 38476 46446 38528 46452
rect 38488 46170 38516 46446
rect 38476 46164 38528 46170
rect 38476 46106 38528 46112
rect 38580 31890 38608 48486
rect 38660 46708 38712 46714
rect 38660 46650 38712 46656
rect 38672 46510 38700 46650
rect 38660 46504 38712 46510
rect 38660 46446 38712 46452
rect 38660 46368 38712 46374
rect 38660 46310 38712 46316
rect 38568 31884 38620 31890
rect 38568 31826 38620 31832
rect 38672 29850 38700 46310
rect 39132 32502 39160 51326
rect 39302 51200 39358 52000
rect 39946 51200 40002 52000
rect 40590 51354 40646 52000
rect 40590 51326 40816 51354
rect 40590 51200 40646 51326
rect 39316 45554 39344 51200
rect 39488 48680 39540 48686
rect 39960 48668 39988 51200
rect 40788 49230 40816 51326
rect 41234 51200 41290 52000
rect 41878 51354 41934 52000
rect 41616 51326 41934 51354
rect 40776 49224 40828 49230
rect 40776 49166 40828 49172
rect 40868 49088 40920 49094
rect 40868 49030 40920 49036
rect 40040 48680 40092 48686
rect 39960 48640 40040 48668
rect 39488 48622 39540 48628
rect 40040 48622 40092 48628
rect 39500 48346 39528 48622
rect 39488 48340 39540 48346
rect 39488 48282 39540 48288
rect 39316 45526 39804 45554
rect 39120 32496 39172 32502
rect 39120 32438 39172 32444
rect 39776 31414 39804 45526
rect 40880 38010 40908 49030
rect 41248 48278 41276 51200
rect 41616 49230 41644 51326
rect 41878 51200 41934 51326
rect 42522 51200 42578 52000
rect 43166 51200 43222 52000
rect 43810 51354 43866 52000
rect 43810 51326 44128 51354
rect 43810 51200 43866 51326
rect 41604 49224 41656 49230
rect 41604 49166 41656 49172
rect 42432 49224 42484 49230
rect 42432 49166 42484 49172
rect 41420 49156 41472 49162
rect 41420 49098 41472 49104
rect 41236 48272 41288 48278
rect 41236 48214 41288 48220
rect 41432 48210 41460 49098
rect 41604 49088 41656 49094
rect 41604 49030 41656 49036
rect 41420 48204 41472 48210
rect 41420 48146 41472 48152
rect 40868 38004 40920 38010
rect 40868 37946 40920 37952
rect 40776 32768 40828 32774
rect 40776 32710 40828 32716
rect 39764 31408 39816 31414
rect 39764 31350 39816 31356
rect 38660 29844 38712 29850
rect 38660 29786 38712 29792
rect 38476 29096 38528 29102
rect 38476 29038 38528 29044
rect 38488 28082 38516 29038
rect 38672 28558 38700 29786
rect 39580 29096 39632 29102
rect 39580 29038 39632 29044
rect 39304 28620 39356 28626
rect 39304 28562 39356 28568
rect 38660 28552 38712 28558
rect 38660 28494 38712 28500
rect 39028 28552 39080 28558
rect 39028 28494 39080 28500
rect 38476 28076 38528 28082
rect 38476 28018 38528 28024
rect 38488 27470 38516 28018
rect 39040 27878 39068 28494
rect 39028 27872 39080 27878
rect 39028 27814 39080 27820
rect 38476 27464 38528 27470
rect 38476 27406 38528 27412
rect 38488 26994 38516 27406
rect 38476 26988 38528 26994
rect 38476 26930 38528 26936
rect 38488 26382 38516 26930
rect 38476 26376 38528 26382
rect 38476 26318 38528 26324
rect 38292 24676 38344 24682
rect 38292 24618 38344 24624
rect 38752 24404 38804 24410
rect 38752 24346 38804 24352
rect 38108 24200 38160 24206
rect 38108 24142 38160 24148
rect 38120 23254 38148 24142
rect 38566 24032 38622 24041
rect 38566 23967 38622 23976
rect 38384 23792 38436 23798
rect 38384 23734 38436 23740
rect 38108 23248 38160 23254
rect 38108 23190 38160 23196
rect 38108 23044 38160 23050
rect 38108 22986 38160 22992
rect 38120 22506 38148 22986
rect 38396 22642 38424 23734
rect 38580 23730 38608 23967
rect 38568 23724 38620 23730
rect 38568 23666 38620 23672
rect 38764 23526 38792 24346
rect 39040 24290 39068 27814
rect 38948 24262 39068 24290
rect 38844 24064 38896 24070
rect 38844 24006 38896 24012
rect 38856 23866 38884 24006
rect 38844 23860 38896 23866
rect 38844 23802 38896 23808
rect 38476 23520 38528 23526
rect 38476 23462 38528 23468
rect 38752 23520 38804 23526
rect 38752 23462 38804 23468
rect 38488 23322 38516 23462
rect 38476 23316 38528 23322
rect 38476 23258 38528 23264
rect 38476 23180 38528 23186
rect 38476 23122 38528 23128
rect 38384 22636 38436 22642
rect 38384 22578 38436 22584
rect 38488 22574 38516 23122
rect 38476 22568 38528 22574
rect 38476 22510 38528 22516
rect 38108 22500 38160 22506
rect 38108 22442 38160 22448
rect 38474 21992 38530 22001
rect 38474 21927 38530 21936
rect 38292 21616 38344 21622
rect 38292 21558 38344 21564
rect 38016 21480 38068 21486
rect 38016 21422 38068 21428
rect 38016 21344 38068 21350
rect 38016 21286 38068 21292
rect 37924 21072 37976 21078
rect 37924 21014 37976 21020
rect 38028 21010 38056 21286
rect 38304 21146 38332 21558
rect 38292 21140 38344 21146
rect 38292 21082 38344 21088
rect 38016 21004 38068 21010
rect 38016 20946 38068 20952
rect 38108 20936 38160 20942
rect 38108 20878 38160 20884
rect 38016 20800 38068 20806
rect 38016 20742 38068 20748
rect 38028 20602 38056 20742
rect 38016 20596 38068 20602
rect 38016 20538 38068 20544
rect 38120 20398 38148 20878
rect 38108 20392 38160 20398
rect 38108 20334 38160 20340
rect 38384 20256 38436 20262
rect 38384 20198 38436 20204
rect 37648 20052 37700 20058
rect 37648 19994 37700 20000
rect 37464 19304 37516 19310
rect 37464 19246 37516 19252
rect 37372 18964 37424 18970
rect 37372 18906 37424 18912
rect 36544 18284 36596 18290
rect 36544 18226 36596 18232
rect 37660 18222 37688 19994
rect 38014 19816 38070 19825
rect 38200 19780 38252 19786
rect 38014 19751 38016 19760
rect 38068 19751 38070 19760
rect 38016 19722 38068 19728
rect 38120 19740 38200 19768
rect 38120 19446 38148 19740
rect 38200 19722 38252 19728
rect 38200 19508 38252 19514
rect 38200 19450 38252 19456
rect 38108 19440 38160 19446
rect 38108 19382 38160 19388
rect 38212 19378 38240 19450
rect 38396 19378 38424 20198
rect 38488 19854 38516 21927
rect 38948 21350 38976 24262
rect 39028 23656 39080 23662
rect 39028 23598 39080 23604
rect 39040 23254 39068 23598
rect 39028 23248 39080 23254
rect 39028 23190 39080 23196
rect 38936 21344 38988 21350
rect 38936 21286 38988 21292
rect 38752 19916 38804 19922
rect 38752 19858 38804 19864
rect 38476 19848 38528 19854
rect 38476 19790 38528 19796
rect 38566 19816 38622 19825
rect 38566 19751 38568 19760
rect 38620 19751 38622 19760
rect 38660 19780 38712 19786
rect 38568 19722 38620 19728
rect 38660 19722 38712 19728
rect 38476 19712 38528 19718
rect 38476 19654 38528 19660
rect 38200 19372 38252 19378
rect 38200 19314 38252 19320
rect 38384 19372 38436 19378
rect 38384 19314 38436 19320
rect 38488 19174 38516 19654
rect 38672 19310 38700 19722
rect 38660 19304 38712 19310
rect 38660 19246 38712 19252
rect 38476 19168 38528 19174
rect 38476 19110 38528 19116
rect 38660 19168 38712 19174
rect 38660 19110 38712 19116
rect 38672 18766 38700 19110
rect 38764 18834 38792 19858
rect 38752 18828 38804 18834
rect 38752 18770 38804 18776
rect 37924 18760 37976 18766
rect 37924 18702 37976 18708
rect 38016 18760 38068 18766
rect 38016 18702 38068 18708
rect 38660 18760 38712 18766
rect 38660 18702 38712 18708
rect 37936 18426 37964 18702
rect 37924 18420 37976 18426
rect 37924 18362 37976 18368
rect 37924 18284 37976 18290
rect 37924 18226 37976 18232
rect 37648 18216 37700 18222
rect 37648 18158 37700 18164
rect 37936 17678 37964 18226
rect 38028 17882 38056 18702
rect 38292 18216 38344 18222
rect 38292 18158 38344 18164
rect 38016 17876 38068 17882
rect 38016 17818 38068 17824
rect 38304 17746 38332 18158
rect 38292 17740 38344 17746
rect 38292 17682 38344 17688
rect 37924 17672 37976 17678
rect 37924 17614 37976 17620
rect 37648 17536 37700 17542
rect 37648 17478 37700 17484
rect 35992 17332 36044 17338
rect 35992 17274 36044 17280
rect 35532 17264 35584 17270
rect 35532 17206 35584 17212
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 35544 16250 35572 17206
rect 36004 16658 36032 17274
rect 36176 17196 36228 17202
rect 36176 17138 36228 17144
rect 35992 16652 36044 16658
rect 35992 16594 36044 16600
rect 35532 16244 35584 16250
rect 35532 16186 35584 16192
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34704 15428 34756 15434
rect 34704 15370 34756 15376
rect 35716 15428 35768 15434
rect 35716 15370 35768 15376
rect 34612 15020 34664 15026
rect 34612 14962 34664 14968
rect 34624 14618 34652 14962
rect 34612 14612 34664 14618
rect 34612 14554 34664 14560
rect 34428 14476 34480 14482
rect 34532 14470 34652 14498
rect 34428 14418 34480 14424
rect 34440 13870 34468 14418
rect 34518 14240 34574 14249
rect 34518 14175 34574 14184
rect 34532 13938 34560 14175
rect 34520 13932 34572 13938
rect 34520 13874 34572 13880
rect 34428 13864 34480 13870
rect 34428 13806 34480 13812
rect 34440 12306 34468 13806
rect 34520 13728 34572 13734
rect 34520 13670 34572 13676
rect 34532 12918 34560 13670
rect 34520 12912 34572 12918
rect 34520 12854 34572 12860
rect 34428 12300 34480 12306
rect 34428 12242 34480 12248
rect 34336 11688 34388 11694
rect 34336 11630 34388 11636
rect 34624 10606 34652 14470
rect 34716 14278 34744 15370
rect 35348 15360 35400 15366
rect 35348 15302 35400 15308
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 35360 14600 35388 15302
rect 35440 15088 35492 15094
rect 35440 15030 35492 15036
rect 35176 14572 35388 14600
rect 34886 14512 34942 14521
rect 34886 14447 34942 14456
rect 34900 14414 34928 14447
rect 35176 14414 35204 14572
rect 35452 14414 35480 15030
rect 35728 14890 35756 15370
rect 35716 14884 35768 14890
rect 35716 14826 35768 14832
rect 34888 14408 34940 14414
rect 34888 14350 34940 14356
rect 35164 14408 35216 14414
rect 35440 14408 35492 14414
rect 35164 14350 35216 14356
rect 35360 14368 35440 14396
rect 34704 14272 34756 14278
rect 34704 14214 34756 14220
rect 35360 14090 35388 14368
rect 35492 14368 35572 14396
rect 35440 14350 35492 14356
rect 35440 14272 35492 14278
rect 35440 14214 35492 14220
rect 35268 14062 35388 14090
rect 35268 13938 35296 14062
rect 35348 14000 35400 14006
rect 35348 13942 35400 13948
rect 35256 13932 35308 13938
rect 35256 13874 35308 13880
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34704 13252 34756 13258
rect 34704 13194 34756 13200
rect 34716 12442 34744 13194
rect 35360 13190 35388 13942
rect 35452 13938 35480 14214
rect 35440 13932 35492 13938
rect 35440 13874 35492 13880
rect 35348 13184 35400 13190
rect 35348 13126 35400 13132
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 34704 12436 34756 12442
rect 34704 12378 34756 12384
rect 35544 12238 35572 14368
rect 35808 13864 35860 13870
rect 35808 13806 35860 13812
rect 35624 13796 35676 13802
rect 35624 13738 35676 13744
rect 35636 12646 35664 13738
rect 35624 12640 35676 12646
rect 35624 12582 35676 12588
rect 35820 12306 35848 13806
rect 35808 12300 35860 12306
rect 35808 12242 35860 12248
rect 36188 12238 36216 17138
rect 37660 17134 37688 17478
rect 37648 17128 37700 17134
rect 37648 17070 37700 17076
rect 37660 16726 37688 17070
rect 37648 16720 37700 16726
rect 37648 16662 37700 16668
rect 37464 16516 37516 16522
rect 37464 16458 37516 16464
rect 37476 16114 37504 16458
rect 37464 16108 37516 16114
rect 37464 16050 37516 16056
rect 38948 16046 38976 21286
rect 39120 19712 39172 19718
rect 39120 19654 39172 19660
rect 39132 19378 39160 19654
rect 39028 19372 39080 19378
rect 39028 19314 39080 19320
rect 39120 19372 39172 19378
rect 39120 19314 39172 19320
rect 39040 18970 39068 19314
rect 39028 18964 39080 18970
rect 39028 18906 39080 18912
rect 39212 16108 39264 16114
rect 39212 16050 39264 16056
rect 38936 16040 38988 16046
rect 38936 15982 38988 15988
rect 38384 15972 38436 15978
rect 38384 15914 38436 15920
rect 37188 15496 37240 15502
rect 37188 15438 37240 15444
rect 36728 15360 36780 15366
rect 36728 15302 36780 15308
rect 36740 14414 36768 15302
rect 36728 14408 36780 14414
rect 36728 14350 36780 14356
rect 35532 12232 35584 12238
rect 35532 12174 35584 12180
rect 35900 12232 35952 12238
rect 35900 12174 35952 12180
rect 36176 12232 36228 12238
rect 36176 12174 36228 12180
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 35912 11082 35940 12174
rect 37200 12102 37228 15438
rect 37924 15428 37976 15434
rect 37924 15370 37976 15376
rect 37936 14958 37964 15370
rect 37924 14952 37976 14958
rect 37924 14894 37976 14900
rect 37936 14618 37964 14894
rect 38396 14890 38424 15914
rect 38948 15638 38976 15982
rect 39224 15706 39252 16050
rect 39212 15700 39264 15706
rect 39212 15642 39264 15648
rect 38936 15632 38988 15638
rect 38936 15574 38988 15580
rect 38844 15428 38896 15434
rect 38844 15370 38896 15376
rect 38384 14884 38436 14890
rect 38384 14826 38436 14832
rect 37924 14612 37976 14618
rect 37924 14554 37976 14560
rect 37462 14512 37518 14521
rect 37462 14447 37464 14456
rect 37516 14447 37518 14456
rect 37464 14418 37516 14424
rect 38396 14414 38424 14826
rect 38856 14822 38884 15370
rect 39028 14952 39080 14958
rect 39028 14894 39080 14900
rect 38844 14816 38896 14822
rect 38844 14758 38896 14764
rect 38384 14408 38436 14414
rect 38384 14350 38436 14356
rect 38292 14340 38344 14346
rect 38292 14282 38344 14288
rect 38304 14249 38332 14282
rect 38476 14272 38528 14278
rect 38290 14240 38346 14249
rect 38476 14214 38528 14220
rect 38290 14175 38346 14184
rect 38488 14006 38516 14214
rect 38476 14000 38528 14006
rect 38476 13942 38528 13948
rect 38856 13870 38884 14758
rect 38844 13864 38896 13870
rect 38844 13806 38896 13812
rect 36084 12096 36136 12102
rect 36084 12038 36136 12044
rect 37188 12096 37240 12102
rect 37188 12038 37240 12044
rect 36096 11898 36124 12038
rect 36084 11892 36136 11898
rect 36084 11834 36136 11840
rect 35900 11076 35952 11082
rect 35900 11018 35952 11024
rect 34612 10600 34664 10606
rect 34612 10542 34664 10548
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 38016 8288 38068 8294
rect 38016 8230 38068 8236
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 35624 6316 35676 6322
rect 35624 6258 35676 6264
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 33968 3732 34020 3738
rect 33968 3674 34020 3680
rect 32956 3392 33008 3398
rect 32956 3334 33008 3340
rect 32968 3126 32996 3334
rect 34992 3194 35388 3210
rect 34980 3188 35388 3194
rect 35032 3182 35388 3188
rect 34980 3130 35032 3136
rect 35360 3126 35388 3182
rect 32956 3120 33008 3126
rect 32956 3062 33008 3068
rect 35348 3120 35400 3126
rect 35348 3062 35400 3068
rect 32772 3052 32824 3058
rect 32772 2994 32824 3000
rect 33508 2984 33560 2990
rect 35440 2984 35492 2990
rect 33508 2926 33560 2932
rect 32864 2440 32916 2446
rect 32864 2382 32916 2388
rect 32876 800 32904 2382
rect 33520 800 33548 2926
rect 34072 2922 34284 2938
rect 35440 2926 35492 2932
rect 34060 2916 34296 2922
rect 34112 2910 34244 2916
rect 34060 2858 34112 2864
rect 34244 2858 34296 2864
rect 34520 2848 34572 2854
rect 34520 2790 34572 2796
rect 35348 2848 35400 2854
rect 35348 2790 35400 2796
rect 34532 2582 34560 2790
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 34520 2576 34572 2582
rect 34520 2518 34572 2524
rect 34152 2440 34204 2446
rect 34152 2382 34204 2388
rect 34796 2440 34848 2446
rect 34796 2382 34848 2388
rect 34164 800 34192 2382
rect 34808 800 34836 2382
rect 35360 1834 35388 2790
rect 35452 2582 35480 2926
rect 35636 2922 35664 6258
rect 36452 4140 36504 4146
rect 36452 4082 36504 4088
rect 36464 4049 36492 4082
rect 36450 4040 36506 4049
rect 36450 3975 36506 3984
rect 36176 3936 36228 3942
rect 36176 3878 36228 3884
rect 37924 3936 37976 3942
rect 37924 3878 37976 3884
rect 36188 3602 36216 3878
rect 37372 3732 37424 3738
rect 37372 3674 37424 3680
rect 36176 3596 36228 3602
rect 36176 3538 36228 3544
rect 36728 3596 36780 3602
rect 36728 3538 36780 3544
rect 35992 3528 36044 3534
rect 35992 3470 36044 3476
rect 36004 3058 36032 3470
rect 35992 3052 36044 3058
rect 35992 2994 36044 3000
rect 35624 2916 35676 2922
rect 35624 2858 35676 2864
rect 35440 2576 35492 2582
rect 35440 2518 35492 2524
rect 36084 2372 36136 2378
rect 36084 2314 36136 2320
rect 35348 1828 35400 1834
rect 35348 1770 35400 1776
rect 36096 800 36124 2314
rect 36740 800 36768 3538
rect 37384 800 37412 3674
rect 37740 3528 37792 3534
rect 37740 3470 37792 3476
rect 37752 3058 37780 3470
rect 37936 3126 37964 3878
rect 37924 3120 37976 3126
rect 37924 3062 37976 3068
rect 37740 3052 37792 3058
rect 37740 2994 37792 3000
rect 38028 800 38056 8230
rect 38752 5160 38804 5166
rect 38752 5102 38804 5108
rect 38764 2582 38792 5102
rect 38752 2576 38804 2582
rect 38752 2518 38804 2524
rect 38660 2440 38712 2446
rect 38660 2382 38712 2388
rect 38672 800 38700 2382
rect 39040 2038 39068 14894
rect 39316 5370 39344 28562
rect 39396 26920 39448 26926
rect 39396 26862 39448 26868
rect 39408 26586 39436 26862
rect 39396 26580 39448 26586
rect 39396 26522 39448 26528
rect 39396 24608 39448 24614
rect 39394 24576 39396 24585
rect 39448 24576 39450 24585
rect 39394 24511 39450 24520
rect 39396 20052 39448 20058
rect 39396 19994 39448 20000
rect 39408 19514 39436 19994
rect 39396 19508 39448 19514
rect 39396 19450 39448 19456
rect 39396 17808 39448 17814
rect 39396 17750 39448 17756
rect 39408 17066 39436 17750
rect 39396 17060 39448 17066
rect 39396 17002 39448 17008
rect 39408 16114 39436 17002
rect 39396 16108 39448 16114
rect 39396 16050 39448 16056
rect 39488 6180 39540 6186
rect 39488 6122 39540 6128
rect 39304 5364 39356 5370
rect 39304 5306 39356 5312
rect 39500 4146 39528 6122
rect 39488 4140 39540 4146
rect 39488 4082 39540 4088
rect 39592 3738 39620 29038
rect 39856 28484 39908 28490
rect 39856 28426 39908 28432
rect 39672 27532 39724 27538
rect 39672 27474 39724 27480
rect 39684 26450 39712 27474
rect 39672 26444 39724 26450
rect 39672 26386 39724 26392
rect 39868 24206 39896 28426
rect 40040 26784 40092 26790
rect 40040 26726 40092 26732
rect 40052 26450 40080 26726
rect 40040 26444 40092 26450
rect 40040 26386 40092 26392
rect 40684 25424 40736 25430
rect 40684 25366 40736 25372
rect 40500 25288 40552 25294
rect 40500 25230 40552 25236
rect 40132 25152 40184 25158
rect 40132 25094 40184 25100
rect 40144 24818 40172 25094
rect 40132 24812 40184 24818
rect 40132 24754 40184 24760
rect 40224 24812 40276 24818
rect 40224 24754 40276 24760
rect 40236 24342 40264 24754
rect 40512 24342 40540 25230
rect 40696 24954 40724 25366
rect 40684 24948 40736 24954
rect 40684 24890 40736 24896
rect 40224 24336 40276 24342
rect 40224 24278 40276 24284
rect 40500 24336 40552 24342
rect 40500 24278 40552 24284
rect 39764 24200 39816 24206
rect 39856 24200 39908 24206
rect 39764 24142 39816 24148
rect 39854 24168 39856 24177
rect 39908 24168 39910 24177
rect 39672 24064 39724 24070
rect 39672 24006 39724 24012
rect 39684 23905 39712 24006
rect 39670 23896 39726 23905
rect 39670 23831 39726 23840
rect 39672 23724 39724 23730
rect 39672 23666 39724 23672
rect 39684 23526 39712 23666
rect 39776 23610 39804 24142
rect 39854 24103 39910 24112
rect 40592 24132 40644 24138
rect 40592 24074 40644 24080
rect 40604 23730 40632 24074
rect 40408 23724 40460 23730
rect 40408 23666 40460 23672
rect 40592 23724 40644 23730
rect 40592 23666 40644 23672
rect 39856 23656 39908 23662
rect 39776 23604 39856 23610
rect 40420 23633 40448 23666
rect 39776 23598 39908 23604
rect 40406 23624 40462 23633
rect 39776 23582 39896 23598
rect 39672 23520 39724 23526
rect 39672 23462 39724 23468
rect 39776 23118 39804 23582
rect 40406 23559 40462 23568
rect 40500 23316 40552 23322
rect 40500 23258 40552 23264
rect 39764 23112 39816 23118
rect 39764 23054 39816 23060
rect 40314 22808 40370 22817
rect 40512 22778 40540 23258
rect 40604 23186 40632 23666
rect 40592 23180 40644 23186
rect 40592 23122 40644 23128
rect 40314 22743 40316 22752
rect 40368 22743 40370 22752
rect 40500 22772 40552 22778
rect 40316 22714 40368 22720
rect 40500 22714 40552 22720
rect 40512 22030 40540 22714
rect 40684 22432 40736 22438
rect 40684 22374 40736 22380
rect 40500 22024 40552 22030
rect 40500 21966 40552 21972
rect 40224 21480 40276 21486
rect 40224 21422 40276 21428
rect 40132 21140 40184 21146
rect 40132 21082 40184 21088
rect 40144 20534 40172 21082
rect 40236 20874 40264 21422
rect 40696 21418 40724 22374
rect 40788 21690 40816 32710
rect 41510 26480 41566 26489
rect 41510 26415 41566 26424
rect 41524 26382 41552 26415
rect 41512 26376 41564 26382
rect 41512 26318 41564 26324
rect 41616 25294 41644 49030
rect 42340 48748 42392 48754
rect 42340 48690 42392 48696
rect 41788 48544 41840 48550
rect 41788 48486 41840 48492
rect 41800 48210 41828 48486
rect 41788 48204 41840 48210
rect 41788 48146 41840 48152
rect 41788 48068 41840 48074
rect 41788 48010 41840 48016
rect 41800 47802 41828 48010
rect 41788 47796 41840 47802
rect 41788 47738 41840 47744
rect 41696 47660 41748 47666
rect 41696 47602 41748 47608
rect 41708 45966 41736 47602
rect 41696 45960 41748 45966
rect 41696 45902 41748 45908
rect 41708 41138 41736 45902
rect 41696 41132 41748 41138
rect 41696 41074 41748 41080
rect 41696 27396 41748 27402
rect 41696 27338 41748 27344
rect 41708 26489 41736 27338
rect 41694 26480 41750 26489
rect 41694 26415 41750 26424
rect 41696 26308 41748 26314
rect 41696 26250 41748 26256
rect 41604 25288 41656 25294
rect 41604 25230 41656 25236
rect 41052 24880 41104 24886
rect 41052 24822 41104 24828
rect 40866 24440 40922 24449
rect 40866 24375 40922 24384
rect 40880 24274 40908 24375
rect 40960 24336 41012 24342
rect 40960 24278 41012 24284
rect 40868 24268 40920 24274
rect 40868 24210 40920 24216
rect 40866 23896 40922 23905
rect 40866 23831 40868 23840
rect 40920 23831 40922 23840
rect 40868 23802 40920 23808
rect 40868 23724 40920 23730
rect 40868 23666 40920 23672
rect 40880 23322 40908 23666
rect 40972 23662 41000 24278
rect 41064 24274 41092 24822
rect 41144 24608 41196 24614
rect 41144 24550 41196 24556
rect 41052 24268 41104 24274
rect 41052 24210 41104 24216
rect 41156 24206 41184 24550
rect 41420 24404 41472 24410
rect 41420 24346 41472 24352
rect 41144 24200 41196 24206
rect 41144 24142 41196 24148
rect 41326 24168 41382 24177
rect 40960 23656 41012 23662
rect 40960 23598 41012 23604
rect 41156 23526 41184 24142
rect 41432 24138 41460 24346
rect 41326 24103 41382 24112
rect 41420 24132 41472 24138
rect 41144 23520 41196 23526
rect 41144 23462 41196 23468
rect 40868 23316 40920 23322
rect 40868 23258 40920 23264
rect 40868 22704 40920 22710
rect 40868 22646 40920 22652
rect 40880 22506 40908 22646
rect 41340 22574 41368 24103
rect 41420 24074 41472 24080
rect 41328 22568 41380 22574
rect 41328 22510 41380 22516
rect 40868 22500 40920 22506
rect 40868 22442 40920 22448
rect 40776 21684 40828 21690
rect 40776 21626 40828 21632
rect 40880 21554 40908 22442
rect 40960 22432 41012 22438
rect 40960 22374 41012 22380
rect 40868 21548 40920 21554
rect 40868 21490 40920 21496
rect 40684 21412 40736 21418
rect 40684 21354 40736 21360
rect 40408 21344 40460 21350
rect 40408 21286 40460 21292
rect 40420 20942 40448 21286
rect 40408 20936 40460 20942
rect 40408 20878 40460 20884
rect 40224 20868 40276 20874
rect 40224 20810 40276 20816
rect 40132 20528 40184 20534
rect 40132 20470 40184 20476
rect 40236 19258 40264 20810
rect 40500 20324 40552 20330
rect 40500 20266 40552 20272
rect 40408 20052 40460 20058
rect 40408 19994 40460 20000
rect 40144 19230 40264 19258
rect 40144 18222 40172 19230
rect 40224 18692 40276 18698
rect 40224 18634 40276 18640
rect 40236 18290 40264 18634
rect 40224 18284 40276 18290
rect 40224 18226 40276 18232
rect 40132 18216 40184 18222
rect 40132 18158 40184 18164
rect 40040 17672 40092 17678
rect 40040 17614 40092 17620
rect 40052 17202 40080 17614
rect 40040 17196 40092 17202
rect 40040 17138 40092 17144
rect 40052 16250 40080 17138
rect 40144 16658 40172 18158
rect 40420 17678 40448 19994
rect 40408 17672 40460 17678
rect 40408 17614 40460 17620
rect 40512 17202 40540 20266
rect 40696 19378 40724 21354
rect 40880 20534 40908 21490
rect 40972 21350 41000 22374
rect 41340 22234 41368 22510
rect 41328 22228 41380 22234
rect 41328 22170 41380 22176
rect 41144 22024 41196 22030
rect 41144 21966 41196 21972
rect 40960 21344 41012 21350
rect 40960 21286 41012 21292
rect 40868 20528 40920 20534
rect 40868 20470 40920 20476
rect 40960 20324 41012 20330
rect 41012 20284 41092 20312
rect 40960 20266 41012 20272
rect 40868 20256 40920 20262
rect 40868 20198 40920 20204
rect 40880 19922 40908 20198
rect 40868 19916 40920 19922
rect 40868 19858 40920 19864
rect 40776 19780 40828 19786
rect 40776 19722 40828 19728
rect 40788 19514 40816 19722
rect 40880 19718 40908 19858
rect 41064 19854 41092 20284
rect 41156 20058 41184 21966
rect 41432 21962 41460 24074
rect 41512 23656 41564 23662
rect 41510 23624 41512 23633
rect 41564 23624 41566 23633
rect 41510 23559 41566 23568
rect 41604 23112 41656 23118
rect 41604 23054 41656 23060
rect 41616 22710 41644 23054
rect 41604 22704 41656 22710
rect 41604 22646 41656 22652
rect 41420 21956 41472 21962
rect 41420 21898 41472 21904
rect 41328 21616 41380 21622
rect 41328 21558 41380 21564
rect 41340 20466 41368 21558
rect 41328 20460 41380 20466
rect 41328 20402 41380 20408
rect 41144 20052 41196 20058
rect 41144 19994 41196 20000
rect 41052 19848 41104 19854
rect 41052 19790 41104 19796
rect 40960 19780 41012 19786
rect 40960 19722 41012 19728
rect 40868 19712 40920 19718
rect 40868 19654 40920 19660
rect 40776 19508 40828 19514
rect 40776 19450 40828 19456
rect 40684 19372 40736 19378
rect 40684 19314 40736 19320
rect 40696 18630 40724 19314
rect 40788 18970 40816 19450
rect 40776 18964 40828 18970
rect 40776 18906 40828 18912
rect 40776 18828 40828 18834
rect 40776 18770 40828 18776
rect 40788 18630 40816 18770
rect 40684 18624 40736 18630
rect 40684 18566 40736 18572
rect 40776 18624 40828 18630
rect 40776 18566 40828 18572
rect 40880 18290 40908 19654
rect 40972 19378 41000 19722
rect 41340 19446 41368 20402
rect 41420 19712 41472 19718
rect 41420 19654 41472 19660
rect 41328 19440 41380 19446
rect 41328 19382 41380 19388
rect 40960 19372 41012 19378
rect 40960 19314 41012 19320
rect 41144 19236 41196 19242
rect 41144 19178 41196 19184
rect 41052 18896 41104 18902
rect 41052 18838 41104 18844
rect 40868 18284 40920 18290
rect 40868 18226 40920 18232
rect 40776 17740 40828 17746
rect 40776 17682 40828 17688
rect 40788 17202 40816 17682
rect 41064 17678 41092 18838
rect 41156 18358 41184 19178
rect 41236 18828 41288 18834
rect 41236 18770 41288 18776
rect 41144 18352 41196 18358
rect 41144 18294 41196 18300
rect 41248 18222 41276 18770
rect 41340 18630 41368 19382
rect 41432 19174 41460 19654
rect 41604 19372 41656 19378
rect 41604 19314 41656 19320
rect 41616 19242 41644 19314
rect 41604 19236 41656 19242
rect 41604 19178 41656 19184
rect 41420 19168 41472 19174
rect 41420 19110 41472 19116
rect 41512 18964 41564 18970
rect 41512 18906 41564 18912
rect 41328 18624 41380 18630
rect 41328 18566 41380 18572
rect 41524 18426 41552 18906
rect 41512 18420 41564 18426
rect 41512 18362 41564 18368
rect 41236 18216 41288 18222
rect 41236 18158 41288 18164
rect 41052 17672 41104 17678
rect 41052 17614 41104 17620
rect 41064 17270 41092 17614
rect 41604 17536 41656 17542
rect 41604 17478 41656 17484
rect 41052 17264 41104 17270
rect 41052 17206 41104 17212
rect 40500 17196 40552 17202
rect 40500 17138 40552 17144
rect 40776 17196 40828 17202
rect 40776 17138 40828 17144
rect 40132 16652 40184 16658
rect 40132 16594 40184 16600
rect 40040 16244 40092 16250
rect 40040 16186 40092 16192
rect 39672 15904 39724 15910
rect 39672 15846 39724 15852
rect 39684 15026 39712 15846
rect 40144 15570 40172 16594
rect 40512 16114 40540 17138
rect 40788 16454 40816 17138
rect 40776 16448 40828 16454
rect 40776 16390 40828 16396
rect 41064 16114 41092 17206
rect 41616 16998 41644 17478
rect 41420 16992 41472 16998
rect 41420 16934 41472 16940
rect 41604 16992 41656 16998
rect 41604 16934 41656 16940
rect 41432 16522 41460 16934
rect 41236 16516 41288 16522
rect 41236 16458 41288 16464
rect 41420 16516 41472 16522
rect 41420 16458 41472 16464
rect 41248 16250 41276 16458
rect 41236 16244 41288 16250
rect 41236 16186 41288 16192
rect 40500 16108 40552 16114
rect 40500 16050 40552 16056
rect 41052 16108 41104 16114
rect 41052 16050 41104 16056
rect 40132 15564 40184 15570
rect 40132 15506 40184 15512
rect 40144 15094 40172 15506
rect 40512 15366 40540 16050
rect 40500 15360 40552 15366
rect 40500 15302 40552 15308
rect 40132 15088 40184 15094
rect 40132 15030 40184 15036
rect 39672 15020 39724 15026
rect 39672 14962 39724 14968
rect 39948 13864 40000 13870
rect 39948 13806 40000 13812
rect 39580 3732 39632 3738
rect 39580 3674 39632 3680
rect 39960 3466 39988 13806
rect 41708 9110 41736 26250
rect 42352 25906 42380 48690
rect 42444 48278 42472 49166
rect 42432 48272 42484 48278
rect 42432 48214 42484 48220
rect 42536 48210 42564 51200
rect 43180 49298 43208 51200
rect 43996 49768 44048 49774
rect 43996 49710 44048 49716
rect 43168 49292 43220 49298
rect 43168 49234 43220 49240
rect 42800 48544 42852 48550
rect 42800 48486 42852 48492
rect 43904 48544 43956 48550
rect 43904 48486 43956 48492
rect 42524 48204 42576 48210
rect 42524 48146 42576 48152
rect 42812 46986 42840 48486
rect 43168 47116 43220 47122
rect 43168 47058 43220 47064
rect 42800 46980 42852 46986
rect 42800 46922 42852 46928
rect 43180 46578 43208 47058
rect 43168 46572 43220 46578
rect 43168 46514 43220 46520
rect 43916 31346 43944 48486
rect 44008 47598 44036 49710
rect 44100 48142 44128 51326
rect 44454 51200 44510 52000
rect 45098 51354 45154 52000
rect 45742 51354 45798 52000
rect 45098 51326 45232 51354
rect 45098 51200 45154 51326
rect 44468 48822 44496 51200
rect 44456 48816 44508 48822
rect 44456 48758 44508 48764
rect 44456 48680 44508 48686
rect 44456 48622 44508 48628
rect 44640 48680 44692 48686
rect 44640 48622 44692 48628
rect 44088 48136 44140 48142
rect 44088 48078 44140 48084
rect 44180 48000 44232 48006
rect 44180 47942 44232 47948
rect 44364 48000 44416 48006
rect 44364 47942 44416 47948
rect 43996 47592 44048 47598
rect 43996 47534 44048 47540
rect 44192 35894 44220 47942
rect 44376 47734 44404 47942
rect 44364 47728 44416 47734
rect 44364 47670 44416 47676
rect 44272 46980 44324 46986
rect 44272 46922 44324 46928
rect 44284 46578 44312 46922
rect 44468 46578 44496 48622
rect 44652 48346 44680 48622
rect 44640 48340 44692 48346
rect 44640 48282 44692 48288
rect 45204 47598 45232 51326
rect 45742 51326 45876 51354
rect 45742 51200 45798 51326
rect 45744 49156 45796 49162
rect 45744 49098 45796 49104
rect 45284 49088 45336 49094
rect 45284 49030 45336 49036
rect 44732 47592 44784 47598
rect 44732 47534 44784 47540
rect 45100 47592 45152 47598
rect 45100 47534 45152 47540
rect 45192 47592 45244 47598
rect 45192 47534 45244 47540
rect 44272 46572 44324 46578
rect 44272 46514 44324 46520
rect 44456 46572 44508 46578
rect 44456 46514 44508 46520
rect 44744 46170 44772 47534
rect 45112 47258 45140 47534
rect 45100 47252 45152 47258
rect 45100 47194 45152 47200
rect 45192 47048 45244 47054
rect 45192 46990 45244 46996
rect 45100 46504 45152 46510
rect 45100 46446 45152 46452
rect 44732 46164 44784 46170
rect 44732 46106 44784 46112
rect 45112 45422 45140 46446
rect 45204 45966 45232 46990
rect 45192 45960 45244 45966
rect 45192 45902 45244 45908
rect 45100 45416 45152 45422
rect 45100 45358 45152 45364
rect 44192 35866 44312 35894
rect 43904 31340 43956 31346
rect 43904 31282 43956 31288
rect 42340 25900 42392 25906
rect 42340 25842 42392 25848
rect 41972 24812 42024 24818
rect 41972 24754 42024 24760
rect 42432 24812 42484 24818
rect 42432 24754 42484 24760
rect 41984 24410 42012 24754
rect 42340 24608 42392 24614
rect 42340 24550 42392 24556
rect 41972 24404 42024 24410
rect 41972 24346 42024 24352
rect 42064 24404 42116 24410
rect 42064 24346 42116 24352
rect 41788 24064 41840 24070
rect 41788 24006 41840 24012
rect 41800 23662 41828 24006
rect 41788 23656 41840 23662
rect 41788 23598 41840 23604
rect 41972 22976 42024 22982
rect 41972 22918 42024 22924
rect 41984 21962 42012 22918
rect 42076 22234 42104 24346
rect 42154 24304 42210 24313
rect 42154 24239 42156 24248
rect 42208 24239 42210 24248
rect 42156 24210 42208 24216
rect 42246 24168 42302 24177
rect 42246 24103 42248 24112
rect 42300 24103 42302 24112
rect 42248 24074 42300 24080
rect 42352 23798 42380 24550
rect 42340 23792 42392 23798
rect 42340 23734 42392 23740
rect 42156 23316 42208 23322
rect 42156 23258 42208 23264
rect 42064 22228 42116 22234
rect 42064 22170 42116 22176
rect 41788 21956 41840 21962
rect 41788 21898 41840 21904
rect 41972 21956 42024 21962
rect 41972 21898 42024 21904
rect 41800 20398 41828 21898
rect 41880 21344 41932 21350
rect 41880 21286 41932 21292
rect 41892 20942 41920 21286
rect 41880 20936 41932 20942
rect 41880 20878 41932 20884
rect 42168 20466 42196 23258
rect 42352 23186 42380 23734
rect 42444 23662 42472 24754
rect 43444 24676 43496 24682
rect 43444 24618 43496 24624
rect 42522 24576 42578 24585
rect 42522 24511 42578 24520
rect 42536 23866 42564 24511
rect 43456 24449 43484 24618
rect 43442 24440 43498 24449
rect 43442 24375 43498 24384
rect 43352 24336 43404 24342
rect 43350 24304 43352 24313
rect 43404 24304 43406 24313
rect 43350 24239 43406 24248
rect 42892 24200 42944 24206
rect 43168 24200 43220 24206
rect 42892 24142 42944 24148
rect 43166 24168 43168 24177
rect 43352 24200 43404 24206
rect 43220 24168 43222 24177
rect 42524 23860 42576 23866
rect 42524 23802 42576 23808
rect 42432 23656 42484 23662
rect 42432 23598 42484 23604
rect 42798 23624 42854 23633
rect 42798 23559 42800 23568
rect 42852 23559 42854 23568
rect 42800 23530 42852 23536
rect 42340 23180 42392 23186
rect 42340 23122 42392 23128
rect 42352 22506 42380 23122
rect 42616 23112 42668 23118
rect 42616 23054 42668 23060
rect 42432 23044 42484 23050
rect 42432 22986 42484 22992
rect 42444 22574 42472 22986
rect 42628 22574 42656 23054
rect 42904 23050 42932 24142
rect 43352 24142 43404 24148
rect 43444 24200 43496 24206
rect 43444 24142 43496 24148
rect 43166 24103 43222 24112
rect 43260 24064 43312 24070
rect 42996 24012 43260 24018
rect 42996 24006 43312 24012
rect 42996 23990 43300 24006
rect 42996 23798 43024 23990
rect 42984 23792 43036 23798
rect 42984 23734 43036 23740
rect 43364 23118 43392 24142
rect 43352 23112 43404 23118
rect 43352 23054 43404 23060
rect 42892 23044 42944 23050
rect 42892 22986 42944 22992
rect 43076 22636 43128 22642
rect 43076 22578 43128 22584
rect 42432 22568 42484 22574
rect 42432 22510 42484 22516
rect 42616 22568 42668 22574
rect 42616 22510 42668 22516
rect 42340 22500 42392 22506
rect 42340 22442 42392 22448
rect 42444 22438 42472 22510
rect 42432 22432 42484 22438
rect 42432 22374 42484 22380
rect 42524 22432 42576 22438
rect 42524 22374 42576 22380
rect 42536 22030 42564 22374
rect 42628 22030 42656 22510
rect 42524 22024 42576 22030
rect 42524 21966 42576 21972
rect 42616 22024 42668 22030
rect 42616 21966 42668 21972
rect 42432 21956 42484 21962
rect 42432 21898 42484 21904
rect 42444 21690 42472 21898
rect 42432 21684 42484 21690
rect 42432 21626 42484 21632
rect 42156 20460 42208 20466
rect 42156 20402 42208 20408
rect 42708 20460 42760 20466
rect 42708 20402 42760 20408
rect 41788 20392 41840 20398
rect 41788 20334 41840 20340
rect 41800 17270 41828 20334
rect 41880 19780 41932 19786
rect 41880 19722 41932 19728
rect 41892 19514 41920 19722
rect 41880 19508 41932 19514
rect 41880 19450 41932 19456
rect 41892 17542 41920 19450
rect 42432 19168 42484 19174
rect 42432 19110 42484 19116
rect 42444 18698 42472 19110
rect 42432 18692 42484 18698
rect 42432 18634 42484 18640
rect 42156 18624 42208 18630
rect 42156 18566 42208 18572
rect 41972 18284 42024 18290
rect 41972 18226 42024 18232
rect 41984 17882 42012 18226
rect 41972 17876 42024 17882
rect 41972 17818 42024 17824
rect 42168 17678 42196 18566
rect 42156 17672 42208 17678
rect 42156 17614 42208 17620
rect 41880 17536 41932 17542
rect 41880 17478 41932 17484
rect 41788 17264 41840 17270
rect 41788 17206 41840 17212
rect 41972 17264 42024 17270
rect 41972 17206 42024 17212
rect 41788 16992 41840 16998
rect 41788 16934 41840 16940
rect 41800 16114 41828 16934
rect 41984 16522 42012 17206
rect 42156 16788 42208 16794
rect 42156 16730 42208 16736
rect 41972 16516 42024 16522
rect 41972 16458 42024 16464
rect 41788 16108 41840 16114
rect 41788 16050 41840 16056
rect 42168 16046 42196 16730
rect 42616 16448 42668 16454
rect 42616 16390 42668 16396
rect 42628 16114 42656 16390
rect 42616 16108 42668 16114
rect 42616 16050 42668 16056
rect 42156 16040 42208 16046
rect 42156 15982 42208 15988
rect 42432 15904 42484 15910
rect 42432 15846 42484 15852
rect 42444 15502 42472 15846
rect 42432 15496 42484 15502
rect 42432 15438 42484 15444
rect 42720 15434 42748 20402
rect 43088 18834 43116 22578
rect 43456 22166 43484 24142
rect 43812 24064 43864 24070
rect 43812 24006 43864 24012
rect 43824 23798 43852 24006
rect 43812 23792 43864 23798
rect 43812 23734 43864 23740
rect 43904 23656 43956 23662
rect 43902 23624 43904 23633
rect 43956 23624 43958 23633
rect 43902 23559 43958 23568
rect 43996 23588 44048 23594
rect 43996 23530 44048 23536
rect 44008 23186 44036 23530
rect 44180 23520 44232 23526
rect 44180 23462 44232 23468
rect 43996 23180 44048 23186
rect 43996 23122 44048 23128
rect 44008 22817 44036 23122
rect 43994 22808 44050 22817
rect 43994 22743 44050 22752
rect 44088 22636 44140 22642
rect 44088 22578 44140 22584
rect 43444 22160 43496 22166
rect 43444 22102 43496 22108
rect 43352 22024 43404 22030
rect 43352 21966 43404 21972
rect 43444 22024 43496 22030
rect 43444 21966 43496 21972
rect 43364 21078 43392 21966
rect 43456 21146 43484 21966
rect 43628 21888 43680 21894
rect 43628 21830 43680 21836
rect 43640 21554 43668 21830
rect 43628 21548 43680 21554
rect 43628 21490 43680 21496
rect 43444 21140 43496 21146
rect 43444 21082 43496 21088
rect 43352 21072 43404 21078
rect 43352 21014 43404 21020
rect 44100 20942 44128 22578
rect 44192 22098 44220 23462
rect 44180 22092 44232 22098
rect 44180 22034 44232 22040
rect 44088 20936 44140 20942
rect 44088 20878 44140 20884
rect 44100 20602 44128 20878
rect 44088 20596 44140 20602
rect 44088 20538 44140 20544
rect 43168 20256 43220 20262
rect 43168 20198 43220 20204
rect 43180 19378 43208 20198
rect 44100 19786 44128 20538
rect 44088 19780 44140 19786
rect 44088 19722 44140 19728
rect 43168 19372 43220 19378
rect 43168 19314 43220 19320
rect 43812 19304 43864 19310
rect 43812 19246 43864 19252
rect 43076 18828 43128 18834
rect 43076 18770 43128 18776
rect 43260 18624 43312 18630
rect 43260 18566 43312 18572
rect 43272 17678 43300 18566
rect 43824 18426 43852 19246
rect 44100 18698 44128 19722
rect 44088 18692 44140 18698
rect 44088 18634 44140 18640
rect 43812 18420 43864 18426
rect 43812 18362 43864 18368
rect 43260 17672 43312 17678
rect 43260 17614 43312 17620
rect 42708 15428 42760 15434
rect 42708 15370 42760 15376
rect 44284 14482 44312 35866
rect 44732 28008 44784 28014
rect 44732 27950 44784 27956
rect 44456 23724 44508 23730
rect 44456 23666 44508 23672
rect 44468 22778 44496 23666
rect 44456 22772 44508 22778
rect 44456 22714 44508 22720
rect 44456 21956 44508 21962
rect 44456 21898 44508 21904
rect 44468 20602 44496 21898
rect 44456 20596 44508 20602
rect 44456 20538 44508 20544
rect 44548 19304 44600 19310
rect 44548 19246 44600 19252
rect 44560 18766 44588 19246
rect 44548 18760 44600 18766
rect 44548 18702 44600 18708
rect 44456 18624 44508 18630
rect 44456 18566 44508 18572
rect 44468 17746 44496 18566
rect 44560 18290 44588 18702
rect 44548 18284 44600 18290
rect 44548 18226 44600 18232
rect 44456 17740 44508 17746
rect 44456 17682 44508 17688
rect 44272 14476 44324 14482
rect 44272 14418 44324 14424
rect 44744 12442 44772 27950
rect 45204 24818 45232 45902
rect 45296 45422 45324 49030
rect 45652 48136 45704 48142
rect 45652 48078 45704 48084
rect 45468 47796 45520 47802
rect 45468 47738 45520 47744
rect 45376 46504 45428 46510
rect 45376 46446 45428 46452
rect 45388 46170 45416 46446
rect 45376 46164 45428 46170
rect 45376 46106 45428 46112
rect 45284 45416 45336 45422
rect 45284 45358 45336 45364
rect 45480 45082 45508 47738
rect 45664 47734 45692 48078
rect 45652 47728 45704 47734
rect 45652 47670 45704 47676
rect 45756 47258 45784 49098
rect 45848 48686 45876 51326
rect 46386 51200 46442 52000
rect 46754 51776 46810 51785
rect 46754 51711 46810 51720
rect 45926 51096 45982 51105
rect 45926 51031 45982 51040
rect 45836 48680 45888 48686
rect 45836 48622 45888 48628
rect 45744 47252 45796 47258
rect 45744 47194 45796 47200
rect 45652 47184 45704 47190
rect 45652 47126 45704 47132
rect 45664 47054 45692 47126
rect 45652 47048 45704 47054
rect 45652 46990 45704 46996
rect 45468 45076 45520 45082
rect 45468 45018 45520 45024
rect 45664 39982 45692 46990
rect 45652 39976 45704 39982
rect 45652 39918 45704 39924
rect 45652 35692 45704 35698
rect 45652 35634 45704 35640
rect 45468 31816 45520 31822
rect 45468 31758 45520 31764
rect 45480 30734 45508 31758
rect 45468 30728 45520 30734
rect 45468 30670 45520 30676
rect 45480 27470 45508 30670
rect 45560 28008 45612 28014
rect 45560 27950 45612 27956
rect 45572 27606 45600 27950
rect 45560 27600 45612 27606
rect 45560 27542 45612 27548
rect 45468 27464 45520 27470
rect 45468 27406 45520 27412
rect 45560 26512 45612 26518
rect 45560 26454 45612 26460
rect 45572 25974 45600 26454
rect 45560 25968 45612 25974
rect 45560 25910 45612 25916
rect 45192 24812 45244 24818
rect 45192 24754 45244 24760
rect 45008 23112 45060 23118
rect 45008 23054 45060 23060
rect 44916 21344 44968 21350
rect 44916 21286 44968 21292
rect 44928 20874 44956 21286
rect 45020 21010 45048 23054
rect 45468 22432 45520 22438
rect 45468 22374 45520 22380
rect 45480 21078 45508 22374
rect 45664 22094 45692 35634
rect 45836 35556 45888 35562
rect 45836 35498 45888 35504
rect 45848 27130 45876 35498
rect 45836 27124 45888 27130
rect 45836 27066 45888 27072
rect 45744 25832 45796 25838
rect 45744 25774 45796 25780
rect 45756 25498 45784 25774
rect 45744 25492 45796 25498
rect 45744 25434 45796 25440
rect 45940 23322 45968 51031
rect 46768 49774 46796 51711
rect 47030 51200 47086 52000
rect 47674 51354 47730 52000
rect 47674 51326 47808 51354
rect 47674 51200 47730 51326
rect 46846 50416 46902 50425
rect 46846 50351 46902 50360
rect 46756 49768 46808 49774
rect 46662 49736 46718 49745
rect 46756 49710 46808 49716
rect 46662 49671 46718 49680
rect 46296 48884 46348 48890
rect 46296 48826 46348 48832
rect 46308 48210 46336 48826
rect 46296 48204 46348 48210
rect 46296 48146 46348 48152
rect 46676 47122 46704 49671
rect 46754 49056 46810 49065
rect 46754 48991 46810 49000
rect 46768 48754 46796 48991
rect 46756 48748 46808 48754
rect 46756 48690 46808 48696
rect 46860 48210 46888 50351
rect 47780 49230 47808 51326
rect 48318 51200 48374 52000
rect 48962 51200 49018 52000
rect 49606 51200 49662 52000
rect 48332 49298 48360 51200
rect 48320 49292 48372 49298
rect 48320 49234 48372 49240
rect 47768 49224 47820 49230
rect 47768 49166 47820 49172
rect 47124 49088 47176 49094
rect 47124 49030 47176 49036
rect 46940 48544 46992 48550
rect 46940 48486 46992 48492
rect 46848 48204 46900 48210
rect 46848 48146 46900 48152
rect 46664 47116 46716 47122
rect 46664 47058 46716 47064
rect 46846 47016 46902 47025
rect 46480 46980 46532 46986
rect 46846 46951 46902 46960
rect 46480 46922 46532 46928
rect 46296 45960 46348 45966
rect 46296 45902 46348 45908
rect 46308 45422 46336 45902
rect 46492 45422 46520 46922
rect 46860 46510 46888 46951
rect 46848 46504 46900 46510
rect 46848 46446 46900 46452
rect 46296 45416 46348 45422
rect 46296 45358 46348 45364
rect 46480 45416 46532 45422
rect 46480 45358 46532 45364
rect 46846 44976 46902 44985
rect 46846 44911 46902 44920
rect 46296 44872 46348 44878
rect 46296 44814 46348 44820
rect 46308 44402 46336 44814
rect 46296 44396 46348 44402
rect 46296 44338 46348 44344
rect 46018 44296 46074 44305
rect 46018 44231 46074 44240
rect 46032 35894 46060 44231
rect 46860 43722 46888 44911
rect 46848 43716 46900 43722
rect 46848 43658 46900 43664
rect 46296 42016 46348 42022
rect 46296 41958 46348 41964
rect 46308 41682 46336 41958
rect 46296 41676 46348 41682
rect 46296 41618 46348 41624
rect 46480 41540 46532 41546
rect 46480 41482 46532 41488
rect 46492 41274 46520 41482
rect 46480 41268 46532 41274
rect 46480 41210 46532 41216
rect 46664 41132 46716 41138
rect 46664 41074 46716 41080
rect 46572 37868 46624 37874
rect 46572 37810 46624 37816
rect 46480 36576 46532 36582
rect 46480 36518 46532 36524
rect 46492 36242 46520 36518
rect 46480 36236 46532 36242
rect 46480 36178 46532 36184
rect 46584 35894 46612 37810
rect 46032 35866 46152 35894
rect 46020 34672 46072 34678
rect 46020 34614 46072 34620
rect 46032 33522 46060 34614
rect 46020 33516 46072 33522
rect 46020 33458 46072 33464
rect 46124 33402 46152 35866
rect 46400 35866 46612 35894
rect 46296 35488 46348 35494
rect 46296 35430 46348 35436
rect 46308 35154 46336 35430
rect 46296 35148 46348 35154
rect 46296 35090 46348 35096
rect 46204 33448 46256 33454
rect 46032 33374 46152 33402
rect 46202 33416 46204 33425
rect 46256 33416 46258 33425
rect 46032 28014 46060 33374
rect 46202 33351 46258 33360
rect 46400 32586 46428 35866
rect 46480 35488 46532 35494
rect 46480 35430 46532 35436
rect 46492 35154 46520 35430
rect 46480 35148 46532 35154
rect 46480 35090 46532 35096
rect 46480 34400 46532 34406
rect 46480 34342 46532 34348
rect 46492 34066 46520 34342
rect 46480 34060 46532 34066
rect 46480 34002 46532 34008
rect 46480 32836 46532 32842
rect 46480 32778 46532 32784
rect 46308 32558 46428 32586
rect 46204 32360 46256 32366
rect 46204 32302 46256 32308
rect 46216 31686 46244 32302
rect 46308 31754 46336 32558
rect 46388 32428 46440 32434
rect 46388 32370 46440 32376
rect 46400 32065 46428 32370
rect 46386 32056 46442 32065
rect 46492 32026 46520 32778
rect 46386 31991 46442 32000
rect 46480 32020 46532 32026
rect 46480 31962 46532 31968
rect 46572 31884 46624 31890
rect 46572 31826 46624 31832
rect 46308 31726 46428 31754
rect 46204 31680 46256 31686
rect 46204 31622 46256 31628
rect 46400 30666 46428 31726
rect 46584 31142 46612 31826
rect 46572 31136 46624 31142
rect 46572 31078 46624 31084
rect 46388 30660 46440 30666
rect 46388 30602 46440 30608
rect 46296 29640 46348 29646
rect 46296 29582 46348 29588
rect 46112 28552 46164 28558
rect 46112 28494 46164 28500
rect 46020 28008 46072 28014
rect 46020 27950 46072 27956
rect 45928 23316 45980 23322
rect 45928 23258 45980 23264
rect 45664 22066 45876 22094
rect 45744 21548 45796 21554
rect 45744 21490 45796 21496
rect 45756 21146 45784 21490
rect 45744 21140 45796 21146
rect 45744 21082 45796 21088
rect 45376 21072 45428 21078
rect 45376 21014 45428 21020
rect 45468 21072 45520 21078
rect 45468 21014 45520 21020
rect 45008 21004 45060 21010
rect 45008 20946 45060 20952
rect 45388 20939 45416 21014
rect 45373 20933 45425 20939
rect 45373 20875 45425 20881
rect 45652 20936 45704 20942
rect 45652 20878 45704 20884
rect 44916 20868 44968 20874
rect 44916 20810 44968 20816
rect 44824 19372 44876 19378
rect 44824 19314 44876 19320
rect 44836 17882 44864 19314
rect 44824 17876 44876 17882
rect 44824 17818 44876 17824
rect 44732 12436 44784 12442
rect 44732 12378 44784 12384
rect 44824 12164 44876 12170
rect 44824 12106 44876 12112
rect 41696 9104 41748 9110
rect 41696 9046 41748 9052
rect 41972 4616 42024 4622
rect 41972 4558 42024 4564
rect 40776 4004 40828 4010
rect 40776 3946 40828 3952
rect 40224 3936 40276 3942
rect 40224 3878 40276 3884
rect 39948 3460 40000 3466
rect 39948 3402 40000 3408
rect 40040 3392 40092 3398
rect 40040 3334 40092 3340
rect 40052 3058 40080 3334
rect 40236 3126 40264 3878
rect 40788 3534 40816 3946
rect 41420 3936 41472 3942
rect 41420 3878 41472 3884
rect 41432 3602 41460 3878
rect 41420 3596 41472 3602
rect 41420 3538 41472 3544
rect 41880 3596 41932 3602
rect 41880 3538 41932 3544
rect 40776 3528 40828 3534
rect 40776 3470 40828 3476
rect 40224 3120 40276 3126
rect 40224 3062 40276 3068
rect 40040 3052 40092 3058
rect 40040 2994 40092 3000
rect 39948 2984 40000 2990
rect 39948 2926 40000 2932
rect 41236 2984 41288 2990
rect 41236 2926 41288 2932
rect 39028 2032 39080 2038
rect 39028 1974 39080 1980
rect 39960 800 39988 2926
rect 41248 800 41276 2926
rect 41892 800 41920 3538
rect 41984 2514 42012 4558
rect 42432 4140 42484 4146
rect 42432 4082 42484 4088
rect 42444 3670 42472 4082
rect 44836 4078 44864 12106
rect 44928 6866 44956 20810
rect 45192 20460 45244 20466
rect 45192 20402 45244 20408
rect 45100 19916 45152 19922
rect 45100 19858 45152 19864
rect 45112 19378 45140 19858
rect 45204 19786 45232 20402
rect 45388 20330 45416 20875
rect 45664 20398 45692 20878
rect 45652 20392 45704 20398
rect 45652 20334 45704 20340
rect 45376 20324 45428 20330
rect 45376 20266 45428 20272
rect 45192 19780 45244 19786
rect 45192 19722 45244 19728
rect 45100 19372 45152 19378
rect 45100 19314 45152 19320
rect 45388 18902 45416 20266
rect 45468 19712 45520 19718
rect 45468 19654 45520 19660
rect 45480 18902 45508 19654
rect 45376 18896 45428 18902
rect 45376 18838 45428 18844
rect 45468 18896 45520 18902
rect 45468 18838 45520 18844
rect 45008 18624 45060 18630
rect 45008 18566 45060 18572
rect 45020 18358 45048 18566
rect 45008 18352 45060 18358
rect 45008 18294 45060 18300
rect 45388 17542 45416 18838
rect 45664 18766 45692 20334
rect 45652 18760 45704 18766
rect 45652 18702 45704 18708
rect 45744 18760 45796 18766
rect 45744 18702 45796 18708
rect 45664 17814 45692 18702
rect 45756 18086 45784 18702
rect 45744 18080 45796 18086
rect 45744 18022 45796 18028
rect 45652 17808 45704 17814
rect 45652 17750 45704 17756
rect 45376 17536 45428 17542
rect 45376 17478 45428 17484
rect 45848 17338 45876 22066
rect 46124 21894 46152 28494
rect 46308 27538 46336 29582
rect 46296 27532 46348 27538
rect 46296 27474 46348 27480
rect 46400 26994 46428 30602
rect 46572 29028 46624 29034
rect 46572 28970 46624 28976
rect 46480 28484 46532 28490
rect 46480 28426 46532 28432
rect 46492 27130 46520 28426
rect 46584 27538 46612 28970
rect 46572 27532 46624 27538
rect 46572 27474 46624 27480
rect 46480 27124 46532 27130
rect 46480 27066 46532 27072
rect 46388 26988 46440 26994
rect 46388 26930 46440 26936
rect 46204 25288 46256 25294
rect 46204 25230 46256 25236
rect 46388 25288 46440 25294
rect 46388 25230 46440 25236
rect 46112 21888 46164 21894
rect 46112 21830 46164 21836
rect 45928 19168 45980 19174
rect 45928 19110 45980 19116
rect 45940 18698 45968 19110
rect 46112 18896 46164 18902
rect 46112 18838 46164 18844
rect 45928 18692 45980 18698
rect 45928 18634 45980 18640
rect 45836 17332 45888 17338
rect 45836 17274 45888 17280
rect 45836 17128 45888 17134
rect 45836 17070 45888 17076
rect 45848 16794 45876 17070
rect 45836 16788 45888 16794
rect 45836 16730 45888 16736
rect 45940 16658 45968 18634
rect 45928 16652 45980 16658
rect 45928 16594 45980 16600
rect 45836 16584 45888 16590
rect 45836 16526 45888 16532
rect 45848 16182 45876 16526
rect 46020 16448 46072 16454
rect 46020 16390 46072 16396
rect 45836 16176 45888 16182
rect 45836 16118 45888 16124
rect 45652 8084 45704 8090
rect 45652 8026 45704 8032
rect 45560 7404 45612 7410
rect 45560 7346 45612 7352
rect 44916 6860 44968 6866
rect 44916 6802 44968 6808
rect 45572 5930 45600 7346
rect 45480 5914 45600 5930
rect 45468 5908 45600 5914
rect 45520 5902 45600 5908
rect 45468 5850 45520 5856
rect 45572 4146 45600 5902
rect 45560 4140 45612 4146
rect 45560 4082 45612 4088
rect 44824 4072 44876 4078
rect 44824 4014 44876 4020
rect 44640 4004 44692 4010
rect 44640 3946 44692 3952
rect 42616 3936 42668 3942
rect 42616 3878 42668 3884
rect 43996 3936 44048 3942
rect 43996 3878 44048 3884
rect 42432 3664 42484 3670
rect 42432 3606 42484 3612
rect 42628 2514 42656 3878
rect 43812 3528 43864 3534
rect 43812 3470 43864 3476
rect 43824 3058 43852 3470
rect 44008 3126 44036 3878
rect 43996 3120 44048 3126
rect 43996 3062 44048 3068
rect 43168 3052 43220 3058
rect 43168 2994 43220 3000
rect 43812 3052 43864 3058
rect 43812 2994 43864 3000
rect 41972 2508 42024 2514
rect 41972 2450 42024 2456
rect 42616 2508 42668 2514
rect 42616 2450 42668 2456
rect 42708 2508 42760 2514
rect 42708 2450 42760 2456
rect 42720 1170 42748 2450
rect 42536 1142 42748 1170
rect 42536 800 42564 1142
rect 43180 800 43208 2994
rect 44456 2984 44508 2990
rect 44456 2926 44508 2932
rect 44468 800 44496 2926
rect 44652 2514 44680 3946
rect 45376 3936 45428 3942
rect 45376 3878 45428 3884
rect 45388 3602 45416 3878
rect 45376 3596 45428 3602
rect 45376 3538 45428 3544
rect 45192 3392 45244 3398
rect 45192 3334 45244 3340
rect 45204 2514 45232 3334
rect 45664 3194 45692 8026
rect 45848 6322 45876 16118
rect 46032 6905 46060 16390
rect 46018 6896 46074 6905
rect 46018 6831 46074 6840
rect 45928 6724 45980 6730
rect 45928 6666 45980 6672
rect 45940 6458 45968 6666
rect 45928 6452 45980 6458
rect 45928 6394 45980 6400
rect 45836 6316 45888 6322
rect 45836 6258 45888 6264
rect 45848 4146 45876 6258
rect 46124 4185 46152 18838
rect 46216 15162 46244 25230
rect 46296 19780 46348 19786
rect 46296 19722 46348 19728
rect 46308 18426 46336 19722
rect 46296 18420 46348 18426
rect 46296 18362 46348 18368
rect 46308 17746 46336 18362
rect 46296 17740 46348 17746
rect 46296 17682 46348 17688
rect 46296 15904 46348 15910
rect 46296 15846 46348 15852
rect 46308 15570 46336 15846
rect 46296 15564 46348 15570
rect 46296 15506 46348 15512
rect 46400 15162 46428 25230
rect 46480 24608 46532 24614
rect 46480 24550 46532 24556
rect 46492 24274 46520 24550
rect 46480 24268 46532 24274
rect 46480 24210 46532 24216
rect 46676 22094 46704 41074
rect 46848 39432 46900 39438
rect 46848 39374 46900 39380
rect 46860 38865 46888 39374
rect 46846 38856 46902 38865
rect 46846 38791 46902 38800
rect 46952 38434 46980 48486
rect 47032 45892 47084 45898
rect 47032 45834 47084 45840
rect 47044 45558 47072 45834
rect 47032 45552 47084 45558
rect 47032 45494 47084 45500
rect 47032 40588 47084 40594
rect 47032 40530 47084 40536
rect 47044 40050 47072 40530
rect 47032 40044 47084 40050
rect 47032 39986 47084 39992
rect 46952 38406 47072 38434
rect 46940 38276 46992 38282
rect 46940 38218 46992 38224
rect 46952 38010 46980 38218
rect 46940 38004 46992 38010
rect 46940 37946 46992 37952
rect 47044 37890 47072 38406
rect 46952 37862 47072 37890
rect 46846 37496 46902 37505
rect 46846 37431 46902 37440
rect 46860 37330 46888 37431
rect 46848 37324 46900 37330
rect 46848 37266 46900 37272
rect 46756 34604 46808 34610
rect 46756 34546 46808 34552
rect 46584 22066 46704 22094
rect 46480 21888 46532 21894
rect 46480 21830 46532 21836
rect 46492 20466 46520 21830
rect 46480 20460 46532 20466
rect 46480 20402 46532 20408
rect 46480 16516 46532 16522
rect 46480 16458 46532 16464
rect 46492 16250 46520 16458
rect 46480 16244 46532 16250
rect 46480 16186 46532 16192
rect 46584 16182 46612 22066
rect 46768 17252 46796 34546
rect 46952 29306 46980 37862
rect 47032 37800 47084 37806
rect 47032 37742 47084 37748
rect 46940 29300 46992 29306
rect 46940 29242 46992 29248
rect 46940 29164 46992 29170
rect 46940 29106 46992 29112
rect 46846 26616 46902 26625
rect 46846 26551 46902 26560
rect 46860 25838 46888 26551
rect 46952 26382 46980 29106
rect 46940 26376 46992 26382
rect 46940 26318 46992 26324
rect 47044 26246 47072 37742
rect 47032 26240 47084 26246
rect 47032 26182 47084 26188
rect 47032 26036 47084 26042
rect 47032 25978 47084 25984
rect 46848 25832 46900 25838
rect 46848 25774 46900 25780
rect 47044 25498 47072 25978
rect 47032 25492 47084 25498
rect 47032 25434 47084 25440
rect 46940 23316 46992 23322
rect 46940 23258 46992 23264
rect 46848 22636 46900 22642
rect 46848 22578 46900 22584
rect 46860 21690 46888 22578
rect 46848 21684 46900 21690
rect 46848 21626 46900 21632
rect 46860 21010 46888 21626
rect 46952 21010 46980 23258
rect 46848 21004 46900 21010
rect 46848 20946 46900 20952
rect 46940 21004 46992 21010
rect 46940 20946 46992 20952
rect 46848 20460 46900 20466
rect 46848 20402 46900 20408
rect 46860 19990 46888 20402
rect 47032 20256 47084 20262
rect 47032 20198 47084 20204
rect 46848 19984 46900 19990
rect 46848 19926 46900 19932
rect 46940 19780 46992 19786
rect 46940 19722 46992 19728
rect 46952 19514 46980 19722
rect 46940 19508 46992 19514
rect 46940 19450 46992 19456
rect 47044 18834 47072 20198
rect 47032 18828 47084 18834
rect 47032 18770 47084 18776
rect 46676 17224 46796 17252
rect 46572 16176 46624 16182
rect 46572 16118 46624 16124
rect 46480 15904 46532 15910
rect 46480 15846 46532 15852
rect 46492 15570 46520 15846
rect 46480 15564 46532 15570
rect 46480 15506 46532 15512
rect 46204 15156 46256 15162
rect 46204 15098 46256 15104
rect 46388 15156 46440 15162
rect 46388 15098 46440 15104
rect 46216 13938 46244 15098
rect 46204 13932 46256 13938
rect 46204 13874 46256 13880
rect 46570 13016 46626 13025
rect 46570 12951 46626 12960
rect 46296 11552 46348 11558
rect 46296 11494 46348 11500
rect 46308 11218 46336 11494
rect 46584 11354 46612 12951
rect 46572 11348 46624 11354
rect 46572 11290 46624 11296
rect 46296 11212 46348 11218
rect 46296 11154 46348 11160
rect 46388 10668 46440 10674
rect 46388 10610 46440 10616
rect 46296 7880 46348 7886
rect 46296 7822 46348 7828
rect 46308 7478 46336 7822
rect 46296 7472 46348 7478
rect 46296 7414 46348 7420
rect 46296 6112 46348 6118
rect 46296 6054 46348 6060
rect 46308 5778 46336 6054
rect 46296 5772 46348 5778
rect 46296 5714 46348 5720
rect 46400 5658 46428 10610
rect 46676 5658 46704 17224
rect 46848 17128 46900 17134
rect 46846 17096 46848 17105
rect 46900 17096 46902 17105
rect 46846 17031 46902 17040
rect 46846 15056 46902 15065
rect 46846 14991 46848 15000
rect 46900 14991 46902 15000
rect 46848 14962 46900 14968
rect 46756 14340 46808 14346
rect 46756 14282 46808 14288
rect 46768 14074 46796 14282
rect 46756 14068 46808 14074
rect 46756 14010 46808 14016
rect 47030 13696 47086 13705
rect 47030 13631 47086 13640
rect 46848 12436 46900 12442
rect 46848 12378 46900 12384
rect 46860 12345 46888 12378
rect 46846 12336 46902 12345
rect 46846 12271 46902 12280
rect 46940 11076 46992 11082
rect 46940 11018 46992 11024
rect 46952 10810 46980 11018
rect 46940 10804 46992 10810
rect 46940 10746 46992 10752
rect 46846 9616 46902 9625
rect 46846 9551 46902 9560
rect 46860 9110 46888 9551
rect 46848 9104 46900 9110
rect 46848 9046 46900 9052
rect 46756 7812 46808 7818
rect 46756 7754 46808 7760
rect 46768 7546 46796 7754
rect 46756 7540 46808 7546
rect 46756 7482 46808 7488
rect 46848 6860 46900 6866
rect 46848 6802 46900 6808
rect 46860 6225 46888 6802
rect 46846 6216 46902 6225
rect 46846 6151 46902 6160
rect 46308 5630 46428 5658
rect 46492 5630 46704 5658
rect 46940 5636 46992 5642
rect 46110 4176 46166 4185
rect 45836 4140 45888 4146
rect 46110 4111 46166 4120
rect 45836 4082 45888 4088
rect 46308 4010 46336 5630
rect 46296 4004 46348 4010
rect 46296 3946 46348 3952
rect 46204 3936 46256 3942
rect 46204 3878 46256 3884
rect 46216 3602 46244 3878
rect 46492 3754 46520 5630
rect 46940 5578 46992 5584
rect 46952 5370 46980 5578
rect 46664 5364 46716 5370
rect 46664 5306 46716 5312
rect 46940 5364 46992 5370
rect 46940 5306 46992 5312
rect 46400 3726 46520 3754
rect 46204 3596 46256 3602
rect 46204 3538 46256 3544
rect 46400 3466 46428 3726
rect 46480 3596 46532 3602
rect 46480 3538 46532 3544
rect 46388 3460 46440 3466
rect 46388 3402 46440 3408
rect 45652 3188 45704 3194
rect 45652 3130 45704 3136
rect 45744 3052 45796 3058
rect 45744 2994 45796 3000
rect 44640 2508 44692 2514
rect 44640 2450 44692 2456
rect 45192 2508 45244 2514
rect 45192 2450 45244 2456
rect 45376 2508 45428 2514
rect 45376 2450 45428 2456
rect 45112 870 45232 898
rect 45112 800 45140 870
rect 11256 734 11560 762
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 23846 0 23902 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 25778 0 25834 800
rect 26422 0 26478 800
rect 27066 0 27122 800
rect 27710 0 27766 800
rect 28354 0 28410 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30286 0 30342 800
rect 30930 0 30986 800
rect 31574 0 31630 800
rect 32218 0 32274 800
rect 32862 0 32918 800
rect 33506 0 33562 800
rect 34150 0 34206 800
rect 34794 0 34850 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 36726 0 36782 800
rect 37370 0 37426 800
rect 38014 0 38070 800
rect 38658 0 38714 800
rect 39946 0 40002 800
rect 40590 0 40646 800
rect 41234 0 41290 800
rect 41878 0 41934 800
rect 42522 0 42578 800
rect 43166 0 43222 800
rect 43810 0 43866 800
rect 44454 0 44510 800
rect 45098 0 45154 800
rect 45204 762 45232 870
rect 45388 762 45416 2450
rect 45756 800 45784 2994
rect 46388 2644 46440 2650
rect 46388 2586 46440 2592
rect 46400 1465 46428 2586
rect 46386 1456 46442 1465
rect 46386 1391 46442 1400
rect 46492 1306 46520 3538
rect 46676 3505 46704 5306
rect 46848 5228 46900 5234
rect 46848 5170 46900 5176
rect 46860 4758 46888 5170
rect 46848 4752 46900 4758
rect 46848 4694 46900 4700
rect 46756 4208 46808 4214
rect 46756 4150 46808 4156
rect 46662 3496 46718 3505
rect 46662 3431 46718 3440
rect 46400 1278 46520 1306
rect 46400 800 46428 1278
rect 45204 734 45416 762
rect 45742 0 45798 800
rect 46386 0 46442 800
rect 46768 105 46796 4150
rect 46860 4146 46888 4694
rect 46940 4548 46992 4554
rect 46940 4490 46992 4496
rect 46952 4146 46980 4490
rect 46848 4140 46900 4146
rect 46848 4082 46900 4088
rect 46940 4140 46992 4146
rect 46940 4082 46992 4088
rect 47044 800 47072 13631
rect 47136 3126 47164 49030
rect 48976 48822 49004 51200
rect 48964 48816 49016 48822
rect 48964 48758 49016 48764
rect 47216 48544 47268 48550
rect 47216 48486 47268 48492
rect 47228 37806 47256 48486
rect 47858 48376 47914 48385
rect 47858 48311 47914 48320
rect 47676 48068 47728 48074
rect 47676 48010 47728 48016
rect 47688 46714 47716 48010
rect 47872 47666 47900 48311
rect 47860 47660 47912 47666
rect 47860 47602 47912 47608
rect 48044 47456 48096 47462
rect 48044 47398 48096 47404
rect 47676 46708 47728 46714
rect 47676 46650 47728 46656
rect 47768 45484 47820 45490
rect 47768 45426 47820 45432
rect 47676 44804 47728 44810
rect 47676 44746 47728 44752
rect 47688 44538 47716 44746
rect 47676 44532 47728 44538
rect 47676 44474 47728 44480
rect 47584 44396 47636 44402
rect 47584 44338 47636 44344
rect 47308 43784 47360 43790
rect 47308 43726 47360 43732
rect 47492 43784 47544 43790
rect 47492 43726 47544 43732
rect 47216 37800 47268 37806
rect 47216 37742 47268 37748
rect 47216 37460 47268 37466
rect 47216 37402 47268 37408
rect 47228 14278 47256 37402
rect 47320 26314 47348 43726
rect 47400 43648 47452 43654
rect 47400 43590 47452 43596
rect 47412 42770 47440 43590
rect 47400 42764 47452 42770
rect 47400 42706 47452 42712
rect 47504 42634 47532 43726
rect 47492 42628 47544 42634
rect 47492 42570 47544 42576
rect 47400 37664 47452 37670
rect 47400 37606 47452 37612
rect 47412 35894 47440 37606
rect 47596 36786 47624 44338
rect 47676 43104 47728 43110
rect 47676 43046 47728 43052
rect 47688 40610 47716 43046
rect 47780 40746 47808 45426
rect 47860 43308 47912 43314
rect 47860 43250 47912 43256
rect 47872 42945 47900 43250
rect 47858 42936 47914 42945
rect 47858 42871 47914 42880
rect 47950 42256 48006 42265
rect 47950 42191 47952 42200
rect 48004 42191 48006 42200
rect 47952 42162 48004 42168
rect 47860 41132 47912 41138
rect 47860 41074 47912 41080
rect 47872 40905 47900 41074
rect 47858 40896 47914 40905
rect 47858 40831 47914 40840
rect 47780 40718 47900 40746
rect 47688 40582 47808 40610
rect 47676 40452 47728 40458
rect 47676 40394 47728 40400
rect 47688 40050 47716 40394
rect 47676 40044 47728 40050
rect 47676 39986 47728 39992
rect 47780 38842 47808 40582
rect 47688 38814 47808 38842
rect 47688 37466 47716 38814
rect 47768 38752 47820 38758
rect 47768 38694 47820 38700
rect 47780 38418 47808 38694
rect 47768 38412 47820 38418
rect 47768 38354 47820 38360
rect 47676 37460 47728 37466
rect 47676 37402 47728 37408
rect 47676 37256 47728 37262
rect 47676 37198 47728 37204
rect 47584 36780 47636 36786
rect 47584 36722 47636 36728
rect 47412 35866 47532 35894
rect 47400 31816 47452 31822
rect 47400 31758 47452 31764
rect 47412 31385 47440 31758
rect 47398 31376 47454 31385
rect 47398 31311 47454 31320
rect 47400 29300 47452 29306
rect 47400 29242 47452 29248
rect 47308 26308 47360 26314
rect 47308 26250 47360 26256
rect 47412 25430 47440 29242
rect 47504 26586 47532 35866
rect 47492 26580 47544 26586
rect 47492 26522 47544 26528
rect 47492 25832 47544 25838
rect 47492 25774 47544 25780
rect 47400 25424 47452 25430
rect 47400 25366 47452 25372
rect 47504 24818 47532 25774
rect 47492 24812 47544 24818
rect 47492 24754 47544 24760
rect 47504 23662 47532 24754
rect 47492 23656 47544 23662
rect 47492 23598 47544 23604
rect 47504 22094 47532 23598
rect 47412 22066 47532 22094
rect 47308 20460 47360 20466
rect 47308 20402 47360 20408
rect 47320 18290 47348 20402
rect 47308 18284 47360 18290
rect 47308 18226 47360 18232
rect 47320 16114 47348 18226
rect 47412 16114 47440 22066
rect 47596 17202 47624 36722
rect 47688 36310 47716 37198
rect 47676 36304 47728 36310
rect 47676 36246 47728 36252
rect 47768 34400 47820 34406
rect 47768 34342 47820 34348
rect 47780 34134 47808 34342
rect 47768 34128 47820 34134
rect 47768 34070 47820 34076
rect 47768 33312 47820 33318
rect 47768 33254 47820 33260
rect 47780 32978 47808 33254
rect 47768 32972 47820 32978
rect 47768 32914 47820 32920
rect 47872 31754 47900 40718
rect 47950 38176 48006 38185
rect 47950 38111 48006 38120
rect 47964 37942 47992 38111
rect 47952 37936 48004 37942
rect 47952 37878 48004 37884
rect 47950 36136 48006 36145
rect 47950 36071 48006 36080
rect 47964 35766 47992 36071
rect 47952 35760 48004 35766
rect 47952 35702 48004 35708
rect 48056 34218 48084 47398
rect 49620 47190 49648 51200
rect 49608 47184 49660 47190
rect 49608 47126 49660 47132
rect 48134 46336 48190 46345
rect 48134 46271 48190 46280
rect 48148 46034 48176 46271
rect 48136 46028 48188 46034
rect 48136 45970 48188 45976
rect 48134 45656 48190 45665
rect 48134 45591 48190 45600
rect 48148 44946 48176 45591
rect 48136 44940 48188 44946
rect 48136 44882 48188 44888
rect 48134 43616 48190 43625
rect 48134 43551 48190 43560
rect 48148 42770 48176 43551
rect 48136 42764 48188 42770
rect 48136 42706 48188 42712
rect 48134 41576 48190 41585
rect 48134 41511 48136 41520
rect 48188 41511 48190 41520
rect 48136 41482 48188 41488
rect 48228 40928 48280 40934
rect 48228 40870 48280 40876
rect 48136 40452 48188 40458
rect 48136 40394 48188 40400
rect 48148 40225 48176 40394
rect 48134 40216 48190 40225
rect 48134 40151 48190 40160
rect 48134 39536 48190 39545
rect 48134 39471 48190 39480
rect 48148 38418 48176 39471
rect 48136 38412 48188 38418
rect 48136 38354 48188 38360
rect 48134 36816 48190 36825
rect 48134 36751 48190 36760
rect 48148 36242 48176 36751
rect 48136 36236 48188 36242
rect 48136 36178 48188 36184
rect 48134 35456 48190 35465
rect 48134 35391 48190 35400
rect 48148 35154 48176 35391
rect 48136 35148 48188 35154
rect 48136 35090 48188 35096
rect 48134 34776 48190 34785
rect 48134 34711 48190 34720
rect 47780 31726 47900 31754
rect 47964 34190 48084 34218
rect 47676 27872 47728 27878
rect 47676 27814 47728 27820
rect 47688 24138 47716 27814
rect 47780 25838 47808 31726
rect 47964 30410 47992 34190
rect 48042 34096 48098 34105
rect 48148 34066 48176 34711
rect 48042 34031 48098 34040
rect 48136 34060 48188 34066
rect 48056 32978 48084 34031
rect 48136 34002 48188 34008
rect 48044 32972 48096 32978
rect 48044 32914 48096 32920
rect 48240 31754 48268 40870
rect 47872 30382 47992 30410
rect 48056 31726 48268 31754
rect 47872 28234 47900 30382
rect 47952 30252 48004 30258
rect 47952 30194 48004 30200
rect 47964 30025 47992 30194
rect 47950 30016 48006 30025
rect 47950 29951 48006 29960
rect 48056 29730 48084 31726
rect 47964 29702 48084 29730
rect 47964 28370 47992 29702
rect 48134 29336 48190 29345
rect 48134 29271 48190 29280
rect 48148 28626 48176 29271
rect 48226 28656 48282 28665
rect 48136 28620 48188 28626
rect 48226 28591 48282 28600
rect 48136 28562 48188 28568
rect 47964 28342 48176 28370
rect 47872 28206 48084 28234
rect 47860 28076 47912 28082
rect 47860 28018 47912 28024
rect 47872 27985 47900 28018
rect 47858 27976 47914 27985
rect 47858 27911 47914 27920
rect 48056 27334 48084 28206
rect 48044 27328 48096 27334
rect 48044 27270 48096 27276
rect 48148 26466 48176 28342
rect 48240 27538 48268 28591
rect 48228 27532 48280 27538
rect 48228 27474 48280 27480
rect 48504 26920 48556 26926
rect 48504 26862 48556 26868
rect 48056 26438 48176 26466
rect 47860 26240 47912 26246
rect 47860 26182 47912 26188
rect 47768 25832 47820 25838
rect 47768 25774 47820 25780
rect 47768 25696 47820 25702
rect 47768 25638 47820 25644
rect 47780 24342 47808 25638
rect 47872 25498 47900 26182
rect 47860 25492 47912 25498
rect 47860 25434 47912 25440
rect 47858 25256 47914 25265
rect 47858 25191 47914 25200
rect 47872 24818 47900 25191
rect 47860 24812 47912 24818
rect 47860 24754 47912 24760
rect 48056 24410 48084 26438
rect 48136 26376 48188 26382
rect 48136 26318 48188 26324
rect 48148 25945 48176 26318
rect 48134 25936 48190 25945
rect 48134 25871 48190 25880
rect 48134 24576 48190 24585
rect 48134 24511 48190 24520
rect 48044 24404 48096 24410
rect 48044 24346 48096 24352
rect 47768 24336 47820 24342
rect 47768 24278 47820 24284
rect 48148 24274 48176 24511
rect 48136 24268 48188 24274
rect 48136 24210 48188 24216
rect 47676 24132 47728 24138
rect 47676 24074 47728 24080
rect 47950 23896 48006 23905
rect 47950 23831 48006 23840
rect 47964 23798 47992 23831
rect 47952 23792 48004 23798
rect 47952 23734 48004 23740
rect 47952 22636 48004 22642
rect 47952 22578 48004 22584
rect 47964 22545 47992 22578
rect 47950 22536 48006 22545
rect 47950 22471 48006 22480
rect 47952 21956 48004 21962
rect 47952 21898 48004 21904
rect 47964 21865 47992 21898
rect 47950 21856 48006 21865
rect 47950 21791 48006 21800
rect 47768 21344 47820 21350
rect 47768 21286 47820 21292
rect 47676 20868 47728 20874
rect 47676 20810 47728 20816
rect 47688 20602 47716 20810
rect 47676 20596 47728 20602
rect 47676 20538 47728 20544
rect 47780 19922 47808 21286
rect 47768 19916 47820 19922
rect 47768 19858 47820 19864
rect 48136 19848 48188 19854
rect 48134 19816 48136 19825
rect 48188 19816 48190 19825
rect 48134 19751 48190 19760
rect 47952 19372 48004 19378
rect 47952 19314 48004 19320
rect 47964 19145 47992 19314
rect 48044 19168 48096 19174
rect 47950 19136 48006 19145
rect 48044 19110 48096 19116
rect 47950 19071 48006 19080
rect 47676 18080 47728 18086
rect 47676 18022 47728 18028
rect 47688 17746 47716 18022
rect 47676 17740 47728 17746
rect 47676 17682 47728 17688
rect 47584 17196 47636 17202
rect 47584 17138 47636 17144
rect 47596 16726 47624 17138
rect 47584 16720 47636 16726
rect 47584 16662 47636 16668
rect 47308 16108 47360 16114
rect 47308 16050 47360 16056
rect 47400 16108 47452 16114
rect 47400 16050 47452 16056
rect 47216 14272 47268 14278
rect 47216 14214 47268 14220
rect 47412 12434 47440 16050
rect 47768 14816 47820 14822
rect 47768 14758 47820 14764
rect 47780 14482 47808 14758
rect 47768 14476 47820 14482
rect 47768 14418 47820 14424
rect 47860 13932 47912 13938
rect 47860 13874 47912 13880
rect 47872 13705 47900 13874
rect 47858 13696 47914 13705
rect 47858 13631 47914 13640
rect 47412 12406 47532 12434
rect 47504 3670 47532 12406
rect 48056 10742 48084 19110
rect 48134 17776 48190 17785
rect 48134 17711 48136 17720
rect 48188 17711 48190 17720
rect 48136 17682 48188 17688
rect 48134 16416 48190 16425
rect 48134 16351 48190 16360
rect 48148 15570 48176 16351
rect 48136 15564 48188 15570
rect 48136 15506 48188 15512
rect 48134 14376 48190 14385
rect 48134 14311 48136 14320
rect 48188 14311 48190 14320
rect 48136 14282 48188 14288
rect 48136 11076 48188 11082
rect 48136 11018 48188 11024
rect 48148 10985 48176 11018
rect 48134 10976 48190 10985
rect 48134 10911 48190 10920
rect 48044 10736 48096 10742
rect 48044 10678 48096 10684
rect 47860 10668 47912 10674
rect 47860 10610 47912 10616
rect 47872 10305 47900 10610
rect 47858 10296 47914 10305
rect 47858 10231 47914 10240
rect 47766 8936 47822 8945
rect 47766 8871 47768 8880
rect 47820 8871 47822 8880
rect 47768 8842 47820 8848
rect 47860 8492 47912 8498
rect 47860 8434 47912 8440
rect 47872 8265 47900 8434
rect 47858 8256 47914 8265
rect 47858 8191 47914 8200
rect 48136 7812 48188 7818
rect 48136 7754 48188 7760
rect 48148 7585 48176 7754
rect 48134 7576 48190 7585
rect 48134 7511 48190 7520
rect 48136 5636 48188 5642
rect 48136 5578 48188 5584
rect 47858 5536 47914 5545
rect 47858 5471 47914 5480
rect 47872 5234 47900 5471
rect 47860 5228 47912 5234
rect 47860 5170 47912 5176
rect 48148 4865 48176 5578
rect 48134 4856 48190 4865
rect 48134 4791 48190 4800
rect 48320 4548 48372 4554
rect 48320 4490 48372 4496
rect 47492 3664 47544 3670
rect 47492 3606 47544 3612
rect 47124 3120 47176 3126
rect 47124 3062 47176 3068
rect 47768 2372 47820 2378
rect 47768 2314 47820 2320
rect 46754 96 46810 105
rect 46754 31 46810 40
rect 47030 0 47086 800
rect 47674 0 47730 800
rect 47780 785 47808 2314
rect 47860 2304 47912 2310
rect 47860 2246 47912 2252
rect 47872 1970 47900 2246
rect 47860 1964 47912 1970
rect 47860 1906 47912 1912
rect 48332 800 48360 4490
rect 47766 776 47822 785
rect 47766 711 47822 720
rect 48318 0 48374 800
rect 48516 762 48544 26862
rect 49608 3052 49660 3058
rect 49608 2994 49660 3000
rect 48884 870 49004 898
rect 48884 762 48912 870
rect 48976 800 49004 870
rect 49620 800 49648 2994
rect 48516 734 48912 762
rect 48962 0 49018 800
rect 49606 0 49662 800
<< via2 >>
rect 3790 51720 3846 51776
rect 1398 45600 1454 45656
rect 1398 44240 1454 44296
rect 1398 43560 1454 43616
rect 1398 40840 1454 40896
rect 1398 37440 1454 37496
rect 3422 51040 3478 51096
rect 2778 49000 2834 49056
rect 4066 50360 4122 50416
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 3882 48320 3938 48376
rect 1858 47660 1914 47696
rect 1858 47640 1860 47660
rect 1860 47640 1912 47660
rect 1912 47640 1914 47660
rect 1398 31340 1454 31376
rect 1398 31320 1400 31340
rect 1400 31320 1452 31340
rect 1452 31320 1454 31340
rect 1398 25900 1454 25936
rect 1398 25880 1400 25900
rect 1400 25880 1452 25900
rect 1452 25880 1454 25900
rect 1398 23840 1454 23896
rect 1858 41520 1914 41576
rect 1858 40160 1914 40216
rect 1858 36760 1914 36816
rect 1858 34720 1914 34776
rect 1858 22480 1914 22536
rect 2778 46960 2834 47016
rect 2778 46280 2834 46336
rect 3054 44920 3110 44976
rect 2778 39500 2834 39536
rect 2778 39480 2780 39500
rect 2780 39480 2832 39500
rect 2832 39480 2834 39500
rect 2778 36080 2834 36136
rect 2778 34040 2834 34096
rect 2778 33396 2780 33416
rect 2780 33396 2832 33416
rect 2832 33396 2834 33416
rect 2778 33360 2834 33396
rect 1858 17040 1914 17096
rect 1858 16360 1914 16416
rect 1398 12280 1454 12336
rect 1398 10920 1454 10976
rect 2778 32680 2834 32736
rect 2870 32000 2926 32056
rect 2778 29960 2834 30016
rect 2778 28620 2834 28656
rect 2778 28600 2780 28620
rect 2780 28600 2832 28620
rect 2832 28600 2834 28620
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 2778 27240 2834 27296
rect 2778 26560 2834 26616
rect 2778 23160 2834 23216
rect 2870 21800 2926 21856
rect 1858 8200 1914 8256
rect 1858 7520 1914 7576
rect 2778 19760 2834 19816
rect 2778 19080 2834 19136
rect 2778 17740 2834 17776
rect 2778 17720 2780 17740
rect 2780 17720 2832 17740
rect 2832 17720 2834 17740
rect 3514 38120 3570 38176
rect 3422 29280 3478 29336
rect 3422 21120 3478 21176
rect 3422 18400 3478 18456
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 2778 13640 2834 13696
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 3054 12960 3110 13016
rect 2778 10240 2834 10296
rect 2778 9560 2834 9616
rect 3146 8880 3202 8936
rect 2778 6840 2834 6896
rect 3422 6160 3478 6216
rect 2778 5480 2834 5536
rect 2778 4800 2834 4856
rect 3422 4120 3478 4176
rect 1858 3440 1914 3496
rect 3422 2080 3478 2136
rect 1398 720 1454 776
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 10414 2352 10470 2408
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19706 34992 19762 35048
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19338 34584 19394 34640
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19338 29960 19394 30016
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 20350 32428 20406 32464
rect 20350 32408 20352 32428
rect 20352 32408 20404 32428
rect 20404 32408 20406 32428
rect 21178 34060 21234 34096
rect 21178 34040 21180 34060
rect 21180 34040 21232 34060
rect 21232 34040 21234 34060
rect 17958 19372 18014 19408
rect 17958 19352 17960 19372
rect 17960 19352 18012 19372
rect 18012 19352 18014 19372
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19798 25236 19800 25256
rect 19800 25236 19852 25256
rect 19852 25236 19854 25256
rect 19798 25200 19854 25236
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19706 24676 19762 24712
rect 19706 24656 19708 24676
rect 19708 24656 19760 24676
rect 19760 24656 19762 24676
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19890 23568 19946 23624
rect 19890 23468 19892 23488
rect 19892 23468 19944 23488
rect 19944 23468 19946 23488
rect 19890 23432 19946 23468
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 18786 19388 18788 19408
rect 18788 19388 18840 19408
rect 18840 19388 18842 19408
rect 18786 19352 18842 19388
rect 19890 22480 19946 22536
rect 20074 21936 20130 21992
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19890 19352 19946 19408
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19890 15988 19892 16008
rect 19892 15988 19944 16008
rect 19944 15988 19946 16008
rect 19890 15952 19946 15988
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19430 14456 19486 14512
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 20074 14764 20076 14784
rect 20076 14764 20128 14784
rect 20128 14764 20130 14784
rect 20074 14728 20130 14764
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19522 9968 19578 10024
rect 19706 10004 19708 10024
rect 19708 10004 19760 10024
rect 19760 10004 19762 10024
rect 19706 9968 19762 10004
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19798 9632 19854 9688
rect 19982 9632 20038 9688
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19982 7248 20038 7304
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 20350 11464 20406 11520
rect 20258 9424 20314 9480
rect 20718 24656 20774 24712
rect 20902 23860 20958 23896
rect 20902 23840 20904 23860
rect 20904 23840 20956 23860
rect 20956 23840 20958 23860
rect 20534 22038 20590 22094
rect 20442 7656 20498 7712
rect 20442 7248 20498 7304
rect 21454 14884 21510 14920
rect 21454 14864 21456 14884
rect 21456 14864 21508 14884
rect 21508 14864 21510 14884
rect 21638 21800 21694 21856
rect 22282 31764 22284 31784
rect 22284 31764 22336 31784
rect 22336 31764 22338 31784
rect 22282 31728 22338 31764
rect 22650 31728 22706 31784
rect 22926 32544 22982 32600
rect 22834 26580 22890 26616
rect 22834 26560 22836 26580
rect 22836 26560 22888 26580
rect 22888 26560 22890 26580
rect 21914 20168 21970 20224
rect 21914 20052 21970 20088
rect 21914 20032 21916 20052
rect 21916 20032 21968 20052
rect 21968 20032 21970 20052
rect 21822 19760 21878 19816
rect 22190 19760 22246 19816
rect 22558 20476 22560 20496
rect 22560 20476 22612 20496
rect 22612 20476 22614 20496
rect 22558 20440 22614 20476
rect 22558 20304 22614 20360
rect 22558 19896 22614 19952
rect 24582 34040 24638 34096
rect 24030 32444 24032 32464
rect 24032 32444 24084 32464
rect 24084 32444 24086 32464
rect 24030 32408 24086 32444
rect 23570 26560 23626 26616
rect 22834 19796 22836 19816
rect 22836 19796 22888 19816
rect 22888 19796 22890 19816
rect 22834 19760 22890 19796
rect 22926 19352 22982 19408
rect 23570 19896 23626 19952
rect 21178 2916 21234 2952
rect 21178 2896 21180 2916
rect 21180 2896 21232 2916
rect 21232 2896 21234 2916
rect 22190 8916 22192 8936
rect 22192 8916 22244 8936
rect 22244 8916 22246 8936
rect 22190 8880 22246 8916
rect 22650 8900 22706 8936
rect 22650 8880 22652 8900
rect 22652 8880 22704 8900
rect 22704 8880 22706 8900
rect 23754 8880 23810 8936
rect 22650 2896 22706 2952
rect 24398 32544 24454 32600
rect 25226 31764 25228 31784
rect 25228 31764 25280 31784
rect 25280 31764 25282 31784
rect 25226 31728 25282 31764
rect 24674 23724 24730 23760
rect 24674 23704 24676 23724
rect 24676 23704 24728 23724
rect 24728 23704 24730 23724
rect 24306 20440 24362 20496
rect 24490 20168 24546 20224
rect 24858 24384 24914 24440
rect 24858 22344 24914 22400
rect 24214 10240 24270 10296
rect 24582 9424 24638 9480
rect 24398 8472 24454 8528
rect 25778 23568 25834 23624
rect 25318 20304 25374 20360
rect 26054 23568 26110 23624
rect 25778 19488 25834 19544
rect 25042 9560 25098 9616
rect 25226 9424 25282 9480
rect 25042 8472 25098 8528
rect 25134 8336 25190 8392
rect 25686 8900 25742 8936
rect 25686 8880 25688 8900
rect 25688 8880 25740 8900
rect 25740 8880 25742 8900
rect 25778 8472 25834 8528
rect 26422 26560 26478 26616
rect 26422 23568 26478 23624
rect 26422 15308 26424 15328
rect 26424 15308 26476 15328
rect 26476 15308 26478 15328
rect 26422 15272 26478 15308
rect 26606 23704 26662 23760
rect 27342 29996 27344 30016
rect 27344 29996 27396 30016
rect 27396 29996 27398 30016
rect 27342 29960 27398 29996
rect 27434 24384 27490 24440
rect 27526 23704 27582 23760
rect 27158 23432 27214 23488
rect 27066 19488 27122 19544
rect 26974 19372 27030 19408
rect 26974 19352 26976 19372
rect 26976 19352 27028 19372
rect 27028 19352 27030 19372
rect 26238 10240 26294 10296
rect 26054 8472 26110 8528
rect 27802 24656 27858 24712
rect 27802 23840 27858 23896
rect 27710 19352 27766 19408
rect 27526 14864 27582 14920
rect 27526 9560 27582 9616
rect 27250 8372 27252 8392
rect 27252 8372 27304 8392
rect 27304 8372 27306 8392
rect 27250 8336 27306 8372
rect 28170 23296 28226 23352
rect 28538 24112 28594 24168
rect 28538 23976 28594 24032
rect 28262 21800 28318 21856
rect 28262 21664 28318 21720
rect 28998 24520 29054 24576
rect 28998 24248 29054 24304
rect 28906 24112 28962 24168
rect 28814 23568 28870 23624
rect 28722 23196 28724 23216
rect 28724 23196 28776 23216
rect 28776 23196 28778 23216
rect 28722 23160 28778 23196
rect 28538 21664 28594 21720
rect 28722 20032 28778 20088
rect 28722 15272 28778 15328
rect 28998 23860 29054 23896
rect 28998 23840 29000 23860
rect 29000 23840 29052 23860
rect 29052 23840 29054 23860
rect 31022 31728 31078 31784
rect 29366 27920 29422 27976
rect 29274 24112 29330 24168
rect 29182 23976 29238 24032
rect 28998 23296 29054 23352
rect 29182 23296 29238 23352
rect 29550 23976 29606 24032
rect 29274 23160 29330 23216
rect 30010 26696 30066 26752
rect 30102 26460 30104 26480
rect 30104 26460 30156 26480
rect 30156 26460 30158 26480
rect 30102 26424 30158 26460
rect 30102 25780 30104 25800
rect 30104 25780 30156 25800
rect 30156 25780 30158 25800
rect 30102 25744 30158 25780
rect 30102 23468 30104 23488
rect 30104 23468 30156 23488
rect 30156 23468 30158 23488
rect 30102 23432 30158 23468
rect 30746 26288 30802 26344
rect 29458 3460 29514 3496
rect 29458 3440 29460 3460
rect 29460 3440 29512 3460
rect 29512 3440 29514 3460
rect 30286 3984 30342 4040
rect 32586 31184 32642 31240
rect 33598 31764 33600 31784
rect 33600 31764 33652 31784
rect 33652 31764 33654 31784
rect 33598 31728 33654 31764
rect 33230 26968 33286 27024
rect 33138 25200 33194 25256
rect 32586 21972 32588 21992
rect 32588 21972 32640 21992
rect 32640 21972 32642 21992
rect 32586 21936 32642 21972
rect 33598 25336 33654 25392
rect 33874 26696 33930 26752
rect 32310 3440 32366 3496
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34426 26732 34428 26752
rect 34428 26732 34480 26752
rect 34480 26732 34482 26752
rect 34426 26696 34482 26732
rect 34518 23840 34574 23896
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 35622 31184 35678 31240
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34702 26188 34704 26208
rect 34704 26188 34756 26208
rect 34756 26188 34758 26208
rect 34702 26152 34758 26188
rect 35530 27920 35586 27976
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 35530 27104 35586 27160
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 35070 26288 35126 26344
rect 35162 26152 35218 26208
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 35346 23704 35402 23760
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 36082 26288 36138 26344
rect 35806 25492 35862 25528
rect 35806 25472 35808 25492
rect 35808 25472 35860 25492
rect 35860 25472 35862 25492
rect 35898 25200 35954 25256
rect 35714 24656 35770 24712
rect 37002 26868 37004 26888
rect 37004 26868 37056 26888
rect 37056 26868 37058 26888
rect 37002 26832 37058 26868
rect 37002 26324 37004 26344
rect 37004 26324 37056 26344
rect 37056 26324 37058 26344
rect 37002 26288 37058 26324
rect 36542 25472 36598 25528
rect 37002 25744 37058 25800
rect 37738 26968 37794 27024
rect 37922 26832 37978 26888
rect 38106 27104 38162 27160
rect 38106 25336 38162 25392
rect 38566 23976 38622 24032
rect 38474 21936 38530 21992
rect 38014 19780 38070 19816
rect 38014 19760 38016 19780
rect 38016 19760 38068 19780
rect 38068 19760 38070 19780
rect 38566 19780 38622 19816
rect 38566 19760 38568 19780
rect 38568 19760 38620 19780
rect 38620 19760 38622 19780
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34518 14184 34574 14240
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34886 14456 34942 14512
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 37462 14476 37518 14512
rect 37462 14456 37464 14476
rect 37464 14456 37516 14476
rect 37516 14456 37518 14476
rect 38290 14184 38346 14240
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 36450 3984 36506 4040
rect 39394 24556 39396 24576
rect 39396 24556 39448 24576
rect 39448 24556 39450 24576
rect 39394 24520 39450 24556
rect 39854 24148 39856 24168
rect 39856 24148 39908 24168
rect 39908 24148 39910 24168
rect 39670 23840 39726 23896
rect 39854 24112 39910 24148
rect 40406 23568 40462 23624
rect 40314 22772 40370 22808
rect 40314 22752 40316 22772
rect 40316 22752 40368 22772
rect 40368 22752 40370 22772
rect 41510 26424 41566 26480
rect 41694 26424 41750 26480
rect 40866 24384 40922 24440
rect 40866 23860 40922 23896
rect 40866 23840 40868 23860
rect 40868 23840 40920 23860
rect 40920 23840 40922 23860
rect 41326 24112 41382 24168
rect 41510 23604 41512 23624
rect 41512 23604 41564 23624
rect 41564 23604 41566 23624
rect 41510 23568 41566 23604
rect 42154 24268 42210 24304
rect 42154 24248 42156 24268
rect 42156 24248 42208 24268
rect 42208 24248 42210 24268
rect 42246 24132 42302 24168
rect 42246 24112 42248 24132
rect 42248 24112 42300 24132
rect 42300 24112 42302 24132
rect 42522 24520 42578 24576
rect 43442 24384 43498 24440
rect 43350 24284 43352 24304
rect 43352 24284 43404 24304
rect 43404 24284 43406 24304
rect 43350 24248 43406 24284
rect 43166 24148 43168 24168
rect 43168 24148 43220 24168
rect 43220 24148 43222 24168
rect 42798 23588 42854 23624
rect 42798 23568 42800 23588
rect 42800 23568 42852 23588
rect 42852 23568 42854 23588
rect 43166 24112 43222 24148
rect 43902 23604 43904 23624
rect 43904 23604 43956 23624
rect 43956 23604 43958 23624
rect 43902 23568 43958 23604
rect 43994 22752 44050 22808
rect 46754 51720 46810 51776
rect 45926 51040 45982 51096
rect 46846 50360 46902 50416
rect 46662 49680 46718 49736
rect 46754 49000 46810 49056
rect 46846 46960 46902 47016
rect 46846 44920 46902 44976
rect 46018 44240 46074 44296
rect 46202 33396 46204 33416
rect 46204 33396 46256 33416
rect 46256 33396 46258 33416
rect 46202 33360 46258 33396
rect 46386 32000 46442 32056
rect 46018 6840 46074 6896
rect 46846 38800 46902 38856
rect 46846 37440 46902 37496
rect 46846 26560 46902 26616
rect 46570 12960 46626 13016
rect 46846 17076 46848 17096
rect 46848 17076 46900 17096
rect 46900 17076 46902 17096
rect 46846 17040 46902 17076
rect 46846 15020 46902 15056
rect 46846 15000 46848 15020
rect 46848 15000 46900 15020
rect 46900 15000 46902 15020
rect 47030 13640 47086 13696
rect 46846 12280 46902 12336
rect 46846 9560 46902 9616
rect 46846 6160 46902 6216
rect 46110 4120 46166 4176
rect 46386 1400 46442 1456
rect 46662 3440 46718 3496
rect 47858 48320 47914 48376
rect 47858 42880 47914 42936
rect 47950 42220 48006 42256
rect 47950 42200 47952 42220
rect 47952 42200 48004 42220
rect 48004 42200 48006 42220
rect 47858 40840 47914 40896
rect 47398 31320 47454 31376
rect 47950 38120 48006 38176
rect 47950 36080 48006 36136
rect 48134 46280 48190 46336
rect 48134 45600 48190 45656
rect 48134 43560 48190 43616
rect 48134 41540 48190 41576
rect 48134 41520 48136 41540
rect 48136 41520 48188 41540
rect 48188 41520 48190 41540
rect 48134 40160 48190 40216
rect 48134 39480 48190 39536
rect 48134 36760 48190 36816
rect 48134 35400 48190 35456
rect 48134 34720 48190 34776
rect 48042 34040 48098 34096
rect 47950 29960 48006 30016
rect 48134 29280 48190 29336
rect 48226 28600 48282 28656
rect 47858 27920 47914 27976
rect 47858 25200 47914 25256
rect 48134 25880 48190 25936
rect 48134 24520 48190 24576
rect 47950 23840 48006 23896
rect 47950 22480 48006 22536
rect 47950 21800 48006 21856
rect 48134 19796 48136 19816
rect 48136 19796 48188 19816
rect 48188 19796 48190 19816
rect 48134 19760 48190 19796
rect 47950 19080 48006 19136
rect 47858 13640 47914 13696
rect 48134 17740 48190 17776
rect 48134 17720 48136 17740
rect 48136 17720 48188 17740
rect 48188 17720 48190 17740
rect 48134 16360 48190 16416
rect 48134 14340 48190 14376
rect 48134 14320 48136 14340
rect 48136 14320 48188 14340
rect 48188 14320 48190 14340
rect 48134 10920 48190 10976
rect 47858 10240 47914 10296
rect 47766 8900 47822 8936
rect 47766 8880 47768 8900
rect 47768 8880 47820 8900
rect 47820 8880 47822 8900
rect 47858 8200 47914 8256
rect 48134 7520 48190 7576
rect 47858 5480 47914 5536
rect 48134 4800 48190 4856
rect 46754 40 46810 96
rect 47766 720 47822 776
<< metal3 >>
rect 0 51778 800 51808
rect 3785 51778 3851 51781
rect 0 51776 3851 51778
rect 0 51720 3790 51776
rect 3846 51720 3851 51776
rect 0 51718 3851 51720
rect 0 51688 800 51718
rect 3785 51715 3851 51718
rect 46749 51778 46815 51781
rect 49200 51778 50000 51808
rect 46749 51776 50000 51778
rect 46749 51720 46754 51776
rect 46810 51720 50000 51776
rect 46749 51718 50000 51720
rect 46749 51715 46815 51718
rect 49200 51688 50000 51718
rect 0 51098 800 51128
rect 3417 51098 3483 51101
rect 0 51096 3483 51098
rect 0 51040 3422 51096
rect 3478 51040 3483 51096
rect 0 51038 3483 51040
rect 0 51008 800 51038
rect 3417 51035 3483 51038
rect 45921 51098 45987 51101
rect 49200 51098 50000 51128
rect 45921 51096 50000 51098
rect 45921 51040 45926 51096
rect 45982 51040 50000 51096
rect 45921 51038 50000 51040
rect 45921 51035 45987 51038
rect 49200 51008 50000 51038
rect 0 50418 800 50448
rect 4061 50418 4127 50421
rect 0 50416 4127 50418
rect 0 50360 4066 50416
rect 4122 50360 4127 50416
rect 0 50358 4127 50360
rect 0 50328 800 50358
rect 4061 50355 4127 50358
rect 46841 50418 46907 50421
rect 49200 50418 50000 50448
rect 46841 50416 50000 50418
rect 46841 50360 46846 50416
rect 46902 50360 50000 50416
rect 46841 50358 50000 50360
rect 46841 50355 46907 50358
rect 49200 50328 50000 50358
rect 0 49648 800 49768
rect 46657 49738 46723 49741
rect 49200 49738 50000 49768
rect 46657 49736 50000 49738
rect 46657 49680 46662 49736
rect 46718 49680 50000 49736
rect 46657 49678 50000 49680
rect 46657 49675 46723 49678
rect 49200 49648 50000 49678
rect 4208 49536 4528 49537
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 49471 4528 49472
rect 34928 49536 35248 49537
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 49471 35248 49472
rect 0 49058 800 49088
rect 2773 49058 2839 49061
rect 0 49056 2839 49058
rect 0 49000 2778 49056
rect 2834 49000 2839 49056
rect 0 48998 2839 49000
rect 0 48968 800 48998
rect 2773 48995 2839 48998
rect 46749 49058 46815 49061
rect 49200 49058 50000 49088
rect 46749 49056 50000 49058
rect 46749 49000 46754 49056
rect 46810 49000 50000 49056
rect 46749 48998 50000 49000
rect 46749 48995 46815 48998
rect 19568 48992 19888 48993
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 49200 48968 50000 48998
rect 19568 48927 19888 48928
rect 4208 48448 4528 48449
rect 0 48378 800 48408
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 48383 4528 48384
rect 34928 48448 35248 48449
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 48383 35248 48384
rect 3877 48378 3943 48381
rect 0 48376 3943 48378
rect 0 48320 3882 48376
rect 3938 48320 3943 48376
rect 0 48318 3943 48320
rect 0 48288 800 48318
rect 3877 48315 3943 48318
rect 47853 48378 47919 48381
rect 49200 48378 50000 48408
rect 47853 48376 50000 48378
rect 47853 48320 47858 48376
rect 47914 48320 50000 48376
rect 47853 48318 50000 48320
rect 47853 48315 47919 48318
rect 49200 48288 50000 48318
rect 19568 47904 19888 47905
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 47839 19888 47840
rect 0 47698 800 47728
rect 1853 47698 1919 47701
rect 0 47696 1919 47698
rect 0 47640 1858 47696
rect 1914 47640 1919 47696
rect 0 47638 1919 47640
rect 0 47608 800 47638
rect 1853 47635 1919 47638
rect 49200 47608 50000 47728
rect 4208 47360 4528 47361
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 47295 4528 47296
rect 34928 47360 35248 47361
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 47295 35248 47296
rect 0 47018 800 47048
rect 2773 47018 2839 47021
rect 0 47016 2839 47018
rect 0 46960 2778 47016
rect 2834 46960 2839 47016
rect 0 46958 2839 46960
rect 0 46928 800 46958
rect 2773 46955 2839 46958
rect 46841 47018 46907 47021
rect 49200 47018 50000 47048
rect 46841 47016 50000 47018
rect 46841 46960 46846 47016
rect 46902 46960 50000 47016
rect 46841 46958 50000 46960
rect 46841 46955 46907 46958
rect 49200 46928 50000 46958
rect 19568 46816 19888 46817
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 46751 19888 46752
rect 0 46338 800 46368
rect 2773 46338 2839 46341
rect 0 46336 2839 46338
rect 0 46280 2778 46336
rect 2834 46280 2839 46336
rect 0 46278 2839 46280
rect 0 46248 800 46278
rect 2773 46275 2839 46278
rect 48129 46338 48195 46341
rect 49200 46338 50000 46368
rect 48129 46336 50000 46338
rect 48129 46280 48134 46336
rect 48190 46280 50000 46336
rect 48129 46278 50000 46280
rect 48129 46275 48195 46278
rect 4208 46272 4528 46273
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 46207 4528 46208
rect 34928 46272 35248 46273
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 49200 46248 50000 46278
rect 34928 46207 35248 46208
rect 19568 45728 19888 45729
rect 0 45658 800 45688
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 45663 19888 45664
rect 1393 45658 1459 45661
rect 0 45656 1459 45658
rect 0 45600 1398 45656
rect 1454 45600 1459 45656
rect 0 45598 1459 45600
rect 0 45568 800 45598
rect 1393 45595 1459 45598
rect 48129 45658 48195 45661
rect 49200 45658 50000 45688
rect 48129 45656 50000 45658
rect 48129 45600 48134 45656
rect 48190 45600 50000 45656
rect 48129 45598 50000 45600
rect 48129 45595 48195 45598
rect 49200 45568 50000 45598
rect 4208 45184 4528 45185
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 45119 4528 45120
rect 34928 45184 35248 45185
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 45119 35248 45120
rect 0 44978 800 45008
rect 3049 44978 3115 44981
rect 0 44976 3115 44978
rect 0 44920 3054 44976
rect 3110 44920 3115 44976
rect 0 44918 3115 44920
rect 0 44888 800 44918
rect 3049 44915 3115 44918
rect 46841 44978 46907 44981
rect 49200 44978 50000 45008
rect 46841 44976 50000 44978
rect 46841 44920 46846 44976
rect 46902 44920 50000 44976
rect 46841 44918 50000 44920
rect 46841 44915 46907 44918
rect 49200 44888 50000 44918
rect 19568 44640 19888 44641
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 44575 19888 44576
rect 0 44298 800 44328
rect 1393 44298 1459 44301
rect 0 44296 1459 44298
rect 0 44240 1398 44296
rect 1454 44240 1459 44296
rect 0 44238 1459 44240
rect 0 44208 800 44238
rect 1393 44235 1459 44238
rect 46013 44298 46079 44301
rect 49200 44298 50000 44328
rect 46013 44296 50000 44298
rect 46013 44240 46018 44296
rect 46074 44240 50000 44296
rect 46013 44238 50000 44240
rect 46013 44235 46079 44238
rect 49200 44208 50000 44238
rect 4208 44096 4528 44097
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 44031 4528 44032
rect 34928 44096 35248 44097
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 44031 35248 44032
rect 0 43618 800 43648
rect 1393 43618 1459 43621
rect 0 43616 1459 43618
rect 0 43560 1398 43616
rect 1454 43560 1459 43616
rect 0 43558 1459 43560
rect 0 43528 800 43558
rect 1393 43555 1459 43558
rect 48129 43618 48195 43621
rect 49200 43618 50000 43648
rect 48129 43616 50000 43618
rect 48129 43560 48134 43616
rect 48190 43560 50000 43616
rect 48129 43558 50000 43560
rect 48129 43555 48195 43558
rect 19568 43552 19888 43553
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 49200 43528 50000 43558
rect 19568 43487 19888 43488
rect 4208 43008 4528 43009
rect 0 42848 800 42968
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 42943 4528 42944
rect 34928 43008 35248 43009
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 42943 35248 42944
rect 47853 42938 47919 42941
rect 49200 42938 50000 42968
rect 47853 42936 50000 42938
rect 47853 42880 47858 42936
rect 47914 42880 50000 42936
rect 47853 42878 50000 42880
rect 47853 42875 47919 42878
rect 49200 42848 50000 42878
rect 19568 42464 19888 42465
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 42399 19888 42400
rect 47945 42258 48011 42261
rect 49200 42258 50000 42288
rect 47945 42256 50000 42258
rect 47945 42200 47950 42256
rect 48006 42200 50000 42256
rect 47945 42198 50000 42200
rect 47945 42195 48011 42198
rect 49200 42168 50000 42198
rect 4208 41920 4528 41921
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 41855 4528 41856
rect 34928 41920 35248 41921
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 41855 35248 41856
rect 0 41578 800 41608
rect 1853 41578 1919 41581
rect 0 41576 1919 41578
rect 0 41520 1858 41576
rect 1914 41520 1919 41576
rect 0 41518 1919 41520
rect 0 41488 800 41518
rect 1853 41515 1919 41518
rect 48129 41578 48195 41581
rect 49200 41578 50000 41608
rect 48129 41576 50000 41578
rect 48129 41520 48134 41576
rect 48190 41520 50000 41576
rect 48129 41518 50000 41520
rect 48129 41515 48195 41518
rect 49200 41488 50000 41518
rect 19568 41376 19888 41377
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 41311 19888 41312
rect 0 40898 800 40928
rect 1393 40898 1459 40901
rect 0 40896 1459 40898
rect 0 40840 1398 40896
rect 1454 40840 1459 40896
rect 0 40838 1459 40840
rect 0 40808 800 40838
rect 1393 40835 1459 40838
rect 47853 40898 47919 40901
rect 49200 40898 50000 40928
rect 47853 40896 50000 40898
rect 47853 40840 47858 40896
rect 47914 40840 50000 40896
rect 47853 40838 50000 40840
rect 47853 40835 47919 40838
rect 4208 40832 4528 40833
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 40767 4528 40768
rect 34928 40832 35248 40833
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 49200 40808 50000 40838
rect 34928 40767 35248 40768
rect 19568 40288 19888 40289
rect 0 40218 800 40248
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 40223 19888 40224
rect 1853 40218 1919 40221
rect 0 40216 1919 40218
rect 0 40160 1858 40216
rect 1914 40160 1919 40216
rect 0 40158 1919 40160
rect 0 40128 800 40158
rect 1853 40155 1919 40158
rect 48129 40218 48195 40221
rect 49200 40218 50000 40248
rect 48129 40216 50000 40218
rect 48129 40160 48134 40216
rect 48190 40160 50000 40216
rect 48129 40158 50000 40160
rect 48129 40155 48195 40158
rect 49200 40128 50000 40158
rect 4208 39744 4528 39745
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 0 39538 800 39568
rect 2773 39538 2839 39541
rect 0 39536 2839 39538
rect 0 39480 2778 39536
rect 2834 39480 2839 39536
rect 0 39478 2839 39480
rect 0 39448 800 39478
rect 2773 39475 2839 39478
rect 48129 39538 48195 39541
rect 49200 39538 50000 39568
rect 48129 39536 50000 39538
rect 48129 39480 48134 39536
rect 48190 39480 50000 39536
rect 48129 39478 50000 39480
rect 48129 39475 48195 39478
rect 49200 39448 50000 39478
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 39135 19888 39136
rect 0 38768 800 38888
rect 46841 38858 46907 38861
rect 49200 38858 50000 38888
rect 46841 38856 50000 38858
rect 46841 38800 46846 38856
rect 46902 38800 50000 38856
rect 46841 38798 50000 38800
rect 46841 38795 46907 38798
rect 49200 38768 50000 38798
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 38591 35248 38592
rect 0 38178 800 38208
rect 3509 38178 3575 38181
rect 0 38176 3575 38178
rect 0 38120 3514 38176
rect 3570 38120 3575 38176
rect 0 38118 3575 38120
rect 0 38088 800 38118
rect 3509 38115 3575 38118
rect 47945 38178 48011 38181
rect 49200 38178 50000 38208
rect 47945 38176 50000 38178
rect 47945 38120 47950 38176
rect 48006 38120 50000 38176
rect 47945 38118 50000 38120
rect 47945 38115 48011 38118
rect 19568 38112 19888 38113
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 49200 38088 50000 38118
rect 19568 38047 19888 38048
rect 4208 37568 4528 37569
rect 0 37498 800 37528
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 1393 37498 1459 37501
rect 0 37496 1459 37498
rect 0 37440 1398 37496
rect 1454 37440 1459 37496
rect 0 37438 1459 37440
rect 0 37408 800 37438
rect 1393 37435 1459 37438
rect 46841 37498 46907 37501
rect 49200 37498 50000 37528
rect 46841 37496 50000 37498
rect 46841 37440 46846 37496
rect 46902 37440 50000 37496
rect 46841 37438 50000 37440
rect 46841 37435 46907 37438
rect 49200 37408 50000 37438
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 0 36818 800 36848
rect 1853 36818 1919 36821
rect 0 36816 1919 36818
rect 0 36760 1858 36816
rect 1914 36760 1919 36816
rect 0 36758 1919 36760
rect 0 36728 800 36758
rect 1853 36755 1919 36758
rect 48129 36818 48195 36821
rect 49200 36818 50000 36848
rect 48129 36816 50000 36818
rect 48129 36760 48134 36816
rect 48190 36760 50000 36816
rect 48129 36758 50000 36760
rect 48129 36755 48195 36758
rect 49200 36728 50000 36758
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 0 36138 800 36168
rect 2773 36138 2839 36141
rect 0 36136 2839 36138
rect 0 36080 2778 36136
rect 2834 36080 2839 36136
rect 0 36078 2839 36080
rect 0 36048 800 36078
rect 2773 36075 2839 36078
rect 47945 36138 48011 36141
rect 49200 36138 50000 36168
rect 47945 36136 50000 36138
rect 47945 36080 47950 36136
rect 48006 36080 50000 36136
rect 47945 36078 50000 36080
rect 47945 36075 48011 36078
rect 49200 36048 50000 36078
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 0 35368 800 35488
rect 48129 35458 48195 35461
rect 49200 35458 50000 35488
rect 48129 35456 50000 35458
rect 48129 35400 48134 35456
rect 48190 35400 50000 35456
rect 48129 35398 50000 35400
rect 48129 35395 48195 35398
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 49200 35368 50000 35398
rect 34928 35327 35248 35328
rect 19701 35050 19767 35053
rect 19382 35048 19767 35050
rect 19382 34992 19706 35048
rect 19762 34992 19767 35048
rect 19382 34990 19767 34992
rect 0 34778 800 34808
rect 1853 34778 1919 34781
rect 0 34776 1919 34778
rect 0 34720 1858 34776
rect 1914 34720 1919 34776
rect 0 34718 1919 34720
rect 0 34688 800 34718
rect 1853 34715 1919 34718
rect 19382 34645 19442 34990
rect 19701 34987 19767 34990
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 48129 34778 48195 34781
rect 49200 34778 50000 34808
rect 48129 34776 50000 34778
rect 48129 34720 48134 34776
rect 48190 34720 50000 34776
rect 48129 34718 50000 34720
rect 48129 34715 48195 34718
rect 49200 34688 50000 34718
rect 19333 34640 19442 34645
rect 19333 34584 19338 34640
rect 19394 34584 19442 34640
rect 19333 34582 19442 34584
rect 19333 34579 19399 34582
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 0 34098 800 34128
rect 2773 34098 2839 34101
rect 0 34096 2839 34098
rect 0 34040 2778 34096
rect 2834 34040 2839 34096
rect 0 34038 2839 34040
rect 0 34008 800 34038
rect 2773 34035 2839 34038
rect 21173 34098 21239 34101
rect 24577 34098 24643 34101
rect 21173 34096 24643 34098
rect 21173 34040 21178 34096
rect 21234 34040 24582 34096
rect 24638 34040 24643 34096
rect 21173 34038 24643 34040
rect 21173 34035 21239 34038
rect 24577 34035 24643 34038
rect 48037 34098 48103 34101
rect 49200 34098 50000 34128
rect 48037 34096 50000 34098
rect 48037 34040 48042 34096
rect 48098 34040 50000 34096
rect 48037 34038 50000 34040
rect 48037 34035 48103 34038
rect 49200 34008 50000 34038
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 0 33418 800 33448
rect 2773 33418 2839 33421
rect 0 33416 2839 33418
rect 0 33360 2778 33416
rect 2834 33360 2839 33416
rect 0 33358 2839 33360
rect 0 33328 800 33358
rect 2773 33355 2839 33358
rect 46197 33418 46263 33421
rect 49200 33418 50000 33448
rect 46197 33416 50000 33418
rect 46197 33360 46202 33416
rect 46258 33360 50000 33416
rect 46197 33358 50000 33360
rect 46197 33355 46263 33358
rect 49200 33328 50000 33358
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 0 32738 800 32768
rect 2773 32738 2839 32741
rect 0 32736 2839 32738
rect 0 32680 2778 32736
rect 2834 32680 2839 32736
rect 0 32678 2839 32680
rect 0 32648 800 32678
rect 2773 32675 2839 32678
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 49200 32648 50000 32768
rect 19568 32607 19888 32608
rect 22921 32602 22987 32605
rect 24393 32602 24459 32605
rect 22921 32600 24459 32602
rect 22921 32544 22926 32600
rect 22982 32544 24398 32600
rect 24454 32544 24459 32600
rect 22921 32542 24459 32544
rect 22921 32539 22987 32542
rect 24393 32539 24459 32542
rect 20345 32466 20411 32469
rect 24025 32466 24091 32469
rect 20345 32464 24091 32466
rect 20345 32408 20350 32464
rect 20406 32408 24030 32464
rect 24086 32408 24091 32464
rect 20345 32406 24091 32408
rect 20345 32403 20411 32406
rect 24025 32403 24091 32406
rect 4208 32128 4528 32129
rect 0 32058 800 32088
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 2865 32058 2931 32061
rect 0 32056 2931 32058
rect 0 32000 2870 32056
rect 2926 32000 2931 32056
rect 0 31998 2931 32000
rect 0 31968 800 31998
rect 2865 31995 2931 31998
rect 46381 32058 46447 32061
rect 49200 32058 50000 32088
rect 46381 32056 50000 32058
rect 46381 32000 46386 32056
rect 46442 32000 50000 32056
rect 46381 31998 50000 32000
rect 46381 31995 46447 31998
rect 49200 31968 50000 31998
rect 22277 31786 22343 31789
rect 22645 31786 22711 31789
rect 25221 31786 25287 31789
rect 22277 31784 25287 31786
rect 22277 31728 22282 31784
rect 22338 31728 22650 31784
rect 22706 31728 25226 31784
rect 25282 31728 25287 31784
rect 22277 31726 25287 31728
rect 22277 31723 22343 31726
rect 22645 31723 22711 31726
rect 25221 31723 25287 31726
rect 31017 31786 31083 31789
rect 33593 31786 33659 31789
rect 31017 31784 33659 31786
rect 31017 31728 31022 31784
rect 31078 31728 33598 31784
rect 33654 31728 33659 31784
rect 31017 31726 33659 31728
rect 31017 31723 31083 31726
rect 33593 31723 33659 31726
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 0 31378 800 31408
rect 1393 31378 1459 31381
rect 0 31376 1459 31378
rect 0 31320 1398 31376
rect 1454 31320 1459 31376
rect 0 31318 1459 31320
rect 0 31288 800 31318
rect 1393 31315 1459 31318
rect 47393 31378 47459 31381
rect 49200 31378 50000 31408
rect 47393 31376 50000 31378
rect 47393 31320 47398 31376
rect 47454 31320 50000 31376
rect 47393 31318 50000 31320
rect 47393 31315 47459 31318
rect 49200 31288 50000 31318
rect 32581 31242 32647 31245
rect 35617 31242 35683 31245
rect 32581 31240 35683 31242
rect 32581 31184 32586 31240
rect 32642 31184 35622 31240
rect 35678 31184 35683 31240
rect 32581 31182 35683 31184
rect 32581 31179 32647 31182
rect 35617 31179 35683 31182
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 0 30608 800 30728
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 0 30018 800 30048
rect 2773 30018 2839 30021
rect 0 30016 2839 30018
rect 0 29960 2778 30016
rect 2834 29960 2839 30016
rect 0 29958 2839 29960
rect 0 29928 800 29958
rect 2773 29955 2839 29958
rect 19333 30018 19399 30021
rect 27337 30018 27403 30021
rect 19333 30016 27403 30018
rect 19333 29960 19338 30016
rect 19394 29960 27342 30016
rect 27398 29960 27403 30016
rect 19333 29958 27403 29960
rect 19333 29955 19399 29958
rect 27337 29955 27403 29958
rect 47945 30018 48011 30021
rect 49200 30018 50000 30048
rect 47945 30016 50000 30018
rect 47945 29960 47950 30016
rect 48006 29960 50000 30016
rect 47945 29958 50000 29960
rect 47945 29955 48011 29958
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 49200 29928 50000 29958
rect 34928 29887 35248 29888
rect 19568 29408 19888 29409
rect 0 29338 800 29368
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 3417 29338 3483 29341
rect 0 29336 3483 29338
rect 0 29280 3422 29336
rect 3478 29280 3483 29336
rect 0 29278 3483 29280
rect 0 29248 800 29278
rect 3417 29275 3483 29278
rect 48129 29338 48195 29341
rect 49200 29338 50000 29368
rect 48129 29336 50000 29338
rect 48129 29280 48134 29336
rect 48190 29280 50000 29336
rect 48129 29278 50000 29280
rect 48129 29275 48195 29278
rect 49200 29248 50000 29278
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 0 28658 800 28688
rect 2773 28658 2839 28661
rect 0 28656 2839 28658
rect 0 28600 2778 28656
rect 2834 28600 2839 28656
rect 0 28598 2839 28600
rect 0 28568 800 28598
rect 2773 28595 2839 28598
rect 48221 28658 48287 28661
rect 49200 28658 50000 28688
rect 48221 28656 50000 28658
rect 48221 28600 48226 28656
rect 48282 28600 50000 28656
rect 48221 28598 50000 28600
rect 48221 28595 48287 28598
rect 49200 28568 50000 28598
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 0 27888 800 28008
rect 29361 27978 29427 27981
rect 35525 27978 35591 27981
rect 29361 27976 35591 27978
rect 29361 27920 29366 27976
rect 29422 27920 35530 27976
rect 35586 27920 35591 27976
rect 29361 27918 35591 27920
rect 29361 27915 29427 27918
rect 35525 27915 35591 27918
rect 47853 27978 47919 27981
rect 49200 27978 50000 28008
rect 47853 27976 50000 27978
rect 47853 27920 47858 27976
rect 47914 27920 50000 27976
rect 47853 27918 50000 27920
rect 47853 27915 47919 27918
rect 49200 27888 50000 27918
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 0 27298 800 27328
rect 2773 27298 2839 27301
rect 0 27296 2839 27298
rect 0 27240 2778 27296
rect 2834 27240 2839 27296
rect 0 27238 2839 27240
rect 0 27208 800 27238
rect 2773 27235 2839 27238
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 49200 27208 50000 27328
rect 19568 27167 19888 27168
rect 35525 27162 35591 27165
rect 38101 27162 38167 27165
rect 35525 27160 38167 27162
rect 35525 27104 35530 27160
rect 35586 27104 38106 27160
rect 38162 27104 38167 27160
rect 35525 27102 38167 27104
rect 35525 27099 35591 27102
rect 38101 27099 38167 27102
rect 33225 27026 33291 27029
rect 37733 27026 37799 27029
rect 33225 27024 37799 27026
rect 33225 26968 33230 27024
rect 33286 26968 37738 27024
rect 37794 26968 37799 27024
rect 33225 26966 37799 26968
rect 33225 26963 33291 26966
rect 37733 26963 37799 26966
rect 36997 26890 37063 26893
rect 37917 26890 37983 26893
rect 36997 26888 37983 26890
rect 36997 26832 37002 26888
rect 37058 26832 37922 26888
rect 37978 26832 37983 26888
rect 36997 26830 37983 26832
rect 36997 26827 37063 26830
rect 37917 26827 37983 26830
rect 30005 26754 30071 26757
rect 33869 26754 33935 26757
rect 34421 26754 34487 26757
rect 30005 26752 34487 26754
rect 30005 26696 30010 26752
rect 30066 26696 33874 26752
rect 33930 26696 34426 26752
rect 34482 26696 34487 26752
rect 30005 26694 34487 26696
rect 30005 26691 30071 26694
rect 33869 26691 33935 26694
rect 34421 26691 34487 26694
rect 4208 26688 4528 26689
rect 0 26618 800 26648
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 2773 26618 2839 26621
rect 0 26616 2839 26618
rect 0 26560 2778 26616
rect 2834 26560 2839 26616
rect 0 26558 2839 26560
rect 0 26528 800 26558
rect 2773 26555 2839 26558
rect 22829 26618 22895 26621
rect 23565 26618 23631 26621
rect 26417 26618 26483 26621
rect 22829 26616 26483 26618
rect 22829 26560 22834 26616
rect 22890 26560 23570 26616
rect 23626 26560 26422 26616
rect 26478 26560 26483 26616
rect 22829 26558 26483 26560
rect 22829 26555 22895 26558
rect 23565 26555 23631 26558
rect 26417 26555 26483 26558
rect 46841 26618 46907 26621
rect 49200 26618 50000 26648
rect 46841 26616 50000 26618
rect 46841 26560 46846 26616
rect 46902 26560 50000 26616
rect 46841 26558 50000 26560
rect 46841 26555 46907 26558
rect 49200 26528 50000 26558
rect 30097 26482 30163 26485
rect 41505 26482 41571 26485
rect 30097 26480 41571 26482
rect 30097 26424 30102 26480
rect 30158 26424 41510 26480
rect 41566 26424 41571 26480
rect 30097 26422 41571 26424
rect 30097 26419 30163 26422
rect 41505 26419 41571 26422
rect 41689 26482 41755 26485
rect 41822 26482 41828 26484
rect 41689 26480 41828 26482
rect 41689 26424 41694 26480
rect 41750 26424 41828 26480
rect 41689 26422 41828 26424
rect 41689 26419 41755 26422
rect 41822 26420 41828 26422
rect 41892 26420 41898 26484
rect 30741 26346 30807 26349
rect 35065 26346 35131 26349
rect 36077 26346 36143 26349
rect 36997 26346 37063 26349
rect 30741 26344 37063 26346
rect 30741 26288 30746 26344
rect 30802 26288 35070 26344
rect 35126 26288 36082 26344
rect 36138 26288 37002 26344
rect 37058 26288 37063 26344
rect 30741 26286 37063 26288
rect 30741 26283 30807 26286
rect 35065 26283 35131 26286
rect 36077 26283 36143 26286
rect 36997 26283 37063 26286
rect 34697 26210 34763 26213
rect 35157 26210 35223 26213
rect 34697 26208 35223 26210
rect 34697 26152 34702 26208
rect 34758 26152 35162 26208
rect 35218 26152 35223 26208
rect 34697 26150 35223 26152
rect 34697 26147 34763 26150
rect 35157 26147 35223 26150
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 0 25938 800 25968
rect 1393 25938 1459 25941
rect 0 25936 1459 25938
rect 0 25880 1398 25936
rect 1454 25880 1459 25936
rect 0 25878 1459 25880
rect 0 25848 800 25878
rect 1393 25875 1459 25878
rect 48129 25938 48195 25941
rect 49200 25938 50000 25968
rect 48129 25936 50000 25938
rect 48129 25880 48134 25936
rect 48190 25880 50000 25936
rect 48129 25878 50000 25880
rect 48129 25875 48195 25878
rect 49200 25848 50000 25878
rect 30097 25802 30163 25805
rect 36997 25802 37063 25805
rect 30097 25800 37063 25802
rect 30097 25744 30102 25800
rect 30158 25744 37002 25800
rect 37058 25744 37063 25800
rect 30097 25742 37063 25744
rect 30097 25739 30163 25742
rect 36997 25739 37063 25742
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 35801 25530 35867 25533
rect 36537 25530 36603 25533
rect 35801 25528 36603 25530
rect 35801 25472 35806 25528
rect 35862 25472 36542 25528
rect 36598 25472 36603 25528
rect 35801 25470 36603 25472
rect 35801 25467 35867 25470
rect 36537 25467 36603 25470
rect 33593 25394 33659 25397
rect 38101 25394 38167 25397
rect 33593 25392 38167 25394
rect 33593 25336 33598 25392
rect 33654 25336 38106 25392
rect 38162 25336 38167 25392
rect 33593 25334 38167 25336
rect 33593 25331 33659 25334
rect 38101 25331 38167 25334
rect 0 25168 800 25288
rect 19793 25258 19859 25261
rect 20110 25258 20116 25260
rect 19793 25256 20116 25258
rect 19793 25200 19798 25256
rect 19854 25200 20116 25256
rect 19793 25198 20116 25200
rect 19793 25195 19859 25198
rect 20110 25196 20116 25198
rect 20180 25196 20186 25260
rect 33133 25258 33199 25261
rect 35893 25258 35959 25261
rect 33133 25256 35959 25258
rect 33133 25200 33138 25256
rect 33194 25200 35898 25256
rect 35954 25200 35959 25256
rect 33133 25198 35959 25200
rect 33133 25195 33199 25198
rect 35893 25195 35959 25198
rect 47853 25258 47919 25261
rect 49200 25258 50000 25288
rect 47853 25256 50000 25258
rect 47853 25200 47858 25256
rect 47914 25200 50000 25256
rect 47853 25198 50000 25200
rect 47853 25195 47919 25198
rect 49200 25168 50000 25198
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 19701 24714 19767 24717
rect 20713 24714 20779 24717
rect 19701 24712 20779 24714
rect 19701 24656 19706 24712
rect 19762 24656 20718 24712
rect 20774 24656 20779 24712
rect 19701 24654 20779 24656
rect 19701 24651 19767 24654
rect 20713 24651 20779 24654
rect 27797 24714 27863 24717
rect 35709 24714 35775 24717
rect 27797 24712 35775 24714
rect 27797 24656 27802 24712
rect 27858 24656 35714 24712
rect 35770 24656 35775 24712
rect 27797 24654 35775 24656
rect 27797 24651 27863 24654
rect 35709 24651 35775 24654
rect 0 24488 800 24608
rect 28993 24578 29059 24581
rect 28950 24576 29059 24578
rect 28950 24520 28998 24576
rect 29054 24520 29059 24576
rect 28950 24515 29059 24520
rect 39389 24578 39455 24581
rect 42517 24578 42583 24581
rect 39389 24576 42583 24578
rect 39389 24520 39394 24576
rect 39450 24520 42522 24576
rect 42578 24520 42583 24576
rect 39389 24518 42583 24520
rect 39389 24515 39455 24518
rect 42517 24515 42583 24518
rect 48129 24578 48195 24581
rect 49200 24578 50000 24608
rect 48129 24576 50000 24578
rect 48129 24520 48134 24576
rect 48190 24520 50000 24576
rect 48129 24518 50000 24520
rect 48129 24515 48195 24518
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 24853 24442 24919 24445
rect 27429 24442 27495 24445
rect 24853 24440 27495 24442
rect 24853 24384 24858 24440
rect 24914 24384 27434 24440
rect 27490 24384 27495 24440
rect 24853 24382 27495 24384
rect 24853 24379 24919 24382
rect 27429 24379 27495 24382
rect 28950 24309 29010 24515
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 49200 24488 50000 24518
rect 34928 24447 35248 24448
rect 40861 24442 40927 24445
rect 43437 24442 43503 24445
rect 40861 24440 43503 24442
rect 40861 24384 40866 24440
rect 40922 24384 43442 24440
rect 43498 24384 43503 24440
rect 40861 24382 43503 24384
rect 40861 24379 40927 24382
rect 43437 24379 43503 24382
rect 28950 24304 29059 24309
rect 28950 24248 28998 24304
rect 29054 24248 29059 24304
rect 28950 24246 29059 24248
rect 28993 24243 29059 24246
rect 42149 24306 42215 24309
rect 43345 24306 43411 24309
rect 42149 24304 43411 24306
rect 42149 24248 42154 24304
rect 42210 24248 43350 24304
rect 43406 24248 43411 24304
rect 42149 24246 43411 24248
rect 42149 24243 42215 24246
rect 43345 24243 43411 24246
rect 28533 24170 28599 24173
rect 28901 24170 28967 24173
rect 28533 24168 28967 24170
rect 28533 24112 28538 24168
rect 28594 24112 28906 24168
rect 28962 24112 28967 24168
rect 28533 24110 28967 24112
rect 28533 24107 28599 24110
rect 28901 24107 28967 24110
rect 29126 24108 29132 24172
rect 29196 24170 29202 24172
rect 29269 24170 29335 24173
rect 29196 24168 29335 24170
rect 29196 24112 29274 24168
rect 29330 24112 29335 24168
rect 29196 24110 29335 24112
rect 29196 24108 29202 24110
rect 29269 24107 29335 24110
rect 39849 24170 39915 24173
rect 41321 24170 41387 24173
rect 42241 24170 42307 24173
rect 43161 24170 43227 24173
rect 39849 24168 43227 24170
rect 39849 24112 39854 24168
rect 39910 24112 41326 24168
rect 41382 24112 42246 24168
rect 42302 24112 43166 24168
rect 43222 24112 43227 24168
rect 39849 24110 43227 24112
rect 39849 24107 39915 24110
rect 41321 24107 41387 24110
rect 42241 24107 42307 24110
rect 43161 24107 43227 24110
rect 28533 24034 28599 24037
rect 29177 24036 29243 24037
rect 28942 24034 28948 24036
rect 28533 24032 28948 24034
rect 28533 23976 28538 24032
rect 28594 23976 28948 24032
rect 28533 23974 28948 23976
rect 28533 23971 28599 23974
rect 28942 23972 28948 23974
rect 29012 23972 29018 24036
rect 29126 24034 29132 24036
rect 29086 23974 29132 24034
rect 29196 24032 29243 24036
rect 29238 23976 29243 24032
rect 29126 23972 29132 23974
rect 29196 23972 29243 23976
rect 29177 23971 29243 23972
rect 29545 24034 29611 24037
rect 38561 24034 38627 24037
rect 29545 24032 38627 24034
rect 29545 23976 29550 24032
rect 29606 23976 38566 24032
rect 38622 23976 38627 24032
rect 29545 23974 38627 23976
rect 29545 23971 29611 23974
rect 38561 23971 38627 23974
rect 19568 23968 19888 23969
rect 0 23898 800 23928
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 1393 23898 1459 23901
rect 0 23896 1459 23898
rect 0 23840 1398 23896
rect 1454 23840 1459 23896
rect 0 23838 1459 23840
rect 0 23808 800 23838
rect 1393 23835 1459 23838
rect 20897 23898 20963 23901
rect 27797 23898 27863 23901
rect 20897 23896 27863 23898
rect 20897 23840 20902 23896
rect 20958 23840 27802 23896
rect 27858 23840 27863 23896
rect 20897 23838 27863 23840
rect 20897 23835 20963 23838
rect 27797 23835 27863 23838
rect 28993 23898 29059 23901
rect 34513 23898 34579 23901
rect 28993 23896 34579 23898
rect 28993 23840 28998 23896
rect 29054 23840 34518 23896
rect 34574 23840 34579 23896
rect 28993 23838 34579 23840
rect 28993 23835 29059 23838
rect 34513 23835 34579 23838
rect 39665 23898 39731 23901
rect 40861 23898 40927 23901
rect 39665 23896 40927 23898
rect 39665 23840 39670 23896
rect 39726 23840 40866 23896
rect 40922 23840 40927 23896
rect 39665 23838 40927 23840
rect 39665 23835 39731 23838
rect 40861 23835 40927 23838
rect 47945 23898 48011 23901
rect 49200 23898 50000 23928
rect 47945 23896 50000 23898
rect 47945 23840 47950 23896
rect 48006 23840 50000 23896
rect 47945 23838 50000 23840
rect 47945 23835 48011 23838
rect 49200 23808 50000 23838
rect 24669 23762 24735 23765
rect 26601 23762 26667 23765
rect 24669 23760 26667 23762
rect 24669 23704 24674 23760
rect 24730 23704 26606 23760
rect 26662 23704 26667 23760
rect 24669 23702 26667 23704
rect 24669 23699 24735 23702
rect 26601 23699 26667 23702
rect 27521 23762 27587 23765
rect 35341 23762 35407 23765
rect 27521 23760 35407 23762
rect 27521 23704 27526 23760
rect 27582 23704 35346 23760
rect 35402 23704 35407 23760
rect 27521 23702 35407 23704
rect 27521 23699 27587 23702
rect 35341 23699 35407 23702
rect 19885 23626 19951 23629
rect 25773 23626 25839 23629
rect 19885 23624 25839 23626
rect 19885 23568 19890 23624
rect 19946 23568 25778 23624
rect 25834 23568 25839 23624
rect 19885 23566 25839 23568
rect 19885 23563 19951 23566
rect 25773 23563 25839 23566
rect 26049 23626 26115 23629
rect 26417 23626 26483 23629
rect 28809 23626 28875 23629
rect 26049 23624 28875 23626
rect 26049 23568 26054 23624
rect 26110 23568 26422 23624
rect 26478 23568 28814 23624
rect 28870 23568 28875 23624
rect 26049 23566 28875 23568
rect 26049 23563 26115 23566
rect 26417 23563 26483 23566
rect 28809 23563 28875 23566
rect 40401 23626 40467 23629
rect 41505 23626 41571 23629
rect 40401 23624 41571 23626
rect 40401 23568 40406 23624
rect 40462 23568 41510 23624
rect 41566 23568 41571 23624
rect 40401 23566 41571 23568
rect 40401 23563 40467 23566
rect 41505 23563 41571 23566
rect 42793 23626 42859 23629
rect 43897 23626 43963 23629
rect 42793 23624 43963 23626
rect 42793 23568 42798 23624
rect 42854 23568 43902 23624
rect 43958 23568 43963 23624
rect 42793 23566 43963 23568
rect 42793 23563 42859 23566
rect 43897 23563 43963 23566
rect 19885 23490 19951 23493
rect 20110 23490 20116 23492
rect 19885 23488 20116 23490
rect 19885 23432 19890 23488
rect 19946 23432 20116 23488
rect 19885 23430 20116 23432
rect 19885 23427 19951 23430
rect 20110 23428 20116 23430
rect 20180 23428 20186 23492
rect 27153 23490 27219 23493
rect 30097 23490 30163 23493
rect 27153 23488 30163 23490
rect 27153 23432 27158 23488
rect 27214 23432 30102 23488
rect 30158 23432 30163 23488
rect 27153 23430 30163 23432
rect 27153 23427 27219 23430
rect 30097 23427 30163 23430
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 28165 23354 28231 23357
rect 28993 23354 29059 23357
rect 29177 23356 29243 23357
rect 28165 23352 29059 23354
rect 28165 23296 28170 23352
rect 28226 23296 28998 23352
rect 29054 23296 29059 23352
rect 28165 23294 29059 23296
rect 28165 23291 28231 23294
rect 28993 23291 29059 23294
rect 29126 23292 29132 23356
rect 29196 23354 29243 23356
rect 29196 23352 29288 23354
rect 29238 23296 29288 23352
rect 29196 23294 29288 23296
rect 29196 23292 29243 23294
rect 29177 23291 29243 23292
rect 0 23218 800 23248
rect 2773 23218 2839 23221
rect 0 23216 2839 23218
rect 0 23160 2778 23216
rect 2834 23160 2839 23216
rect 0 23158 2839 23160
rect 0 23128 800 23158
rect 2773 23155 2839 23158
rect 28717 23218 28783 23221
rect 29269 23218 29335 23221
rect 28717 23216 29335 23218
rect 28717 23160 28722 23216
rect 28778 23160 29274 23216
rect 29330 23160 29335 23216
rect 28717 23158 29335 23160
rect 28717 23155 28783 23158
rect 29269 23155 29335 23158
rect 49200 23128 50000 23248
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 40309 22810 40375 22813
rect 43989 22810 44055 22813
rect 40309 22808 44055 22810
rect 40309 22752 40314 22808
rect 40370 22752 43994 22808
rect 44050 22752 44055 22808
rect 40309 22750 44055 22752
rect 40309 22747 40375 22750
rect 43989 22747 44055 22750
rect 0 22538 800 22568
rect 1853 22538 1919 22541
rect 0 22536 1919 22538
rect 0 22480 1858 22536
rect 1914 22480 1919 22536
rect 0 22478 1919 22480
rect 0 22448 800 22478
rect 1853 22475 1919 22478
rect 19885 22538 19951 22541
rect 20110 22538 20116 22540
rect 19885 22536 20116 22538
rect 19885 22480 19890 22536
rect 19946 22480 20116 22536
rect 19885 22478 20116 22480
rect 19885 22475 19951 22478
rect 20110 22476 20116 22478
rect 20180 22476 20186 22540
rect 47945 22538 48011 22541
rect 49200 22538 50000 22568
rect 47945 22536 50000 22538
rect 47945 22480 47950 22536
rect 48006 22480 50000 22536
rect 47945 22478 50000 22480
rect 47945 22475 48011 22478
rect 49200 22448 50000 22478
rect 24853 22404 24919 22405
rect 24853 22400 24900 22404
rect 24964 22402 24970 22404
rect 24853 22344 24858 22400
rect 24853 22340 24900 22344
rect 24964 22342 25010 22402
rect 24964 22340 24970 22342
rect 24853 22339 24919 22340
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 20529 22096 20595 22099
rect 20486 22094 20595 22096
rect 20486 22038 20534 22094
rect 20590 22038 20595 22094
rect 20486 22033 20595 22038
rect 20069 21994 20135 21997
rect 20486 21994 20546 22033
rect 20069 21992 20546 21994
rect 20069 21936 20074 21992
rect 20130 21936 20546 21992
rect 20069 21934 20546 21936
rect 32581 21994 32647 21997
rect 38469 21994 38535 21997
rect 32581 21992 38535 21994
rect 32581 21936 32586 21992
rect 32642 21936 38474 21992
rect 38530 21936 38535 21992
rect 32581 21934 38535 21936
rect 20069 21931 20135 21934
rect 32581 21931 32647 21934
rect 38469 21931 38535 21934
rect 0 21858 800 21888
rect 2865 21858 2931 21861
rect 0 21856 2931 21858
rect 0 21800 2870 21856
rect 2926 21800 2931 21856
rect 0 21798 2931 21800
rect 0 21768 800 21798
rect 2865 21795 2931 21798
rect 21633 21858 21699 21861
rect 28257 21858 28323 21861
rect 21633 21856 28323 21858
rect 21633 21800 21638 21856
rect 21694 21800 28262 21856
rect 28318 21800 28323 21856
rect 21633 21798 28323 21800
rect 21633 21795 21699 21798
rect 28257 21795 28323 21798
rect 47945 21858 48011 21861
rect 49200 21858 50000 21888
rect 47945 21856 50000 21858
rect 47945 21800 47950 21856
rect 48006 21800 50000 21856
rect 47945 21798 50000 21800
rect 47945 21795 48011 21798
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 49200 21768 50000 21798
rect 19568 21727 19888 21728
rect 28257 21722 28323 21725
rect 28533 21722 28599 21725
rect 28257 21720 28599 21722
rect 28257 21664 28262 21720
rect 28318 21664 28538 21720
rect 28594 21664 28599 21720
rect 28257 21662 28599 21664
rect 28257 21659 28323 21662
rect 28533 21659 28599 21662
rect 4208 21248 4528 21249
rect 0 21178 800 21208
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 3417 21178 3483 21181
rect 0 21176 3483 21178
rect 0 21120 3422 21176
rect 3478 21120 3483 21176
rect 0 21118 3483 21120
rect 0 21088 800 21118
rect 3417 21115 3483 21118
rect 49200 21088 50000 21208
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 0 20408 800 20528
rect 22553 20498 22619 20501
rect 24301 20498 24367 20501
rect 22553 20496 24367 20498
rect 22553 20440 22558 20496
rect 22614 20440 24306 20496
rect 24362 20440 24367 20496
rect 22553 20438 24367 20440
rect 22553 20435 22619 20438
rect 24301 20435 24367 20438
rect 49200 20408 50000 20528
rect 22553 20362 22619 20365
rect 25313 20362 25379 20365
rect 22553 20360 25379 20362
rect 22553 20304 22558 20360
rect 22614 20304 25318 20360
rect 25374 20304 25379 20360
rect 22553 20302 25379 20304
rect 22553 20299 22619 20302
rect 25313 20299 25379 20302
rect 21909 20226 21975 20229
rect 24485 20226 24551 20229
rect 21909 20224 24551 20226
rect 21909 20168 21914 20224
rect 21970 20168 24490 20224
rect 24546 20168 24551 20224
rect 21909 20166 24551 20168
rect 21909 20163 21975 20166
rect 24485 20163 24551 20166
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 21909 20090 21975 20093
rect 28717 20090 28783 20093
rect 21909 20088 28783 20090
rect 21909 20032 21914 20088
rect 21970 20032 28722 20088
rect 28778 20032 28783 20088
rect 21909 20030 28783 20032
rect 21909 20027 21975 20030
rect 28717 20027 28783 20030
rect 22553 19954 22619 19957
rect 23565 19954 23631 19957
rect 22553 19952 23631 19954
rect 22553 19896 22558 19952
rect 22614 19896 23570 19952
rect 23626 19896 23631 19952
rect 22553 19894 23631 19896
rect 22553 19891 22619 19894
rect 23565 19891 23631 19894
rect 0 19818 800 19848
rect 2773 19818 2839 19821
rect 0 19816 2839 19818
rect 0 19760 2778 19816
rect 2834 19760 2839 19816
rect 0 19758 2839 19760
rect 0 19728 800 19758
rect 2773 19755 2839 19758
rect 21817 19818 21883 19821
rect 22185 19818 22251 19821
rect 21817 19816 22251 19818
rect 21817 19760 21822 19816
rect 21878 19760 22190 19816
rect 22246 19760 22251 19816
rect 21817 19758 22251 19760
rect 21817 19755 21883 19758
rect 22185 19755 22251 19758
rect 22829 19818 22895 19821
rect 38009 19818 38075 19821
rect 38561 19818 38627 19821
rect 22829 19816 22938 19818
rect 22829 19760 22834 19816
rect 22890 19760 22938 19816
rect 22829 19755 22938 19760
rect 38009 19816 38627 19818
rect 38009 19760 38014 19816
rect 38070 19760 38566 19816
rect 38622 19760 38627 19816
rect 38009 19758 38627 19760
rect 38009 19755 38075 19758
rect 38561 19755 38627 19758
rect 48129 19818 48195 19821
rect 49200 19818 50000 19848
rect 48129 19816 50000 19818
rect 48129 19760 48134 19816
rect 48190 19760 50000 19816
rect 48129 19758 50000 19760
rect 48129 19755 48195 19758
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 22878 19413 22938 19755
rect 49200 19728 50000 19758
rect 25773 19546 25839 19549
rect 27061 19546 27127 19549
rect 25773 19544 27127 19546
rect 25773 19488 25778 19544
rect 25834 19488 27066 19544
rect 27122 19488 27127 19544
rect 25773 19486 27127 19488
rect 25773 19483 25839 19486
rect 27061 19483 27127 19486
rect 17953 19410 18019 19413
rect 18781 19410 18847 19413
rect 17953 19408 18847 19410
rect 17953 19352 17958 19408
rect 18014 19352 18786 19408
rect 18842 19352 18847 19408
rect 17953 19350 18847 19352
rect 17953 19347 18019 19350
rect 18781 19347 18847 19350
rect 19885 19410 19951 19413
rect 20110 19410 20116 19412
rect 19885 19408 20116 19410
rect 19885 19352 19890 19408
rect 19946 19352 20116 19408
rect 19885 19350 20116 19352
rect 19885 19347 19951 19350
rect 20110 19348 20116 19350
rect 20180 19348 20186 19412
rect 22878 19408 22987 19413
rect 22878 19352 22926 19408
rect 22982 19352 22987 19408
rect 22878 19350 22987 19352
rect 22921 19347 22987 19350
rect 26969 19410 27035 19413
rect 27705 19410 27771 19413
rect 26969 19408 27771 19410
rect 26969 19352 26974 19408
rect 27030 19352 27710 19408
rect 27766 19352 27771 19408
rect 26969 19350 27771 19352
rect 26969 19347 27035 19350
rect 27705 19347 27771 19350
rect 0 19138 800 19168
rect 2773 19138 2839 19141
rect 0 19136 2839 19138
rect 0 19080 2778 19136
rect 2834 19080 2839 19136
rect 0 19078 2839 19080
rect 0 19048 800 19078
rect 2773 19075 2839 19078
rect 47945 19138 48011 19141
rect 49200 19138 50000 19168
rect 47945 19136 50000 19138
rect 47945 19080 47950 19136
rect 48006 19080 50000 19136
rect 47945 19078 50000 19080
rect 47945 19075 48011 19078
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 49200 19048 50000 19078
rect 34928 19007 35248 19008
rect 19568 18528 19888 18529
rect 0 18458 800 18488
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 3417 18458 3483 18461
rect 0 18456 3483 18458
rect 0 18400 3422 18456
rect 3478 18400 3483 18456
rect 0 18398 3483 18400
rect 0 18368 800 18398
rect 3417 18395 3483 18398
rect 49200 18368 50000 18488
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 0 17778 800 17808
rect 2773 17778 2839 17781
rect 0 17776 2839 17778
rect 0 17720 2778 17776
rect 2834 17720 2839 17776
rect 0 17718 2839 17720
rect 0 17688 800 17718
rect 2773 17715 2839 17718
rect 48129 17778 48195 17781
rect 49200 17778 50000 17808
rect 48129 17776 50000 17778
rect 48129 17720 48134 17776
rect 48190 17720 50000 17776
rect 48129 17718 50000 17720
rect 48129 17715 48195 17718
rect 49200 17688 50000 17718
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 0 17098 800 17128
rect 1853 17098 1919 17101
rect 0 17096 1919 17098
rect 0 17040 1858 17096
rect 1914 17040 1919 17096
rect 0 17038 1919 17040
rect 0 17008 800 17038
rect 1853 17035 1919 17038
rect 46841 17098 46907 17101
rect 49200 17098 50000 17128
rect 46841 17096 50000 17098
rect 46841 17040 46846 17096
rect 46902 17040 50000 17096
rect 46841 17038 50000 17040
rect 46841 17035 46907 17038
rect 49200 17008 50000 17038
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 0 16418 800 16448
rect 1853 16418 1919 16421
rect 0 16416 1919 16418
rect 0 16360 1858 16416
rect 1914 16360 1919 16416
rect 0 16358 1919 16360
rect 0 16328 800 16358
rect 1853 16355 1919 16358
rect 48129 16418 48195 16421
rect 49200 16418 50000 16448
rect 48129 16416 50000 16418
rect 48129 16360 48134 16416
rect 48190 16360 50000 16416
rect 48129 16358 50000 16360
rect 48129 16355 48195 16358
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 49200 16328 50000 16358
rect 19568 16287 19888 16288
rect 19885 16010 19951 16013
rect 20110 16010 20116 16012
rect 19885 16008 20116 16010
rect 19885 15952 19890 16008
rect 19946 15952 20116 16008
rect 19885 15950 20116 15952
rect 19885 15947 19951 15950
rect 20110 15948 20116 15950
rect 20180 15948 20186 16012
rect 4208 15808 4528 15809
rect 0 15648 800 15768
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 49200 15648 50000 15768
rect 26417 15330 26483 15333
rect 28717 15330 28783 15333
rect 26417 15328 28783 15330
rect 26417 15272 26422 15328
rect 26478 15272 28722 15328
rect 28778 15272 28783 15328
rect 26417 15270 28783 15272
rect 26417 15267 26483 15270
rect 28717 15267 28783 15270
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 0 14968 800 15088
rect 46841 15058 46907 15061
rect 49200 15058 50000 15088
rect 46841 15056 50000 15058
rect 46841 15000 46846 15056
rect 46902 15000 50000 15056
rect 46841 14998 50000 15000
rect 46841 14995 46907 14998
rect 49200 14968 50000 14998
rect 21449 14922 21515 14925
rect 27521 14922 27587 14925
rect 21449 14920 27587 14922
rect 21449 14864 21454 14920
rect 21510 14864 27526 14920
rect 27582 14864 27587 14920
rect 21449 14862 27587 14864
rect 21449 14859 21515 14862
rect 27521 14859 27587 14862
rect 20069 14786 20135 14789
rect 20294 14786 20300 14788
rect 20069 14784 20300 14786
rect 20069 14728 20074 14784
rect 20130 14728 20300 14784
rect 20069 14726 20300 14728
rect 20069 14723 20135 14726
rect 20294 14724 20300 14726
rect 20364 14724 20370 14788
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 19425 14516 19491 14517
rect 19374 14452 19380 14516
rect 19444 14514 19491 14516
rect 34881 14514 34947 14517
rect 37457 14514 37523 14517
rect 19444 14512 19536 14514
rect 19486 14456 19536 14512
rect 19444 14454 19536 14456
rect 34881 14512 37523 14514
rect 34881 14456 34886 14512
rect 34942 14456 37462 14512
rect 37518 14456 37523 14512
rect 34881 14454 37523 14456
rect 19444 14452 19491 14454
rect 19425 14451 19491 14452
rect 34881 14451 34947 14454
rect 37457 14451 37523 14454
rect 0 14288 800 14408
rect 48129 14378 48195 14381
rect 49200 14378 50000 14408
rect 48129 14376 50000 14378
rect 48129 14320 48134 14376
rect 48190 14320 50000 14376
rect 48129 14318 50000 14320
rect 48129 14315 48195 14318
rect 49200 14288 50000 14318
rect 34513 14242 34579 14245
rect 38285 14242 38351 14245
rect 34513 14240 38351 14242
rect 34513 14184 34518 14240
rect 34574 14184 38290 14240
rect 38346 14184 38351 14240
rect 34513 14182 38351 14184
rect 34513 14179 34579 14182
rect 38285 14179 38351 14182
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 0 13698 800 13728
rect 2773 13698 2839 13701
rect 0 13696 2839 13698
rect 0 13640 2778 13696
rect 2834 13640 2839 13696
rect 0 13638 2839 13640
rect 0 13608 800 13638
rect 2773 13635 2839 13638
rect 41822 13636 41828 13700
rect 41892 13698 41898 13700
rect 47025 13698 47091 13701
rect 41892 13696 47091 13698
rect 41892 13640 47030 13696
rect 47086 13640 47091 13696
rect 41892 13638 47091 13640
rect 41892 13636 41898 13638
rect 47025 13635 47091 13638
rect 47853 13698 47919 13701
rect 49200 13698 50000 13728
rect 47853 13696 50000 13698
rect 47853 13640 47858 13696
rect 47914 13640 50000 13696
rect 47853 13638 50000 13640
rect 47853 13635 47919 13638
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 49200 13608 50000 13638
rect 34928 13567 35248 13568
rect 19568 13088 19888 13089
rect 0 13018 800 13048
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 3049 13018 3115 13021
rect 0 13016 3115 13018
rect 0 12960 3054 13016
rect 3110 12960 3115 13016
rect 0 12958 3115 12960
rect 0 12928 800 12958
rect 3049 12955 3115 12958
rect 46565 13018 46631 13021
rect 49200 13018 50000 13048
rect 46565 13016 50000 13018
rect 46565 12960 46570 13016
rect 46626 12960 50000 13016
rect 46565 12958 50000 12960
rect 46565 12955 46631 12958
rect 49200 12928 50000 12958
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 0 12338 800 12368
rect 1393 12338 1459 12341
rect 0 12336 1459 12338
rect 0 12280 1398 12336
rect 1454 12280 1459 12336
rect 0 12278 1459 12280
rect 0 12248 800 12278
rect 1393 12275 1459 12278
rect 46841 12338 46907 12341
rect 49200 12338 50000 12368
rect 46841 12336 50000 12338
rect 46841 12280 46846 12336
rect 46902 12280 50000 12336
rect 46841 12278 50000 12280
rect 46841 12275 46907 12278
rect 49200 12248 50000 12278
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 0 11568 800 11688
rect 49200 11568 50000 11688
rect 19374 11460 19380 11524
rect 19444 11522 19450 11524
rect 20345 11522 20411 11525
rect 19444 11520 20411 11522
rect 19444 11464 20350 11520
rect 20406 11464 20411 11520
rect 19444 11462 20411 11464
rect 19444 11460 19450 11462
rect 20345 11459 20411 11462
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 0 10978 800 11008
rect 1393 10978 1459 10981
rect 0 10976 1459 10978
rect 0 10920 1398 10976
rect 1454 10920 1459 10976
rect 0 10918 1459 10920
rect 0 10888 800 10918
rect 1393 10915 1459 10918
rect 48129 10978 48195 10981
rect 49200 10978 50000 11008
rect 48129 10976 50000 10978
rect 48129 10920 48134 10976
rect 48190 10920 50000 10976
rect 48129 10918 50000 10920
rect 48129 10915 48195 10918
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 49200 10888 50000 10918
rect 19568 10847 19888 10848
rect 4208 10368 4528 10369
rect 0 10298 800 10328
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 2773 10298 2839 10301
rect 0 10296 2839 10298
rect 0 10240 2778 10296
rect 2834 10240 2839 10296
rect 0 10238 2839 10240
rect 0 10208 800 10238
rect 2773 10235 2839 10238
rect 24209 10298 24275 10301
rect 26233 10298 26299 10301
rect 24209 10296 26299 10298
rect 24209 10240 24214 10296
rect 24270 10240 26238 10296
rect 26294 10240 26299 10296
rect 24209 10238 26299 10240
rect 24209 10235 24275 10238
rect 26233 10235 26299 10238
rect 47853 10298 47919 10301
rect 49200 10298 50000 10328
rect 47853 10296 50000 10298
rect 47853 10240 47858 10296
rect 47914 10240 50000 10296
rect 47853 10238 50000 10240
rect 47853 10235 47919 10238
rect 49200 10208 50000 10238
rect 19517 10026 19583 10029
rect 19382 10024 19583 10026
rect 19382 9968 19522 10024
rect 19578 9968 19583 10024
rect 19382 9966 19583 9968
rect 19382 9690 19442 9966
rect 19517 9963 19583 9966
rect 19701 10026 19767 10029
rect 19701 10024 20040 10026
rect 19701 9968 19706 10024
rect 19762 9968 20040 10024
rect 19701 9966 20040 9968
rect 19701 9963 19767 9966
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 19980 9693 20040 9966
rect 20294 9754 20300 9756
rect 20118 9694 20300 9754
rect 19793 9690 19859 9693
rect 19382 9688 19859 9690
rect 0 9618 800 9648
rect 19382 9632 19798 9688
rect 19854 9632 19859 9688
rect 19382 9630 19859 9632
rect 19793 9627 19859 9630
rect 19977 9688 20043 9693
rect 19977 9632 19982 9688
rect 20038 9632 20043 9688
rect 19977 9627 20043 9632
rect 2773 9618 2839 9621
rect 0 9616 2839 9618
rect 0 9560 2778 9616
rect 2834 9560 2839 9616
rect 0 9558 2839 9560
rect 20118 9618 20178 9694
rect 20294 9692 20300 9694
rect 20364 9692 20370 9756
rect 25037 9618 25103 9621
rect 27521 9618 27587 9621
rect 20118 9558 20316 9618
rect 0 9528 800 9558
rect 2773 9555 2839 9558
rect 20256 9485 20316 9558
rect 25037 9616 27587 9618
rect 25037 9560 25042 9616
rect 25098 9560 27526 9616
rect 27582 9560 27587 9616
rect 25037 9558 27587 9560
rect 25037 9555 25103 9558
rect 27521 9555 27587 9558
rect 46841 9618 46907 9621
rect 49200 9618 50000 9648
rect 46841 9616 50000 9618
rect 46841 9560 46846 9616
rect 46902 9560 50000 9616
rect 46841 9558 50000 9560
rect 46841 9555 46907 9558
rect 49200 9528 50000 9558
rect 20253 9480 20319 9485
rect 20253 9424 20258 9480
rect 20314 9424 20319 9480
rect 20253 9419 20319 9424
rect 24577 9482 24643 9485
rect 25221 9482 25287 9485
rect 24577 9480 25287 9482
rect 24577 9424 24582 9480
rect 24638 9424 25226 9480
rect 25282 9424 25287 9480
rect 24577 9422 25287 9424
rect 24577 9419 24643 9422
rect 25221 9419 25287 9422
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 0 8938 800 8968
rect 3141 8938 3207 8941
rect 0 8936 3207 8938
rect 0 8880 3146 8936
rect 3202 8880 3207 8936
rect 0 8878 3207 8880
rect 0 8848 800 8878
rect 3141 8875 3207 8878
rect 22185 8938 22251 8941
rect 22645 8938 22711 8941
rect 22185 8936 22711 8938
rect 22185 8880 22190 8936
rect 22246 8880 22650 8936
rect 22706 8880 22711 8936
rect 22185 8878 22711 8880
rect 22185 8875 22251 8878
rect 22645 8875 22711 8878
rect 23749 8938 23815 8941
rect 25681 8938 25747 8941
rect 23749 8936 25747 8938
rect 23749 8880 23754 8936
rect 23810 8880 25686 8936
rect 25742 8880 25747 8936
rect 23749 8878 25747 8880
rect 23749 8875 23815 8878
rect 25681 8875 25747 8878
rect 47761 8938 47827 8941
rect 49200 8938 50000 8968
rect 47761 8936 50000 8938
rect 47761 8880 47766 8936
rect 47822 8880 50000 8936
rect 47761 8878 50000 8880
rect 47761 8875 47827 8878
rect 49200 8848 50000 8878
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 24393 8530 24459 8533
rect 25037 8530 25103 8533
rect 25773 8530 25839 8533
rect 26049 8530 26115 8533
rect 24393 8528 26115 8530
rect 24393 8472 24398 8528
rect 24454 8472 25042 8528
rect 25098 8472 25778 8528
rect 25834 8472 26054 8528
rect 26110 8472 26115 8528
rect 24393 8470 26115 8472
rect 24393 8467 24459 8470
rect 25037 8467 25103 8470
rect 25773 8467 25839 8470
rect 26049 8467 26115 8470
rect 25129 8394 25195 8397
rect 27245 8394 27311 8397
rect 25129 8392 27311 8394
rect 25129 8336 25134 8392
rect 25190 8336 27250 8392
rect 27306 8336 27311 8392
rect 25129 8334 27311 8336
rect 25129 8331 25195 8334
rect 27245 8331 27311 8334
rect 0 8258 800 8288
rect 1853 8258 1919 8261
rect 0 8256 1919 8258
rect 0 8200 1858 8256
rect 1914 8200 1919 8256
rect 0 8198 1919 8200
rect 0 8168 800 8198
rect 1853 8195 1919 8198
rect 47853 8258 47919 8261
rect 49200 8258 50000 8288
rect 47853 8256 50000 8258
rect 47853 8200 47858 8256
rect 47914 8200 50000 8256
rect 47853 8198 50000 8200
rect 47853 8195 47919 8198
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 49200 8168 50000 8198
rect 34928 8127 35248 8128
rect 20437 7714 20503 7717
rect 20437 7712 20546 7714
rect 20437 7656 20442 7712
rect 20498 7656 20546 7712
rect 20437 7651 20546 7656
rect 19568 7648 19888 7649
rect 0 7578 800 7608
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 1853 7578 1919 7581
rect 0 7576 1919 7578
rect 0 7520 1858 7576
rect 1914 7520 1919 7576
rect 0 7518 1919 7520
rect 0 7488 800 7518
rect 1853 7515 1919 7518
rect 20486 7309 20546 7651
rect 48129 7578 48195 7581
rect 49200 7578 50000 7608
rect 48129 7576 50000 7578
rect 48129 7520 48134 7576
rect 48190 7520 50000 7576
rect 48129 7518 50000 7520
rect 48129 7515 48195 7518
rect 49200 7488 50000 7518
rect 19977 7306 20043 7309
rect 20110 7306 20116 7308
rect 19977 7304 20116 7306
rect 19977 7248 19982 7304
rect 20038 7248 20116 7304
rect 19977 7246 20116 7248
rect 19977 7243 20043 7246
rect 20110 7244 20116 7246
rect 20180 7244 20186 7308
rect 20437 7304 20546 7309
rect 20437 7248 20442 7304
rect 20498 7248 20546 7304
rect 20437 7246 20546 7248
rect 20437 7243 20503 7246
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 0 6898 800 6928
rect 2773 6898 2839 6901
rect 0 6896 2839 6898
rect 0 6840 2778 6896
rect 2834 6840 2839 6896
rect 0 6838 2839 6840
rect 0 6808 800 6838
rect 2773 6835 2839 6838
rect 46013 6898 46079 6901
rect 49200 6898 50000 6928
rect 46013 6896 50000 6898
rect 46013 6840 46018 6896
rect 46074 6840 50000 6896
rect 46013 6838 50000 6840
rect 46013 6835 46079 6838
rect 49200 6808 50000 6838
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 0 6218 800 6248
rect 3417 6218 3483 6221
rect 0 6216 3483 6218
rect 0 6160 3422 6216
rect 3478 6160 3483 6216
rect 0 6158 3483 6160
rect 0 6128 800 6158
rect 3417 6155 3483 6158
rect 46841 6218 46907 6221
rect 49200 6218 50000 6248
rect 46841 6216 50000 6218
rect 46841 6160 46846 6216
rect 46902 6160 50000 6216
rect 46841 6158 50000 6160
rect 46841 6155 46907 6158
rect 49200 6128 50000 6158
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 0 5538 800 5568
rect 2773 5538 2839 5541
rect 0 5536 2839 5538
rect 0 5480 2778 5536
rect 2834 5480 2839 5536
rect 0 5478 2839 5480
rect 0 5448 800 5478
rect 2773 5475 2839 5478
rect 47853 5538 47919 5541
rect 49200 5538 50000 5568
rect 47853 5536 50000 5538
rect 47853 5480 47858 5536
rect 47914 5480 50000 5536
rect 47853 5478 50000 5480
rect 47853 5475 47919 5478
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 49200 5448 50000 5478
rect 19568 5407 19888 5408
rect 4208 4928 4528 4929
rect 0 4858 800 4888
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 2773 4858 2839 4861
rect 0 4856 2839 4858
rect 0 4800 2778 4856
rect 2834 4800 2839 4856
rect 0 4798 2839 4800
rect 0 4768 800 4798
rect 2773 4795 2839 4798
rect 48129 4858 48195 4861
rect 49200 4858 50000 4888
rect 48129 4856 50000 4858
rect 48129 4800 48134 4856
rect 48190 4800 50000 4856
rect 48129 4798 50000 4800
rect 48129 4795 48195 4798
rect 49200 4768 50000 4798
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 0 4178 800 4208
rect 3417 4178 3483 4181
rect 0 4176 3483 4178
rect 0 4120 3422 4176
rect 3478 4120 3483 4176
rect 0 4118 3483 4120
rect 0 4088 800 4118
rect 3417 4115 3483 4118
rect 46105 4178 46171 4181
rect 49200 4178 50000 4208
rect 46105 4176 50000 4178
rect 46105 4120 46110 4176
rect 46166 4120 50000 4176
rect 46105 4118 50000 4120
rect 46105 4115 46171 4118
rect 49200 4088 50000 4118
rect 30281 4042 30347 4045
rect 36445 4042 36511 4045
rect 30281 4040 36511 4042
rect 30281 3984 30286 4040
rect 30342 3984 36450 4040
rect 36506 3984 36511 4040
rect 30281 3982 36511 3984
rect 30281 3979 30347 3982
rect 36445 3979 36511 3982
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 0 3498 800 3528
rect 1853 3498 1919 3501
rect 0 3496 1919 3498
rect 0 3440 1858 3496
rect 1914 3440 1919 3496
rect 0 3438 1919 3440
rect 0 3408 800 3438
rect 1853 3435 1919 3438
rect 29453 3498 29519 3501
rect 32305 3498 32371 3501
rect 29453 3496 32371 3498
rect 29453 3440 29458 3496
rect 29514 3440 32310 3496
rect 32366 3440 32371 3496
rect 29453 3438 32371 3440
rect 29453 3435 29519 3438
rect 32305 3435 32371 3438
rect 46657 3498 46723 3501
rect 49200 3498 50000 3528
rect 46657 3496 50000 3498
rect 46657 3440 46662 3496
rect 46718 3440 50000 3496
rect 46657 3438 50000 3440
rect 46657 3435 46723 3438
rect 49200 3408 50000 3438
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 21173 2954 21239 2957
rect 22645 2954 22711 2957
rect 21173 2952 22711 2954
rect 21173 2896 21178 2952
rect 21234 2896 22650 2952
rect 22706 2896 22711 2952
rect 21173 2894 22711 2896
rect 21173 2891 21239 2894
rect 22645 2891 22711 2894
rect 0 2728 800 2848
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 49200 2728 50000 2848
rect 34928 2687 35248 2688
rect 10409 2410 10475 2413
rect 24894 2410 24900 2412
rect 10409 2408 24900 2410
rect 10409 2352 10414 2408
rect 10470 2352 24900 2408
rect 10409 2350 24900 2352
rect 10409 2347 10475 2350
rect 24894 2348 24900 2350
rect 24964 2348 24970 2412
rect 19568 2208 19888 2209
rect 0 2138 800 2168
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 3417 2138 3483 2141
rect 0 2136 3483 2138
rect 0 2080 3422 2136
rect 3478 2080 3483 2136
rect 0 2078 3483 2080
rect 0 2048 800 2078
rect 3417 2075 3483 2078
rect 49200 2048 50000 2168
rect 0 1368 800 1488
rect 46381 1458 46447 1461
rect 49200 1458 50000 1488
rect 46381 1456 50000 1458
rect 46381 1400 46386 1456
rect 46442 1400 50000 1456
rect 46381 1398 50000 1400
rect 46381 1395 46447 1398
rect 49200 1368 50000 1398
rect 0 778 800 808
rect 1393 778 1459 781
rect 0 776 1459 778
rect 0 720 1398 776
rect 1454 720 1459 776
rect 0 718 1459 720
rect 0 688 800 718
rect 1393 715 1459 718
rect 47761 778 47827 781
rect 49200 778 50000 808
rect 47761 776 50000 778
rect 47761 720 47766 776
rect 47822 720 50000 776
rect 47761 718 50000 720
rect 47761 715 47827 718
rect 49200 688 50000 718
rect 46749 98 46815 101
rect 49200 98 50000 128
rect 46749 96 50000 98
rect 46749 40 46754 96
rect 46810 40 50000 96
rect 46749 38 50000 40
rect 46749 35 46815 38
rect 49200 8 50000 38
<< via3 >>
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 41828 26420 41892 26484
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 20116 25196 20180 25260
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 29132 24108 29196 24172
rect 28948 23972 29012 24036
rect 29132 24032 29196 24036
rect 29132 23976 29182 24032
rect 29182 23976 29196 24032
rect 29132 23972 29196 23976
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 20116 23428 20180 23492
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 29132 23352 29196 23356
rect 29132 23296 29182 23352
rect 29182 23296 29196 23352
rect 29132 23292 29196 23296
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 20116 22476 20180 22540
rect 24900 22400 24964 22404
rect 24900 22344 24914 22400
rect 24914 22344 24964 22400
rect 24900 22340 24964 22344
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 20116 19348 20180 19412
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 20116 15948 20180 16012
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 20300 14724 20364 14788
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19380 14512 19444 14516
rect 19380 14456 19430 14512
rect 19430 14456 19444 14512
rect 19380 14452 19444 14456
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 41828 13636 41892 13700
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 19380 11460 19444 11524
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 20300 9692 20364 9756
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 20116 7244 20180 7308
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 24900 2348 24964 2412
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 49536 4528 49552
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 19568 48992 19888 49552
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 34928 49536 35248 49552
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 41827 26484 41893 26485
rect 41827 26420 41828 26484
rect 41892 26420 41893 26484
rect 41827 26419 41893 26420
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 20115 25260 20181 25261
rect 20115 25196 20116 25260
rect 20180 25196 20181 25260
rect 20115 25195 20181 25196
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 20118 23493 20178 25195
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 29131 24172 29197 24173
rect 29131 24170 29132 24172
rect 28950 24110 29132 24170
rect 28950 24037 29010 24110
rect 29131 24108 29132 24110
rect 29196 24108 29197 24172
rect 29131 24107 29197 24108
rect 28947 24036 29013 24037
rect 28947 23972 28948 24036
rect 29012 23972 29013 24036
rect 28947 23971 29013 23972
rect 29131 24036 29197 24037
rect 29131 23972 29132 24036
rect 29196 23972 29197 24036
rect 29131 23971 29197 23972
rect 20115 23492 20181 23493
rect 20115 23428 20116 23492
rect 20180 23428 20181 23492
rect 20115 23427 20181 23428
rect 29134 23357 29194 23971
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 29131 23356 29197 23357
rect 29131 23292 29132 23356
rect 29196 23292 29197 23356
rect 29131 23291 29197 23292
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 20115 22540 20181 22541
rect 20115 22476 20116 22540
rect 20180 22476 20181 22540
rect 20115 22475 20181 22476
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 20118 19413 20178 22475
rect 24899 22404 24965 22405
rect 24899 22340 24900 22404
rect 24964 22340 24965 22404
rect 24899 22339 24965 22340
rect 20115 19412 20181 19413
rect 20115 19348 20116 19412
rect 20180 19348 20181 19412
rect 20115 19347 20181 19348
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 20115 16012 20181 16013
rect 20115 15948 20116 16012
rect 20180 15948 20181 16012
rect 20115 15947 20181 15948
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19379 14516 19445 14517
rect 19379 14452 19380 14516
rect 19444 14452 19445 14516
rect 19379 14451 19445 14452
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 19382 11525 19442 14451
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19379 11524 19445 11525
rect 19379 11460 19380 11524
rect 19444 11460 19445 11524
rect 19379 11459 19445 11460
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 20118 7309 20178 15947
rect 20299 14788 20365 14789
rect 20299 14724 20300 14788
rect 20364 14724 20365 14788
rect 20299 14723 20365 14724
rect 20302 9757 20362 14723
rect 20299 9756 20365 9757
rect 20299 9692 20300 9756
rect 20364 9692 20365 9756
rect 20299 9691 20365 9692
rect 20115 7308 20181 7309
rect 20115 7244 20116 7308
rect 20180 7244 20181 7308
rect 20115 7243 20181 7244
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 24902 2413 24962 22339
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 41830 13701 41890 26419
rect 41827 13700 41893 13701
rect 41827 13636 41828 13700
rect 41892 13636 41893 13700
rect 41827 13635 41893 13636
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 24899 2412 24965 2413
rect 24899 2348 24900 2412
rect 24964 2348 24965 2412
rect 24899 2347 24965 2348
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28980 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1644511149
transform -1 0 15640 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1644511149
transform -1 0 32016 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1644511149
transform 1 0 20148 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1644511149
transform -1 0 30728 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1644511149
transform 1 0 47104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1644511149
transform 1 0 30636 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1644511149
transform 1 0 28428 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1644511149
transform 1 0 35512 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15
timestamp 1644511149
transform 1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5152 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65
timestamp 1644511149
transform 1 0 7084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76
timestamp 1644511149
transform 1 0 8096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_95
timestamp 1644511149
transform 1 0 9844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_103
timestamp 1644511149
transform 1 0 10580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1644511149
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1644511149
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_149
timestamp 1644511149
transform 1 0 14812 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_161
timestamp 1644511149
transform 1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1644511149
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177
timestamp 1644511149
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_188
timestamp 1644511149
transform 1 0 18400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_205
timestamp 1644511149
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_210
timestamp 1644511149
transform 1 0 20424 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1644511149
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_233
timestamp 1644511149
transform 1 0 22540 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_238
timestamp 1644511149
transform 1 0 23000 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_245
timestamp 1644511149
transform 1 0 23644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1644511149
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_257
timestamp 1644511149
transform 1 0 24748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_261
timestamp 1644511149
transform 1 0 25116 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_266
timestamp 1644511149
transform 1 0 25576 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1644511149
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_287
timestamp 1644511149
transform 1 0 27508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_295
timestamp 1644511149
transform 1 0 28244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1644511149
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_309
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_320
timestamp 1644511149
transform 1 0 30544 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_332
timestamp 1644511149
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_345
timestamp 1644511149
transform 1 0 32844 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_350
timestamp 1644511149
transform 1 0 33304 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_356
timestamp 1644511149
transform 1 0 33856 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_360
timestamp 1644511149
transform 1 0 34224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_370
timestamp 1644511149
transform 1 0 35144 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_378 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_385
timestamp 1644511149
transform 1 0 36524 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1644511149
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_393
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_405
timestamp 1644511149
transform 1 0 38364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_412
timestamp 1644511149
transform 1 0 39008 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_421
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_433
timestamp 1644511149
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1644511149
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_470
timestamp 1644511149
transform 1 0 44344 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_498
timestamp 1644511149
transform 1 0 46920 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_505
timestamp 1644511149
transform 1 0 47564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_512
timestamp 1644511149
transform 1 0 48208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_28
timestamp 1644511149
transform 1 0 3680 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_35
timestamp 1644511149
transform 1 0 4324 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_43
timestamp 1644511149
transform 1 0 5060 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_48
timestamp 1644511149
transform 1 0 5520 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_78
timestamp 1644511149
transform 1 0 8280 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1644511149
transform 1 0 9016 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1644511149
transform 1 0 10120 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1644511149
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_117
timestamp 1644511149
transform 1 0 11868 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_139
timestamp 1644511149
transform 1 0 13892 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1644511149
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_202
timestamp 1644511149
transform 1 0 19688 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_209
timestamp 1644511149
transform 1 0 20332 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_215
timestamp 1644511149
transform 1 0 20884 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_219
timestamp 1644511149
transform 1 0 21252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1644511149
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_237
timestamp 1644511149
transform 1 0 22908 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_264
timestamp 1644511149
transform 1 0 25392 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_268
timestamp 1644511149
transform 1 0 25760 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_272
timestamp 1644511149
transform 1 0 26128 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_293
timestamp 1644511149
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_305
timestamp 1644511149
transform 1 0 29164 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_332
timestamp 1644511149
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_343
timestamp 1644511149
transform 1 0 32660 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_365
timestamp 1644511149
transform 1 0 34684 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_378
timestamp 1644511149
transform 1 0 35880 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1644511149
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1644511149
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_397
timestamp 1644511149
transform 1 0 37628 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_419
timestamp 1644511149
transform 1 0 39652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_444
timestamp 1644511149
transform 1 0 41952 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_449
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_453
timestamp 1644511149
transform 1 0 42780 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_460
timestamp 1644511149
transform 1 0 43424 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_485
timestamp 1644511149
transform 1 0 45724 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_495
timestamp 1644511149
transform 1 0 46644 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1644511149
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_505
timestamp 1644511149
transform 1 0 47564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_512
timestamp 1644511149
transform 1 0 48208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1644511149
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_50
timestamp 1644511149
transform 1 0 5704 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_54
timestamp 1644511149
transform 1 0 6072 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_76
timestamp 1644511149
transform 1 0 8096 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_97
timestamp 1644511149
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_109
timestamp 1644511149
transform 1 0 11132 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_113
timestamp 1644511149
transform 1 0 11500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_117
timestamp 1644511149
transform 1 0 11868 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_124
timestamp 1644511149
transform 1 0 12512 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_128
timestamp 1644511149
transform 1 0 12880 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_132
timestamp 1644511149
transform 1 0 13248 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_148
timestamp 1644511149
transform 1 0 14720 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_155
timestamp 1644511149
transform 1 0 15364 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_167
timestamp 1644511149
transform 1 0 16468 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_182
timestamp 1644511149
transform 1 0 17848 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1644511149
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1644511149
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_205
timestamp 1644511149
transform 1 0 19964 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_228
timestamp 1644511149
transform 1 0 22080 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_232
timestamp 1644511149
transform 1 0 22448 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_236
timestamp 1644511149
transform 1 0 22816 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_243
timestamp 1644511149
transform 1 0 23460 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1644511149
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_265
timestamp 1644511149
transform 1 0 25484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_290
timestamp 1644511149
transform 1 0 27784 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_298
timestamp 1644511149
transform 1 0 28520 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_304
timestamp 1644511149
transform 1 0 29072 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_312
timestamp 1644511149
transform 1 0 29808 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_339
timestamp 1644511149
transform 1 0 32292 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_347
timestamp 1644511149
transform 1 0 33028 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_351
timestamp 1644511149
transform 1 0 33396 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1644511149
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_400
timestamp 1644511149
transform 1 0 37904 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_408
timestamp 1644511149
transform 1 0 38640 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_412
timestamp 1644511149
transform 1 0 39008 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_421
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_427
timestamp 1644511149
transform 1 0 40388 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_434
timestamp 1644511149
transform 1 0 41032 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_459
timestamp 1644511149
transform 1 0 43332 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_463
timestamp 1644511149
transform 1 0 43700 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_467
timestamp 1644511149
transform 1 0 44068 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1644511149
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_480
timestamp 1644511149
transform 1 0 45264 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_509
timestamp 1644511149
transform 1 0 47932 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_515
timestamp 1644511149
transform 1 0 48484 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_8
timestamp 1644511149
transform 1 0 1840 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_15
timestamp 1644511149
transform 1 0 2484 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_24
timestamp 1644511149
transform 1 0 3312 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_31
timestamp 1644511149
transform 1 0 3956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_43
timestamp 1644511149
transform 1 0 5060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1644511149
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_60
timestamp 1644511149
transform 1 0 6624 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_67
timestamp 1644511149
transform 1 0 7268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_79
timestamp 1644511149
transform 1 0 8372 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_91
timestamp 1644511149
transform 1 0 9476 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_103
timestamp 1644511149
transform 1 0 10580 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1644511149
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_120
timestamp 1644511149
transform 1 0 12144 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_127
timestamp 1644511149
transform 1 0 12788 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_152
timestamp 1644511149
transform 1 0 15088 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1644511149
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_181
timestamp 1644511149
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_193
timestamp 1644511149
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_205
timestamp 1644511149
transform 1 0 19964 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_211
timestamp 1644511149
transform 1 0 20516 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_218
timestamp 1644511149
transform 1 0 21160 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_246
timestamp 1644511149
transform 1 0 23736 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_258
timestamp 1644511149
transform 1 0 24840 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_270
timestamp 1644511149
transform 1 0 25944 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1644511149
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_309
timestamp 1644511149
transform 1 0 29532 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_313
timestamp 1644511149
transform 1 0 29900 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_319
timestamp 1644511149
transform 1 0 30452 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_323
timestamp 1644511149
transform 1 0 30820 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_330
timestamp 1644511149
transform 1 0 31464 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_343
timestamp 1644511149
transform 1 0 32660 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_347
timestamp 1644511149
transform 1 0 33028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_359
timestamp 1644511149
transform 1 0 34132 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_371
timestamp 1644511149
transform 1 0 35236 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_386
timestamp 1644511149
transform 1 0 36616 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_404
timestamp 1644511149
transform 1 0 38272 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_416
timestamp 1644511149
transform 1 0 39376 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_420
timestamp 1644511149
transform 1 0 39744 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_432
timestamp 1644511149
transform 1 0 40848 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_438
timestamp 1644511149
transform 1 0 41400 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_442
timestamp 1644511149
transform 1 0 41768 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_452
timestamp 1644511149
transform 1 0 42688 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_460
timestamp 1644511149
transform 1 0 43424 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_464
timestamp 1644511149
transform 1 0 43792 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_471
timestamp 1644511149
transform 1 0 44436 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_482
timestamp 1644511149
transform 1 0 45448 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_489
timestamp 1644511149
transform 1 0 46092 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_500
timestamp 1644511149
transform 1 0 47104 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_505
timestamp 1644511149
transform 1 0 47564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_512
timestamp 1644511149
transform 1 0 48208 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1644511149
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_59
timestamp 1644511149
transform 1 0 6532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_71
timestamp 1644511149
transform 1 0 7636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_109
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_121
timestamp 1644511149
transform 1 0 12236 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_129
timestamp 1644511149
transform 1 0 12972 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_134
timestamp 1644511149
transform 1 0 13432 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_221
timestamp 1644511149
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_233
timestamp 1644511149
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1644511149
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1644511149
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1644511149
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_338
timestamp 1644511149
transform 1 0 32200 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_350
timestamp 1644511149
transform 1 0 33304 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_362
timestamp 1644511149
transform 1 0 34408 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_401
timestamp 1644511149
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1644511149
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1644511149
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_421
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_433
timestamp 1644511149
transform 1 0 40940 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_441
timestamp 1644511149
transform 1 0 41676 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_445
timestamp 1644511149
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_457
timestamp 1644511149
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1644511149
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1644511149
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_477
timestamp 1644511149
transform 1 0 44988 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_483
timestamp 1644511149
transform 1 0 45540 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_487
timestamp 1644511149
transform 1 0 45908 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_512
timestamp 1644511149
transform 1 0 48208 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_28
timestamp 1644511149
transform 1 0 3680 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_40
timestamp 1644511149
transform 1 0 4784 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1644511149
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_205
timestamp 1644511149
transform 1 0 19964 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_211
timestamp 1644511149
transform 1 0 20516 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_220
timestamp 1644511149
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_241
timestamp 1644511149
transform 1 0 23276 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_250
timestamp 1644511149
transform 1 0 24104 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_262
timestamp 1644511149
transform 1 0 25208 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_274
timestamp 1644511149
transform 1 0 26312 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_297
timestamp 1644511149
transform 1 0 28428 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_309
timestamp 1644511149
transform 1 0 29532 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_321
timestamp 1644511149
transform 1 0 30636 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_333
timestamp 1644511149
transform 1 0 31740 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1644511149
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_405
timestamp 1644511149
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_417
timestamp 1644511149
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_429
timestamp 1644511149
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1644511149
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1644511149
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_449
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_461
timestamp 1644511149
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_473
timestamp 1644511149
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_485
timestamp 1644511149
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_500
timestamp 1644511149
transform 1 0 47104 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_505
timestamp 1644511149
transform 1 0 47564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_512
timestamp 1644511149
transform 1 0 48208 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_8
timestamp 1644511149
transform 1 0 1840 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_22
timestamp 1644511149
transform 1 0 3128 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_228
timestamp 1644511149
transform 1 0 22080 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_240
timestamp 1644511149
transform 1 0 23184 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_269
timestamp 1644511149
transform 1 0 25852 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_281
timestamp 1644511149
transform 1 0 26956 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_299
timestamp 1644511149
transform 1 0 28612 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1644511149
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1644511149
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_433
timestamp 1644511149
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_445
timestamp 1644511149
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_457
timestamp 1644511149
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1644511149
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1644511149
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_477
timestamp 1644511149
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_489
timestamp 1644511149
transform 1 0 46092 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_512
timestamp 1644511149
transform 1 0 48208 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_6
timestamp 1644511149
transform 1 0 1656 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_31
timestamp 1644511149
transform 1 0 3956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_43
timestamp 1644511149
transform 1 0 5060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_213
timestamp 1644511149
transform 1 0 20700 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_219
timestamp 1644511149
transform 1 0 21252 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_241
timestamp 1644511149
transform 1 0 23276 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_250
timestamp 1644511149
transform 1 0 24104 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_262
timestamp 1644511149
transform 1 0 25208 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_274
timestamp 1644511149
transform 1 0 26312 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_287
timestamp 1644511149
transform 1 0 27508 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1644511149
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1644511149
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_461
timestamp 1644511149
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_473
timestamp 1644511149
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_485
timestamp 1644511149
transform 1 0 45724 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_489
timestamp 1644511149
transform 1 0 46092 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_501
timestamp 1644511149
transform 1 0 47196 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_508
timestamp 1644511149
transform 1 0 47840 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_19
timestamp 1644511149
transform 1 0 2852 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_23
timestamp 1644511149
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_201
timestamp 1644511149
transform 1 0 19596 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_213
timestamp 1644511149
transform 1 0 20700 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_220
timestamp 1644511149
transform 1 0 21344 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_232
timestamp 1644511149
transform 1 0 22448 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_244
timestamp 1644511149
transform 1 0 23552 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_330
timestamp 1644511149
transform 1 0 31464 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_342
timestamp 1644511149
transform 1 0 32568 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_354
timestamp 1644511149
transform 1 0 33672 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_362
timestamp 1644511149
transform 1 0 34408 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_401
timestamp 1644511149
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1644511149
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1644511149
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_433
timestamp 1644511149
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_445
timestamp 1644511149
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_457
timestamp 1644511149
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1644511149
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1644511149
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_477
timestamp 1644511149
transform 1 0 44988 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_483
timestamp 1644511149
transform 1 0 45540 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_505
timestamp 1644511149
transform 1 0 47564 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_513
timestamp 1644511149
transform 1 0 48300 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_14
timestamp 1644511149
transform 1 0 2392 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_26
timestamp 1644511149
transform 1 0 3496 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_38
timestamp 1644511149
transform 1 0 4600 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_50
timestamp 1644511149
transform 1 0 5704 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_187
timestamp 1644511149
transform 1 0 18308 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_191
timestamp 1644511149
transform 1 0 18676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_197
timestamp 1644511149
transform 1 0 19228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_206
timestamp 1644511149
transform 1 0 20056 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_218
timestamp 1644511149
transform 1 0 21160 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_259
timestamp 1644511149
transform 1 0 24932 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_271
timestamp 1644511149
transform 1 0 26036 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_299
timestamp 1644511149
transform 1 0 28612 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_319
timestamp 1644511149
transform 1 0 30452 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_326
timestamp 1644511149
transform 1 0 31096 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_334
timestamp 1644511149
transform 1 0 31832 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_417
timestamp 1644511149
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_429
timestamp 1644511149
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1644511149
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1644511149
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_461
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_473
timestamp 1644511149
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_485
timestamp 1644511149
transform 1 0 45724 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_493
timestamp 1644511149
transform 1 0 46460 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_498
timestamp 1644511149
transform 1 0 46920 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_508
timestamp 1644511149
transform 1 0 47840 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_13
timestamp 1644511149
transform 1 0 2300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1644511149
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_185
timestamp 1644511149
transform 1 0 18124 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_192
timestamp 1644511149
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_218
timestamp 1644511149
transform 1 0 21160 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_226
timestamp 1644511149
transform 1 0 21896 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_237
timestamp 1644511149
transform 1 0 22908 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_249
timestamp 1644511149
transform 1 0 24012 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_261
timestamp 1644511149
transform 1 0 25116 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_278
timestamp 1644511149
transform 1 0 26680 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_290
timestamp 1644511149
transform 1 0 27784 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_302
timestamp 1644511149
transform 1 0 28888 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_315
timestamp 1644511149
transform 1 0 30084 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_340
timestamp 1644511149
transform 1 0 32384 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_352
timestamp 1644511149
transform 1 0 33488 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1644511149
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1644511149
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1644511149
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_457
timestamp 1644511149
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1644511149
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1644511149
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_477
timestamp 1644511149
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_489
timestamp 1644511149
transform 1 0 46092 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_512
timestamp 1644511149
transform 1 0 48208 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_13
timestamp 1644511149
transform 1 0 2300 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_25
timestamp 1644511149
transform 1 0 3404 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_37
timestamp 1644511149
transform 1 0 4508 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_49
timestamp 1644511149
transform 1 0 5612 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_177
timestamp 1644511149
transform 1 0 17388 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_195
timestamp 1644511149
transform 1 0 19044 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_220
timestamp 1644511149
transform 1 0 21344 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_241
timestamp 1644511149
transform 1 0 23276 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_258
timestamp 1644511149
transform 1 0 24840 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_268
timestamp 1644511149
transform 1 0 25760 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_292
timestamp 1644511149
transform 1 0 27968 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_312
timestamp 1644511149
transform 1 0 29808 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_332
timestamp 1644511149
transform 1 0 31648 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_342
timestamp 1644511149
transform 1 0 32568 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_354
timestamp 1644511149
transform 1 0 33672 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_366
timestamp 1644511149
transform 1 0 34776 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_378
timestamp 1644511149
transform 1 0 35880 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_390
timestamp 1644511149
transform 1 0 36984 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_417
timestamp 1644511149
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1644511149
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1644511149
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_449
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_461
timestamp 1644511149
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_473
timestamp 1644511149
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_485
timestamp 1644511149
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1644511149
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1644511149
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_505
timestamp 1644511149
transform 1 0 47564 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_512
timestamp 1644511149
transform 1 0 48208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_14
timestamp 1644511149
transform 1 0 2392 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1644511149
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_192
timestamp 1644511149
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_213
timestamp 1644511149
transform 1 0 20700 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_223
timestamp 1644511149
transform 1 0 21620 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_236
timestamp 1644511149
transform 1 0 22816 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_248
timestamp 1644511149
transform 1 0 23920 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_262
timestamp 1644511149
transform 1 0 25208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_273
timestamp 1644511149
transform 1 0 26220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_282
timestamp 1644511149
transform 1 0 27048 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_302
timestamp 1644511149
transform 1 0 28888 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_329
timestamp 1644511149
transform 1 0 31372 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_341
timestamp 1644511149
transform 1 0 32476 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_353
timestamp 1644511149
transform 1 0 33580 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_361
timestamp 1644511149
transform 1 0 34316 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_445
timestamp 1644511149
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_457
timestamp 1644511149
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1644511149
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1644511149
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_477
timestamp 1644511149
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_489
timestamp 1644511149
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_501
timestamp 1644511149
transform 1 0 47196 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_505
timestamp 1644511149
transform 1 0 47564 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_512
timestamp 1644511149
transform 1 0 48208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_28
timestamp 1644511149
transform 1 0 3680 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_40
timestamp 1644511149
transform 1 0 4784 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_52
timestamp 1644511149
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_180
timestamp 1644511149
transform 1 0 17664 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_189
timestamp 1644511149
transform 1 0 18492 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_197
timestamp 1644511149
transform 1 0 19228 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_207
timestamp 1644511149
transform 1 0 20148 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_219
timestamp 1644511149
transform 1 0 21252 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_235
timestamp 1644511149
transform 1 0 22724 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_243
timestamp 1644511149
transform 1 0 23460 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_260
timestamp 1644511149
transform 1 0 25024 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_266
timestamp 1644511149
transform 1 0 25576 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_276
timestamp 1644511149
transform 1 0 26496 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_292
timestamp 1644511149
transform 1 0 27968 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_304
timestamp 1644511149
transform 1 0 29072 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_316
timestamp 1644511149
transform 1 0 30176 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_332
timestamp 1644511149
transform 1 0 31648 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_342
timestamp 1644511149
transform 1 0 32568 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_354
timestamp 1644511149
transform 1 0 33672 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_366
timestamp 1644511149
transform 1 0 34776 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_378
timestamp 1644511149
transform 1 0 35880 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_390
timestamp 1644511149
transform 1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_417
timestamp 1644511149
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_429
timestamp 1644511149
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1644511149
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1644511149
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_461
timestamp 1644511149
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_473
timestamp 1644511149
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_485
timestamp 1644511149
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1644511149
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1644511149
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_505
timestamp 1644511149
transform 1 0 47564 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_513
timestamp 1644511149
transform 1 0 48300 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_7
timestamp 1644511149
transform 1 0 1748 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_11
timestamp 1644511149
transform 1 0 2116 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_23
timestamp 1644511149
transform 1 0 3220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_187
timestamp 1644511149
transform 1 0 18308 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_203
timestamp 1644511149
transform 1 0 19780 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_215
timestamp 1644511149
transform 1 0 20884 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_223
timestamp 1644511149
transform 1 0 21620 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_230
timestamp 1644511149
transform 1 0 22264 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_236
timestamp 1644511149
transform 1 0 22816 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_240
timestamp 1644511149
transform 1 0 23184 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_248
timestamp 1644511149
transform 1 0 23920 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_258
timestamp 1644511149
transform 1 0 24840 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_269
timestamp 1644511149
transform 1 0 25852 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_279
timestamp 1644511149
transform 1 0 26772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_287
timestamp 1644511149
transform 1 0 27508 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_304
timestamp 1644511149
transform 1 0 29072 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_325
timestamp 1644511149
transform 1 0 31004 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_347
timestamp 1644511149
transform 1 0 33028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_359
timestamp 1644511149
transform 1 0 34132 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1644511149
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1644511149
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_433
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_445
timestamp 1644511149
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_457
timestamp 1644511149
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1644511149
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1644511149
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_477
timestamp 1644511149
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_489
timestamp 1644511149
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_501
timestamp 1644511149
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_513
timestamp 1644511149
transform 1 0 48300 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_7
timestamp 1644511149
transform 1 0 1748 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_14
timestamp 1644511149
transform 1 0 2392 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_26
timestamp 1644511149
transform 1 0 3496 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_38
timestamp 1644511149
transform 1 0 4600 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_50
timestamp 1644511149
transform 1 0 5704 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_197
timestamp 1644511149
transform 1 0 19228 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_209
timestamp 1644511149
transform 1 0 20332 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_221
timestamp 1644511149
transform 1 0 21436 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_233
timestamp 1644511149
transform 1 0 22540 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_243
timestamp 1644511149
transform 1 0 23460 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_251
timestamp 1644511149
transform 1 0 24196 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_266
timestamp 1644511149
transform 1 0 25576 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_270
timestamp 1644511149
transform 1 0 25944 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_275
timestamp 1644511149
transform 1 0 26404 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_284
timestamp 1644511149
transform 1 0 27232 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_296
timestamp 1644511149
transform 1 0 28336 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_308
timestamp 1644511149
transform 1 0 29440 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_320
timestamp 1644511149
transform 1 0 30544 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_332
timestamp 1644511149
transform 1 0 31648 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_341
timestamp 1644511149
transform 1 0 32476 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_345
timestamp 1644511149
transform 1 0 32844 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_370
timestamp 1644511149
transform 1 0 35144 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_382
timestamp 1644511149
transform 1 0 36248 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_390
timestamp 1644511149
transform 1 0 36984 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_417
timestamp 1644511149
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_429
timestamp 1644511149
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1644511149
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1644511149
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_461
timestamp 1644511149
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_473
timestamp 1644511149
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_485
timestamp 1644511149
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_500
timestamp 1644511149
transform 1 0 47104 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_505
timestamp 1644511149
transform 1 0 47564 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_512
timestamp 1644511149
transform 1 0 48208 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_24
timestamp 1644511149
transform 1 0 3312 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1644511149
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_202
timestamp 1644511149
transform 1 0 19688 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_226
timestamp 1644511149
transform 1 0 21896 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_230
timestamp 1644511149
transform 1 0 22264 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_247
timestamp 1644511149
transform 1 0 23828 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_260
timestamp 1644511149
transform 1 0 25024 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_270
timestamp 1644511149
transform 1 0 25944 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_278
timestamp 1644511149
transform 1 0 26680 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_293
timestamp 1644511149
transform 1 0 28060 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1644511149
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_317
timestamp 1644511149
transform 1 0 30268 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_329
timestamp 1644511149
transform 1 0 31372 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_346
timestamp 1644511149
transform 1 0 32936 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_358
timestamp 1644511149
transform 1 0 34040 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1644511149
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1644511149
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_433
timestamp 1644511149
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_445
timestamp 1644511149
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_457
timestamp 1644511149
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1644511149
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1644511149
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_477
timestamp 1644511149
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_489
timestamp 1644511149
transform 1 0 46092 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_512
timestamp 1644511149
transform 1 0 48208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_9
timestamp 1644511149
transform 1 0 1932 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_13
timestamp 1644511149
transform 1 0 2300 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_25
timestamp 1644511149
transform 1 0 3404 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_37
timestamp 1644511149
transform 1 0 4508 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_49
timestamp 1644511149
transform 1 0 5612 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_197
timestamp 1644511149
transform 1 0 19228 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_209
timestamp 1644511149
transform 1 0 20332 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_221
timestamp 1644511149
transform 1 0 21436 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_234
timestamp 1644511149
transform 1 0 22632 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_244
timestamp 1644511149
transform 1 0 23552 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_256
timestamp 1644511149
transform 1 0 24656 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_264
timestamp 1644511149
transform 1 0 25392 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_271
timestamp 1644511149
transform 1 0 26036 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_289
timestamp 1644511149
transform 1 0 27692 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_306
timestamp 1644511149
transform 1 0 29256 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_314
timestamp 1644511149
transform 1 0 29992 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_320
timestamp 1644511149
transform 1 0 30544 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_332
timestamp 1644511149
transform 1 0 31648 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_342
timestamp 1644511149
transform 1 0 32568 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_369
timestamp 1644511149
transform 1 0 35052 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_381
timestamp 1644511149
transform 1 0 36156 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_389
timestamp 1644511149
transform 1 0 36892 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_417
timestamp 1644511149
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_429
timestamp 1644511149
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1644511149
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1644511149
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_449
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_461
timestamp 1644511149
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_473
timestamp 1644511149
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_485
timestamp 1644511149
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1644511149
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1644511149
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_508
timestamp 1644511149
transform 1 0 47840 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_183
timestamp 1644511149
transform 1 0 17940 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_192
timestamp 1644511149
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_218
timestamp 1644511149
transform 1 0 21160 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_222
timestamp 1644511149
transform 1 0 21528 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_232
timestamp 1644511149
transform 1 0 22448 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_243
timestamp 1644511149
transform 1 0 23460 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_259
timestamp 1644511149
transform 1 0 24932 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_270
timestamp 1644511149
transform 1 0 25944 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_282
timestamp 1644511149
transform 1 0 27048 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_293
timestamp 1644511149
transform 1 0 28060 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_305
timestamp 1644511149
transform 1 0 29164 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_317
timestamp 1644511149
transform 1 0 30268 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_322
timestamp 1644511149
transform 1 0 30728 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_336
timestamp 1644511149
transform 1 0 32016 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_345
timestamp 1644511149
transform 1 0 32844 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_352
timestamp 1644511149
transform 1 0 33488 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_373
timestamp 1644511149
transform 1 0 35420 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_382
timestamp 1644511149
transform 1 0 36248 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_394
timestamp 1644511149
transform 1 0 37352 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_406
timestamp 1644511149
transform 1 0 38456 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_418
timestamp 1644511149
transform 1 0 39560 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_421
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_433
timestamp 1644511149
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_445
timestamp 1644511149
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_457
timestamp 1644511149
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1644511149
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1644511149
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_477
timestamp 1644511149
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_489
timestamp 1644511149
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_501
timestamp 1644511149
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_513
timestamp 1644511149
transform 1 0 48300 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_7
timestamp 1644511149
transform 1 0 1748 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_19
timestamp 1644511149
transform 1 0 2852 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_31
timestamp 1644511149
transform 1 0 3956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_43
timestamp 1644511149
transform 1 0 5060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1644511149
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_190
timestamp 1644511149
transform 1 0 18584 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_208
timestamp 1644511149
transform 1 0 20240 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_215
timestamp 1644511149
transform 1 0 20884 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1644511149
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_231
timestamp 1644511149
transform 1 0 22356 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_249
timestamp 1644511149
transform 1 0 24012 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_257
timestamp 1644511149
transform 1 0 24748 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_267
timestamp 1644511149
transform 1 0 25668 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_275
timestamp 1644511149
transform 1 0 26404 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_288
timestamp 1644511149
transform 1 0 27600 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_294
timestamp 1644511149
transform 1 0 28152 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_311
timestamp 1644511149
transform 1 0 29716 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_328
timestamp 1644511149
transform 1 0 31280 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_353
timestamp 1644511149
transform 1 0 33580 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_378
timestamp 1644511149
transform 1 0 35880 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_390
timestamp 1644511149
transform 1 0 36984 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_417
timestamp 1644511149
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_429
timestamp 1644511149
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1644511149
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1644511149
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_461
timestamp 1644511149
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_473
timestamp 1644511149
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_485
timestamp 1644511149
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1644511149
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1644511149
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_505
timestamp 1644511149
transform 1 0 47564 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_513
timestamp 1644511149
transform 1 0 48300 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_9
timestamp 1644511149
transform 1 0 1932 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_13
timestamp 1644511149
transform 1 0 2300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_25
timestamp 1644511149
transform 1 0 3404 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_165
timestamp 1644511149
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_177
timestamp 1644511149
transform 1 0 17388 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_183
timestamp 1644511149
transform 1 0 17940 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_192
timestamp 1644511149
transform 1 0 18768 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_207
timestamp 1644511149
transform 1 0 20148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_224
timestamp 1644511149
transform 1 0 21712 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_236
timestamp 1644511149
transform 1 0 22816 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1644511149
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_262
timestamp 1644511149
transform 1 0 25208 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_274
timestamp 1644511149
transform 1 0 26312 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_282
timestamp 1644511149
transform 1 0 27048 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_295
timestamp 1644511149
transform 1 0 28244 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_304
timestamp 1644511149
transform 1 0 29072 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_317
timestamp 1644511149
transform 1 0 30268 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_322
timestamp 1644511149
transform 1 0 30728 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_330
timestamp 1644511149
transform 1 0 31464 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_335
timestamp 1644511149
transform 1 0 31924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_360
timestamp 1644511149
transform 1 0 34224 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_381
timestamp 1644511149
transform 1 0 36156 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_393
timestamp 1644511149
transform 1 0 37260 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_405
timestamp 1644511149
transform 1 0 38364 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_417
timestamp 1644511149
transform 1 0 39468 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_433
timestamp 1644511149
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_445
timestamp 1644511149
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_457
timestamp 1644511149
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1644511149
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1644511149
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_477
timestamp 1644511149
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_489
timestamp 1644511149
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_501
timestamp 1644511149
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_513
timestamp 1644511149
transform 1 0 48300 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_28
timestamp 1644511149
transform 1 0 3680 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_40
timestamp 1644511149
transform 1 0 4784 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp 1644511149
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1644511149
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1644511149
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_172
timestamp 1644511149
transform 1 0 16928 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_192
timestamp 1644511149
transform 1 0 18768 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_202
timestamp 1644511149
transform 1 0 19688 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_209
timestamp 1644511149
transform 1 0 20332 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_220
timestamp 1644511149
transform 1 0 21344 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_234
timestamp 1644511149
transform 1 0 22632 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_242
timestamp 1644511149
transform 1 0 23368 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_250
timestamp 1644511149
transform 1 0 24104 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_256
timestamp 1644511149
transform 1 0 24656 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_266
timestamp 1644511149
transform 1 0 25576 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_276
timestamp 1644511149
transform 1 0 26496 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_294
timestamp 1644511149
transform 1 0 28152 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_300
timestamp 1644511149
transform 1 0 28704 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_305
timestamp 1644511149
transform 1 0 29164 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_313
timestamp 1644511149
transform 1 0 29900 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_325
timestamp 1644511149
transform 1 0 31004 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_333
timestamp 1644511149
transform 1 0 31740 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_340
timestamp 1644511149
transform 1 0 32384 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_348
timestamp 1644511149
transform 1 0 33120 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_357
timestamp 1644511149
transform 1 0 33948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_369
timestamp 1644511149
transform 1 0 35052 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_378
timestamp 1644511149
transform 1 0 35880 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_390
timestamp 1644511149
transform 1 0 36984 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_401
timestamp 1644511149
transform 1 0 37996 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_425
timestamp 1644511149
transform 1 0 40204 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_437
timestamp 1644511149
transform 1 0 41308 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_445
timestamp 1644511149
transform 1 0 42044 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_461
timestamp 1644511149
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_473
timestamp 1644511149
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_485
timestamp 1644511149
transform 1 0 45724 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_493
timestamp 1644511149
transform 1 0 46460 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_498
timestamp 1644511149
transform 1 0 46920 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_21_505
timestamp 1644511149
transform 1 0 47564 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_512
timestamp 1644511149
transform 1 0 48208 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_7
timestamp 1644511149
transform 1 0 1748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_11
timestamp 1644511149
transform 1 0 2116 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_23
timestamp 1644511149
transform 1 0 3220 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_153
timestamp 1644511149
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_165
timestamp 1644511149
transform 1 0 16284 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_169
timestamp 1644511149
transform 1 0 16652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_176
timestamp 1644511149
transform 1 0 17296 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_192
timestamp 1644511149
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_213
timestamp 1644511149
transform 1 0 20700 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_217
timestamp 1644511149
transform 1 0 21068 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_222
timestamp 1644511149
transform 1 0 21528 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_226
timestamp 1644511149
transform 1 0 21896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_236
timestamp 1644511149
transform 1 0 22816 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_248
timestamp 1644511149
transform 1 0 23920 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_260
timestamp 1644511149
transform 1 0 25024 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_271
timestamp 1644511149
transform 1 0 26036 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_282
timestamp 1644511149
transform 1 0 27048 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_286
timestamp 1644511149
transform 1 0 27416 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_296
timestamp 1644511149
transform 1 0 28336 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_321
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_325
timestamp 1644511149
transform 1 0 31004 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_331
timestamp 1644511149
transform 1 0 31556 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_339
timestamp 1644511149
transform 1 0 32292 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_344
timestamp 1644511149
transform 1 0 32752 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_360
timestamp 1644511149
transform 1 0 34224 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_373
timestamp 1644511149
transform 1 0 35420 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_381
timestamp 1644511149
transform 1 0 36156 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_400
timestamp 1644511149
transform 1 0 37904 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_404
timestamp 1644511149
transform 1 0 38272 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_408
timestamp 1644511149
transform 1 0 38640 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_433
timestamp 1644511149
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_445
timestamp 1644511149
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_457
timestamp 1644511149
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1644511149
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1644511149
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_477
timestamp 1644511149
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_489
timestamp 1644511149
transform 1 0 46092 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_512
timestamp 1644511149
transform 1 0 48208 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1644511149
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1644511149
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1644511149
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_164
timestamp 1644511149
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_190
timestamp 1644511149
transform 1 0 18584 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_214
timestamp 1644511149
transform 1 0 20792 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1644511149
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_232
timestamp 1644511149
transform 1 0 22448 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_242
timestamp 1644511149
transform 1 0 23368 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_248
timestamp 1644511149
transform 1 0 23920 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_253
timestamp 1644511149
transform 1 0 24380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_261
timestamp 1644511149
transform 1 0 25116 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_269
timestamp 1644511149
transform 1 0 25852 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_276
timestamp 1644511149
transform 1 0 26496 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_285
timestamp 1644511149
transform 1 0 27324 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_295
timestamp 1644511149
transform 1 0 28244 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_318
timestamp 1644511149
transform 1 0 30360 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_322
timestamp 1644511149
transform 1 0 30728 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_332
timestamp 1644511149
transform 1 0 31648 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_353
timestamp 1644511149
transform 1 0 33580 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_377
timestamp 1644511149
transform 1 0 35788 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_388
timestamp 1644511149
transform 1 0 36800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_414
timestamp 1644511149
transform 1 0 39192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_434
timestamp 1644511149
transform 1 0 41032 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_446
timestamp 1644511149
transform 1 0 42136 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_461
timestamp 1644511149
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_473
timestamp 1644511149
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_485
timestamp 1644511149
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_500
timestamp 1644511149
transform 1 0 47104 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_508
timestamp 1644511149
transform 1 0 47840 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1644511149
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1644511149
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_144
timestamp 1644511149
transform 1 0 14352 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_152
timestamp 1644511149
transform 1 0 15088 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_158
timestamp 1644511149
transform 1 0 15640 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_166
timestamp 1644511149
transform 1 0 16376 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_191
timestamp 1644511149
transform 1 0 18676 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1644511149
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_214
timestamp 1644511149
transform 1 0 20792 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_222
timestamp 1644511149
transform 1 0 21528 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_228
timestamp 1644511149
transform 1 0 22080 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_248
timestamp 1644511149
transform 1 0 23920 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_258
timestamp 1644511149
transform 1 0 24840 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_265
timestamp 1644511149
transform 1 0 25484 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_269
timestamp 1644511149
transform 1 0 25852 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_279
timestamp 1644511149
transform 1 0 26772 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_287
timestamp 1644511149
transform 1 0 27508 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_304
timestamp 1644511149
transform 1 0 29072 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_317
timestamp 1644511149
transform 1 0 30268 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_336
timestamp 1644511149
transform 1 0 32016 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_348
timestamp 1644511149
transform 1 0 33120 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_360
timestamp 1644511149
transform 1 0 34224 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_370
timestamp 1644511149
transform 1 0 35144 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_382
timestamp 1644511149
transform 1 0 36248 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_394
timestamp 1644511149
transform 1 0 37352 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_403
timestamp 1644511149
transform 1 0 38180 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_407
timestamp 1644511149
transform 1 0 38548 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1644511149
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1644511149
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_425
timestamp 1644511149
transform 1 0 40204 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_443
timestamp 1644511149
transform 1 0 41860 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_455
timestamp 1644511149
transform 1 0 42964 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_467
timestamp 1644511149
transform 1 0 44068 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1644511149
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_477
timestamp 1644511149
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_489
timestamp 1644511149
transform 1 0 46092 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_512
timestamp 1644511149
transform 1 0 48208 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_14
timestamp 1644511149
transform 1 0 2392 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_26
timestamp 1644511149
transform 1 0 3496 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_38
timestamp 1644511149
transform 1 0 4600 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_50
timestamp 1644511149
transform 1 0 5704 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_137
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1644511149
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1644511149
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_192
timestamp 1644511149
transform 1 0 18768 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_208
timestamp 1644511149
transform 1 0 20240 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_215
timestamp 1644511149
transform 1 0 20884 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_234
timestamp 1644511149
transform 1 0 22632 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_240
timestamp 1644511149
transform 1 0 23184 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_246
timestamp 1644511149
transform 1 0 23736 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_255
timestamp 1644511149
transform 1 0 24564 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_262
timestamp 1644511149
transform 1 0 25208 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_274
timestamp 1644511149
transform 1 0 26312 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_305
timestamp 1644511149
transform 1 0 29164 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_311
timestamp 1644511149
transform 1 0 29716 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_325
timestamp 1644511149
transform 1 0 31004 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_333
timestamp 1644511149
transform 1 0 31740 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_345
timestamp 1644511149
transform 1 0 32844 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_355
timestamp 1644511149
transform 1 0 33764 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_375
timestamp 1644511149
transform 1 0 35604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_387
timestamp 1644511149
transform 1 0 36708 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_399
timestamp 1644511149
transform 1 0 37812 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_407
timestamp 1644511149
transform 1 0 38548 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_417
timestamp 1644511149
transform 1 0 39468 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_425
timestamp 1644511149
transform 1 0 40204 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_432
timestamp 1644511149
transform 1 0 40848 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_439
timestamp 1644511149
transform 1 0 41492 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1644511149
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_452
timestamp 1644511149
transform 1 0 42688 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_464
timestamp 1644511149
transform 1 0 43792 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_476
timestamp 1644511149
transform 1 0 44896 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_484
timestamp 1644511149
transform 1 0 45632 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_488
timestamp 1644511149
transform 1 0 46000 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_495
timestamp 1644511149
transform 1 0 46644 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1644511149
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_508
timestamp 1644511149
transform 1 0 47840 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1644511149
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_121
timestamp 1644511149
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1644511149
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1644511149
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_153
timestamp 1644511149
transform 1 0 15180 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_164
timestamp 1644511149
transform 1 0 16192 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_188
timestamp 1644511149
transform 1 0 18400 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_203
timestamp 1644511149
transform 1 0 19780 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_207
timestamp 1644511149
transform 1 0 20148 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_224
timestamp 1644511149
transform 1 0 21712 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_231
timestamp 1644511149
transform 1 0 22356 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_244
timestamp 1644511149
transform 1 0 23552 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_263
timestamp 1644511149
transform 1 0 25300 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_274
timestamp 1644511149
transform 1 0 26312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_282
timestamp 1644511149
transform 1 0 27048 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_292
timestamp 1644511149
transform 1 0 27968 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_304
timestamp 1644511149
transform 1 0 29072 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_321
timestamp 1644511149
transform 1 0 30636 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_327
timestamp 1644511149
transform 1 0 31188 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_347
timestamp 1644511149
transform 1 0 33028 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_359
timestamp 1644511149
transform 1 0 34132 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_403
timestamp 1644511149
transform 1 0 38180 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_416
timestamp 1644511149
transform 1 0 39376 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_421
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_440
timestamp 1644511149
transform 1 0 41584 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_449
timestamp 1644511149
transform 1 0 42412 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_461
timestamp 1644511149
transform 1 0 43516 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_473
timestamp 1644511149
transform 1 0 44620 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_477
timestamp 1644511149
transform 1 0 44988 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_483
timestamp 1644511149
transform 1 0 45540 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_487
timestamp 1644511149
transform 1 0 45908 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_512
timestamp 1644511149
transform 1 0 48208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_11
timestamp 1644511149
transform 1 0 2116 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_18
timestamp 1644511149
transform 1 0 2760 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_30
timestamp 1644511149
transform 1 0 3864 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_42
timestamp 1644511149
transform 1 0 4968 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1644511149
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_137
timestamp 1644511149
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_149
timestamp 1644511149
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_164
timestamp 1644511149
transform 1 0 16192 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_190
timestamp 1644511149
transform 1 0 18584 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_210
timestamp 1644511149
transform 1 0 20424 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1644511149
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_233
timestamp 1644511149
transform 1 0 22540 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_240
timestamp 1644511149
transform 1 0 23184 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_244
timestamp 1644511149
transform 1 0 23552 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_249
timestamp 1644511149
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_261
timestamp 1644511149
transform 1 0 25116 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_268
timestamp 1644511149
transform 1 0 25760 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_276
timestamp 1644511149
transform 1 0 26496 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_287
timestamp 1644511149
transform 1 0 27508 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_294
timestamp 1644511149
transform 1 0 28152 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_306
timestamp 1644511149
transform 1 0 29256 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_319
timestamp 1644511149
transform 1 0 30452 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_327
timestamp 1644511149
transform 1 0 31188 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1644511149
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_355
timestamp 1644511149
transform 1 0 33764 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_361
timestamp 1644511149
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_373
timestamp 1644511149
transform 1 0 35420 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_381
timestamp 1644511149
transform 1 0 36156 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_389
timestamp 1644511149
transform 1 0 36892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_401
timestamp 1644511149
transform 1 0 37996 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_413
timestamp 1644511149
transform 1 0 39100 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_425
timestamp 1644511149
transform 1 0 40204 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_434
timestamp 1644511149
transform 1 0 41032 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_443
timestamp 1644511149
transform 1 0 41860 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1644511149
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_449
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_461
timestamp 1644511149
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_473
timestamp 1644511149
transform 1 0 44620 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_500
timestamp 1644511149
transform 1 0 47104 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_508
timestamp 1644511149
transform 1 0 47840 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1644511149
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1644511149
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1644511149
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_153
timestamp 1644511149
transform 1 0 15180 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_162
timestamp 1644511149
transform 1 0 16008 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_174
timestamp 1644511149
transform 1 0 17112 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_183
timestamp 1644511149
transform 1 0 17940 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1644511149
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_214
timestamp 1644511149
transform 1 0 20792 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_226
timestamp 1644511149
transform 1 0 21896 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_236
timestamp 1644511149
transform 1 0 22816 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_246
timestamp 1644511149
transform 1 0 23736 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_261
timestamp 1644511149
transform 1 0 25116 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_269
timestamp 1644511149
transform 1 0 25852 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_277
timestamp 1644511149
transform 1 0 26588 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_285
timestamp 1644511149
transform 1 0 27324 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_290
timestamp 1644511149
transform 1 0 27784 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_298
timestamp 1644511149
transform 1 0 28520 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_304
timestamp 1644511149
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_325
timestamp 1644511149
transform 1 0 31004 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_339
timestamp 1644511149
transform 1 0 32292 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_347
timestamp 1644511149
transform 1 0 33028 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_360
timestamp 1644511149
transform 1 0 34224 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_389
timestamp 1644511149
transform 1 0 36892 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_397
timestamp 1644511149
transform 1 0 37628 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_403
timestamp 1644511149
transform 1 0 38180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_415
timestamp 1644511149
transform 1 0 39284 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1644511149
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_421
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_432
timestamp 1644511149
transform 1 0 40848 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_439
timestamp 1644511149
transform 1 0 41492 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_443
timestamp 1644511149
transform 1 0 41860 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_447
timestamp 1644511149
transform 1 0 42228 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_455
timestamp 1644511149
transform 1 0 42964 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_459
timestamp 1644511149
transform 1 0 43332 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_471
timestamp 1644511149
transform 1 0 44436 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1644511149
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_485
timestamp 1644511149
transform 1 0 45724 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_512
timestamp 1644511149
transform 1 0 48208 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_9
timestamp 1644511149
transform 1 0 1932 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_13
timestamp 1644511149
transform 1 0 2300 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_20
timestamp 1644511149
transform 1 0 2944 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_32
timestamp 1644511149
transform 1 0 4048 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_44
timestamp 1644511149
transform 1 0 5152 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_125
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_137
timestamp 1644511149
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_149
timestamp 1644511149
transform 1 0 14812 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_162
timestamp 1644511149
transform 1 0 16008 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_186
timestamp 1644511149
transform 1 0 18216 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_198
timestamp 1644511149
transform 1 0 19320 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_206
timestamp 1644511149
transform 1 0 20056 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1644511149
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1644511149
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_233
timestamp 1644511149
transform 1 0 22540 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_243
timestamp 1644511149
transform 1 0 23460 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_251
timestamp 1644511149
transform 1 0 24196 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_263
timestamp 1644511149
transform 1 0 25300 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_276
timestamp 1644511149
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_292
timestamp 1644511149
transform 1 0 27968 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_300
timestamp 1644511149
transform 1 0 28704 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_317
timestamp 1644511149
transform 1 0 30268 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_323
timestamp 1644511149
transform 1 0 30820 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_332
timestamp 1644511149
transform 1 0 31648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_342
timestamp 1644511149
transform 1 0 32568 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_354
timestamp 1644511149
transform 1 0 33672 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_373
timestamp 1644511149
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1644511149
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1644511149
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_400
timestamp 1644511149
transform 1 0 37904 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_409
timestamp 1644511149
transform 1 0 38732 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_421
timestamp 1644511149
transform 1 0 39836 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_433
timestamp 1644511149
transform 1 0 40940 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_440
timestamp 1644511149
transform 1 0 41584 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_465
timestamp 1644511149
transform 1 0 43884 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_477
timestamp 1644511149
transform 1 0 44988 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_494
timestamp 1644511149
transform 1 0 46552 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_502
timestamp 1644511149
transform 1 0 47288 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_508
timestamp 1644511149
transform 1 0 47840 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_24
timestamp 1644511149
transform 1 0 3312 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_121
timestamp 1644511149
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1644511149
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_153
timestamp 1644511149
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_181
timestamp 1644511149
transform 1 0 17756 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_190
timestamp 1644511149
transform 1 0 18584 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_214
timestamp 1644511149
transform 1 0 20792 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_232
timestamp 1644511149
transform 1 0 22448 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1644511149
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1644511149
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_259
timestamp 1644511149
transform 1 0 24932 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_273
timestamp 1644511149
transform 1 0 26220 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_282
timestamp 1644511149
transform 1 0 27048 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_302
timestamp 1644511149
transform 1 0 28888 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_321
timestamp 1644511149
transform 1 0 30636 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_342
timestamp 1644511149
transform 1 0 32568 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_30_358
timestamp 1644511149
transform 1 0 34040 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_382
timestamp 1644511149
transform 1 0 36248 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_394
timestamp 1644511149
transform 1 0 37352 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_404
timestamp 1644511149
transform 1 0 38272 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_415
timestamp 1644511149
transform 1 0 39284 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1644511149
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_421
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_430
timestamp 1644511149
transform 1 0 40664 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_441
timestamp 1644511149
transform 1 0 41676 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_461
timestamp 1644511149
transform 1 0 43516 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_472
timestamp 1644511149
transform 1 0 44528 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_485
timestamp 1644511149
transform 1 0 45724 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_512
timestamp 1644511149
transform 1 0 48208 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_8
timestamp 1644511149
transform 1 0 1840 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1644511149
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1644511149
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1644511149
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1644511149
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1644511149
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_125
timestamp 1644511149
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_137
timestamp 1644511149
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_149
timestamp 1644511149
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1644511149
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1644511149
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_173
timestamp 1644511149
transform 1 0 17020 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_179
timestamp 1644511149
transform 1 0 17572 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_191
timestamp 1644511149
transform 1 0 18676 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_206
timestamp 1644511149
transform 1 0 20056 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_218
timestamp 1644511149
transform 1 0 21160 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_231
timestamp 1644511149
transform 1 0 22356 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_244
timestamp 1644511149
transform 1 0 23552 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_256
timestamp 1644511149
transform 1 0 24656 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_260
timestamp 1644511149
transform 1 0 25024 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_270
timestamp 1644511149
transform 1 0 25944 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1644511149
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_285
timestamp 1644511149
transform 1 0 27324 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_297
timestamp 1644511149
transform 1 0 28428 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_303
timestamp 1644511149
transform 1 0 28980 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_308
timestamp 1644511149
transform 1 0 29440 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_320
timestamp 1644511149
transform 1 0 30544 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_326
timestamp 1644511149
transform 1 0 31096 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_334
timestamp 1644511149
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_337
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_345
timestamp 1644511149
transform 1 0 32844 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_356
timestamp 1644511149
transform 1 0 33856 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_365
timestamp 1644511149
transform 1 0 34684 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_377
timestamp 1644511149
transform 1 0 35788 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_389
timestamp 1644511149
transform 1 0 36892 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_397
timestamp 1644511149
transform 1 0 37628 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_409
timestamp 1644511149
transform 1 0 38732 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_417
timestamp 1644511149
transform 1 0 39468 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_430
timestamp 1644511149
transform 1 0 40664 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1644511149
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1644511149
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_452
timestamp 1644511149
transform 1 0 42688 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_466
timestamp 1644511149
transform 1 0 43976 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_488
timestamp 1644511149
transform 1 0 46000 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_496
timestamp 1644511149
transform 1 0 46736 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_500
timestamp 1644511149
transform 1 0 47104 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_505
timestamp 1644511149
transform 1 0 47564 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_512
timestamp 1644511149
transform 1 0 48208 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1644511149
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_109
timestamp 1644511149
transform 1 0 11132 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_115
timestamp 1644511149
transform 1 0 11684 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_119
timestamp 1644511149
transform 1 0 12052 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_131
timestamp 1644511149
transform 1 0 13156 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1644511149
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_153
timestamp 1644511149
transform 1 0 15180 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_175
timestamp 1644511149
transform 1 0 17204 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_191
timestamp 1644511149
transform 1 0 18676 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1644511149
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_200
timestamp 1644511149
transform 1 0 19504 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_228
timestamp 1644511149
transform 1 0 22080 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_232
timestamp 1644511149
transform 1 0 22448 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_239
timestamp 1644511149
transform 1 0 23092 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1644511149
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_265
timestamp 1644511149
transform 1 0 25484 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_270
timestamp 1644511149
transform 1 0 25944 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_278
timestamp 1644511149
transform 1 0 26680 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_290
timestamp 1644511149
transform 1 0 27784 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_296
timestamp 1644511149
transform 1 0 28336 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1644511149
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1644511149
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_320
timestamp 1644511149
transform 1 0 30544 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_328
timestamp 1644511149
transform 1 0 31280 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_334
timestamp 1644511149
transform 1 0 31832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_340
timestamp 1644511149
transform 1 0 32384 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_352
timestamp 1644511149
transform 1 0 33488 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_385
timestamp 1644511149
transform 1 0 36524 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_395
timestamp 1644511149
transform 1 0 37444 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_406
timestamp 1644511149
transform 1 0 38456 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_418
timestamp 1644511149
transform 1 0 39560 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_421
timestamp 1644511149
transform 1 0 39836 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_429
timestamp 1644511149
transform 1 0 40572 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_437
timestamp 1644511149
transform 1 0 41308 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_446
timestamp 1644511149
transform 1 0 42136 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_458
timestamp 1644511149
transform 1 0 43240 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_470
timestamp 1644511149
transform 1 0 44344 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_477
timestamp 1644511149
transform 1 0 44988 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_483
timestamp 1644511149
transform 1 0 45540 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_512
timestamp 1644511149
transform 1 0 48208 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1644511149
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_136
timestamp 1644511149
transform 1 0 13616 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_151
timestamp 1644511149
transform 1 0 14996 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_164
timestamp 1644511149
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_173
timestamp 1644511149
transform 1 0 17020 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_181
timestamp 1644511149
transform 1 0 17756 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_191
timestamp 1644511149
transform 1 0 18676 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_195
timestamp 1644511149
transform 1 0 19044 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_206
timestamp 1644511149
transform 1 0 20056 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_218
timestamp 1644511149
transform 1 0 21160 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_233
timestamp 1644511149
transform 1 0 22540 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_242
timestamp 1644511149
transform 1 0 23368 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_252
timestamp 1644511149
transform 1 0 24288 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_263
timestamp 1644511149
transform 1 0 25300 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_275
timestamp 1644511149
transform 1 0 26404 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1644511149
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_293
timestamp 1644511149
transform 1 0 28060 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_303
timestamp 1644511149
transform 1 0 28980 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_311
timestamp 1644511149
transform 1 0 29716 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_321
timestamp 1644511149
transform 1 0 30636 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_332
timestamp 1644511149
transform 1 0 31648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_358
timestamp 1644511149
transform 1 0 34040 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_370
timestamp 1644511149
transform 1 0 35144 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_388
timestamp 1644511149
transform 1 0 36800 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_400
timestamp 1644511149
transform 1 0 37904 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_407
timestamp 1644511149
transform 1 0 38548 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_419
timestamp 1644511149
transform 1 0 39652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_427
timestamp 1644511149
transform 1 0 40388 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1644511149
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1644511149
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_449
timestamp 1644511149
transform 1 0 42412 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_457
timestamp 1644511149
transform 1 0 43148 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_461
timestamp 1644511149
transform 1 0 43516 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_469
timestamp 1644511149
transform 1 0 44252 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_479
timestamp 1644511149
transform 1 0 45172 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_488
timestamp 1644511149
transform 1 0 46000 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_496
timestamp 1644511149
transform 1 0 46736 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_500
timestamp 1644511149
transform 1 0 47104 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_508
timestamp 1644511149
transform 1 0 47840 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_109
timestamp 1644511149
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_121
timestamp 1644511149
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1644511149
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1644511149
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_158
timestamp 1644511149
transform 1 0 15640 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_183
timestamp 1644511149
transform 1 0 17940 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_192
timestamp 1644511149
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_205
timestamp 1644511149
transform 1 0 19964 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_213
timestamp 1644511149
transform 1 0 20700 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_220
timestamp 1644511149
transform 1 0 21344 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_232
timestamp 1644511149
transform 1 0 22448 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1644511149
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1644511149
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_256
timestamp 1644511149
transform 1 0 24656 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_268
timestamp 1644511149
transform 1 0 25760 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_277
timestamp 1644511149
transform 1 0 26588 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_286
timestamp 1644511149
transform 1 0 27416 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_294
timestamp 1644511149
transform 1 0 28152 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_300
timestamp 1644511149
transform 1 0 28704 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_325
timestamp 1644511149
transform 1 0 31004 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_339
timestamp 1644511149
transform 1 0 32292 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_343
timestamp 1644511149
transform 1 0 32660 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_360
timestamp 1644511149
transform 1 0 34224 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_370
timestamp 1644511149
transform 1 0 35144 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_382
timestamp 1644511149
transform 1 0 36248 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_403
timestamp 1644511149
transform 1 0 38180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_415
timestamp 1644511149
transform 1 0 39284 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1644511149
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_437
timestamp 1644511149
transform 1 0 41308 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_444
timestamp 1644511149
transform 1 0 41952 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_450
timestamp 1644511149
transform 1 0 42504 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_461
timestamp 1644511149
transform 1 0 43516 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_472
timestamp 1644511149
transform 1 0 44528 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_485
timestamp 1644511149
transform 1 0 45724 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_512
timestamp 1644511149
transform 1 0 48208 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_23
timestamp 1644511149
transform 1 0 3220 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_45
timestamp 1644511149
transform 1 0 5244 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp 1644511149
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_137
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_141
timestamp 1644511149
transform 1 0 14076 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_147
timestamp 1644511149
transform 1 0 14628 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_164
timestamp 1644511149
transform 1 0 16192 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_193
timestamp 1644511149
transform 1 0 18860 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_213
timestamp 1644511149
transform 1 0 20700 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_221
timestamp 1644511149
transform 1 0 21436 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_241
timestamp 1644511149
transform 1 0 23276 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_251
timestamp 1644511149
transform 1 0 24196 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_259
timestamp 1644511149
transform 1 0 24932 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_276
timestamp 1644511149
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_301
timestamp 1644511149
transform 1 0 28796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_310
timestamp 1644511149
transform 1 0 29624 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_314
timestamp 1644511149
transform 1 0 29992 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_332
timestamp 1644511149
transform 1 0 31648 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_340
timestamp 1644511149
transform 1 0 32384 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_352
timestamp 1644511149
transform 1 0 33488 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_372
timestamp 1644511149
transform 1 0 35328 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_384
timestamp 1644511149
transform 1 0 36432 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_402
timestamp 1644511149
transform 1 0 38088 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_410
timestamp 1644511149
transform 1 0 38824 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_422
timestamp 1644511149
transform 1 0 39928 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_428
timestamp 1644511149
transform 1 0 40480 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_436
timestamp 1644511149
transform 1 0 41216 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_449
timestamp 1644511149
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_477
timestamp 1644511149
transform 1 0 44988 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_481
timestamp 1644511149
transform 1 0 45356 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_498
timestamp 1644511149
transform 1 0 46920 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_508
timestamp 1644511149
transform 1 0 47840 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_24
timestamp 1644511149
transform 1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_50
timestamp 1644511149
transform 1 0 5704 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_62
timestamp 1644511149
transform 1 0 6808 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_74
timestamp 1644511149
transform 1 0 7912 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1644511149
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_109
timestamp 1644511149
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_121
timestamp 1644511149
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1644511149
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_162
timestamp 1644511149
transform 1 0 16008 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_170
timestamp 1644511149
transform 1 0 16744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_187
timestamp 1644511149
transform 1 0 18308 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1644511149
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_202
timestamp 1644511149
transform 1 0 19688 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_214
timestamp 1644511149
transform 1 0 20792 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_226
timestamp 1644511149
transform 1 0 21896 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_238
timestamp 1644511149
transform 1 0 23000 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1644511149
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_272
timestamp 1644511149
transform 1 0 26128 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_280
timestamp 1644511149
transform 1 0 26864 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_289
timestamp 1644511149
transform 1 0 27692 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_293
timestamp 1644511149
transform 1 0 28060 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_304
timestamp 1644511149
transform 1 0 29072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_317
timestamp 1644511149
transform 1 0 30268 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_339
timestamp 1644511149
transform 1 0 32292 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_360
timestamp 1644511149
transform 1 0 34224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_377
timestamp 1644511149
transform 1 0 35788 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_384
timestamp 1644511149
transform 1 0 36432 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_398
timestamp 1644511149
transform 1 0 37720 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_410
timestamp 1644511149
transform 1 0 38824 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_418
timestamp 1644511149
transform 1 0 39560 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_421
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_425
timestamp 1644511149
transform 1 0 40204 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_430
timestamp 1644511149
transform 1 0 40664 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_434
timestamp 1644511149
transform 1 0 41032 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_438
timestamp 1644511149
transform 1 0 41400 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_442
timestamp 1644511149
transform 1 0 41768 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_448
timestamp 1644511149
transform 1 0 42320 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_454
timestamp 1644511149
transform 1 0 42872 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_463
timestamp 1644511149
transform 1 0 43700 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1644511149
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_477
timestamp 1644511149
transform 1 0 44988 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_494
timestamp 1644511149
transform 1 0 46552 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_506
timestamp 1644511149
transform 1 0 47656 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_512
timestamp 1644511149
transform 1 0 48208 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_11
timestamp 1644511149
transform 1 0 2116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_23
timestamp 1644511149
transform 1 0 3220 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_28
timestamp 1644511149
transform 1 0 3680 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_40
timestamp 1644511149
transform 1 0 4784 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_52
timestamp 1644511149
transform 1 0 5888 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_125
timestamp 1644511149
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_137
timestamp 1644511149
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_149
timestamp 1644511149
transform 1 0 14812 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_164
timestamp 1644511149
transform 1 0 16192 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_173
timestamp 1644511149
transform 1 0 17020 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_182
timestamp 1644511149
transform 1 0 17848 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_194
timestamp 1644511149
transform 1 0 18952 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_200
timestamp 1644511149
transform 1 0 19504 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_207
timestamp 1644511149
transform 1 0 20148 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_219
timestamp 1644511149
transform 1 0 21252 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1644511149
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_237
timestamp 1644511149
transform 1 0 22908 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_244
timestamp 1644511149
transform 1 0 23552 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_252
timestamp 1644511149
transform 1 0 24288 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_263
timestamp 1644511149
transform 1 0 25300 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_275
timestamp 1644511149
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1644511149
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_285
timestamp 1644511149
transform 1 0 27324 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_291
timestamp 1644511149
transform 1 0 27876 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_304
timestamp 1644511149
transform 1 0 29072 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_311
timestamp 1644511149
transform 1 0 29716 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_323
timestamp 1644511149
transform 1 0 30820 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_332
timestamp 1644511149
transform 1 0 31648 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_346
timestamp 1644511149
transform 1 0 32936 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_358
timestamp 1644511149
transform 1 0 34040 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_370
timestamp 1644511149
transform 1 0 35144 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_376
timestamp 1644511149
transform 1 0 35696 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_382
timestamp 1644511149
transform 1 0 36248 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_390
timestamp 1644511149
transform 1 0 36984 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_398
timestamp 1644511149
transform 1 0 37720 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_406
timestamp 1644511149
transform 1 0 38456 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_418
timestamp 1644511149
transform 1 0 39560 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_431
timestamp 1644511149
transform 1 0 40756 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_444
timestamp 1644511149
transform 1 0 41952 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_455
timestamp 1644511149
transform 1 0 42964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_467
timestamp 1644511149
transform 1 0 44068 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_479
timestamp 1644511149
transform 1 0 45172 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_485
timestamp 1644511149
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1644511149
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1644511149
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_505
timestamp 1644511149
transform 1 0 47564 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_512
timestamp 1644511149
transform 1 0 48208 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_121
timestamp 1644511149
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1644511149
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_153
timestamp 1644511149
transform 1 0 15180 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_161
timestamp 1644511149
transform 1 0 15916 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_180
timestamp 1644511149
transform 1 0 17664 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_187
timestamp 1644511149
transform 1 0 18308 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1644511149
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_203
timestamp 1644511149
transform 1 0 19780 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_210
timestamp 1644511149
transform 1 0 20424 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_222
timestamp 1644511149
transform 1 0 21528 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_234
timestamp 1644511149
transform 1 0 22632 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_240
timestamp 1644511149
transform 1 0 23184 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_246
timestamp 1644511149
transform 1 0 23736 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_265
timestamp 1644511149
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_277
timestamp 1644511149
transform 1 0 26588 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_285
timestamp 1644511149
transform 1 0 27324 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_290
timestamp 1644511149
transform 1 0 27784 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_299
timestamp 1644511149
transform 1 0 28612 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1644511149
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_317
timestamp 1644511149
transform 1 0 30268 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_328
timestamp 1644511149
transform 1 0 31280 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_336
timestamp 1644511149
transform 1 0 32016 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_342
timestamp 1644511149
transform 1 0 32568 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_354
timestamp 1644511149
transform 1 0 33672 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_362
timestamp 1644511149
transform 1 0 34408 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_372
timestamp 1644511149
transform 1 0 35328 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_382
timestamp 1644511149
transform 1 0 36248 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_390
timestamp 1644511149
transform 1 0 36984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_397
timestamp 1644511149
transform 1 0 37628 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_410
timestamp 1644511149
transform 1 0 38824 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_418
timestamp 1644511149
transform 1 0 39560 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_426
timestamp 1644511149
transform 1 0 40296 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_434
timestamp 1644511149
transform 1 0 41032 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_444
timestamp 1644511149
transform 1 0 41952 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_458
timestamp 1644511149
transform 1 0 43240 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_472
timestamp 1644511149
transform 1 0 44528 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_477
timestamp 1644511149
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_489
timestamp 1644511149
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_501
timestamp 1644511149
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_513
timestamp 1644511149
transform 1 0 48300 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_28
timestamp 1644511149
transform 1 0 3680 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_40
timestamp 1644511149
transform 1 0 4784 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_52
timestamp 1644511149
transform 1 0 5888 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_137
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_149
timestamp 1644511149
transform 1 0 14812 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_157
timestamp 1644511149
transform 1 0 15548 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_164
timestamp 1644511149
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_39_193
timestamp 1644511149
transform 1 0 18860 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_201
timestamp 1644511149
transform 1 0 19596 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_208
timestamp 1644511149
transform 1 0 20240 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_218
timestamp 1644511149
transform 1 0 21160 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_248
timestamp 1644511149
transform 1 0 23920 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_255
timestamp 1644511149
transform 1 0 24564 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_267
timestamp 1644511149
transform 1 0 25668 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_276
timestamp 1644511149
transform 1 0 26496 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_289
timestamp 1644511149
transform 1 0 27692 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_301
timestamp 1644511149
transform 1 0 28796 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_305
timestamp 1644511149
transform 1 0 29164 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_312
timestamp 1644511149
transform 1 0 29808 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_320
timestamp 1644511149
transform 1 0 30544 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_332
timestamp 1644511149
transform 1 0 31648 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_343
timestamp 1644511149
transform 1 0 32660 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_349
timestamp 1644511149
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_361
timestamp 1644511149
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_373
timestamp 1644511149
transform 1 0 35420 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_379
timestamp 1644511149
transform 1 0 35972 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_387
timestamp 1644511149
transform 1 0 36708 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1644511149
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_398
timestamp 1644511149
transform 1 0 37720 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_415
timestamp 1644511149
transform 1 0 39284 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_425
timestamp 1644511149
transform 1 0 40204 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_434
timestamp 1644511149
transform 1 0 41032 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_443
timestamp 1644511149
transform 1 0 41860 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1644511149
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_449
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_453
timestamp 1644511149
transform 1 0 42780 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_470
timestamp 1644511149
transform 1 0 44344 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_482
timestamp 1644511149
transform 1 0 45448 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_494
timestamp 1644511149
transform 1 0 46552 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_502
timestamp 1644511149
transform 1 0 47288 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_505
timestamp 1644511149
transform 1 0 47564 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_512
timestamp 1644511149
transform 1 0 48208 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_13
timestamp 1644511149
transform 1 0 2300 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_20
timestamp 1644511149
transform 1 0 2944 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_121
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1644511149
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_153
timestamp 1644511149
transform 1 0 15180 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_160
timestamp 1644511149
transform 1 0 15824 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_167
timestamp 1644511149
transform 1 0 16468 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1644511149
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_201
timestamp 1644511149
transform 1 0 19596 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_208
timestamp 1644511149
transform 1 0 20240 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_218
timestamp 1644511149
transform 1 0 21160 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_40_242
timestamp 1644511149
transform 1 0 23368 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1644511149
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_257
timestamp 1644511149
transform 1 0 24748 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_279
timestamp 1644511149
transform 1 0 26772 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_292
timestamp 1644511149
transform 1 0 27968 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_304
timestamp 1644511149
transform 1 0 29072 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_317
timestamp 1644511149
transform 1 0 30268 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_328
timestamp 1644511149
transform 1 0 31280 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_340
timestamp 1644511149
transform 1 0 32384 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_360
timestamp 1644511149
transform 1 0 34224 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_381
timestamp 1644511149
transform 1 0 36156 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_389
timestamp 1644511149
transform 1 0 36892 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_395
timestamp 1644511149
transform 1 0 37444 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_405
timestamp 1644511149
transform 1 0 38364 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_415
timestamp 1644511149
transform 1 0 39284 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1644511149
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_421
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_429
timestamp 1644511149
transform 1 0 40572 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_436
timestamp 1644511149
transform 1 0 41216 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_445
timestamp 1644511149
transform 1 0 42044 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_453
timestamp 1644511149
transform 1 0 42780 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_460
timestamp 1644511149
transform 1 0 43424 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_467
timestamp 1644511149
transform 1 0 44068 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1644511149
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_477
timestamp 1644511149
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_489
timestamp 1644511149
transform 1 0 46092 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_512
timestamp 1644511149
transform 1 0 48208 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_14
timestamp 1644511149
transform 1 0 2392 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_26
timestamp 1644511149
transform 1 0 3496 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_38
timestamp 1644511149
transform 1 0 4600 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_50
timestamp 1644511149
transform 1 0 5704 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_137
timestamp 1644511149
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_149
timestamp 1644511149
transform 1 0 14812 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_157
timestamp 1644511149
transform 1 0 15548 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_164
timestamp 1644511149
transform 1 0 16192 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_185
timestamp 1644511149
transform 1 0 18124 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_191
timestamp 1644511149
transform 1 0 18676 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_198
timestamp 1644511149
transform 1 0 19320 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_208
timestamp 1644511149
transform 1 0 20240 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_218
timestamp 1644511149
transform 1 0 21160 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_239
timestamp 1644511149
transform 1 0 23092 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_246
timestamp 1644511149
transform 1 0 23736 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_258
timestamp 1644511149
transform 1 0 24840 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_276
timestamp 1644511149
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_289
timestamp 1644511149
transform 1 0 27692 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_298
timestamp 1644511149
transform 1 0 28520 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_312
timestamp 1644511149
transform 1 0 29808 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_332
timestamp 1644511149
transform 1 0 31648 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_345
timestamp 1644511149
transform 1 0 32844 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_365
timestamp 1644511149
transform 1 0 34684 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_377
timestamp 1644511149
transform 1 0 35788 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_389
timestamp 1644511149
transform 1 0 36892 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_433
timestamp 1644511149
transform 1 0 40940 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_444
timestamp 1644511149
transform 1 0 41952 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_465
timestamp 1644511149
transform 1 0 43884 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_477
timestamp 1644511149
transform 1 0 44988 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_489
timestamp 1644511149
transform 1 0 46092 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_500
timestamp 1644511149
transform 1 0 47104 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_505
timestamp 1644511149
transform 1 0 47564 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_512
timestamp 1644511149
transform 1 0 48208 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1644511149
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_97
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_109
timestamp 1644511149
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_121
timestamp 1644511149
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1644511149
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1644511149
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_149
timestamp 1644511149
transform 1 0 14812 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_163
timestamp 1644511149
transform 1 0 16100 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_183
timestamp 1644511149
transform 1 0 17940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1644511149
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_201
timestamp 1644511149
transform 1 0 19596 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_208
timestamp 1644511149
transform 1 0 20240 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_212
timestamp 1644511149
transform 1 0 20608 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_219
timestamp 1644511149
transform 1 0 21252 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_231
timestamp 1644511149
transform 1 0 22356 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_243
timestamp 1644511149
transform 1 0 23460 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1644511149
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_259
timestamp 1644511149
transform 1 0 24932 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_268
timestamp 1644511149
transform 1 0 25760 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_280
timestamp 1644511149
transform 1 0 26864 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_296
timestamp 1644511149
transform 1 0 28336 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_304
timestamp 1644511149
transform 1 0 29072 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_323
timestamp 1644511149
transform 1 0 30820 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_332
timestamp 1644511149
transform 1 0 31648 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_344
timestamp 1644511149
transform 1 0 32752 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_356
timestamp 1644511149
transform 1 0 33856 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_378
timestamp 1644511149
transform 1 0 35880 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_398
timestamp 1644511149
transform 1 0 37720 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_410
timestamp 1644511149
transform 1 0 38824 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_418
timestamp 1644511149
transform 1 0 39560 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_421
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_427
timestamp 1644511149
transform 1 0 40388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_439
timestamp 1644511149
transform 1 0 41492 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_451
timestamp 1644511149
transform 1 0 42596 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_463
timestamp 1644511149
transform 1 0 43700 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1644511149
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_477
timestamp 1644511149
transform 1 0 44988 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_483
timestamp 1644511149
transform 1 0 45540 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_487
timestamp 1644511149
transform 1 0 45908 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_499
timestamp 1644511149
transform 1 0 47012 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_502
timestamp 1644511149
transform 1 0 47288 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_511
timestamp 1644511149
transform 1 0 48116 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_515
timestamp 1644511149
transform 1 0 48484 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_13
timestamp 1644511149
transform 1 0 2300 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_20
timestamp 1644511149
transform 1 0 2944 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_32
timestamp 1644511149
transform 1 0 4048 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_44
timestamp 1644511149
transform 1 0 5152 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_125
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_137
timestamp 1644511149
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_149
timestamp 1644511149
transform 1 0 14812 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_155
timestamp 1644511149
transform 1 0 15364 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_158
timestamp 1644511149
transform 1 0 15640 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1644511149
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_185
timestamp 1644511149
transform 1 0 18124 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_197
timestamp 1644511149
transform 1 0 19228 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_214
timestamp 1644511149
transform 1 0 20792 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1644511149
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_237
timestamp 1644511149
transform 1 0 22908 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_241
timestamp 1644511149
transform 1 0 23276 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_247
timestamp 1644511149
transform 1 0 23828 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_259
timestamp 1644511149
transform 1 0 24932 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_271
timestamp 1644511149
transform 1 0 26036 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1644511149
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_293
timestamp 1644511149
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_305
timestamp 1644511149
transform 1 0 29164 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_309
timestamp 1644511149
transform 1 0 29532 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_315
timestamp 1644511149
transform 1 0 30084 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_323
timestamp 1644511149
transform 1 0 30820 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1644511149
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_345
timestamp 1644511149
transform 1 0 32844 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_354
timestamp 1644511149
transform 1 0 33672 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_366
timestamp 1644511149
transform 1 0 34776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_371
timestamp 1644511149
transform 1 0 35236 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_379
timestamp 1644511149
transform 1 0 35972 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_388
timestamp 1644511149
transform 1 0 36800 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_405
timestamp 1644511149
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_417
timestamp 1644511149
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_429
timestamp 1644511149
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1644511149
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1644511149
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_449
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_461
timestamp 1644511149
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_473
timestamp 1644511149
transform 1 0 44620 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_500
timestamp 1644511149
transform 1 0 47104 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_508
timestamp 1644511149
transform 1 0 47840 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_24
timestamp 1644511149
transform 1 0 3312 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_121
timestamp 1644511149
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_153
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_157
timestamp 1644511149
transform 1 0 15548 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_179
timestamp 1644511149
transform 1 0 17572 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_185
timestamp 1644511149
transform 1 0 18124 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_191
timestamp 1644511149
transform 1 0 18676 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1644511149
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_205
timestamp 1644511149
transform 1 0 19964 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_44_215
timestamp 1644511149
transform 1 0 20884 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_227
timestamp 1644511149
transform 1 0 21988 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_231
timestamp 1644511149
transform 1 0 22356 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_248
timestamp 1644511149
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_261
timestamp 1644511149
transform 1 0 25116 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_273
timestamp 1644511149
transform 1 0 26220 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_285
timestamp 1644511149
transform 1 0 27324 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_297
timestamp 1644511149
transform 1 0 28428 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_305
timestamp 1644511149
transform 1 0 29164 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_315
timestamp 1644511149
transform 1 0 30084 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_333
timestamp 1644511149
transform 1 0 31740 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_341
timestamp 1644511149
transform 1 0 32476 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_353
timestamp 1644511149
transform 1 0 33580 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_359
timestamp 1644511149
transform 1 0 34132 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1644511149
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_373
timestamp 1644511149
transform 1 0 35420 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_381
timestamp 1644511149
transform 1 0 36156 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_400
timestamp 1644511149
transform 1 0 37904 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_412
timestamp 1644511149
transform 1 0 39008 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_416
timestamp 1644511149
transform 1 0 39376 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_442
timestamp 1644511149
transform 1 0 41768 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_454
timestamp 1644511149
transform 1 0 42872 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_466
timestamp 1644511149
transform 1 0 43976 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_474
timestamp 1644511149
transform 1 0 44712 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_477
timestamp 1644511149
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_489
timestamp 1644511149
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_501
timestamp 1644511149
transform 1 0 47196 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_512
timestamp 1644511149
transform 1 0 48208 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_28
timestamp 1644511149
transform 1 0 3680 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_40
timestamp 1644511149
transform 1 0 4784 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_52
timestamp 1644511149
transform 1 0 5888 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_137
timestamp 1644511149
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_149
timestamp 1644511149
transform 1 0 14812 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_157
timestamp 1644511149
transform 1 0 15548 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_162
timestamp 1644511149
transform 1 0 16008 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_181
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_185
timestamp 1644511149
transform 1 0 18124 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_207
timestamp 1644511149
transform 1 0 20148 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_220
timestamp 1644511149
transform 1 0 21344 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_241
timestamp 1644511149
transform 1 0 23276 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_45_263
timestamp 1644511149
transform 1 0 25300 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1644511149
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1644511149
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_285
timestamp 1644511149
transform 1 0 27324 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_291
timestamp 1644511149
transform 1 0 27876 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_298
timestamp 1644511149
transform 1 0 28520 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_310
timestamp 1644511149
transform 1 0 29624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_319
timestamp 1644511149
transform 1 0 30452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_331
timestamp 1644511149
transform 1 0 31556 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1644511149
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_366
timestamp 1644511149
transform 1 0 34776 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_370
timestamp 1644511149
transform 1 0 35144 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_376
timestamp 1644511149
transform 1 0 35696 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_388
timestamp 1644511149
transform 1 0 36800 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_401
timestamp 1644511149
transform 1 0 37996 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_410
timestamp 1644511149
transform 1 0 38824 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_435
timestamp 1644511149
transform 1 0 41124 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1644511149
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_461
timestamp 1644511149
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_473
timestamp 1644511149
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_485
timestamp 1644511149
transform 1 0 45724 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_45_496
timestamp 1644511149
transform 1 0 46736 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_45_505
timestamp 1644511149
transform 1 0 47564 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_513
timestamp 1644511149
transform 1 0 48300 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_8
timestamp 1644511149
transform 1 0 1840 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_22
timestamp 1644511149
transform 1 0 3128 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_121
timestamp 1644511149
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1644511149
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_153
timestamp 1644511149
transform 1 0 15180 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_177
timestamp 1644511149
transform 1 0 17388 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_183
timestamp 1644511149
transform 1 0 17940 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1644511149
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_216
timestamp 1644511149
transform 1 0 20976 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_228
timestamp 1644511149
transform 1 0 22080 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_236
timestamp 1644511149
transform 1 0 22816 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_248
timestamp 1644511149
transform 1 0 23920 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_258
timestamp 1644511149
transform 1 0 24840 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_266
timestamp 1644511149
transform 1 0 25576 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_275
timestamp 1644511149
transform 1 0 26404 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_295
timestamp 1644511149
transform 1 0 28244 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_303
timestamp 1644511149
transform 1 0 28980 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1644511149
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_313
timestamp 1644511149
transform 1 0 29900 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_325
timestamp 1644511149
transform 1 0 31004 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_343
timestamp 1644511149
transform 1 0 32660 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_351
timestamp 1644511149
transform 1 0 33396 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_359
timestamp 1644511149
transform 1 0 34132 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1644511149
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_369
timestamp 1644511149
transform 1 0 35052 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_375
timestamp 1644511149
transform 1 0 35604 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_396
timestamp 1644511149
transform 1 0 37536 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_408
timestamp 1644511149
transform 1 0 38640 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_412
timestamp 1644511149
transform 1 0 39008 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_416
timestamp 1644511149
transform 1 0 39376 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_442
timestamp 1644511149
transform 1 0 41768 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_454
timestamp 1644511149
transform 1 0 42872 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_466
timestamp 1644511149
transform 1 0 43976 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_474
timestamp 1644511149
transform 1 0 44712 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_477
timestamp 1644511149
transform 1 0 44988 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_481
timestamp 1644511149
transform 1 0 45356 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_485
timestamp 1644511149
transform 1 0 45724 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_512
timestamp 1644511149
transform 1 0 48208 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_11
timestamp 1644511149
transform 1 0 2116 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_128
timestamp 1644511149
transform 1 0 12880 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_140
timestamp 1644511149
transform 1 0 13984 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_152
timestamp 1644511149
transform 1 0 15088 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_164
timestamp 1644511149
transform 1 0 16192 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_175
timestamp 1644511149
transform 1 0 17204 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_192
timestamp 1644511149
transform 1 0 18768 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_204
timestamp 1644511149
transform 1 0 19872 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_213
timestamp 1644511149
transform 1 0 20700 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_221
timestamp 1644511149
transform 1 0 21436 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_229
timestamp 1644511149
transform 1 0 22172 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_238
timestamp 1644511149
transform 1 0 23000 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_250
timestamp 1644511149
transform 1 0 24104 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_258
timestamp 1644511149
transform 1 0 24840 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_276
timestamp 1644511149
transform 1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_293
timestamp 1644511149
transform 1 0 28060 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_303
timestamp 1644511149
transform 1 0 28980 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_47_327
timestamp 1644511149
transform 1 0 31188 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1644511149
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_340
timestamp 1644511149
transform 1 0 32384 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_352
timestamp 1644511149
transform 1 0 33488 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_363
timestamp 1644511149
transform 1 0 34500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_375
timestamp 1644511149
transform 1 0 35604 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_383
timestamp 1644511149
transform 1 0 36340 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_387
timestamp 1644511149
transform 1 0 36708 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1644511149
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_398
timestamp 1644511149
transform 1 0 37720 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_406
timestamp 1644511149
transform 1 0 38456 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_410
timestamp 1644511149
transform 1 0 38824 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_435
timestamp 1644511149
transform 1 0 41124 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1644511149
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_449
timestamp 1644511149
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_461
timestamp 1644511149
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_473
timestamp 1644511149
transform 1 0 44620 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_500
timestamp 1644511149
transform 1 0 47104 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_47_505
timestamp 1644511149
transform 1 0 47564 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_512
timestamp 1644511149
transform 1 0 48208 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_24
timestamp 1644511149
transform 1 0 3312 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1644511149
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_153
timestamp 1644511149
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_165
timestamp 1644511149
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_177
timestamp 1644511149
transform 1 0 17388 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_185
timestamp 1644511149
transform 1 0 18124 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_193
timestamp 1644511149
transform 1 0 18860 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_200
timestamp 1644511149
transform 1 0 19504 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_212
timestamp 1644511149
transform 1 0 20608 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_224
timestamp 1644511149
transform 1 0 21712 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_232
timestamp 1644511149
transform 1 0 22448 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_240
timestamp 1644511149
transform 1 0 23184 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_246
timestamp 1644511149
transform 1 0 23736 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_261
timestamp 1644511149
transform 1 0 25116 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_270
timestamp 1644511149
transform 1 0 25944 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_278
timestamp 1644511149
transform 1 0 26680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_284
timestamp 1644511149
transform 1 0 27232 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_293
timestamp 1644511149
transform 1 0 28060 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_303
timestamp 1644511149
transform 1 0 28980 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1644511149
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_321
timestamp 1644511149
transform 1 0 30636 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_329
timestamp 1644511149
transform 1 0 31372 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_339
timestamp 1644511149
transform 1 0 32292 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_48_348
timestamp 1644511149
transform 1 0 33120 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_360
timestamp 1644511149
transform 1 0 34224 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_372
timestamp 1644511149
transform 1 0 35328 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_405
timestamp 1644511149
transform 1 0 38364 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1644511149
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1644511149
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_421
timestamp 1644511149
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_433
timestamp 1644511149
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_445
timestamp 1644511149
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_457
timestamp 1644511149
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1644511149
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1644511149
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_477
timestamp 1644511149
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_489
timestamp 1644511149
transform 1 0 46092 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_512
timestamp 1644511149
transform 1 0 48208 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_7
timestamp 1644511149
transform 1 0 1748 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_11
timestamp 1644511149
transform 1 0 2116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_23
timestamp 1644511149
transform 1 0 3220 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_35
timestamp 1644511149
transform 1 0 4324 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_47
timestamp 1644511149
transform 1 0 5428 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_137
timestamp 1644511149
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_149
timestamp 1644511149
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1644511149
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1644511149
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_177
timestamp 1644511149
transform 1 0 17388 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_186
timestamp 1644511149
transform 1 0 18216 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_198
timestamp 1644511149
transform 1 0 19320 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_210
timestamp 1644511149
transform 1 0 20424 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_222
timestamp 1644511149
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_235
timestamp 1644511149
transform 1 0 22724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_247
timestamp 1644511149
transform 1 0 23828 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_251
timestamp 1644511149
transform 1 0 24196 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_260
timestamp 1644511149
transform 1 0 25024 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_272
timestamp 1644511149
transform 1 0 26128 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_289
timestamp 1644511149
transform 1 0 27692 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_49_302
timestamp 1644511149
transform 1 0 28888 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_310
timestamp 1644511149
transform 1 0 29624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_316
timestamp 1644511149
transform 1 0 30176 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_328
timestamp 1644511149
transform 1 0 31280 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_345
timestamp 1644511149
transform 1 0 32844 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_369
timestamp 1644511149
transform 1 0 35052 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_379
timestamp 1644511149
transform 1 0 35972 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_388
timestamp 1644511149
transform 1 0 36800 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_414
timestamp 1644511149
transform 1 0 39192 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_426
timestamp 1644511149
transform 1 0 40296 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_438
timestamp 1644511149
transform 1 0 41400 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_446
timestamp 1644511149
transform 1 0 42136 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_449
timestamp 1644511149
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_461
timestamp 1644511149
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_473
timestamp 1644511149
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_485
timestamp 1644511149
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1644511149
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1644511149
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_508
timestamp 1644511149
transform 1 0 47840 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_24
timestamp 1644511149
transform 1 0 3312 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_153
timestamp 1644511149
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_165
timestamp 1644511149
transform 1 0 16284 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_169
timestamp 1644511149
transform 1 0 16652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_186
timestamp 1644511149
transform 1 0 18216 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_194
timestamp 1644511149
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_205
timestamp 1644511149
transform 1 0 19964 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_223
timestamp 1644511149
transform 1 0 21620 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1644511149
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1644511149
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_275
timestamp 1644511149
transform 1 0 26404 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_283
timestamp 1644511149
transform 1 0 27140 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_289
timestamp 1644511149
transform 1 0 27692 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_299
timestamp 1644511149
transform 1 0 28612 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1644511149
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_319
timestamp 1644511149
transform 1 0 30452 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_327
timestamp 1644511149
transform 1 0 31188 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_335
timestamp 1644511149
transform 1 0 31924 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_340
timestamp 1644511149
transform 1 0 32384 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_360
timestamp 1644511149
transform 1 0 34224 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_370
timestamp 1644511149
transform 1 0 35144 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_382
timestamp 1644511149
transform 1 0 36248 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_390
timestamp 1644511149
transform 1 0 36984 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_409
timestamp 1644511149
transform 1 0 38732 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_417
timestamp 1644511149
transform 1 0 39468 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_421
timestamp 1644511149
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_433
timestamp 1644511149
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_445
timestamp 1644511149
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_457
timestamp 1644511149
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1644511149
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1644511149
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_477
timestamp 1644511149
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_489
timestamp 1644511149
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_501
timestamp 1644511149
transform 1 0 47196 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_507
timestamp 1644511149
transform 1 0 47748 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_515
timestamp 1644511149
transform 1 0 48484 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_7
timestamp 1644511149
transform 1 0 1748 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_14
timestamp 1644511149
transform 1 0 2392 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_26
timestamp 1644511149
transform 1 0 3496 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_38
timestamp 1644511149
transform 1 0 4600 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_50
timestamp 1644511149
transform 1 0 5704 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_149
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1644511149
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1644511149
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_177
timestamp 1644511149
transform 1 0 17388 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_194
timestamp 1644511149
transform 1 0 18952 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_207
timestamp 1644511149
transform 1 0 20148 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_220
timestamp 1644511149
transform 1 0 21344 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_230
timestamp 1644511149
transform 1 0 22264 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_51_245
timestamp 1644511149
transform 1 0 23644 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_253
timestamp 1644511149
transform 1 0 24380 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_261
timestamp 1644511149
transform 1 0 25116 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_269
timestamp 1644511149
transform 1 0 25852 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_277
timestamp 1644511149
transform 1 0 26588 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_289
timestamp 1644511149
transform 1 0 27692 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_297
timestamp 1644511149
transform 1 0 28428 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_306
timestamp 1644511149
transform 1 0 29256 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_312
timestamp 1644511149
transform 1 0 29808 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1644511149
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1644511149
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_349
timestamp 1644511149
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_361
timestamp 1644511149
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_373
timestamp 1644511149
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1644511149
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1644511149
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_397
timestamp 1644511149
transform 1 0 37628 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_409
timestamp 1644511149
transform 1 0 38732 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_421
timestamp 1644511149
transform 1 0 39836 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_433
timestamp 1644511149
transform 1 0 40940 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_445
timestamp 1644511149
transform 1 0 42044 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_449
timestamp 1644511149
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_461
timestamp 1644511149
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_473
timestamp 1644511149
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_485
timestamp 1644511149
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1644511149
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1644511149
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_505
timestamp 1644511149
transform 1 0 47564 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_512
timestamp 1644511149
transform 1 0 48208 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_7
timestamp 1644511149
transform 1 0 1748 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_11
timestamp 1644511149
transform 1 0 2116 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_23
timestamp 1644511149
transform 1 0 3220 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_165
timestamp 1644511149
transform 1 0 16284 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_184
timestamp 1644511149
transform 1 0 18032 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_202
timestamp 1644511149
transform 1 0 19688 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_210
timestamp 1644511149
transform 1 0 20424 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_219
timestamp 1644511149
transform 1 0 21252 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_232
timestamp 1644511149
transform 1 0 22448 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_240
timestamp 1644511149
transform 1 0 23184 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_269
timestamp 1644511149
transform 1 0 25852 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_281
timestamp 1644511149
transform 1 0 26956 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_287
timestamp 1644511149
transform 1 0 27508 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_304
timestamp 1644511149
transform 1 0 29072 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_329
timestamp 1644511149
transform 1 0 31372 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_341
timestamp 1644511149
transform 1 0 32476 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_353
timestamp 1644511149
transform 1 0 33580 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_361
timestamp 1644511149
transform 1 0 34316 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_373
timestamp 1644511149
transform 1 0 35420 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_380
timestamp 1644511149
transform 1 0 36064 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_393
timestamp 1644511149
transform 1 0 37260 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_399
timestamp 1644511149
transform 1 0 37812 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_403
timestamp 1644511149
transform 1 0 38180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_415
timestamp 1644511149
transform 1 0 39284 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1644511149
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_421
timestamp 1644511149
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_433
timestamp 1644511149
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_445
timestamp 1644511149
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_457
timestamp 1644511149
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1644511149
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1644511149
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_477
timestamp 1644511149
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_489
timestamp 1644511149
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_501
timestamp 1644511149
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_513
timestamp 1644511149
transform 1 0 48300 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_13
timestamp 1644511149
transform 1 0 2300 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_20
timestamp 1644511149
transform 1 0 2944 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_32
timestamp 1644511149
transform 1 0 4048 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_44
timestamp 1644511149
transform 1 0 5152 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_149
timestamp 1644511149
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1644511149
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_179
timestamp 1644511149
transform 1 0 17572 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_187
timestamp 1644511149
transform 1 0 18308 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_198
timestamp 1644511149
transform 1 0 19320 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_206
timestamp 1644511149
transform 1 0 20056 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_209
timestamp 1644511149
transform 1 0 20332 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_216
timestamp 1644511149
transform 1 0 20976 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_233
timestamp 1644511149
transform 1 0 22540 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_243
timestamp 1644511149
transform 1 0 23460 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_255
timestamp 1644511149
transform 1 0 24564 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_262
timestamp 1644511149
transform 1 0 25208 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_274
timestamp 1644511149
transform 1 0 26312 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_289
timestamp 1644511149
transform 1 0 27692 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_295
timestamp 1644511149
transform 1 0 28244 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_299
timestamp 1644511149
transform 1 0 28612 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_306
timestamp 1644511149
transform 1 0 29256 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_317
timestamp 1644511149
transform 1 0 30268 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_325
timestamp 1644511149
transform 1 0 31004 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_332
timestamp 1644511149
transform 1 0 31648 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_348
timestamp 1644511149
transform 1 0 33120 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_360
timestamp 1644511149
transform 1 0 34224 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_372
timestamp 1644511149
transform 1 0 35328 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_376
timestamp 1644511149
transform 1 0 35696 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_388
timestamp 1644511149
transform 1 0 36800 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_396
timestamp 1644511149
transform 1 0 37536 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_421
timestamp 1644511149
transform 1 0 39836 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_433
timestamp 1644511149
transform 1 0 40940 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_445
timestamp 1644511149
transform 1 0 42044 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_449
timestamp 1644511149
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_461
timestamp 1644511149
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_473
timestamp 1644511149
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_485
timestamp 1644511149
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1644511149
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1644511149
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_505
timestamp 1644511149
transform 1 0 47564 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_513
timestamp 1644511149
transform 1 0 48300 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_24
timestamp 1644511149
transform 1 0 3312 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_153
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_170
timestamp 1644511149
transform 1 0 16744 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_190
timestamp 1644511149
transform 1 0 18584 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_54_219
timestamp 1644511149
transform 1 0 21252 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_227
timestamp 1644511149
transform 1 0 21988 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_232
timestamp 1644511149
transform 1 0 22448 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_244
timestamp 1644511149
transform 1 0 23552 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_261
timestamp 1644511149
transform 1 0 25116 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_265
timestamp 1644511149
transform 1 0 25484 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_270
timestamp 1644511149
transform 1 0 25944 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_278
timestamp 1644511149
transform 1 0 26680 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_290
timestamp 1644511149
transform 1 0 27784 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_299
timestamp 1644511149
transform 1 0 28612 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1644511149
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_321
timestamp 1644511149
transform 1 0 30636 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_329
timestamp 1644511149
transform 1 0 31372 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_336
timestamp 1644511149
transform 1 0 32016 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_348
timestamp 1644511149
transform 1 0 33120 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_356
timestamp 1644511149
transform 1 0 33856 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_373
timestamp 1644511149
transform 1 0 35420 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_378
timestamp 1644511149
transform 1 0 35880 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_388
timestamp 1644511149
transform 1 0 36800 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1644511149
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1644511149
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_421
timestamp 1644511149
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_433
timestamp 1644511149
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_445
timestamp 1644511149
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_457
timestamp 1644511149
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1644511149
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1644511149
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_477
timestamp 1644511149
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_489
timestamp 1644511149
transform 1 0 46092 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_498
timestamp 1644511149
transform 1 0 46920 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_512
timestamp 1644511149
transform 1 0 48208 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_30
timestamp 1644511149
transform 1 0 3864 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_42
timestamp 1644511149
transform 1 0 4968 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_54
timestamp 1644511149
transform 1 0 6072 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_55_160
timestamp 1644511149
transform 1 0 15824 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_181
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_185
timestamp 1644511149
transform 1 0 18124 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_191
timestamp 1644511149
transform 1 0 18676 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_203
timestamp 1644511149
transform 1 0 19780 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_215
timestamp 1644511149
transform 1 0 20884 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1644511149
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_228
timestamp 1644511149
transform 1 0 22080 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_236
timestamp 1644511149
transform 1 0 22816 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_248
timestamp 1644511149
transform 1 0 23920 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_261
timestamp 1644511149
transform 1 0 25116 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_269
timestamp 1644511149
transform 1 0 25852 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_276
timestamp 1644511149
transform 1 0 26496 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_301
timestamp 1644511149
transform 1 0 28796 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_313
timestamp 1644511149
transform 1 0 29900 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_321
timestamp 1644511149
transform 1 0 30636 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_332
timestamp 1644511149
transform 1 0 31648 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_341
timestamp 1644511149
transform 1 0 32476 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_358
timestamp 1644511149
transform 1 0 34040 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_370
timestamp 1644511149
transform 1 0 35144 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_388
timestamp 1644511149
transform 1 0 36800 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_414
timestamp 1644511149
transform 1 0 39192 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_426
timestamp 1644511149
transform 1 0 40296 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_438
timestamp 1644511149
transform 1 0 41400 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_446
timestamp 1644511149
transform 1 0 42136 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_449
timestamp 1644511149
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_461
timestamp 1644511149
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_473
timestamp 1644511149
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_485
timestamp 1644511149
transform 1 0 45724 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_500
timestamp 1644511149
transform 1 0 47104 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_505
timestamp 1644511149
transform 1 0 47564 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_513
timestamp 1644511149
transform 1 0 48300 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_6
timestamp 1644511149
transform 1 0 1656 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_13
timestamp 1644511149
transform 1 0 2300 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_20
timestamp 1644511149
transform 1 0 2944 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_178
timestamp 1644511149
transform 1 0 17480 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_190
timestamp 1644511149
transform 1 0 18584 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_56_197
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_204
timestamp 1644511149
transform 1 0 19872 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_214
timestamp 1644511149
transform 1 0 20792 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_228
timestamp 1644511149
transform 1 0 22080 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_239
timestamp 1644511149
transform 1 0 23092 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_248
timestamp 1644511149
transform 1 0 23920 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_269
timestamp 1644511149
transform 1 0 25852 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_277
timestamp 1644511149
transform 1 0 26588 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_287
timestamp 1644511149
transform 1 0 27508 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_304
timestamp 1644511149
transform 1 0 29072 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_56_320
timestamp 1644511149
transform 1 0 30544 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_56_335
timestamp 1644511149
transform 1 0 31924 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_341
timestamp 1644511149
transform 1 0 32476 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_358
timestamp 1644511149
transform 1 0 34040 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_377
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_384
timestamp 1644511149
transform 1 0 36432 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_396
timestamp 1644511149
transform 1 0 37536 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_408
timestamp 1644511149
transform 1 0 38640 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_421
timestamp 1644511149
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_433
timestamp 1644511149
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_445
timestamp 1644511149
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_457
timestamp 1644511149
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1644511149
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1644511149
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_477
timestamp 1644511149
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_489
timestamp 1644511149
transform 1 0 46092 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_512
timestamp 1644511149
transform 1 0 48208 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_28
timestamp 1644511149
transform 1 0 3680 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_40
timestamp 1644511149
transform 1 0 4784 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_52
timestamp 1644511149
transform 1 0 5888 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1644511149
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_200
timestamp 1644511149
transform 1 0 19504 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_208
timestamp 1644511149
transform 1 0 20240 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_220
timestamp 1644511149
transform 1 0 21344 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_233
timestamp 1644511149
transform 1 0 22540 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_242
timestamp 1644511149
transform 1 0 23368 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_250
timestamp 1644511149
transform 1 0 24104 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_261
timestamp 1644511149
transform 1 0 25116 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_269
timestamp 1644511149
transform 1 0 25852 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_276
timestamp 1644511149
transform 1 0 26496 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_297
timestamp 1644511149
transform 1 0 28428 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_305
timestamp 1644511149
transform 1 0 29164 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_317
timestamp 1644511149
transform 1 0 30268 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_323
timestamp 1644511149
transform 1 0 30820 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_328
timestamp 1644511149
transform 1 0 31280 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_342
timestamp 1644511149
transform 1 0 32568 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_354
timestamp 1644511149
transform 1 0 33672 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_366
timestamp 1644511149
transform 1 0 34776 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_378
timestamp 1644511149
transform 1 0 35880 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_390
timestamp 1644511149
transform 1 0 36984 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_417
timestamp 1644511149
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_429
timestamp 1644511149
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1644511149
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1644511149
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_449
timestamp 1644511149
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_461
timestamp 1644511149
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_473
timestamp 1644511149
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_485
timestamp 1644511149
transform 1 0 45724 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_489
timestamp 1644511149
transform 1 0 46092 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_500
timestamp 1644511149
transform 1 0 47104 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_508
timestamp 1644511149
transform 1 0 47840 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_7
timestamp 1644511149
transform 1 0 1748 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_11
timestamp 1644511149
transform 1 0 2116 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_23
timestamp 1644511149
transform 1 0 3220 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_165
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_177
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1644511149
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_206
timestamp 1644511149
transform 1 0 20056 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_219
timestamp 1644511149
transform 1 0 21252 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_58_235
timestamp 1644511149
transform 1 0 22724 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_248
timestamp 1644511149
transform 1 0 23920 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_259
timestamp 1644511149
transform 1 0 24932 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_273
timestamp 1644511149
transform 1 0 26220 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_277
timestamp 1644511149
transform 1 0 26588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_283
timestamp 1644511149
transform 1 0 27140 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_296
timestamp 1644511149
transform 1 0 28336 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_325
timestamp 1644511149
transform 1 0 31004 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_343
timestamp 1644511149
transform 1 0 32660 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_355
timestamp 1644511149
transform 1 0 33764 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1644511149
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_377
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_389
timestamp 1644511149
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_401
timestamp 1644511149
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1644511149
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1644511149
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_421
timestamp 1644511149
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_433
timestamp 1644511149
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_445
timestamp 1644511149
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_457
timestamp 1644511149
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1644511149
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1644511149
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_477
timestamp 1644511149
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_489
timestamp 1644511149
transform 1 0 46092 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_512
timestamp 1644511149
transform 1 0 48208 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_28
timestamp 1644511149
transform 1 0 3680 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_40
timestamp 1644511149
transform 1 0 4784 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_52
timestamp 1644511149
transform 1 0 5888 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_181
timestamp 1644511149
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_193
timestamp 1644511149
transform 1 0 18860 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_205
timestamp 1644511149
transform 1 0 19964 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_214
timestamp 1644511149
transform 1 0 20792 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_222
timestamp 1644511149
transform 1 0 21528 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_245
timestamp 1644511149
transform 1 0 23644 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_258
timestamp 1644511149
transform 1 0 24840 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_264
timestamp 1644511149
transform 1 0 25392 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_271
timestamp 1644511149
transform 1 0 26036 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1644511149
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_293
timestamp 1644511149
transform 1 0 28060 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_301
timestamp 1644511149
transform 1 0 28796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_315
timestamp 1644511149
transform 1 0 30084 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_326
timestamp 1644511149
transform 1 0 31096 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_334
timestamp 1644511149
transform 1 0 31832 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_344
timestamp 1644511149
transform 1 0 32752 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_356
timestamp 1644511149
transform 1 0 33856 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_368
timestamp 1644511149
transform 1 0 34960 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_380
timestamp 1644511149
transform 1 0 36064 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_417
timestamp 1644511149
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_429
timestamp 1644511149
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1644511149
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1644511149
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_449
timestamp 1644511149
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_461
timestamp 1644511149
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_473
timestamp 1644511149
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_485
timestamp 1644511149
transform 1 0 45724 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_493
timestamp 1644511149
transform 1 0 46460 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_499
timestamp 1644511149
transform 1 0 47012 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1644511149
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_508
timestamp 1644511149
transform 1 0 47840 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_11
timestamp 1644511149
transform 1 0 2116 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_18
timestamp 1644511149
transform 1 0 2760 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_26
timestamp 1644511149
transform 1 0 3496 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_177
timestamp 1644511149
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1644511149
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1644511149
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_208
timestamp 1644511149
transform 1 0 20240 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_218
timestamp 1644511149
transform 1 0 21160 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_226
timestamp 1644511149
transform 1 0 21896 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_238
timestamp 1644511149
transform 1 0 23000 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_250
timestamp 1644511149
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_259
timestamp 1644511149
transform 1 0 24932 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_267
timestamp 1644511149
transform 1 0 25668 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_279
timestamp 1644511149
transform 1 0 26772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_291
timestamp 1644511149
transform 1 0 27876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_303
timestamp 1644511149
transform 1 0 28980 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1644511149
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_314
timestamp 1644511149
transform 1 0 29992 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_323
timestamp 1644511149
transform 1 0 30820 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_342
timestamp 1644511149
transform 1 0 32568 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_354
timestamp 1644511149
transform 1 0 33672 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_362
timestamp 1644511149
transform 1 0 34408 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_401
timestamp 1644511149
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1644511149
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1644511149
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_421
timestamp 1644511149
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_433
timestamp 1644511149
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_445
timestamp 1644511149
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_457
timestamp 1644511149
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1644511149
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1644511149
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_477
timestamp 1644511149
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_489
timestamp 1644511149
transform 1 0 46092 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_512
timestamp 1644511149
transform 1 0 48208 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_30
timestamp 1644511149
transform 1 0 3864 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_42
timestamp 1644511149
transform 1 0 4968 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1644511149
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_201
timestamp 1644511149
transform 1 0 19596 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_205
timestamp 1644511149
transform 1 0 19964 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_214
timestamp 1644511149
transform 1 0 20792 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_222
timestamp 1644511149
transform 1 0 21528 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_237
timestamp 1644511149
transform 1 0 22908 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_245
timestamp 1644511149
transform 1 0 23644 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_253
timestamp 1644511149
transform 1 0 24380 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_263
timestamp 1644511149
transform 1 0 25300 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_276
timestamp 1644511149
transform 1 0 26496 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_290
timestamp 1644511149
transform 1 0 27784 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_298
timestamp 1644511149
transform 1 0 28520 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_302
timestamp 1644511149
transform 1 0 28888 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_309
timestamp 1644511149
transform 1 0 29532 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_322
timestamp 1644511149
transform 1 0 30728 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_334
timestamp 1644511149
transform 1 0 31832 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_353
timestamp 1644511149
transform 1 0 33580 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_365
timestamp 1644511149
transform 1 0 34684 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_377
timestamp 1644511149
transform 1 0 35788 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_389
timestamp 1644511149
transform 1 0 36892 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_417
timestamp 1644511149
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_429
timestamp 1644511149
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1644511149
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1644511149
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_449
timestamp 1644511149
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_461
timestamp 1644511149
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_473
timestamp 1644511149
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_485
timestamp 1644511149
transform 1 0 45724 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_492
timestamp 1644511149
transform 1 0 46368 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_499
timestamp 1644511149
transform 1 0 47012 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1644511149
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_61_505
timestamp 1644511149
transform 1 0 47564 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_512
timestamp 1644511149
transform 1 0 48208 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_15
timestamp 1644511149
transform 1 0 2484 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_62_21
timestamp 1644511149
transform 1 0 3036 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1644511149
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_165
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_177
timestamp 1644511149
transform 1 0 17388 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_183
timestamp 1644511149
transform 1 0 17940 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_192
timestamp 1644511149
transform 1 0 18768 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_202
timestamp 1644511149
transform 1 0 19688 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_210
timestamp 1644511149
transform 1 0 20424 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_228
timestamp 1644511149
transform 1 0 22080 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_241
timestamp 1644511149
transform 1 0 23276 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_249
timestamp 1644511149
transform 1 0 24012 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_253
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_273
timestamp 1644511149
transform 1 0 26220 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_287
timestamp 1644511149
transform 1 0 27508 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_299
timestamp 1644511149
transform 1 0 28612 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1644511149
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_309
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_319
timestamp 1644511149
transform 1 0 30452 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_323
timestamp 1644511149
transform 1 0 30820 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_330
timestamp 1644511149
transform 1 0 31464 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_334
timestamp 1644511149
transform 1 0 31832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_342
timestamp 1644511149
transform 1 0 32568 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_354
timestamp 1644511149
transform 1 0 33672 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_362
timestamp 1644511149
transform 1 0 34408 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_401
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1644511149
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1644511149
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_421
timestamp 1644511149
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_433
timestamp 1644511149
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_445
timestamp 1644511149
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_457
timestamp 1644511149
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1644511149
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1644511149
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_477
timestamp 1644511149
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_489
timestamp 1644511149
transform 1 0 46092 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_512
timestamp 1644511149
transform 1 0 48208 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_9
timestamp 1644511149
transform 1 0 1932 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_13
timestamp 1644511149
transform 1 0 2300 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_25
timestamp 1644511149
transform 1 0 3404 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_37
timestamp 1644511149
transform 1 0 4508 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_49
timestamp 1644511149
transform 1 0 5612 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1644511149
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_200
timestamp 1644511149
transform 1 0 19504 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_208
timestamp 1644511149
transform 1 0 20240 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_215
timestamp 1644511149
transform 1 0 20884 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1644511149
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_230
timestamp 1644511149
transform 1 0 22264 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_242
timestamp 1644511149
transform 1 0 23368 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_254
timestamp 1644511149
transform 1 0 24472 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_265
timestamp 1644511149
transform 1 0 25484 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_276
timestamp 1644511149
transform 1 0 26496 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_287
timestamp 1644511149
transform 1 0 27508 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_297
timestamp 1644511149
transform 1 0 28428 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_306
timestamp 1644511149
transform 1 0 29256 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_310
timestamp 1644511149
transform 1 0 29624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_327
timestamp 1644511149
transform 1 0 31188 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1644511149
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_353
timestamp 1644511149
transform 1 0 33580 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_365
timestamp 1644511149
transform 1 0 34684 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_377
timestamp 1644511149
transform 1 0 35788 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_389
timestamp 1644511149
transform 1 0 36892 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_417
timestamp 1644511149
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_429
timestamp 1644511149
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1644511149
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1644511149
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_449
timestamp 1644511149
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_461
timestamp 1644511149
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_473
timestamp 1644511149
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_485
timestamp 1644511149
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1644511149
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1644511149
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_508
timestamp 1644511149
transform 1 0 47840 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_11
timestamp 1644511149
transform 1 0 2116 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_23
timestamp 1644511149
transform 1 0 3220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_183
timestamp 1644511149
transform 1 0 17940 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_192
timestamp 1644511149
transform 1 0 18768 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_210
timestamp 1644511149
transform 1 0 20424 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_230
timestamp 1644511149
transform 1 0 22264 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_242
timestamp 1644511149
transform 1 0 23368 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_250
timestamp 1644511149
transform 1 0 24104 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_64_268
timestamp 1644511149
transform 1 0 25760 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_276
timestamp 1644511149
transform 1 0 26496 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_286
timestamp 1644511149
transform 1 0 27416 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_299
timestamp 1644511149
transform 1 0 28612 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1644511149
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_325
timestamp 1644511149
transform 1 0 31004 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_333
timestamp 1644511149
transform 1 0 31740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_336
timestamp 1644511149
transform 1 0 32016 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_343
timestamp 1644511149
transform 1 0 32660 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_355
timestamp 1644511149
transform 1 0 33764 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1644511149
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_377
timestamp 1644511149
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_389
timestamp 1644511149
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_401
timestamp 1644511149
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1644511149
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1644511149
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_421
timestamp 1644511149
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_433
timestamp 1644511149
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_445
timestamp 1644511149
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_457
timestamp 1644511149
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1644511149
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1644511149
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_477
timestamp 1644511149
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_489
timestamp 1644511149
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_501
timestamp 1644511149
transform 1 0 47196 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_507
timestamp 1644511149
transform 1 0 47748 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_515
timestamp 1644511149
transform 1 0 48484 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_13
timestamp 1644511149
transform 1 0 2300 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_25
timestamp 1644511149
transform 1 0 3404 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_37
timestamp 1644511149
transform 1 0 4508 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_49
timestamp 1644511149
transform 1 0 5612 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_149
timestamp 1644511149
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1644511149
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1644511149
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_181
timestamp 1644511149
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_193
timestamp 1644511149
transform 1 0 18860 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_197
timestamp 1644511149
transform 1 0 19228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_203
timestamp 1644511149
transform 1 0 19780 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_211
timestamp 1644511149
transform 1 0 20516 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_220
timestamp 1644511149
transform 1 0 21344 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_234
timestamp 1644511149
transform 1 0 22632 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_246
timestamp 1644511149
transform 1 0 23736 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_257
timestamp 1644511149
transform 1 0 24748 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_266
timestamp 1644511149
transform 1 0 25576 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_275
timestamp 1644511149
transform 1 0 26404 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1644511149
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_281
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_65_303
timestamp 1644511149
transform 1 0 28980 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_311
timestamp 1644511149
transform 1 0 29716 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_65_318
timestamp 1644511149
transform 1 0 30360 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_330
timestamp 1644511149
transform 1 0 31464 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_65_337
timestamp 1644511149
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_349
timestamp 1644511149
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_361
timestamp 1644511149
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_373
timestamp 1644511149
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1644511149
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1644511149
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_393
timestamp 1644511149
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_405
timestamp 1644511149
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_417
timestamp 1644511149
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_429
timestamp 1644511149
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1644511149
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1644511149
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_449
timestamp 1644511149
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_461
timestamp 1644511149
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_473
timestamp 1644511149
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_485
timestamp 1644511149
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_500
timestamp 1644511149
transform 1 0 47104 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_65_505
timestamp 1644511149
transform 1 0 47564 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_512
timestamp 1644511149
transform 1 0 48208 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1644511149
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1644511149
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1644511149
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_165
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_177
timestamp 1644511149
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1644511149
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1644511149
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_197
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_209
timestamp 1644511149
transform 1 0 20332 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_218
timestamp 1644511149
transform 1 0 21160 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_238
timestamp 1644511149
transform 1 0 23000 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_250
timestamp 1644511149
transform 1 0 24104 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_269
timestamp 1644511149
transform 1 0 25852 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_297
timestamp 1644511149
transform 1 0 28428 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_305
timestamp 1644511149
transform 1 0 29164 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_309
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_321
timestamp 1644511149
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_333
timestamp 1644511149
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_345
timestamp 1644511149
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1644511149
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1644511149
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_365
timestamp 1644511149
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_377
timestamp 1644511149
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_389
timestamp 1644511149
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_401
timestamp 1644511149
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1644511149
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1644511149
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_421
timestamp 1644511149
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_433
timestamp 1644511149
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_445
timestamp 1644511149
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_457
timestamp 1644511149
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1644511149
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1644511149
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_477
timestamp 1644511149
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_489
timestamp 1644511149
transform 1 0 46092 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_512
timestamp 1644511149
transform 1 0 48208 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_9
timestamp 1644511149
transform 1 0 1932 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_13
timestamp 1644511149
transform 1 0 2300 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_25
timestamp 1644511149
transform 1 0 3404 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_37
timestamp 1644511149
transform 1 0 4508 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_49
timestamp 1644511149
transform 1 0 5612 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1644511149
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1644511149
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_149
timestamp 1644511149
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1644511149
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1644511149
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_181
timestamp 1644511149
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_193
timestamp 1644511149
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_205
timestamp 1644511149
transform 1 0 19964 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_213
timestamp 1644511149
transform 1 0 20700 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_220
timestamp 1644511149
transform 1 0 21344 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_225
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_237
timestamp 1644511149
transform 1 0 22908 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_245
timestamp 1644511149
transform 1 0 23644 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_264
timestamp 1644511149
transform 1 0 25392 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_276
timestamp 1644511149
transform 1 0 26496 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_281
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_293
timestamp 1644511149
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_305
timestamp 1644511149
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_317
timestamp 1644511149
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1644511149
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1644511149
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_337
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_349
timestamp 1644511149
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_361
timestamp 1644511149
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_373
timestamp 1644511149
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1644511149
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1644511149
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_393
timestamp 1644511149
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_405
timestamp 1644511149
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_417
timestamp 1644511149
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_429
timestamp 1644511149
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1644511149
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1644511149
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_449
timestamp 1644511149
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_461
timestamp 1644511149
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_473
timestamp 1644511149
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_485
timestamp 1644511149
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1644511149
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1644511149
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_508
timestamp 1644511149
transform 1 0 47840 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_24
timestamp 1644511149
transform 1 0 3312 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_41
timestamp 1644511149
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_53
timestamp 1644511149
transform 1 0 5980 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_59
timestamp 1644511149
transform 1 0 6532 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_63
timestamp 1644511149
transform 1 0 6900 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_68_72
timestamp 1644511149
transform 1 0 7728 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_109
timestamp 1644511149
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_121
timestamp 1644511149
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1644511149
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1644511149
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1644511149
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_165
timestamp 1644511149
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_177
timestamp 1644511149
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1644511149
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1644511149
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_197
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_209
timestamp 1644511149
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_221
timestamp 1644511149
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_233
timestamp 1644511149
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1644511149
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1644511149
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_261
timestamp 1644511149
transform 1 0 25116 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_273
timestamp 1644511149
transform 1 0 26220 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_285
timestamp 1644511149
transform 1 0 27324 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_297
timestamp 1644511149
transform 1 0 28428 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_305
timestamp 1644511149
transform 1 0 29164 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_321
timestamp 1644511149
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_333
timestamp 1644511149
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_345
timestamp 1644511149
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1644511149
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1644511149
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_365
timestamp 1644511149
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_377
timestamp 1644511149
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_389
timestamp 1644511149
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_401
timestamp 1644511149
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1644511149
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1644511149
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_421
timestamp 1644511149
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_433
timestamp 1644511149
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_445
timestamp 1644511149
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_457
timestamp 1644511149
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1644511149
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1644511149
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_477
timestamp 1644511149
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_489
timestamp 1644511149
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_501
timestamp 1644511149
transform 1 0 47196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_512
timestamp 1644511149
transform 1 0 48208 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_7
timestamp 1644511149
transform 1 0 1748 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_11
timestamp 1644511149
transform 1 0 2116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_23
timestamp 1644511149
transform 1 0 3220 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_35
timestamp 1644511149
transform 1 0 4324 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_47
timestamp 1644511149
transform 1 0 5428 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1644511149
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1644511149
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1644511149
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_93
timestamp 1644511149
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1644511149
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1644511149
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_113
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_125
timestamp 1644511149
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_137
timestamp 1644511149
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_149
timestamp 1644511149
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1644511149
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1644511149
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_169
timestamp 1644511149
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_181
timestamp 1644511149
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_193
timestamp 1644511149
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_205
timestamp 1644511149
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1644511149
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1644511149
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_225
timestamp 1644511149
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_237
timestamp 1644511149
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_249
timestamp 1644511149
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_261
timestamp 1644511149
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1644511149
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1644511149
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_281
timestamp 1644511149
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_293
timestamp 1644511149
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_305
timestamp 1644511149
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_317
timestamp 1644511149
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1644511149
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1644511149
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_337
timestamp 1644511149
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_349
timestamp 1644511149
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_361
timestamp 1644511149
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_373
timestamp 1644511149
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1644511149
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1644511149
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_393
timestamp 1644511149
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_405
timestamp 1644511149
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_417
timestamp 1644511149
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_429
timestamp 1644511149
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1644511149
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1644511149
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_449
timestamp 1644511149
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_461
timestamp 1644511149
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_473
timestamp 1644511149
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_485
timestamp 1644511149
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_500
timestamp 1644511149
transform 1 0 47104 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_508
timestamp 1644511149
transform 1 0 47840 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_3
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_11
timestamp 1644511149
transform 1 0 2116 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_23
timestamp 1644511149
transform 1 0 3220 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1644511149
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1644511149
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1644511149
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1644511149
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1644511149
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1644511149
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_97
timestamp 1644511149
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_109
timestamp 1644511149
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_121
timestamp 1644511149
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1644511149
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1644511149
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_153
timestamp 1644511149
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_165
timestamp 1644511149
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_177
timestamp 1644511149
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1644511149
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1644511149
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_197
timestamp 1644511149
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_209
timestamp 1644511149
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_221
timestamp 1644511149
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_233
timestamp 1644511149
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1644511149
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1644511149
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_253
timestamp 1644511149
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_265
timestamp 1644511149
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_277
timestamp 1644511149
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_289
timestamp 1644511149
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1644511149
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1644511149
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_309
timestamp 1644511149
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_321
timestamp 1644511149
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_333
timestamp 1644511149
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_345
timestamp 1644511149
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1644511149
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1644511149
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_365
timestamp 1644511149
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_377
timestamp 1644511149
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_389
timestamp 1644511149
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_401
timestamp 1644511149
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1644511149
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1644511149
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_421
timestamp 1644511149
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_433
timestamp 1644511149
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_445
timestamp 1644511149
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_457
timestamp 1644511149
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1644511149
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1644511149
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_477
timestamp 1644511149
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_489
timestamp 1644511149
transform 1 0 46092 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_512
timestamp 1644511149
transform 1 0 48208 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_7
timestamp 1644511149
transform 1 0 1748 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_14
timestamp 1644511149
transform 1 0 2392 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_26
timestamp 1644511149
transform 1 0 3496 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_38
timestamp 1644511149
transform 1 0 4600 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_50
timestamp 1644511149
transform 1 0 5704 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1644511149
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_93
timestamp 1644511149
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1644511149
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1644511149
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_125
timestamp 1644511149
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_137
timestamp 1644511149
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_149
timestamp 1644511149
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1644511149
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1644511149
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_169
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_181
timestamp 1644511149
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_193
timestamp 1644511149
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_205
timestamp 1644511149
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1644511149
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1644511149
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_225
timestamp 1644511149
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_237
timestamp 1644511149
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_249
timestamp 1644511149
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_261
timestamp 1644511149
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1644511149
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1644511149
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_281
timestamp 1644511149
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_293
timestamp 1644511149
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_305
timestamp 1644511149
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_317
timestamp 1644511149
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1644511149
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1644511149
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_337
timestamp 1644511149
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_349
timestamp 1644511149
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_361
timestamp 1644511149
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_373
timestamp 1644511149
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1644511149
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1644511149
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_393
timestamp 1644511149
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_405
timestamp 1644511149
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_417
timestamp 1644511149
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_429
timestamp 1644511149
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1644511149
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1644511149
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_449
timestamp 1644511149
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_461
timestamp 1644511149
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_473
timestamp 1644511149
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_485
timestamp 1644511149
transform 1 0 45724 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_493
timestamp 1644511149
transform 1 0 46460 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_499
timestamp 1644511149
transform 1 0 47012 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1644511149
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_71_505
timestamp 1644511149
transform 1 0 47564 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_512
timestamp 1644511149
transform 1 0 48208 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_24
timestamp 1644511149
transform 1 0 3312 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1644511149
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1644511149
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1644511149
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1644511149
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1644511149
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1644511149
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_97
timestamp 1644511149
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_109
timestamp 1644511149
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_121
timestamp 1644511149
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1644511149
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1644511149
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1644511149
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_153
timestamp 1644511149
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_165
timestamp 1644511149
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_177
timestamp 1644511149
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1644511149
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1644511149
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_197
timestamp 1644511149
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_209
timestamp 1644511149
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_221
timestamp 1644511149
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_233
timestamp 1644511149
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1644511149
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1644511149
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_253
timestamp 1644511149
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_265
timestamp 1644511149
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_277
timestamp 1644511149
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_289
timestamp 1644511149
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1644511149
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1644511149
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_309
timestamp 1644511149
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_321
timestamp 1644511149
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_333
timestamp 1644511149
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_345
timestamp 1644511149
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1644511149
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1644511149
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_365
timestamp 1644511149
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_377
timestamp 1644511149
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_389
timestamp 1644511149
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_401
timestamp 1644511149
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1644511149
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1644511149
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_421
timestamp 1644511149
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_433
timestamp 1644511149
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_445
timestamp 1644511149
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_457
timestamp 1644511149
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1644511149
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1644511149
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_477
timestamp 1644511149
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_489
timestamp 1644511149
transform 1 0 46092 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_512
timestamp 1644511149
transform 1 0 48208 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_3
timestamp 1644511149
transform 1 0 1380 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_7
timestamp 1644511149
transform 1 0 1748 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_11
timestamp 1644511149
transform 1 0 2116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_23
timestamp 1644511149
transform 1 0 3220 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_35
timestamp 1644511149
transform 1 0 4324 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_47
timestamp 1644511149
transform 1 0 5428 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1644511149
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1644511149
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_93
timestamp 1644511149
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1644511149
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1644511149
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1644511149
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1644511149
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_137
timestamp 1644511149
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_149
timestamp 1644511149
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1644511149
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1644511149
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_169
timestamp 1644511149
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_181
timestamp 1644511149
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_193
timestamp 1644511149
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_205
timestamp 1644511149
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1644511149
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1644511149
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_225
timestamp 1644511149
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_237
timestamp 1644511149
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_249
timestamp 1644511149
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_261
timestamp 1644511149
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1644511149
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1644511149
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_281
timestamp 1644511149
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_293
timestamp 1644511149
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_305
timestamp 1644511149
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_317
timestamp 1644511149
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1644511149
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1644511149
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_337
timestamp 1644511149
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_349
timestamp 1644511149
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_361
timestamp 1644511149
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_373
timestamp 1644511149
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1644511149
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1644511149
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_393
timestamp 1644511149
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_405
timestamp 1644511149
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_417
timestamp 1644511149
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_429
timestamp 1644511149
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1644511149
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1644511149
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_449
timestamp 1644511149
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_461
timestamp 1644511149
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_473
timestamp 1644511149
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_485
timestamp 1644511149
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_500
timestamp 1644511149
transform 1 0 47104 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_73_505
timestamp 1644511149
transform 1 0 47564 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_512
timestamp 1644511149
transform 1 0 48208 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1644511149
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1644511149
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1644511149
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1644511149
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1644511149
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_53
timestamp 1644511149
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_65
timestamp 1644511149
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1644511149
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1644511149
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_85
timestamp 1644511149
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_97
timestamp 1644511149
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_109
timestamp 1644511149
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_121
timestamp 1644511149
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1644511149
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1644511149
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1644511149
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_153
timestamp 1644511149
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_165
timestamp 1644511149
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_177
timestamp 1644511149
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1644511149
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1644511149
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_197
timestamp 1644511149
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_209
timestamp 1644511149
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_221
timestamp 1644511149
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_233
timestamp 1644511149
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1644511149
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1644511149
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_253
timestamp 1644511149
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_265
timestamp 1644511149
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_277
timestamp 1644511149
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_289
timestamp 1644511149
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1644511149
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1644511149
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_309
timestamp 1644511149
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_321
timestamp 1644511149
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_333
timestamp 1644511149
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_345
timestamp 1644511149
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1644511149
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1644511149
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_365
timestamp 1644511149
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_377
timestamp 1644511149
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_389
timestamp 1644511149
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_401
timestamp 1644511149
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1644511149
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1644511149
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_421
timestamp 1644511149
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_433
timestamp 1644511149
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_445
timestamp 1644511149
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_457
timestamp 1644511149
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1644511149
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1644511149
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_477
timestamp 1644511149
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_489
timestamp 1644511149
transform 1 0 46092 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_512
timestamp 1644511149
transform 1 0 48208 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_3
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_15
timestamp 1644511149
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_27
timestamp 1644511149
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_39
timestamp 1644511149
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1644511149
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1644511149
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1644511149
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1644511149
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_93
timestamp 1644511149
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1644511149
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1644511149
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_113
timestamp 1644511149
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_125
timestamp 1644511149
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_137
timestamp 1644511149
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_149
timestamp 1644511149
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1644511149
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1644511149
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_169
timestamp 1644511149
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_181
timestamp 1644511149
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_193
timestamp 1644511149
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_205
timestamp 1644511149
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1644511149
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1644511149
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_225
timestamp 1644511149
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_237
timestamp 1644511149
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_249
timestamp 1644511149
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_261
timestamp 1644511149
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1644511149
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1644511149
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_281
timestamp 1644511149
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_293
timestamp 1644511149
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_305
timestamp 1644511149
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_317
timestamp 1644511149
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1644511149
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1644511149
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_337
timestamp 1644511149
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_349
timestamp 1644511149
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_361
timestamp 1644511149
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_373
timestamp 1644511149
transform 1 0 35420 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_381
timestamp 1644511149
transform 1 0 36156 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_387
timestamp 1644511149
transform 1 0 36708 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1644511149
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_393
timestamp 1644511149
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_405
timestamp 1644511149
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_417
timestamp 1644511149
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_429
timestamp 1644511149
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1644511149
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1644511149
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_449
timestamp 1644511149
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_461
timestamp 1644511149
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_473
timestamp 1644511149
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_485
timestamp 1644511149
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1644511149
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1644511149
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_75_505
timestamp 1644511149
transform 1 0 47564 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_512
timestamp 1644511149
transform 1 0 48208 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_9
timestamp 1644511149
transform 1 0 1932 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_17
timestamp 1644511149
transform 1 0 2668 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_76_22
timestamp 1644511149
transform 1 0 3128 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1644511149
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1644511149
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1644511149
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_65
timestamp 1644511149
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1644511149
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1644511149
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_85
timestamp 1644511149
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_97
timestamp 1644511149
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_109
timestamp 1644511149
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_121
timestamp 1644511149
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1644511149
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1644511149
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_141
timestamp 1644511149
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_153
timestamp 1644511149
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_165
timestamp 1644511149
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_177
timestamp 1644511149
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1644511149
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1644511149
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_197
timestamp 1644511149
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_209
timestamp 1644511149
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_221
timestamp 1644511149
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_233
timestamp 1644511149
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1644511149
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1644511149
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_253
timestamp 1644511149
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_265
timestamp 1644511149
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_277
timestamp 1644511149
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_289
timestamp 1644511149
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1644511149
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1644511149
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_309
timestamp 1644511149
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_321
timestamp 1644511149
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_333
timestamp 1644511149
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_345
timestamp 1644511149
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1644511149
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1644511149
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_365
timestamp 1644511149
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_377
timestamp 1644511149
transform 1 0 35788 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_404
timestamp 1644511149
transform 1 0 38272 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_416
timestamp 1644511149
transform 1 0 39376 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_421
timestamp 1644511149
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_433
timestamp 1644511149
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_445
timestamp 1644511149
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_457
timestamp 1644511149
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1644511149
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1644511149
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_477
timestamp 1644511149
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_489
timestamp 1644511149
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_501
timestamp 1644511149
transform 1 0 47196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_505
timestamp 1644511149
transform 1 0 47564 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_512
timestamp 1644511149
transform 1 0 48208 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_3
timestamp 1644511149
transform 1 0 1380 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_9
timestamp 1644511149
transform 1 0 1932 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_31
timestamp 1644511149
transform 1 0 3956 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_43
timestamp 1644511149
transform 1 0 5060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1644511149
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1644511149
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1644511149
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1644511149
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_93
timestamp 1644511149
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1644511149
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1644511149
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_113
timestamp 1644511149
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_125
timestamp 1644511149
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_137
timestamp 1644511149
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_149
timestamp 1644511149
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1644511149
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1644511149
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_169
timestamp 1644511149
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_181
timestamp 1644511149
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_193
timestamp 1644511149
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_205
timestamp 1644511149
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1644511149
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1644511149
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_225
timestamp 1644511149
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_237
timestamp 1644511149
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_249
timestamp 1644511149
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_261
timestamp 1644511149
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1644511149
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1644511149
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_281
timestamp 1644511149
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_293
timestamp 1644511149
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_305
timestamp 1644511149
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_317
timestamp 1644511149
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1644511149
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1644511149
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_337
timestamp 1644511149
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_349
timestamp 1644511149
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_361
timestamp 1644511149
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_373
timestamp 1644511149
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1644511149
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1644511149
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_393
timestamp 1644511149
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_405
timestamp 1644511149
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_417
timestamp 1644511149
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_429
timestamp 1644511149
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1644511149
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1644511149
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_449
timestamp 1644511149
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_461
timestamp 1644511149
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_473
timestamp 1644511149
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_485
timestamp 1644511149
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_500
timestamp 1644511149
transform 1 0 47104 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_508
timestamp 1644511149
transform 1 0 47840 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_78_7
timestamp 1644511149
transform 1 0 1748 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_14
timestamp 1644511149
transform 1 0 2392 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_21
timestamp 1644511149
transform 1 0 3036 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1644511149
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1644511149
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_41
timestamp 1644511149
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_53
timestamp 1644511149
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_65
timestamp 1644511149
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1644511149
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1644511149
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_85
timestamp 1644511149
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_97
timestamp 1644511149
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_109
timestamp 1644511149
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_121
timestamp 1644511149
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1644511149
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1644511149
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1644511149
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_153
timestamp 1644511149
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_165
timestamp 1644511149
transform 1 0 16284 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_177
timestamp 1644511149
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1644511149
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1644511149
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_197
timestamp 1644511149
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_209
timestamp 1644511149
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_221
timestamp 1644511149
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_233
timestamp 1644511149
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1644511149
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1644511149
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_253
timestamp 1644511149
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_265
timestamp 1644511149
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_277
timestamp 1644511149
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_289
timestamp 1644511149
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1644511149
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1644511149
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_309
timestamp 1644511149
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_321
timestamp 1644511149
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_78_333
timestamp 1644511149
transform 1 0 31740 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_78_356
timestamp 1644511149
transform 1 0 33856 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_365
timestamp 1644511149
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_377
timestamp 1644511149
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_389
timestamp 1644511149
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_401
timestamp 1644511149
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1644511149
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1644511149
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_421
timestamp 1644511149
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_433
timestamp 1644511149
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_445
timestamp 1644511149
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_457
timestamp 1644511149
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1644511149
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1644511149
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_78_477
timestamp 1644511149
transform 1 0 44988 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_483
timestamp 1644511149
transform 1 0 45540 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_487
timestamp 1644511149
transform 1 0 45908 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_512
timestamp 1644511149
transform 1 0 48208 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_7
timestamp 1644511149
transform 1 0 1748 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_11
timestamp 1644511149
transform 1 0 2116 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_16
timestamp 1644511149
transform 1 0 2576 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_28
timestamp 1644511149
transform 1 0 3680 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_40
timestamp 1644511149
transform 1 0 4784 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_52
timestamp 1644511149
transform 1 0 5888 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1644511149
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1644511149
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_81
timestamp 1644511149
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_93
timestamp 1644511149
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1644511149
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1644511149
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_113
timestamp 1644511149
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_125
timestamp 1644511149
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_137
timestamp 1644511149
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_149
timestamp 1644511149
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1644511149
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1644511149
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_169
timestamp 1644511149
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_181
timestamp 1644511149
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_193
timestamp 1644511149
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_205
timestamp 1644511149
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1644511149
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1644511149
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_225
timestamp 1644511149
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_237
timestamp 1644511149
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_249
timestamp 1644511149
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_261
timestamp 1644511149
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1644511149
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1644511149
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_281
timestamp 1644511149
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_293
timestamp 1644511149
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_305
timestamp 1644511149
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_317
timestamp 1644511149
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1644511149
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1644511149
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_337
timestamp 1644511149
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_349
timestamp 1644511149
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_361
timestamp 1644511149
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_373
timestamp 1644511149
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1644511149
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1644511149
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_393
timestamp 1644511149
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_405
timestamp 1644511149
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_417
timestamp 1644511149
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_429
timestamp 1644511149
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1644511149
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1644511149
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_449
timestamp 1644511149
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_461
timestamp 1644511149
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_473
timestamp 1644511149
transform 1 0 44620 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_479
timestamp 1644511149
transform 1 0 45172 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_486
timestamp 1644511149
transform 1 0 45816 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_493
timestamp 1644511149
transform 1 0 46460 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_500
timestamp 1644511149
transform 1 0 47104 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_508
timestamp 1644511149
transform 1 0 47840 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_80_24
timestamp 1644511149
transform 1 0 3312 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_29
timestamp 1644511149
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_41
timestamp 1644511149
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_53
timestamp 1644511149
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_65
timestamp 1644511149
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1644511149
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1644511149
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_85
timestamp 1644511149
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_97
timestamp 1644511149
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_120
timestamp 1644511149
transform 1 0 12144 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_132
timestamp 1644511149
transform 1 0 13248 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_141
timestamp 1644511149
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_153
timestamp 1644511149
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_165
timestamp 1644511149
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_177
timestamp 1644511149
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1644511149
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1644511149
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_197
timestamp 1644511149
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_209
timestamp 1644511149
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_221
timestamp 1644511149
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_233
timestamp 1644511149
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1644511149
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1644511149
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_253
timestamp 1644511149
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_265
timestamp 1644511149
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_277
timestamp 1644511149
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_289
timestamp 1644511149
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1644511149
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1644511149
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_309
timestamp 1644511149
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_321
timestamp 1644511149
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_333
timestamp 1644511149
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_345
timestamp 1644511149
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1644511149
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1644511149
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_365
timestamp 1644511149
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_377
timestamp 1644511149
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_389
timestamp 1644511149
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_401
timestamp 1644511149
transform 1 0 37996 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_408
timestamp 1644511149
transform 1 0 38640 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_421
timestamp 1644511149
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_433
timestamp 1644511149
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_445
timestamp 1644511149
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_457
timestamp 1644511149
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_472
timestamp 1644511149
transform 1 0 44528 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_477
timestamp 1644511149
transform 1 0 44988 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_80_482
timestamp 1644511149
transform 1 0 45448 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_490
timestamp 1644511149
transform 1 0 46184 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_512
timestamp 1644511149
transform 1 0 48208 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_3
timestamp 1644511149
transform 1 0 1380 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_28
timestamp 1644511149
transform 1 0 3680 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_35
timestamp 1644511149
transform 1 0 4324 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_47
timestamp 1644511149
transform 1 0 5428 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1644511149
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1644511149
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_69
timestamp 1644511149
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_81
timestamp 1644511149
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_93
timestamp 1644511149
transform 1 0 9660 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_101
timestamp 1644511149
transform 1 0 10396 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_108
timestamp 1644511149
transform 1 0 11040 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_113
timestamp 1644511149
transform 1 0 11500 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_137
timestamp 1644511149
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_149
timestamp 1644511149
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1644511149
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1644511149
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_169
timestamp 1644511149
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_181
timestamp 1644511149
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_193
timestamp 1644511149
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_205
timestamp 1644511149
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1644511149
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1644511149
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_225
timestamp 1644511149
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_237
timestamp 1644511149
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_249
timestamp 1644511149
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_261
timestamp 1644511149
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1644511149
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1644511149
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_281
timestamp 1644511149
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_293
timestamp 1644511149
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_305
timestamp 1644511149
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_317
timestamp 1644511149
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1644511149
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1644511149
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_337
timestamp 1644511149
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_349
timestamp 1644511149
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_361
timestamp 1644511149
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_373
timestamp 1644511149
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1644511149
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1644511149
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_393
timestamp 1644511149
transform 1 0 37260 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_401
timestamp 1644511149
transform 1 0 37996 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_423
timestamp 1644511149
transform 1 0 40020 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_435
timestamp 1644511149
transform 1 0 41124 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1644511149
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_449
timestamp 1644511149
transform 1 0 42412 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_81_458
timestamp 1644511149
transform 1 0 43240 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_467
timestamp 1644511149
transform 1 0 44068 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_474
timestamp 1644511149
transform 1 0 44712 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_478
timestamp 1644511149
transform 1 0 45080 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_500
timestamp 1644511149
transform 1 0 47104 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_508
timestamp 1644511149
transform 1 0 47840 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_3
timestamp 1644511149
transform 1 0 1380 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_8
timestamp 1644511149
transform 1 0 1840 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_15
timestamp 1644511149
transform 1 0 2484 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_22
timestamp 1644511149
transform 1 0 3128 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_82_32
timestamp 1644511149
transform 1 0 4048 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_61
timestamp 1644511149
transform 1 0 6716 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_73
timestamp 1644511149
transform 1 0 7820 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_81
timestamp 1644511149
transform 1 0 8556 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_85
timestamp 1644511149
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_97
timestamp 1644511149
transform 1 0 10028 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_105
timestamp 1644511149
transform 1 0 10764 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_129
timestamp 1644511149
transform 1 0 12972 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_137
timestamp 1644511149
transform 1 0 13708 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_141
timestamp 1644511149
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_153
timestamp 1644511149
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_165
timestamp 1644511149
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_177
timestamp 1644511149
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1644511149
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1644511149
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_197
timestamp 1644511149
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_209
timestamp 1644511149
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_221
timestamp 1644511149
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_233
timestamp 1644511149
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1644511149
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1644511149
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_253
timestamp 1644511149
transform 1 0 24380 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_261
timestamp 1644511149
transform 1 0 25116 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_267
timestamp 1644511149
transform 1 0 25668 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_274
timestamp 1644511149
transform 1 0 26312 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_281
timestamp 1644511149
transform 1 0 26956 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_289
timestamp 1644511149
transform 1 0 27692 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_293
timestamp 1644511149
transform 1 0 28060 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_300
timestamp 1644511149
transform 1 0 28704 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_82_312
timestamp 1644511149
transform 1 0 29808 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_316
timestamp 1644511149
transform 1 0 30176 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_320
timestamp 1644511149
transform 1 0 30544 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_332
timestamp 1644511149
transform 1 0 31648 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_344
timestamp 1644511149
transform 1 0 32752 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_356
timestamp 1644511149
transform 1 0 33856 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_365
timestamp 1644511149
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_377
timestamp 1644511149
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_389
timestamp 1644511149
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_401
timestamp 1644511149
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1644511149
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1644511149
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_421
timestamp 1644511149
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_433
timestamp 1644511149
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_445
timestamp 1644511149
transform 1 0 42044 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_472
timestamp 1644511149
transform 1 0 44528 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_480
timestamp 1644511149
transform 1 0 45264 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_487
timestamp 1644511149
transform 1 0 45908 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_512
timestamp 1644511149
transform 1 0 48208 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_3
timestamp 1644511149
transform 1 0 1380 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_11
timestamp 1644511149
transform 1 0 2116 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_18
timestamp 1644511149
transform 1 0 2760 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_83_25
timestamp 1644511149
transform 1 0 3404 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_31
timestamp 1644511149
transform 1 0 3956 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_83_35
timestamp 1644511149
transform 1 0 4324 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_83_44
timestamp 1644511149
transform 1 0 5152 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1644511149
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1644511149
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_57
timestamp 1644511149
transform 1 0 6348 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_64
timestamp 1644511149
transform 1 0 6992 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_83_89
timestamp 1644511149
transform 1 0 9292 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_97
timestamp 1644511149
transform 1 0 10028 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_101
timestamp 1644511149
transform 1 0 10396 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_108
timestamp 1644511149
transform 1 0 11040 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_83_125
timestamp 1644511149
transform 1 0 12604 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_131
timestamp 1644511149
transform 1 0 13156 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_135
timestamp 1644511149
transform 1 0 13524 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_83_146
timestamp 1644511149
transform 1 0 14536 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_83_157
timestamp 1644511149
transform 1 0 15548 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_83_165
timestamp 1644511149
transform 1 0 16284 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_83_169
timestamp 1644511149
transform 1 0 16652 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_177
timestamp 1644511149
transform 1 0 17388 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_83_182
timestamp 1644511149
transform 1 0 17848 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_188
timestamp 1644511149
transform 1 0 18400 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_192
timestamp 1644511149
transform 1 0 18768 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_204
timestamp 1644511149
transform 1 0 19872 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_216
timestamp 1644511149
transform 1 0 20976 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_83_225
timestamp 1644511149
transform 1 0 21804 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_232
timestamp 1644511149
transform 1 0 22448 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_83_239
timestamp 1644511149
transform 1 0 23092 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_83_247
timestamp 1644511149
transform 1 0 23828 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_83_253
timestamp 1644511149
transform 1 0 24380 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_83_268
timestamp 1644511149
transform 1 0 25760 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_272
timestamp 1644511149
transform 1 0 26128 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_276
timestamp 1644511149
transform 1 0 26496 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_83_281
timestamp 1644511149
transform 1 0 26956 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_83_287
timestamp 1644511149
transform 1 0 27508 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_293
timestamp 1644511149
transform 1 0 28060 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_315
timestamp 1644511149
transform 1 0 30084 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_322
timestamp 1644511149
transform 1 0 30728 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 1644511149
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1644511149
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_340
timestamp 1644511149
transform 1 0 32384 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_344
timestamp 1644511149
transform 1 0 32752 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_348
timestamp 1644511149
transform 1 0 33120 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_373
timestamp 1644511149
transform 1 0 35420 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_380
timestamp 1644511149
transform 1 0 36064 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_387
timestamp 1644511149
transform 1 0 36708 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1644511149
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_393
timestamp 1644511149
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_405
timestamp 1644511149
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_417
timestamp 1644511149
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_429
timestamp 1644511149
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_444
timestamp 1644511149
transform 1 0 41952 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_470
timestamp 1644511149
transform 1 0 44344 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_83_495
timestamp 1644511149
transform 1 0 46644 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1644511149
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_83_505
timestamp 1644511149
transform 1 0 47564 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_83_512
timestamp 1644511149
transform 1 0 48208 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_24
timestamp 1644511149
transform 1 0 3312 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_84_32
timestamp 1644511149
transform 1 0 4048 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_38
timestamp 1644511149
transform 1 0 4600 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_60
timestamp 1644511149
transform 1 0 6624 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_67
timestamp 1644511149
transform 1 0 7268 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_84_74
timestamp 1644511149
transform 1 0 7912 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_82
timestamp 1644511149
transform 1 0 8648 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_85
timestamp 1644511149
transform 1 0 8924 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_84_90
timestamp 1644511149
transform 1 0 9384 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_84_119
timestamp 1644511149
transform 1 0 12052 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_127
timestamp 1644511149
transform 1 0 12788 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1644511149
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1644511149
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_141
timestamp 1644511149
transform 1 0 14076 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_166
timestamp 1644511149
transform 1 0 16376 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_84_173
timestamp 1644511149
transform 1 0 17020 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_185
timestamp 1644511149
transform 1 0 18124 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_84_193
timestamp 1644511149
transform 1 0 18860 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_84_200
timestamp 1644511149
transform 1 0 19504 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_212
timestamp 1644511149
transform 1 0 20608 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_84_221
timestamp 1644511149
transform 1 0 21436 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_84_246
timestamp 1644511149
transform 1 0 23736 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_84_274
timestamp 1644511149
transform 1 0 26312 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_282
timestamp 1644511149
transform 1 0 27048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_304
timestamp 1644511149
transform 1 0 29072 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_330
timestamp 1644511149
transform 1 0 31464 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_84_355
timestamp 1644511149
transform 1 0 33764 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 1644511149
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_84_365
timestamp 1644511149
transform 1 0 34684 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_84_375
timestamp 1644511149
transform 1 0 35604 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_84_400
timestamp 1644511149
transform 1 0 37904 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_412
timestamp 1644511149
transform 1 0 39008 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_84_424
timestamp 1644511149
transform 1 0 40112 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_84_432
timestamp 1644511149
transform 1 0 40848 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_84_438
timestamp 1644511149
transform 1 0 41400 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_463
timestamp 1644511149
transform 1 0 43700 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_471
timestamp 1644511149
transform 1 0 44436 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1644511149
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_480
timestamp 1644511149
transform 1 0 45264 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_487
timestamp 1644511149
transform 1 0 45908 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_512
timestamp 1644511149
transform 1 0 48208 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_9
timestamp 1644511149
transform 1 0 1932 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_17
timestamp 1644511149
transform 1 0 2668 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_21
timestamp 1644511149
transform 1 0 3036 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_43
timestamp 1644511149
transform 1 0 5060 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1644511149
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1644511149
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_57
timestamp 1644511149
transform 1 0 6348 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_82
timestamp 1644511149
transform 1 0 8648 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_86
timestamp 1644511149
transform 1 0 9016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_108
timestamp 1644511149
transform 1 0 11040 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_113
timestamp 1644511149
transform 1 0 11500 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_118
timestamp 1644511149
transform 1 0 11960 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_143
timestamp 1644511149
transform 1 0 14260 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_85_151
timestamp 1644511149
transform 1 0 14996 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_85_159
timestamp 1644511149
transform 1 0 15732 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_85_164
timestamp 1644511149
transform 1 0 16192 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_85_190
timestamp 1644511149
transform 1 0 18584 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_196
timestamp 1644511149
transform 1 0 19136 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_85_218
timestamp 1644511149
transform 1 0 21160 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_225
timestamp 1644511149
transform 1 0 21804 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_229
timestamp 1644511149
transform 1 0 22172 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_85_254
timestamp 1644511149
transform 1 0 24472 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_85_262
timestamp 1644511149
transform 1 0 25208 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_266
timestamp 1644511149
transform 1 0 25576 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_85_274
timestamp 1644511149
transform 1 0 26312 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_85_281
timestamp 1644511149
transform 1 0 26956 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_285
timestamp 1644511149
transform 1 0 27324 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_307
timestamp 1644511149
transform 1 0 29348 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_332
timestamp 1644511149
transform 1 0 31648 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_85_358
timestamp 1644511149
transform 1 0 34040 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_85_366
timestamp 1644511149
transform 1 0 34776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_388
timestamp 1644511149
transform 1 0 36800 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_393
timestamp 1644511149
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_85_405
timestamp 1644511149
transform 1 0 38364 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_85_411
timestamp 1644511149
transform 1 0 38916 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_436
timestamp 1644511149
transform 1 0 41216 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_440
timestamp 1644511149
transform 1 0 41584 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_444
timestamp 1644511149
transform 1 0 41952 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_452
timestamp 1644511149
transform 1 0 42688 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_459
timestamp 1644511149
transform 1 0 43332 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_467
timestamp 1644511149
transform 1 0 44068 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_492
timestamp 1644511149
transform 1 0 46368 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_500
timestamp 1644511149
transform 1 0 47104 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_85_505
timestamp 1644511149
transform 1 0 47564 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_85_512
timestamp 1644511149
transform 1 0 48208 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_24
timestamp 1644511149
transform 1 0 3312 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_29
timestamp 1644511149
transform 1 0 3772 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_39
timestamp 1644511149
transform 1 0 4692 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_49
timestamp 1644511149
transform 1 0 5612 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_55
timestamp 1644511149
transform 1 0 6164 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_86_57
timestamp 1644511149
transform 1 0 6348 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_86_63
timestamp 1644511149
transform 1 0 6900 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_70
timestamp 1644511149
transform 1 0 7544 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1644511149
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1644511149
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_85
timestamp 1644511149
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_97
timestamp 1644511149
transform 1 0 10028 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_101
timestamp 1644511149
transform 1 0 10396 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_108
timestamp 1644511149
transform 1 0 11040 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_134
timestamp 1644511149
transform 1 0 13432 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_86_141
timestamp 1644511149
transform 1 0 14076 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_86_153
timestamp 1644511149
transform 1 0 15180 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_86_160
timestamp 1644511149
transform 1 0 15824 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_86_169
timestamp 1644511149
transform 1 0 16652 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_177
timestamp 1644511149
transform 1 0 17388 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_181
timestamp 1644511149
transform 1 0 17756 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_192
timestamp 1644511149
transform 1 0 18768 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_197
timestamp 1644511149
transform 1 0 19228 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_202
timestamp 1644511149
transform 1 0 19688 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_86_210
timestamp 1644511149
transform 1 0 20424 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_86_222
timestamp 1644511149
transform 1 0 21528 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_225
timestamp 1644511149
transform 1 0 21804 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_86_237
timestamp 1644511149
transform 1 0 22908 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_86_248
timestamp 1644511149
transform 1 0 23920 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_86_263
timestamp 1644511149
transform 1 0 25300 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_271
timestamp 1644511149
transform 1 0 26036 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_86_276
timestamp 1644511149
transform 1 0 26496 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_302
timestamp 1644511149
transform 1 0 28888 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_86_309
timestamp 1644511149
transform 1 0 29532 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_317
timestamp 1644511149
transform 1 0 30268 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_86_326
timestamp 1644511149
transform 1 0 31096 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_334
timestamp 1644511149
transform 1 0 31832 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_86_340
timestamp 1644511149
transform 1 0 32384 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_352
timestamp 1644511149
transform 1 0 33488 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_356
timestamp 1644511149
transform 1 0 33856 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_86_365
timestamp 1644511149
transform 1 0 34684 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_86_376
timestamp 1644511149
transform 1 0 35696 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_86_383
timestamp 1644511149
transform 1 0 36340 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_391
timestamp 1644511149
transform 1 0 37076 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_393
timestamp 1644511149
transform 1 0 37260 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_401
timestamp 1644511149
transform 1 0 37996 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_406
timestamp 1644511149
transform 1 0 38456 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_86_418
timestamp 1644511149
transform 1 0 39560 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_86_421
timestamp 1644511149
transform 1 0 39836 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_429
timestamp 1644511149
transform 1 0 40572 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_86_434
timestamp 1644511149
transform 1 0 41032 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_86_444
timestamp 1644511149
transform 1 0 41952 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_470
timestamp 1644511149
transform 1 0 44344 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_86_477
timestamp 1644511149
transform 1 0 44988 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_86_500
timestamp 1644511149
transform 1 0 47104 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_505
timestamp 1644511149
transform 1 0 47564 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_512
timestamp 1644511149
transform 1 0 48208 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 48852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 48852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 48852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 48852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 48852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 48852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 48852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 48852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 48852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 48852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 48852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 48852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 48852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 48852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 48852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 48852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 48852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 48852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 48852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 48852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 48852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 48852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 48852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 48852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 48852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 48852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 48852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 48852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 48852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 48852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 48852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 48852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 48852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 48852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 48852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 48852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 48852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 48852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 48852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 48852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 48852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 48852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 48852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 48852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 48852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 48852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 48852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 48852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 48852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 48852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 48852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 48852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 48852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 48852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 48852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 48852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 48852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 48852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 48852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 48852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 48852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 48852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 48852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 48852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 48852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 48852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 48852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 48852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 48852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 48852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 48852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 48852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 48852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 48852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 48852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 48852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1644511149
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1644511149
transform -1 0 48852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1644511149
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1644511149
transform -1 0 48852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1644511149
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1644511149
transform -1 0 48852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1644511149
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1644511149
transform -1 0 48852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1644511149
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1644511149
transform -1 0 48852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1644511149
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1644511149
transform -1 0 48852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1644511149
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1644511149
transform -1 0 48852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1644511149
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1644511149
transform -1 0 48852 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1644511149
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1644511149
transform -1 0 48852 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1644511149
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1644511149
transform -1 0 48852 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1644511149
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1644511149
transform -1 0 48852 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1644511149
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1644511149
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1644511149
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1644511149
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1644511149
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1644511149
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1644511149
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1644511149
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1644511149
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1644511149
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1644511149
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1644511149
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1644511149
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1644511149
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1644511149
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1644511149
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1644511149
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1644511149
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1644511149
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1644511149
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1644511149
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1644511149
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1644511149
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1644511149
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1644511149
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1644511149
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1644511149
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1644511149
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1644511149
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1644511149
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1644511149
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1644511149
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1644511149
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1644511149
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1644511149
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1644511149
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1644511149
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1644511149
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1644511149
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1644511149
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1644511149
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1644511149
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1644511149
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1644511149
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1644511149
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1644511149
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1644511149
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1644511149
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1644511149
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1644511149
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1644511149
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1644511149
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1644511149
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1644511149
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1644511149
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1644511149
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1644511149
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1644511149
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1644511149
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1644511149
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1644511149
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1644511149
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1644511149
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1644511149
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1644511149
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1644511149
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1644511149
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1644511149
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1644511149
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1644511149
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1644511149
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1644511149
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1644511149
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1644511149
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1644511149
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1644511149
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1644511149
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1644511149
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1644511149
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1644511149
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1644511149
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1644511149
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1644511149
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1644511149
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1644511149
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1644511149
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1644511149
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1644511149
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1644511149
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1644511149
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1644511149
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1644511149
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1644511149
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1644511149
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1644511149
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1644511149
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1644511149
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1644511149
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1644511149
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1644511149
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1644511149
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1644511149
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1644511149
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1644511149
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1644511149
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1644511149
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1644511149
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1644511149
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1644511149
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1644511149
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1644511149
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1644511149
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1644511149
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1644511149
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1644511149
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1644511149
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1644511149
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1644511149
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1644511149
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1644511149
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1644511149
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1644511149
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1644511149
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1644511149
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1644511149
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1644511149
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1644511149
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1644511149
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1644511149
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1644511149
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1644511149
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1644511149
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1644511149
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1644511149
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1644511149
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1644511149
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1644511149
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1644511149
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1644511149
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1644511149
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1644511149
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1644511149
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1644511149
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1644511149
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1644511149
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1644511149
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1644511149
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1644511149
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1644511149
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1644511149
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1644511149
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1644511149
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1644511149
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1644511149
transform 1 0 6256 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1644511149
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1644511149
transform 1 0 11408 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1644511149
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1644511149
transform 1 0 16560 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1644511149
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1644511149
transform 1 0 21712 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1644511149
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1644511149
transform 1 0 26864 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1644511149
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1644511149
transform 1 0 32016 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1644511149
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1644511149
transform 1 0 37168 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1644511149
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1644511149
transform 1 0 42320 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1644511149
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1644511149
transform 1 0 47472 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0855_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5520 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0856_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15824 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _0857_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15640 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  _0858_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16560 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _0859_
timestamp 1644511149
transform 1 0 47564 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0860_
timestamp 1644511149
transform 1 0 2852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0861_
timestamp 1644511149
transform 1 0 47564 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0862_
timestamp 1644511149
transform 1 0 20884 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0863_
timestamp 1644511149
transform 1 0 47564 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0864_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15640 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  _0865_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0866_
timestamp 1644511149
transform 1 0 47564 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0867_
timestamp 1644511149
transform 1 0 47564 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0868_
timestamp 1644511149
transform 1 0 46828 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0869_
timestamp 1644511149
transform 1 0 44988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0870_
timestamp 1644511149
transform 1 0 6992 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _0871_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16468 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0872_
timestamp 1644511149
transform 1 0 46828 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0873_
timestamp 1644511149
transform 1 0 6716 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0874_
timestamp 1644511149
transform 1 0 47288 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0875_
timestamp 1644511149
transform 1 0 46828 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0876_
timestamp 1644511149
transform 1 0 2944 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _0877_
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0878_
timestamp 1644511149
transform 1 0 2116 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0879_
timestamp 1644511149
transform 1 0 36340 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0880_
timestamp 1644511149
transform 1 0 45172 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0881_
timestamp 1644511149
transform 1 0 2116 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0882_
timestamp 1644511149
transform 1 0 44988 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0883_
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0884_
timestamp 1644511149
transform 1 0 2668 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0885_
timestamp 1644511149
transform 1 0 45632 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0886_
timestamp 1644511149
transform 1 0 24104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0887_
timestamp 1644511149
transform 1 0 2116 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0888_
timestamp 1644511149
transform 1 0 47564 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _0889_
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0890_
timestamp 1644511149
transform 1 0 2484 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0891_
timestamp 1644511149
transform 1 0 11592 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0892_
timestamp 1644511149
transform 1 0 42412 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0893_
timestamp 1644511149
transform 1 0 2208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0894_
timestamp 1644511149
transform 1 0 33120 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0895_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16008 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  _0896_
timestamp 1644511149
transform 1 0 17664 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0897_
timestamp 1644511149
transform 1 0 22172 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0898_
timestamp 1644511149
transform 1 0 2024 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0899_
timestamp 1644511149
transform 1 0 2024 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0900_
timestamp 1644511149
transform 1 0 37996 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0901_
timestamp 1644511149
transform 1 0 2024 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0902_
timestamp 1644511149
transform 1 0 16744 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0903_
timestamp 1644511149
transform 1 0 18032 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0904_
timestamp 1644511149
transform 1 0 19320 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0905_
timestamp 1644511149
transform 1 0 20608 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0906_
timestamp 1644511149
transform 1 0 17388 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0907_
timestamp 1644511149
transform 1 0 18400 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0908_
timestamp 1644511149
transform 1 0 19136 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0909_
timestamp 1644511149
transform 1 0 28336 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0910_
timestamp 1644511149
transform 1 0 32568 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0911_
timestamp 1644511149
transform 1 0 30820 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0912_
timestamp 1644511149
transform 1 0 33212 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0913_
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0914_
timestamp 1644511149
transform 1 0 17664 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0915_
timestamp 1644511149
transform 1 0 45632 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0916_
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0917_
timestamp 1644511149
transform 1 0 46644 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0918_
timestamp 1644511149
transform 1 0 23184 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0919_
timestamp 1644511149
transform 1 0 13248 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _0920_
timestamp 1644511149
transform 1 0 18952 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _0921_
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0922_
timestamp 1644511149
transform 1 0 20056 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0923_
timestamp 1644511149
transform 1 0 40756 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0924_
timestamp 1644511149
transform 1 0 46736 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0925_
timestamp 1644511149
transform 1 0 4048 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0926_
timestamp 1644511149
transform 1 0 17388 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  _0927_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 38548 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0928_
timestamp 1644511149
transform 1 0 41676 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0929_
timestamp 1644511149
transform 1 0 46736 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0930_
timestamp 1644511149
transform 1 0 45816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0931_
timestamp 1644511149
transform 1 0 38364 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0932_
timestamp 1644511149
transform 1 0 45816 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0933_
timestamp 1644511149
transform 1 0 37444 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0934_
timestamp 1644511149
transform 1 0 47564 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0935_
timestamp 1644511149
transform 1 0 47564 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0936_
timestamp 1644511149
transform 1 0 46368 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0937_
timestamp 1644511149
transform 1 0 38364 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0938_
timestamp 1644511149
transform 1 0 36524 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _0939_
timestamp 1644511149
transform 1 0 36340 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _0940_
timestamp 1644511149
transform 1 0 12236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0941_
timestamp 1644511149
transform 1 0 46736 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0942_
timestamp 1644511149
transform 1 0 6992 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0943_
timestamp 1644511149
transform 1 0 15732 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0944_
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0945_
timestamp 1644511149
transform 1 0 19136 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0946_
timestamp 1644511149
transform 1 0 16744 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0947_
timestamp 1644511149
transform 1 0 27232 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0948_
timestamp 1644511149
transform 1 0 30452 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0949_
timestamp 1644511149
transform 1 0 3036 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0950_
timestamp 1644511149
transform 1 0 2668 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0951_
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0952_
timestamp 1644511149
transform 1 0 16744 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0953_
timestamp 1644511149
transform 1 0 15916 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0954_
timestamp 1644511149
transform 1 0 29624 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0955_
timestamp 1644511149
transform 1 0 14720 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0956_
timestamp 1644511149
transform 1 0 15364 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0957_
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _0958_
timestamp 1644511149
transform 1 0 14812 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0959_
timestamp 1644511149
transform 1 0 1564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0960_
timestamp 1644511149
transform 1 0 2116 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0961_
timestamp 1644511149
transform 1 0 17572 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0962_
timestamp 1644511149
transform 1 0 18492 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0963_
timestamp 1644511149
transform 1 0 15088 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _0964_
timestamp 1644511149
transform 1 0 14720 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0965_
timestamp 1644511149
transform 1 0 30544 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0966_
timestamp 1644511149
transform 1 0 2668 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0967_
timestamp 1644511149
transform 1 0 46828 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0968_
timestamp 1644511149
transform 1 0 31096 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0969_
timestamp 1644511149
transform 1 0 2116 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _0970_
timestamp 1644511149
transform 1 0 17020 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1644511149
transform 1 0 22816 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0972_
timestamp 1644511149
transform 1 0 2208 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0973_
timestamp 1644511149
transform 1 0 47564 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0974_
timestamp 1644511149
transform 1 0 3128 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0975_
timestamp 1644511149
transform 1 0 46828 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0976_
timestamp 1644511149
transform 1 0 15364 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0977_
timestamp 1644511149
transform 1 0 2024 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0978_
timestamp 1644511149
transform 1 0 15916 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0979_
timestamp 1644511149
transform 1 0 2116 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0980_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17020 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0981_
timestamp 1644511149
transform 1 0 2024 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0982_
timestamp 1644511149
transform 1 0 15364 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0983_
timestamp 1644511149
transform 1 0 13800 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0984_
timestamp 1644511149
transform 1 0 10764 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0985_
timestamp 1644511149
transform 1 0 11776 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0986_
timestamp 1644511149
transform 1 0 32108 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0987_
timestamp 1644511149
transform 1 0 31372 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0988_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35880 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__buf_6  _0989_
timestamp 1644511149
transform 1 0 36432 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0990_
timestamp 1644511149
transform 1 0 46460 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0991_
timestamp 1644511149
transform 1 0 46828 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0992_
timestamp 1644511149
transform 1 0 2760 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0993_
timestamp 1644511149
transform 1 0 3036 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0994_
timestamp 1644511149
transform 1 0 3404 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0995_
timestamp 1644511149
transform 1 0 36248 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0996_
timestamp 1644511149
transform 1 0 36432 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0997_
timestamp 1644511149
transform 1 0 44988 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0998_
timestamp 1644511149
transform 1 0 39836 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0999_
timestamp 1644511149
transform 1 0 35236 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1000_
timestamp 1644511149
transform 1 0 36432 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1001_
timestamp 1644511149
transform 1 0 36248 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _1002_
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1003_
timestamp 1644511149
transform 1 0 37904 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1004_
timestamp 1644511149
transform 1 0 46644 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1005_
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1006_
timestamp 1644511149
transform 1 0 45448 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1007_
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1008_
timestamp 1644511149
transform 1 0 38548 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1009_
timestamp 1644511149
transform 1 0 39100 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1010_
timestamp 1644511149
transform 1 0 39100 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1011_
timestamp 1644511149
transform 1 0 38548 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1012_
timestamp 1644511149
transform 1 0 36524 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1013_
timestamp 1644511149
transform 1 0 35512 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1014_
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1015_
timestamp 1644511149
transform 1 0 35604 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1016_
timestamp 1644511149
transform 1 0 15548 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1017_
timestamp 1644511149
transform 1 0 36432 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1018_
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1019_
timestamp 1644511149
transform 1 0 10672 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _1020_
timestamp 1644511149
transform 1 0 10212 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1021_
timestamp 1644511149
transform 1 0 4876 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1022_
timestamp 1644511149
transform 1 0 32844 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1023_
timestamp 1644511149
transform 1 0 14260 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1024_
timestamp 1644511149
transform 1 0 2208 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1025_
timestamp 1644511149
transform 1 0 2208 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  _1026_
timestamp 1644511149
transform 1 0 11132 0 1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _1027_
timestamp 1644511149
transform 1 0 2208 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1028_
timestamp 1644511149
transform 1 0 46644 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1029_
timestamp 1644511149
transform 1 0 44160 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1030_
timestamp 1644511149
transform 1 0 2208 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1031_
timestamp 1644511149
transform 1 0 27784 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _1032_
timestamp 1644511149
transform 1 0 11868 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _1033_
timestamp 1644511149
transform 1 0 46828 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1034_
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1035_
timestamp 1644511149
transform 1 0 46828 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1036_
timestamp 1644511149
transform 1 0 10120 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1037_
timestamp 1644511149
transform 1 0 12972 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _1038_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11132 0 1 45696
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _1039_
timestamp 1644511149
transform 1 0 26220 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1040_
timestamp 1644511149
transform 1 0 45632 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1041_
timestamp 1644511149
transform 1 0 7452 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1042_
timestamp 1644511149
transform 1 0 35788 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1043_
timestamp 1644511149
transform 1 0 47564 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1044_
timestamp 1644511149
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1045_
timestamp 1644511149
transform 1 0 2208 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1046_
timestamp 1644511149
transform 1 0 39468 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1047_
timestamp 1644511149
transform 1 0 2852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1048_
timestamp 1644511149
transform 1 0 28428 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1049_
timestamp 1644511149
transform 1 0 29532 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1050_
timestamp 1644511149
transform 1 0 15916 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1051_
timestamp 1644511149
transform 1 0 15732 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1052_
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1053_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24932 0 -1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1054_
timestamp 1644511149
transform 1 0 24932 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1055_
timestamp 1644511149
transform 1 0 24012 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1056_
timestamp 1644511149
transform 1 0 28612 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1057_
timestamp 1644511149
transform 1 0 27968 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1058_
timestamp 1644511149
transform 1 0 23460 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1059_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22540 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1060_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24288 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1061_
timestamp 1644511149
transform 1 0 24656 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1062_
timestamp 1644511149
transform 1 0 24288 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1063_
timestamp 1644511149
transform 1 0 25576 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1064_
timestamp 1644511149
transform 1 0 23828 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1065_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25208 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1066_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22080 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1067_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23184 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1068_
timestamp 1644511149
transform 1 0 28612 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1069_
timestamp 1644511149
transform 1 0 22908 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1070_
timestamp 1644511149
transform 1 0 23184 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1071_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23184 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1072_
timestamp 1644511149
transform 1 0 34224 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1073_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1074_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27600 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1075_
timestamp 1644511149
transform 1 0 28244 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1076_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28428 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1077_
timestamp 1644511149
transform 1 0 30820 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1078_
timestamp 1644511149
transform 1 0 32108 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _1079_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1080_
timestamp 1644511149
transform 1 0 33028 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1081_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28428 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1082_
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1083_
timestamp 1644511149
transform 1 0 23184 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1084_
timestamp 1644511149
transform 1 0 25484 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1085_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24932 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1086_
timestamp 1644511149
transform 1 0 23368 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1087_
timestamp 1644511149
transform 1 0 26220 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1088_
timestamp 1644511149
transform 1 0 28704 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _1089_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23276 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1090_
timestamp 1644511149
transform 1 0 23276 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_1  _1091_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22724 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1092_
timestamp 1644511149
transform 1 0 40020 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1093_
timestamp 1644511149
transform 1 0 43608 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1094_
timestamp 1644511149
transform 1 0 42320 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1095_
timestamp 1644511149
transform 1 0 40940 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1096_
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1097_
timestamp 1644511149
transform 1 0 39928 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1098_
timestamp 1644511149
transform 1 0 43056 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1099_
timestamp 1644511149
transform 1 0 43056 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1100_
timestamp 1644511149
transform 1 0 40756 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1101_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 41124 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1102_
timestamp 1644511149
transform 1 0 17480 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1103_
timestamp 1644511149
transform 1 0 29440 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1104_
timestamp 1644511149
transform 1 0 25944 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1105_
timestamp 1644511149
transform 1 0 19688 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1106_
timestamp 1644511149
transform 1 0 19688 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1107_
timestamp 1644511149
transform 1 0 20332 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_2  _1108_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 47472 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1109_
timestamp 1644511149
transform 1 0 28336 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _1110_
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1111_
timestamp 1644511149
transform 1 0 28152 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1112_
timestamp 1644511149
transform 1 0 20516 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _1113_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35052 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1114_
timestamp 1644511149
transform 1 0 19688 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1115_
timestamp 1644511149
transform 1 0 19872 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1116_
timestamp 1644511149
transform 1 0 20608 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_4  _1117_
timestamp 1644511149
transform 1 0 27140 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1118_
timestamp 1644511149
transform 1 0 27416 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1119_
timestamp 1644511149
transform 1 0 29900 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1120_
timestamp 1644511149
transform 1 0 30176 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1121_
timestamp 1644511149
transform 1 0 27416 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1122_
timestamp 1644511149
transform 1 0 24472 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1123_
timestamp 1644511149
transform 1 0 24932 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1124_
timestamp 1644511149
transform 1 0 27600 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1125_
timestamp 1644511149
transform 1 0 27968 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1126_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24932 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1127_
timestamp 1644511149
transform 1 0 34960 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1128_
timestamp 1644511149
transform 1 0 28244 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1129_
timestamp 1644511149
transform 1 0 29716 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1130_
timestamp 1644511149
transform 1 0 30820 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1131_
timestamp 1644511149
transform 1 0 31648 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1132_
timestamp 1644511149
transform 1 0 35604 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1133_
timestamp 1644511149
transform 1 0 32752 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1134_
timestamp 1644511149
transform 1 0 33120 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1135_
timestamp 1644511149
transform 1 0 32384 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1136_
timestamp 1644511149
transform 1 0 32936 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1137_
timestamp 1644511149
transform 1 0 31188 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1138_
timestamp 1644511149
transform 1 0 30084 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1139_
timestamp 1644511149
transform 1 0 30452 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1140_
timestamp 1644511149
transform 1 0 37076 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1141_
timestamp 1644511149
transform 1 0 28152 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1142_
timestamp 1644511149
transform 1 0 28888 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1143_
timestamp 1644511149
transform 1 0 35420 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1144_
timestamp 1644511149
transform 1 0 28704 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1145_
timestamp 1644511149
transform 1 0 36064 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1146_
timestamp 1644511149
transform 1 0 35236 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1147_
timestamp 1644511149
transform 1 0 36064 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1148_
timestamp 1644511149
transform 1 0 29624 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1149_
timestamp 1644511149
transform 1 0 29716 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1150_
timestamp 1644511149
transform 1 0 35144 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1151_
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1152_
timestamp 1644511149
transform 1 0 33672 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1153_
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1154_
timestamp 1644511149
transform 1 0 29900 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1155_
timestamp 1644511149
transform 1 0 28520 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1156_
timestamp 1644511149
transform 1 0 20792 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1157_
timestamp 1644511149
transform 1 0 28428 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1158_
timestamp 1644511149
transform 1 0 22448 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1159_
timestamp 1644511149
transform 1 0 27600 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1160_
timestamp 1644511149
transform 1 0 27692 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1161_
timestamp 1644511149
transform 1 0 29808 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1162_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29808 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1163_
timestamp 1644511149
transform 1 0 20884 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1164_
timestamp 1644511149
transform 1 0 20608 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1165_
timestamp 1644511149
transform 1 0 23644 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1166_
timestamp 1644511149
transform 1 0 23368 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1167_
timestamp 1644511149
transform 1 0 28612 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1168_
timestamp 1644511149
transform 1 0 29808 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1169_
timestamp 1644511149
transform 1 0 30360 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1170_
timestamp 1644511149
transform 1 0 30084 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1171_
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1172_
timestamp 1644511149
transform 1 0 27416 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1173_
timestamp 1644511149
transform 1 0 29348 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1174_
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1175_
timestamp 1644511149
transform 1 0 33488 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1176_
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1177_
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1178_
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1179_
timestamp 1644511149
transform 1 0 31096 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1180_
timestamp 1644511149
transform 1 0 30912 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1181_
timestamp 1644511149
transform 1 0 29900 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1182_
timestamp 1644511149
transform 1 0 30268 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1183_
timestamp 1644511149
transform 1 0 26036 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1184_
timestamp 1644511149
transform 1 0 25852 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1185_
timestamp 1644511149
transform 1 0 25024 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1186_
timestamp 1644511149
transform 1 0 26128 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1187_
timestamp 1644511149
transform 1 0 25024 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1188_
timestamp 1644511149
transform 1 0 24840 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1189_
timestamp 1644511149
transform 1 0 24564 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1190_
timestamp 1644511149
transform 1 0 26956 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1191_
timestamp 1644511149
transform 1 0 26956 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _1192_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27968 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1193_
timestamp 1644511149
transform 1 0 27968 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1194_
timestamp 1644511149
transform 1 0 29348 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1195_
timestamp 1644511149
transform 1 0 18768 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1196_
timestamp 1644511149
transform 1 0 19688 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1197_
timestamp 1644511149
transform 1 0 20608 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1198_
timestamp 1644511149
transform 1 0 19596 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1199_
timestamp 1644511149
transform 1 0 20608 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1200_
timestamp 1644511149
transform 1 0 20700 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1201_
timestamp 1644511149
transform 1 0 16192 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1202_
timestamp 1644511149
transform 1 0 28336 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1203_
timestamp 1644511149
transform 1 0 26128 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1204_
timestamp 1644511149
transform 1 0 23644 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _1205_
timestamp 1644511149
transform 1 0 24104 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1206_
timestamp 1644511149
transform 1 0 22448 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1207_
timestamp 1644511149
transform 1 0 22816 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1208_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21988 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1209_
timestamp 1644511149
transform 1 0 22080 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1210_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1211_
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1212_
timestamp 1644511149
transform 1 0 21068 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1213_
timestamp 1644511149
transform 1 0 22816 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1214_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1215_
timestamp 1644511149
transform 1 0 19964 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1216_
timestamp 1644511149
transform 1 0 20056 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1217_
timestamp 1644511149
transform 1 0 24564 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1218_
timestamp 1644511149
transform 1 0 21620 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1219_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1220_
timestamp 1644511149
transform 1 0 25208 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1221_
timestamp 1644511149
transform 1 0 27140 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1222_
timestamp 1644511149
transform 1 0 21252 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1223_
timestamp 1644511149
transform 1 0 23092 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__or3b_1  _1224_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22816 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1225_
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1226_
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1227_
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1228_
timestamp 1644511149
transform 1 0 24564 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1229_
timestamp 1644511149
transform 1 0 26312 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1230_
timestamp 1644511149
transform 1 0 23828 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1231_
timestamp 1644511149
transform 1 0 22908 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1232_
timestamp 1644511149
transform 1 0 23000 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1233_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22816 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1234_
timestamp 1644511149
transform 1 0 22080 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1235_
timestamp 1644511149
transform 1 0 22356 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1236_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21252 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1237_
timestamp 1644511149
transform 1 0 21988 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1238_
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1239_
timestamp 1644511149
transform 1 0 23368 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1240_
timestamp 1644511149
transform 1 0 26220 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1241_
timestamp 1644511149
transform 1 0 24380 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1242_
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1243_
timestamp 1644511149
transform 1 0 26680 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1244_
timestamp 1644511149
transform 1 0 24748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1245_
timestamp 1644511149
transform 1 0 27140 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1246_
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1247_
timestamp 1644511149
transform 1 0 26036 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1248_
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1249_
timestamp 1644511149
transform 1 0 27140 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1250_
timestamp 1644511149
transform 1 0 25668 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or4_2  _1251_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25208 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1252_
timestamp 1644511149
transform 1 0 23736 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1253_
timestamp 1644511149
transform 1 0 25576 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1254_
timestamp 1644511149
transform 1 0 25392 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1255_
timestamp 1644511149
transform 1 0 24932 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1256_
timestamp 1644511149
transform 1 0 27232 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1257_
timestamp 1644511149
transform 1 0 25484 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1258_
timestamp 1644511149
transform 1 0 25300 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1259_
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1260_
timestamp 1644511149
transform 1 0 27232 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1261_
timestamp 1644511149
transform 1 0 27324 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1262_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26404 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1263_
timestamp 1644511149
transform 1 0 28612 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1264_
timestamp 1644511149
transform 1 0 27416 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1265_
timestamp 1644511149
transform 1 0 27416 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1266_
timestamp 1644511149
transform 1 0 25944 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1267_
timestamp 1644511149
transform 1 0 26036 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1268_
timestamp 1644511149
transform 1 0 26404 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1269_
timestamp 1644511149
transform 1 0 27508 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1270_
timestamp 1644511149
transform 1 0 25944 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_1  _1271_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25392 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1272_
timestamp 1644511149
transform 1 0 25024 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1273_
timestamp 1644511149
transform 1 0 25024 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1274_
timestamp 1644511149
transform 1 0 25484 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1275_
timestamp 1644511149
transform 1 0 25668 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1276_
timestamp 1644511149
transform 1 0 19964 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1277_
timestamp 1644511149
transform 1 0 20608 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1278_
timestamp 1644511149
transform 1 0 25300 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1279_
timestamp 1644511149
transform 1 0 25668 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1280_
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1281_
timestamp 1644511149
transform 1 0 26312 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1282_
timestamp 1644511149
transform 1 0 27140 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1283_
timestamp 1644511149
transform 1 0 25116 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1284_
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1285_
timestamp 1644511149
transform 1 0 26588 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1286_
timestamp 1644511149
transform 1 0 24932 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1287_
timestamp 1644511149
transform 1 0 25208 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1288_
timestamp 1644511149
transform 1 0 20240 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1289_
timestamp 1644511149
transform 1 0 19780 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1290_
timestamp 1644511149
transform 1 0 22724 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1291_
timestamp 1644511149
transform 1 0 21896 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _1292_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22540 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1293_
timestamp 1644511149
transform 1 0 22816 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1294_
timestamp 1644511149
transform 1 0 21988 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1295_
timestamp 1644511149
transform 1 0 28428 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1296_
timestamp 1644511149
transform 1 0 22816 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1297_
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1298_
timestamp 1644511149
transform 1 0 23736 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _1299_
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1300_
timestamp 1644511149
transform 1 0 23644 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1301_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22724 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1302_
timestamp 1644511149
transform 1 0 21896 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1303_
timestamp 1644511149
transform 1 0 35420 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1304_
timestamp 1644511149
transform 1 0 30084 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1305_
timestamp 1644511149
transform 1 0 28980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1306_
timestamp 1644511149
transform 1 0 28244 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1307_
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1308_
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1309_
timestamp 1644511149
transform 1 0 20240 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1310_
timestamp 1644511149
transform 1 0 22908 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1311_
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1312_
timestamp 1644511149
transform 1 0 25484 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_2  _1313_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25300 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1314_
timestamp 1644511149
transform 1 0 22448 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1315_
timestamp 1644511149
transform 1 0 25852 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1316_
timestamp 1644511149
transform 1 0 25668 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1317_
timestamp 1644511149
transform 1 0 33672 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1318_
timestamp 1644511149
transform 1 0 39836 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1319_
timestamp 1644511149
transform 1 0 40296 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1320_
timestamp 1644511149
transform 1 0 35696 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1321_
timestamp 1644511149
transform 1 0 36800 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__xor2_1  _1322_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 36800 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1323_
timestamp 1644511149
transform 1 0 38640 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1324_
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1325_
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1326_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 37996 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1327_
timestamp 1644511149
transform 1 0 36248 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1328_
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1329_
timestamp 1644511149
transform 1 0 38272 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1330_
timestamp 1644511149
transform 1 0 39100 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1331_
timestamp 1644511149
transform 1 0 38180 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1332_
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1333_
timestamp 1644511149
transform 1 0 37904 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1334_
timestamp 1644511149
transform 1 0 38272 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1335_
timestamp 1644511149
transform 1 0 35788 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1336_
timestamp 1644511149
transform 1 0 36156 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1337_
timestamp 1644511149
transform 1 0 37628 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1338_
timestamp 1644511149
transform 1 0 38456 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1339_
timestamp 1644511149
transform 1 0 38732 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1340_
timestamp 1644511149
transform 1 0 39652 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1341_
timestamp 1644511149
transform 1 0 38180 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1342_
timestamp 1644511149
transform 1 0 38456 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1343_
timestamp 1644511149
transform 1 0 36340 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1344_
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1345_
timestamp 1644511149
transform 1 0 38088 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1346_
timestamp 1644511149
transform 1 0 37076 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _1347_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 37352 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o41a_1  _1348_
timestamp 1644511149
transform 1 0 37444 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1349_
timestamp 1644511149
transform 1 0 40756 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1350_
timestamp 1644511149
transform 1 0 37996 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1351_
timestamp 1644511149
transform 1 0 40572 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1352_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 39928 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1353_
timestamp 1644511149
transform 1 0 40112 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1354_
timestamp 1644511149
transform 1 0 43148 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1355_
timestamp 1644511149
transform 1 0 41400 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1356_
timestamp 1644511149
transform 1 0 41584 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1357_
timestamp 1644511149
transform 1 0 41676 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1358_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 42412 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1359_
timestamp 1644511149
transform 1 0 41308 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1360_
timestamp 1644511149
transform 1 0 41860 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1361_
timestamp 1644511149
transform 1 0 43792 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1362_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 40112 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1363_
timestamp 1644511149
transform 1 0 41308 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1364_
timestamp 1644511149
transform 1 0 40572 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1365_
timestamp 1644511149
transform 1 0 41676 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1366_
timestamp 1644511149
transform 1 0 40204 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1367_
timestamp 1644511149
transform 1 0 41676 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1368_
timestamp 1644511149
transform 1 0 41032 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1369_
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1370_
timestamp 1644511149
transform 1 0 40204 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1371_
timestamp 1644511149
transform 1 0 41124 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1372_
timestamp 1644511149
transform 1 0 41032 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1373_
timestamp 1644511149
transform 1 0 41952 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1374_
timestamp 1644511149
transform 1 0 41216 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1375_
timestamp 1644511149
transform 1 0 40572 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1376_
timestamp 1644511149
transform 1 0 41400 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1377_
timestamp 1644511149
transform 1 0 41216 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1378_
timestamp 1644511149
transform 1 0 40296 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1379_
timestamp 1644511149
transform 1 0 39836 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1380_
timestamp 1644511149
transform 1 0 41952 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1381_
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1382_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26772 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1383_
timestamp 1644511149
transform 1 0 26312 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1384_
timestamp 1644511149
transform 1 0 25576 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1385_
timestamp 1644511149
transform 1 0 27324 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1386_
timestamp 1644511149
transform 1 0 27324 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1387_
timestamp 1644511149
transform 1 0 23092 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1388_
timestamp 1644511149
transform 1 0 18124 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1389_
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1390_
timestamp 1644511149
transform 1 0 22172 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1391_
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1392_
timestamp 1644511149
transform 1 0 19320 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1393_
timestamp 1644511149
transform 1 0 17756 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1394_
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1395_
timestamp 1644511149
transform 1 0 22816 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1396_
timestamp 1644511149
transform 1 0 18492 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1397_
timestamp 1644511149
transform 1 0 18216 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1398_
timestamp 1644511149
transform 1 0 16836 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1399_
timestamp 1644511149
transform 1 0 20516 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1400_
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1401_
timestamp 1644511149
transform 1 0 20516 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1402_
timestamp 1644511149
transform 1 0 22816 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1403_
timestamp 1644511149
transform 1 0 21988 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1404_
timestamp 1644511149
transform 1 0 21988 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1405_
timestamp 1644511149
transform 1 0 21528 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1406_
timestamp 1644511149
transform 1 0 23276 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1407_
timestamp 1644511149
transform 1 0 19412 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1408_
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1409_
timestamp 1644511149
transform 1 0 20792 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1410_
timestamp 1644511149
transform 1 0 18032 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1411_
timestamp 1644511149
transform 1 0 22448 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1412_
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1413_
timestamp 1644511149
transform 1 0 20424 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1414_
timestamp 1644511149
transform 1 0 21160 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1415_
timestamp 1644511149
transform 1 0 22080 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1416_
timestamp 1644511149
transform 1 0 20424 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1417_
timestamp 1644511149
transform 1 0 20056 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1418_
timestamp 1644511149
transform 1 0 19596 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1419_
timestamp 1644511149
transform 1 0 19320 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1420_
timestamp 1644511149
transform 1 0 18032 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1421_
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1422_
timestamp 1644511149
transform 1 0 20884 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1423_
timestamp 1644511149
transform 1 0 20608 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1424_
timestamp 1644511149
transform 1 0 22080 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1425_
timestamp 1644511149
transform 1 0 24564 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1426_
timestamp 1644511149
transform 1 0 20424 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1427_
timestamp 1644511149
transform 1 0 20332 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1428_
timestamp 1644511149
transform 1 0 19504 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1429_
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1430_
timestamp 1644511149
transform 1 0 20516 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1431_
timestamp 1644511149
transform 1 0 19596 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1432_
timestamp 1644511149
transform 1 0 20148 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1433_
timestamp 1644511149
transform 1 0 26220 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1434_
timestamp 1644511149
transform 1 0 24288 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1435_
timestamp 1644511149
transform 1 0 23460 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1436_
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1437_
timestamp 1644511149
transform 1 0 24288 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1438_
timestamp 1644511149
transform 1 0 22632 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1439_
timestamp 1644511149
transform 1 0 23184 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1440_
timestamp 1644511149
transform 1 0 24012 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1441_
timestamp 1644511149
transform 1 0 23460 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1442_
timestamp 1644511149
transform 1 0 21988 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1443_
timestamp 1644511149
transform 1 0 26588 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1444_
timestamp 1644511149
transform 1 0 25300 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1445_
timestamp 1644511149
transform 1 0 24656 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1446_
timestamp 1644511149
transform 1 0 25116 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1447_
timestamp 1644511149
transform 1 0 27600 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1448_
timestamp 1644511149
transform 1 0 28152 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1449_
timestamp 1644511149
transform 1 0 24012 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1450_
timestamp 1644511149
transform 1 0 24932 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1451_
timestamp 1644511149
transform 1 0 25944 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1452_
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1453_
timestamp 1644511149
transform 1 0 26220 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1454_
timestamp 1644511149
transform 1 0 27600 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1455_
timestamp 1644511149
transform 1 0 28796 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1456_
timestamp 1644511149
transform 1 0 26680 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1457_
timestamp 1644511149
transform 1 0 27784 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1458_
timestamp 1644511149
transform 1 0 26036 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1459_
timestamp 1644511149
transform 1 0 27876 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1460_
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1461_
timestamp 1644511149
transform 1 0 26036 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1462_
timestamp 1644511149
transform 1 0 24564 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1463_
timestamp 1644511149
transform 1 0 28244 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1464_
timestamp 1644511149
transform 1 0 28152 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1465_
timestamp 1644511149
transform 1 0 36064 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1466_
timestamp 1644511149
transform 1 0 27048 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1467_
timestamp 1644511149
transform 1 0 27508 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1468_
timestamp 1644511149
transform 1 0 26680 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1469_
timestamp 1644511149
transform 1 0 26772 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1470_
timestamp 1644511149
transform 1 0 31096 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1471_
timestamp 1644511149
transform 1 0 31556 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1472_
timestamp 1644511149
transform 1 0 32384 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1473_
timestamp 1644511149
transform 1 0 30820 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1474_
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1475_
timestamp 1644511149
transform 1 0 32384 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1476_
timestamp 1644511149
transform 1 0 29348 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1477_
timestamp 1644511149
transform 1 0 29164 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1478_
timestamp 1644511149
transform 1 0 31740 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1479_
timestamp 1644511149
transform 1 0 32292 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1480_
timestamp 1644511149
transform 1 0 31924 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1481_
timestamp 1644511149
transform 1 0 32200 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1482_
timestamp 1644511149
transform 1 0 31924 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1483_
timestamp 1644511149
transform 1 0 29900 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1484_
timestamp 1644511149
transform 1 0 29808 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1485_
timestamp 1644511149
transform 1 0 31004 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1486_
timestamp 1644511149
transform 1 0 30084 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1487_
timestamp 1644511149
transform 1 0 30360 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1488_
timestamp 1644511149
transform 1 0 30452 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1489_
timestamp 1644511149
transform 1 0 28612 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1490_
timestamp 1644511149
transform 1 0 28796 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1491_
timestamp 1644511149
transform 1 0 28612 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1492_
timestamp 1644511149
transform 1 0 29716 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1493_
timestamp 1644511149
transform 1 0 29808 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1494_
timestamp 1644511149
transform 1 0 27784 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1495_
timestamp 1644511149
transform 1 0 29624 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1496_
timestamp 1644511149
transform 1 0 20976 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1497_
timestamp 1644511149
transform 1 0 17664 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1498_
timestamp 1644511149
transform 1 0 18032 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1499_
timestamp 1644511149
transform 1 0 23000 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1500_
timestamp 1644511149
transform 1 0 18216 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1501_
timestamp 1644511149
transform 1 0 19136 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1502_
timestamp 1644511149
transform 1 0 20240 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1503_
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1504_
timestamp 1644511149
transform 1 0 20884 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1505_
timestamp 1644511149
transform 1 0 21344 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1506_
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1507_
timestamp 1644511149
transform 1 0 23368 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1508_
timestamp 1644511149
transform 1 0 23368 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1509_
timestamp 1644511149
transform 1 0 22264 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1510_
timestamp 1644511149
transform 1 0 25484 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1511_
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1512_
timestamp 1644511149
transform 1 0 24656 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1513_
timestamp 1644511149
transform 1 0 24288 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1514_
timestamp 1644511149
transform 1 0 38732 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1515_
timestamp 1644511149
transform 1 0 37444 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1516_
timestamp 1644511149
transform 1 0 42596 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1517_
timestamp 1644511149
transform 1 0 43240 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1518_
timestamp 1644511149
transform 1 0 44068 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1519_
timestamp 1644511149
transform 1 0 42964 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1520_
timestamp 1644511149
transform 1 0 45264 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1521_
timestamp 1644511149
transform 1 0 37628 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1522_
timestamp 1644511149
transform 1 0 44988 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1523_
timestamp 1644511149
transform 1 0 45080 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1524_
timestamp 1644511149
transform 1 0 44988 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1525_
timestamp 1644511149
transform 1 0 44068 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1526_
timestamp 1644511149
transform 1 0 44988 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1527_
timestamp 1644511149
transform 1 0 45540 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1528_
timestamp 1644511149
transform 1 0 44436 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1529_
timestamp 1644511149
transform 1 0 38640 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1530_
timestamp 1644511149
transform 1 0 38732 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1531_
timestamp 1644511149
transform 1 0 37720 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1532_
timestamp 1644511149
transform 1 0 35880 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1533_
timestamp 1644511149
transform 1 0 36616 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1534_
timestamp 1644511149
transform 1 0 32844 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _1535_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31556 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1536_
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1537_
timestamp 1644511149
transform 1 0 29164 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1538_
timestamp 1644511149
transform 1 0 28612 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1539_
timestamp 1644511149
transform 1 0 19320 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_4  _1540_
timestamp 1644511149
transform 1 0 28244 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1541_
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1542_
timestamp 1644511149
transform 1 0 18308 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1543_
timestamp 1644511149
transform 1 0 18032 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1544_
timestamp 1644511149
transform 1 0 19320 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1545_
timestamp 1644511149
transform 1 0 19412 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1546_
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1547_
timestamp 1644511149
transform 1 0 19596 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1548_
timestamp 1644511149
transform 1 0 18032 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1549_
timestamp 1644511149
transform 1 0 18492 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1550_
timestamp 1644511149
transform 1 0 18308 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1551_
timestamp 1644511149
transform 1 0 30176 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1552_
timestamp 1644511149
transform 1 0 19320 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1553_
timestamp 1644511149
transform 1 0 30360 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1554_
timestamp 1644511149
transform 1 0 30360 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1555_
timestamp 1644511149
transform 1 0 29624 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1556_
timestamp 1644511149
transform 1 0 29072 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1557_
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1558_
timestamp 1644511149
transform 1 0 30912 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1559_
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1560_
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1561_
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1562_
timestamp 1644511149
transform 1 0 30912 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1563_
timestamp 1644511149
transform 1 0 32384 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1564_
timestamp 1644511149
transform 1 0 30728 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1565_
timestamp 1644511149
transform 1 0 31280 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1566_
timestamp 1644511149
transform 1 0 30820 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1567_
timestamp 1644511149
transform 1 0 31372 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1568_
timestamp 1644511149
transform 1 0 33856 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1569_
timestamp 1644511149
transform 1 0 33396 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1570_
timestamp 1644511149
transform 1 0 30728 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1571_
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1572_
timestamp 1644511149
transform 1 0 34224 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1573_
timestamp 1644511149
transform 1 0 33304 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1574_
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1575_
timestamp 1644511149
transform 1 0 30912 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1576_
timestamp 1644511149
transform 1 0 33764 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1577_
timestamp 1644511149
transform 1 0 30912 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1578_
timestamp 1644511149
transform 1 0 33120 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1579_
timestamp 1644511149
transform 1 0 31372 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1580_
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1581_
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1582_
timestamp 1644511149
transform 1 0 32752 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1583_
timestamp 1644511149
transform 1 0 30820 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1584_
timestamp 1644511149
transform 1 0 30912 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1585_
timestamp 1644511149
transform 1 0 32108 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1586_
timestamp 1644511149
transform 1 0 32200 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1587_
timestamp 1644511149
transform 1 0 31924 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1588_
timestamp 1644511149
transform 1 0 33304 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1589_
timestamp 1644511149
transform 1 0 30084 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1590_
timestamp 1644511149
transform 1 0 29072 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1591_
timestamp 1644511149
transform 1 0 29900 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1592_
timestamp 1644511149
transform 1 0 19136 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1593_
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1594_
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1595_
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1596_
timestamp 1644511149
transform 1 0 17112 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1597_
timestamp 1644511149
transform 1 0 17940 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1598_
timestamp 1644511149
transform 1 0 18124 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1599_
timestamp 1644511149
transform 1 0 17940 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1600_
timestamp 1644511149
transform 1 0 18308 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1601_
timestamp 1644511149
transform 1 0 17940 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1602_
timestamp 1644511149
transform 1 0 17388 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1603_
timestamp 1644511149
transform 1 0 18216 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1604_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15272 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1605_
timestamp 1644511149
transform 1 0 32752 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1606_
timestamp 1644511149
transform 1 0 29716 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1607_
timestamp 1644511149
transform 1 0 21896 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1608_
timestamp 1644511149
transform 1 0 22448 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1609_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22356 0 -1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1610_
timestamp 1644511149
transform 1 0 24932 0 -1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1611_
timestamp 1644511149
transform 1 0 32752 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1612_
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1613_
timestamp 1644511149
transform 1 0 33212 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1614_
timestamp 1644511149
transform 1 0 30176 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1615_
timestamp 1644511149
transform 1 0 36248 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1616_
timestamp 1644511149
transform 1 0 36340 0 1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1617_
timestamp 1644511149
transform 1 0 30176 0 1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1618_
timestamp 1644511149
transform 1 0 35972 0 1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1619_
timestamp 1644511149
transform 1 0 33212 0 -1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1620_
timestamp 1644511149
transform 1 0 20608 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1621_
timestamp 1644511149
transform 1 0 27140 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1622_
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1623_
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1624_
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1625_
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1626_
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1627_
timestamp 1644511149
transform 1 0 34408 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1628_
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1629_
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1630_
timestamp 1644511149
transform 1 0 30544 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1631_
timestamp 1644511149
transform 1 0 25300 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1632_
timestamp 1644511149
transform 1 0 25024 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1633_
timestamp 1644511149
transform 1 0 24656 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1634_
timestamp 1644511149
transform 1 0 27324 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1635_
timestamp 1644511149
transform 1 0 16192 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1636_
timestamp 1644511149
transform 1 0 20240 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1637_
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1638_
timestamp 1644511149
transform 1 0 20424 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1639_
timestamp 1644511149
transform 1 0 22356 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1640_
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1641_
timestamp 1644511149
transform 1 0 23460 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1642_
timestamp 1644511149
transform 1 0 27416 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1643_
timestamp 1644511149
transform 1 0 25208 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1644_
timestamp 1644511149
transform 1 0 27784 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1645_
timestamp 1644511149
transform 1 0 28244 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1646_
timestamp 1644511149
transform 1 0 27600 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1647_
timestamp 1644511149
transform 1 0 18952 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1648_
timestamp 1644511149
transform 1 0 27416 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1649_
timestamp 1644511149
transform 1 0 19320 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1650_
timestamp 1644511149
transform 1 0 20608 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1651_
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1652_
timestamp 1644511149
transform 1 0 33580 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1653_
timestamp 1644511149
transform 1 0 26772 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1654_
timestamp 1644511149
transform 1 0 39468 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1655_
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1656_
timestamp 1644511149
transform 1 0 42872 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1657_
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1658_
timestamp 1644511149
transform 1 0 42044 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1659_
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1660_
timestamp 1644511149
transform 1 0 40112 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1661_
timestamp 1644511149
transform 1 0 40296 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1662_
timestamp 1644511149
transform 1 0 16560 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1663_
timestamp 1644511149
transform 1 0 16744 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1664_
timestamp 1644511149
transform 1 0 17112 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1665_
timestamp 1644511149
transform 1 0 20148 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1666_
timestamp 1644511149
transform 1 0 22172 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1667_
timestamp 1644511149
transform 1 0 18124 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1668_
timestamp 1644511149
transform 1 0 21528 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1669_
timestamp 1644511149
transform 1 0 20608 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1670_
timestamp 1644511149
transform 1 0 18032 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1671_
timestamp 1644511149
transform 1 0 20792 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1672_
timestamp 1644511149
transform 1 0 18032 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1673_
timestamp 1644511149
transform 1 0 19780 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1674_
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1675_
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1676_
timestamp 1644511149
transform 1 0 22172 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1677_
timestamp 1644511149
transform 1 0 23920 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1678_
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1679_
timestamp 1644511149
transform 1 0 26956 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1680_
timestamp 1644511149
transform 1 0 27508 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1681_
timestamp 1644511149
transform 1 0 24748 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1682_
timestamp 1644511149
transform 1 0 27324 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1683_
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1684_
timestamp 1644511149
transform 1 0 32568 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1685_
timestamp 1644511149
transform 1 0 32568 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1686_
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1687_
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1688_
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1689_
timestamp 1644511149
transform 1 0 29716 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1690_
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1691_
timestamp 1644511149
transform 1 0 27600 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1692_
timestamp 1644511149
transform 1 0 29900 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1693_
timestamp 1644511149
transform 1 0 29900 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1694_
timestamp 1644511149
transform 1 0 15916 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1695_
timestamp 1644511149
transform 1 0 17296 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1696_
timestamp 1644511149
transform 1 0 19412 0 1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1697_
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1698_
timestamp 1644511149
transform 1 0 23828 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1699_
timestamp 1644511149
transform 1 0 22448 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1700_
timestamp 1644511149
transform 1 0 25024 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1701_
timestamp 1644511149
transform 1 0 24932 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1702_
timestamp 1644511149
transform 1 0 37260 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1703_
timestamp 1644511149
transform 1 0 43516 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1704_
timestamp 1644511149
transform 1 0 45448 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1705_
timestamp 1644511149
transform 1 0 45080 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1706_
timestamp 1644511149
transform 1 0 44528 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1707_
timestamp 1644511149
transform 1 0 45080 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1708_
timestamp 1644511149
transform 1 0 39560 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1709_
timestamp 1644511149
transform 1 0 36432 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1710_
timestamp 1644511149
transform 1 0 31096 0 1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1711_
timestamp 1644511149
transform 1 0 16468 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1712_
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1713_
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1714_
timestamp 1644511149
transform 1 0 16836 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1715_
timestamp 1644511149
transform 1 0 17572 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1716_
timestamp 1644511149
transform 1 0 28980 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1717_
timestamp 1644511149
transform 1 0 31556 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1718_
timestamp 1644511149
transform 1 0 30176 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1719_
timestamp 1644511149
transform 1 0 31464 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1720_
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1721_
timestamp 1644511149
transform 1 0 34132 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1722_
timestamp 1644511149
transform 1 0 31556 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1723_
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1724_
timestamp 1644511149
transform 1 0 31004 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1725_
timestamp 1644511149
transform 1 0 33948 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1726_
timestamp 1644511149
transform 1 0 33856 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1727_
timestamp 1644511149
transform 1 0 30084 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1728_
timestamp 1644511149
transform 1 0 32660 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1729_
timestamp 1644511149
transform 1 0 32752 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1730_
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1731_
timestamp 1644511149
transform 1 0 19228 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1732_
timestamp 1644511149
transform 1 0 16284 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1733_
timestamp 1644511149
transform 1 0 16744 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1734_
timestamp 1644511149
transform 1 0 15732 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1735_
timestamp 1644511149
transform 1 0 16836 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1736__200 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 40112 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1737__201
timestamp 1644511149
transform 1 0 32108 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1738__202
timestamp 1644511149
transform 1 0 10120 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1739__203
timestamp 1644511149
transform 1 0 1840 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1740__96
timestamp 1644511149
transform 1 0 4048 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1741__97
timestamp 1644511149
transform 1 0 26220 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1742__98
timestamp 1644511149
transform 1 0 15916 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1743__99
timestamp 1644511149
transform 1 0 25852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1744__100
timestamp 1644511149
transform 1 0 36064 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1745__101
timestamp 1644511149
transform 1 0 2024 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1746__102
timestamp 1644511149
transform 1 0 47564 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1747__103
timestamp 1644511149
transform 1 0 1564 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1748__104
timestamp 1644511149
transform 1 0 1564 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1749__105
timestamp 1644511149
transform 1 0 2116 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1750__106
timestamp 1644511149
transform 1 0 31188 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1751__107
timestamp 1644511149
transform 1 0 15548 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1752__108
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1753__109
timestamp 1644511149
transform 1 0 30820 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1754__110
timestamp 1644511149
transform 1 0 5244 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1755__111
timestamp 1644511149
transform 1 0 47564 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1756__112
timestamp 1644511149
transform 1 0 22540 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1757__113
timestamp 1644511149
transform 1 0 15548 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1758__114
timestamp 1644511149
transform 1 0 28796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1759__115
timestamp 1644511149
transform 1 0 20240 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1760__116
timestamp 1644511149
transform 1 0 41492 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1761__117
timestamp 1644511149
transform 1 0 47564 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1762__118
timestamp 1644511149
transform 1 0 3772 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1763__119
timestamp 1644511149
transform 1 0 41676 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1764__120
timestamp 1644511149
transform 1 0 2852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1765__121
timestamp 1644511149
transform 1 0 1472 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1766__122
timestamp 1644511149
transform 1 0 18216 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1767__123
timestamp 1644511149
transform 1 0 19228 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1768__124
timestamp 1644511149
transform 1 0 14444 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1769__125
timestamp 1644511149
transform 1 0 30268 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1770__126
timestamp 1644511149
transform 1 0 1840 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1771__127
timestamp 1644511149
transform 1 0 47564 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1772__128
timestamp 1644511149
transform 1 0 30268 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1773__129
timestamp 1644511149
transform 1 0 2484 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1774__130
timestamp 1644511149
transform 1 0 21896 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1775__131
timestamp 1644511149
transform 1 0 1840 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1776__132
timestamp 1644511149
transform 1 0 43056 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1777__133
timestamp 1644511149
transform 1 0 1564 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1778__134
timestamp 1644511149
transform 1 0 46828 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1779__135
timestamp 1644511149
transform 1 0 45172 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1780__136
timestamp 1644511149
transform 1 0 46828 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1781__137
timestamp 1644511149
transform 1 0 2852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1782__138
timestamp 1644511149
transform 1 0 35420 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1783__139
timestamp 1644511149
transform 1 0 12512 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1784__140
timestamp 1644511149
transform 1 0 46092 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1785__141
timestamp 1644511149
transform 1 0 44436 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1786__142
timestamp 1644511149
transform 1 0 38640 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1787__143
timestamp 1644511149
transform 1 0 10764 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1788__144
timestamp 1644511149
transform 1 0 7268 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1789__145
timestamp 1644511149
transform 1 0 47564 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1790__146
timestamp 1644511149
transform 1 0 33580 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1791__147
timestamp 1644511149
transform 1 0 15272 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1792__148
timestamp 1644511149
transform 1 0 4048 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1793__149
timestamp 1644511149
transform 1 0 2484 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1794__150
timestamp 1644511149
transform 1 0 1564 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1795__151
timestamp 1644511149
transform 1 0 47564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1796__152
timestamp 1644511149
transform 1 0 43792 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1797__153
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1798__154
timestamp 1644511149
transform 1 0 25300 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1799__155
timestamp 1644511149
transform 1 0 46184 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1800__156
timestamp 1644511149
transform 1 0 41768 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1801__157
timestamp 1644511149
transform 1 0 47564 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1802__158
timestamp 1644511149
transform 1 0 9108 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1803__159
timestamp 1644511149
transform 1 0 13156 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1804__160
timestamp 1644511149
transform 1 0 26680 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1805__161
timestamp 1644511149
transform 1 0 45540 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1806__162
timestamp 1644511149
transform 1 0 6624 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1807__163
timestamp 1644511149
transform 1 0 41124 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1808__164
timestamp 1644511149
transform 1 0 7912 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1809__165
timestamp 1644511149
transform 1 0 46828 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1810__166
timestamp 1644511149
transform 1 0 2760 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1811__167
timestamp 1644511149
transform 1 0 47472 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1812__168
timestamp 1644511149
transform 1 0 20976 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1813__169
timestamp 1644511149
transform 1 0 45632 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1814__170
timestamp 1644511149
transform 1 0 43792 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1815__171
timestamp 1644511149
transform 1 0 45724 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1816__172
timestamp 1644511149
transform 1 0 47564 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1817__173
timestamp 1644511149
transform 1 0 43516 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1818__174
timestamp 1644511149
transform 1 0 6256 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1819__175
timestamp 1644511149
transform 1 0 45632 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1820__176
timestamp 1644511149
transform 1 0 7636 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1821__177
timestamp 1644511149
transform 1 0 47932 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1822__178
timestamp 1644511149
transform 1 0 47564 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1823__179
timestamp 1644511149
transform 1 0 2116 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1824__180
timestamp 1644511149
transform 1 0 1840 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1825__181
timestamp 1644511149
transform 1 0 36248 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1826__182
timestamp 1644511149
transform 1 0 44896 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1827__183
timestamp 1644511149
transform 1 0 1840 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1828__184
timestamp 1644511149
transform 1 0 44252 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1829__185
timestamp 1644511149
transform 1 0 2852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1830__186
timestamp 1644511149
transform 1 0 45632 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1831__187
timestamp 1644511149
transform 1 0 23644 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1832__188
timestamp 1644511149
transform 1 0 2668 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1833__189
timestamp 1644511149
transform 1 0 47472 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1834__190
timestamp 1644511149
transform 1 0 3772 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1835__191
timestamp 1644511149
transform 1 0 11868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1836__192
timestamp 1644511149
transform 1 0 42964 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1837__193
timestamp 1644511149
transform 1 0 3680 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1838__194
timestamp 1644511149
transform 1 0 32752 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1839__195
timestamp 1644511149
transform 1 0 21160 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1840__196
timestamp 1644511149
transform 1 0 2668 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1841__197
timestamp 1644511149
transform 1 0 1840 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1842__198
timestamp 1644511149
transform 1 0 38732 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1843__199
timestamp 1644511149
transform 1 0 1840 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1844_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16836 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1845_
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1846_
timestamp 1644511149
transform 1 0 19412 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1847_
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1848_
timestamp 1644511149
transform 1 0 16836 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1849_
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1850_
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1851_
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1852_
timestamp 1644511149
transform 1 0 30452 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1853_
timestamp 1644511149
transform 1 0 33120 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1854_
timestamp 1644511149
transform 1 0 32292 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1855_
timestamp 1644511149
transform 1 0 45172 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1856_
timestamp 1644511149
transform 1 0 13984 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1857_
timestamp 1644511149
transform 1 0 36340 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1858_
timestamp 1644511149
transform 1 0 31924 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1859_
timestamp 1644511149
transform 1 0 46276 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1860_
timestamp 1644511149
transform 1 0 37904 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1861_
timestamp 1644511149
transform 1 0 3312 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1862_
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1863_
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1864_
timestamp 1644511149
transform 1 0 11684 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1865_
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1866_
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1867_
timestamp 1644511149
transform 1 0 16744 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1868_
timestamp 1644511149
transform 1 0 16008 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1869_
timestamp 1644511149
transform 1 0 16836 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1870_
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1871_
timestamp 1644511149
transform 1 0 27416 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1872_
timestamp 1644511149
transform 1 0 16652 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1873_
timestamp 1644511149
transform 1 0 25852 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1874_
timestamp 1644511149
transform 1 0 35972 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1875_
timestamp 1644511149
transform 1 0 1932 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1876_
timestamp 1644511149
transform 1 0 46276 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_2  _1877_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15180 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_8  _1878_
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1879_
timestamp 1644511149
transform 1 0 29532 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1880_
timestamp 1644511149
transform 1 0 28152 0 -1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1881_
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1882_
timestamp 1644511149
transform 1 0 40020 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1883_
timestamp 1644511149
transform 1 0 32108 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1884_
timestamp 1644511149
transform 1 0 10120 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1885_
timestamp 1644511149
transform 1 0 1748 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1886_
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1887_
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1888_
timestamp 1644511149
transform 1 0 30360 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1889_
timestamp 1644511149
transform 1 0 16928 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1890_
timestamp 1644511149
transform 1 0 1932 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1891_
timestamp 1644511149
transform 1 0 29716 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1892_
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1893_
timestamp 1644511149
transform 1 0 46276 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1894_
timestamp 1644511149
transform 1 0 23460 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1895_
timestamp 1644511149
transform 1 0 12328 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1896_
timestamp 1644511149
transform 1 0 29716 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1897_
timestamp 1644511149
transform 1 0 20148 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1898_
timestamp 1644511149
transform 1 0 41400 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1899_
timestamp 1644511149
transform 1 0 46276 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1900_
timestamp 1644511149
transform 1 0 3128 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1901_
timestamp 1644511149
transform 1 0 41768 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1902_
timestamp 1644511149
transform 1 0 1748 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1903_
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1904_
timestamp 1644511149
transform 1 0 17756 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1905_
timestamp 1644511149
transform 1 0 19228 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1906_
timestamp 1644511149
transform 1 0 14260 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1907_
timestamp 1644511149
transform 1 0 30268 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1908_
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1909_
timestamp 1644511149
transform 1 0 46276 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1910_
timestamp 1644511149
transform 1 0 31832 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1911_
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1912_
timestamp 1644511149
transform 1 0 22540 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1913_
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1914_
timestamp 1644511149
transform 1 0 46276 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1915_
timestamp 1644511149
transform 1 0 1380 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1916_
timestamp 1644511149
transform 1 0 46276 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1917_
timestamp 1644511149
transform 1 0 46000 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1918_
timestamp 1644511149
transform 1 0 46276 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1919_
timestamp 1644511149
transform 1 0 1748 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1920_
timestamp 1644511149
transform 1 0 38088 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1921_
timestamp 1644511149
transform 1 0 45632 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1922_
timestamp 1644511149
transform 1 0 46276 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1923_
timestamp 1644511149
transform 1 0 46276 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1924_
timestamp 1644511149
transform 1 0 46276 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1925_
timestamp 1644511149
transform 1 0 46276 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1926_
timestamp 1644511149
transform 1 0 38272 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1927_
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1928_
timestamp 1644511149
transform 1 0 34868 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1929_
timestamp 1644511149
transform 1 0 11960 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1930_
timestamp 1644511149
transform 1 0 46276 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1931_
timestamp 1644511149
transform 1 0 44436 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1932_
timestamp 1644511149
transform 1 0 39284 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1933_
timestamp 1644511149
transform 1 0 11500 0 1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1934_
timestamp 1644511149
transform 1 0 6716 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1935_
timestamp 1644511149
transform 1 0 46276 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1936_
timestamp 1644511149
transform 1 0 15640 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1937_
timestamp 1644511149
transform 1 0 18216 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1938_
timestamp 1644511149
transform 1 0 45172 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1939_
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1940_
timestamp 1644511149
transform 1 0 39192 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1941_
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1942_
timestamp 1644511149
transform 1 0 39192 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1943_
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1944_
timestamp 1644511149
transform 1 0 37168 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1945_
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1946_
timestamp 1644511149
transform 1 0 15548 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1947_
timestamp 1644511149
transform 1 0 36432 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1948_
timestamp 1644511149
transform 1 0 11776 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1949_
timestamp 1644511149
transform 1 0 4784 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1950_
timestamp 1644511149
transform 1 0 33488 0 -1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1951_
timestamp 1644511149
transform 1 0 14444 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1952_
timestamp 1644511149
transform 1 0 1380 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1953_
timestamp 1644511149
transform 1 0 1748 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1954_
timestamp 1644511149
transform 1 0 1748 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1955_
timestamp 1644511149
transform 1 0 46276 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1956_
timestamp 1644511149
transform 1 0 43792 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1957_
timestamp 1644511149
transform 1 0 1748 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1958_
timestamp 1644511149
transform 1 0 27140 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1959_
timestamp 1644511149
transform 1 0 46276 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1960_
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1961_
timestamp 1644511149
transform 1 0 46276 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1962_
timestamp 1644511149
transform 1 0 9108 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1963_
timestamp 1644511149
transform 1 0 13156 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1964_
timestamp 1644511149
transform 1 0 26956 0 1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1965_
timestamp 1644511149
transform 1 0 45172 0 1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1966_
timestamp 1644511149
transform 1 0 6624 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1967_
timestamp 1644511149
transform 1 0 42412 0 1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1968_
timestamp 1644511149
transform 1 0 4692 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1969_
timestamp 1644511149
transform 1 0 46276 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1970_
timestamp 1644511149
transform 1 0 2024 0 -1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1971_
timestamp 1644511149
transform 1 0 46276 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1972_
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1973_
timestamp 1644511149
transform 1 0 45172 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1974_
timestamp 1644511149
transform 1 0 46276 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1975_
timestamp 1644511149
transform 1 0 46276 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1976_
timestamp 1644511149
transform 1 0 46276 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1977_
timestamp 1644511149
transform 1 0 44988 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1978_
timestamp 1644511149
transform 1 0 6164 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1979_
timestamp 1644511149
transform 1 0 46276 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1980_
timestamp 1644511149
transform 1 0 7360 0 -1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1981_
timestamp 1644511149
transform 1 0 46276 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1982_
timestamp 1644511149
transform 1 0 46276 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1983_
timestamp 1644511149
transform 1 0 2024 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1984_
timestamp 1644511149
transform 1 0 1380 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1985_
timestamp 1644511149
transform 1 0 35972 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1986_
timestamp 1644511149
transform 1 0 45172 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1987_
timestamp 1644511149
transform 1 0 1748 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1988_
timestamp 1644511149
transform 1 0 44712 0 -1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1989_
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1990_
timestamp 1644511149
transform 1 0 42412 0 -1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1991_
timestamp 1644511149
transform 1 0 24380 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1992_
timestamp 1644511149
transform 1 0 1748 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1993_
timestamp 1644511149
transform 1 0 46276 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1994_
timestamp 1644511149
transform 1 0 1380 0 1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1995_
timestamp 1644511149
transform 1 0 11684 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1996_
timestamp 1644511149
transform 1 0 42596 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1997_
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1998_
timestamp 1644511149
transform 1 0 32752 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1999_
timestamp 1644511149
transform 1 0 21804 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2000_
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2001_
timestamp 1644511149
transform 1 0 1748 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2002_
timestamp 1644511149
transform 1 0 37720 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2003_
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i
timestamp 1644511149
transform 1 0 30452 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 28796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 27324 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 26036 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 32384 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 25484 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 32476 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 24472 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 23000 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 32752 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 33396 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_4_0_wb_clk_i
timestamp 1644511149
transform 1 0 22080 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_5_0_wb_clk_i
timestamp 1644511149
transform 1 0 19412 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_6_0_wb_clk_i
timestamp 1644511149
transform 1 0 33764 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_7_0_wb_clk_i
timestamp 1644511149
transform 1 0 31280 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 21896 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 23552 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 21160 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 21712 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_4_0_wb_clk_i
timestamp 1644511149
transform 1 0 31556 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_5_0_wb_clk_i
timestamp 1644511149
transform 1 0 33856 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_6_0_wb_clk_i
timestamp 1644511149
transform 1 0 32660 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_7_0_wb_clk_i
timestamp 1644511149
transform 1 0 35788 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_8_0_wb_clk_i
timestamp 1644511149
transform 1 0 20516 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_9_0_wb_clk_i
timestamp 1644511149
transform 1 0 24748 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_10_0_wb_clk_i
timestamp 1644511149
transform 1 0 19596 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_11_0_wb_clk_i
timestamp 1644511149
transform 1 0 25484 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_12_0_wb_clk_i
timestamp 1644511149
transform 1 0 32108 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_13_0_wb_clk_i
timestamp 1644511149
transform 1 0 34868 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_14_0_wb_clk_i
timestamp 1644511149
transform 1 0 30912 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_15_0_wb_clk_i
timestamp 1644511149
transform 1 0 33488 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  input1
timestamp 1644511149
transform 1 0 46276 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  input2
timestamp 1644511149
transform 1 0 1748 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1644511149
transform 1 0 14628 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1644511149
transform 1 0 22632 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1644511149
transform 1 0 1748 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input6
timestamp 1644511149
transform 1 0 47656 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input7
timestamp 1644511149
transform 1 0 47840 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1644511149
transform 1 0 21988 0 1 48960
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1644511149
transform 1 0 12972 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1644511149
transform 1 0 17848 0 1 48960
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input11
timestamp 1644511149
transform 1 0 27140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input12
timestamp 1644511149
transform 1 0 32936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1644511149
transform 1 0 1748 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input14
timestamp 1644511149
transform 1 0 8648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input15
timestamp 1644511149
transform 1 0 1748 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1644511149
transform 1 0 17020 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 1644511149
transform 1 0 47840 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1644511149
transform 1 0 47288 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp 1644511149
transform 1 0 46184 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20
timestamp 1644511149
transform 1 0 47288 0 1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1644511149
transform 1 0 24380 0 1 48960
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1644511149
transform 1 0 1748 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input23
timestamp 1644511149
transform 1 0 2300 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1644511149
transform 1 0 47840 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1644511149
transform 1 0 1748 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input26
timestamp 1644511149
transform 1 0 47840 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1644511149
transform 1 0 14812 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1644511149
transform 1 0 47840 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1644511149
transform 1 0 47840 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1644511149
transform 1 0 1748 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1644511149
transform 1 0 5428 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input32
timestamp 1644511149
transform 1 0 20056 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1644511149
transform 1 0 40664 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1644511149
transform 1 0 26036 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input36
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input37
timestamp 1644511149
transform 1 0 38088 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1644511149
transform 1 0 20056 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input40
timestamp 1644511149
transform 1 0 6532 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input41
timestamp 1644511149
transform 1 0 47840 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input42
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1644511149
transform 1 0 27876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input44
timestamp 1644511149
transform 1 0 1380 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1644511149
transform 1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input46
timestamp 1644511149
transform 1 0 42872 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input47
timestamp 1644511149
transform 1 0 43700 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input48
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1644511149
transform 1 0 25208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1644511149
transform 1 0 36156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input51
timestamp 1644511149
transform 1 0 47840 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input52
timestamp 1644511149
transform 1 0 19320 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input53
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input54
timestamp 1644511149
transform 1 0 4600 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1644511149
transform 1 0 29900 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input56
timestamp 1644511149
transform 1 0 47840 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input57
timestamp 1644511149
transform 1 0 47840 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input58
timestamp 1644511149
transform 1 0 17480 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1644511149
transform 1 0 47840 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1644511149
transform 1 0 46828 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1644511149
transform 1 0 34868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input62
timestamp 1644511149
transform 1 0 47656 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1644511149
transform 1 0 33948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 1644511149
transform 1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input65
timestamp 1644511149
transform 1 0 1380 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input66
timestamp 1644511149
transform 1 0 46092 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input67
timestamp 1644511149
transform 1 0 47656 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1644511149
transform 1 0 25392 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1644511149
transform 1 0 47840 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input70
timestamp 1644511149
transform 1 0 1380 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input71
timestamp 1644511149
transform 1 0 4140 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input72
timestamp 1644511149
transform 1 0 5060 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input73
timestamp 1644511149
transform 1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input74
timestamp 1644511149
transform 1 0 10212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input75
timestamp 1644511149
transform 1 0 47840 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input76
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input77
timestamp 1644511149
transform 1 0 41584 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input78
timestamp 1644511149
transform 1 0 46736 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input79
timestamp 1644511149
transform 1 0 11592 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input80
timestamp 1644511149
transform 1 0 7176 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1644511149
transform 1 0 47932 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input82
timestamp 1644511149
transform 1 0 47840 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input83
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input84
timestamp 1644511149
transform 1 0 47840 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input85
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1644511149
transform 1 0 38732 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input87
timestamp 1644511149
transform 1 0 47840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input88
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1644511149
transform 1 0 23368 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input90
timestamp 1644511149
transform 1 0 47840 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input91
timestamp 1644511149
transform 1 0 44068 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input92
timestamp 1644511149
transform 1 0 47840 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input93
timestamp 1644511149
transform 1 0 47840 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input94
timestamp 1644511149
transform 1 0 1380 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input95
timestamp 1644511149
transform 1 0 47840 0 -1 25024
box -38 -48 406 592
<< labels >>
rlabel metal3 s 49200 31968 50000 32088 6 active
port 0 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 25134 51200 25190 52000 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 49200 15648 50000 15768 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 21270 51200 21326 52000 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 49200 2048 50000 2168 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 io_in[18]
port 10 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 49200 18368 50000 18488 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 0 30608 800 30728 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 49200 21088 50000 21208 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 49200 32648 50000 32768 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 49200 23128 50000 23248 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 2594 51200 2650 52000 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 46386 51200 46442 52000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 9034 51200 9090 52000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 31574 51200 31630 52000 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 49200 47608 50000 47728 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 49200 20408 50000 20528 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 35438 51200 35494 52000 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 49200 2728 50000 2848 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 3882 51200 3938 52000 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 io_oeb[0]
port 39 nsew signal tristate
rlabel metal3 s 49200 24488 50000 24608 6 io_oeb[10]
port 40 nsew signal tristate
rlabel metal2 s 45098 0 45154 800 6 io_oeb[11]
port 41 nsew signal tristate
rlabel metal2 s 5814 0 5870 800 6 io_oeb[12]
port 42 nsew signal tristate
rlabel metal2 s 48318 0 48374 800 6 io_oeb[13]
port 43 nsew signal tristate
rlabel metal2 s 7746 51200 7802 52000 6 io_oeb[14]
port 44 nsew signal tristate
rlabel metal3 s 49200 43528 50000 43648 6 io_oeb[15]
port 45 nsew signal tristate
rlabel metal3 s 49200 4768 50000 4888 6 io_oeb[16]
port 46 nsew signal tristate
rlabel metal3 s 0 6808 800 6928 6 io_oeb[17]
port 47 nsew signal tristate
rlabel metal3 s 0 41488 800 41608 6 io_oeb[18]
port 48 nsew signal tristate
rlabel metal2 s 36726 0 36782 800 6 io_oeb[19]
port 49 nsew signal tristate
rlabel metal2 s 43166 51200 43222 52000 6 io_oeb[1]
port 50 nsew signal tristate
rlabel metal3 s 49200 46928 50000 47048 6 io_oeb[20]
port 51 nsew signal tristate
rlabel metal3 s 0 9528 800 9648 6 io_oeb[21]
port 52 nsew signal tristate
rlabel metal2 s 45098 51200 45154 52000 6 io_oeb[22]
port 53 nsew signal tristate
rlabel metal3 s 0 26528 800 26648 6 io_oeb[23]
port 54 nsew signal tristate
rlabel metal3 s 49200 51688 50000 51808 6 io_oeb[24]
port 55 nsew signal tristate
rlabel metal2 s 24490 51200 24546 52000 6 io_oeb[25]
port 56 nsew signal tristate
rlabel metal3 s 0 23128 800 23248 6 io_oeb[26]
port 57 nsew signal tristate
rlabel metal3 s 49200 28568 50000 28688 6 io_oeb[27]
port 58 nsew signal tristate
rlabel metal2 s 1306 51200 1362 52000 6 io_oeb[28]
port 59 nsew signal tristate
rlabel metal2 s 12254 0 12310 800 6 io_oeb[29]
port 60 nsew signal tristate
rlabel metal3 s 0 51688 800 51808 6 io_oeb[2]
port 61 nsew signal tristate
rlabel metal2 s 49606 51200 49662 52000 6 io_oeb[30]
port 62 nsew signal tristate
rlabel metal3 s 0 3408 800 3528 6 io_oeb[31]
port 63 nsew signal tristate
rlabel metal2 s 33506 0 33562 800 6 io_oeb[32]
port 64 nsew signal tristate
rlabel metal2 s 22558 51200 22614 52000 6 io_oeb[33]
port 65 nsew signal tristate
rlabel metal3 s 0 17688 800 17808 6 io_oeb[34]
port 66 nsew signal tristate
rlabel metal3 s 0 13608 800 13728 6 io_oeb[35]
port 67 nsew signal tristate
rlabel metal2 s 39946 0 40002 800 6 io_oeb[36]
port 68 nsew signal tristate
rlabel metal3 s 0 39448 800 39568 6 io_oeb[37]
port 69 nsew signal tristate
rlabel metal3 s 49200 45568 50000 45688 6 io_oeb[3]
port 70 nsew signal tristate
rlabel metal3 s 0 44888 800 45008 6 io_oeb[4]
port 71 nsew signal tristate
rlabel metal3 s 49200 36728 50000 36848 6 io_oeb[5]
port 72 nsew signal tristate
rlabel metal2 s 21270 0 21326 800 6 io_oeb[6]
port 73 nsew signal tristate
rlabel metal3 s 49200 17008 50000 17128 6 io_oeb[7]
port 74 nsew signal tristate
rlabel metal3 s 49200 49648 50000 49768 6 io_oeb[8]
port 75 nsew signal tristate
rlabel metal3 s 49200 16328 50000 16448 6 io_oeb[9]
port 76 nsew signal tristate
rlabel metal2 s 36082 51200 36138 52000 6 io_out[0]
port 77 nsew signal tristate
rlabel metal3 s 49200 44208 50000 44328 6 io_out[10]
port 78 nsew signal tristate
rlabel metal3 s 49200 9528 50000 9648 6 io_out[11]
port 79 nsew signal tristate
rlabel metal2 s 48962 0 49018 800 6 io_out[12]
port 80 nsew signal tristate
rlabel metal2 s 47030 0 47086 800 6 io_out[13]
port 81 nsew signal tristate
rlabel metal3 s 49200 12248 50000 12368 6 io_out[14]
port 82 nsew signal tristate
rlabel metal2 s 37370 0 37426 800 6 io_out[15]
port 83 nsew signal tristate
rlabel metal2 s 37370 51200 37426 52000 6 io_out[16]
port 84 nsew signal tristate
rlabel metal2 s 38658 51200 38714 52000 6 io_out[17]
port 85 nsew signal tristate
rlabel metal2 s 15474 51200 15530 52000 6 io_out[18]
port 86 nsew signal tristate
rlabel metal3 s 49200 3408 50000 3528 6 io_out[19]
port 87 nsew signal tristate
rlabel metal2 s 12898 0 12954 800 6 io_out[1]
port 88 nsew signal tristate
rlabel metal2 s 11610 0 11666 800 6 io_out[20]
port 89 nsew signal tristate
rlabel metal3 s 0 48288 800 48408 6 io_out[21]
port 90 nsew signal tristate
rlabel metal2 s 34794 51200 34850 52000 6 io_out[22]
port 91 nsew signal tristate
rlabel metal2 s 14830 51200 14886 52000 6 io_out[23]
port 92 nsew signal tristate
rlabel metal3 s 0 46248 800 46368 6 io_out[24]
port 93 nsew signal tristate
rlabel metal3 s 0 34008 800 34128 6 io_out[25]
port 94 nsew signal tristate
rlabel metal3 s 0 27208 800 27328 6 io_out[26]
port 95 nsew signal tristate
rlabel metal3 s 49200 7488 50000 7608 6 io_out[27]
port 96 nsew signal tristate
rlabel metal2 s 44454 0 44510 800 6 io_out[28]
port 97 nsew signal tristate
rlabel metal3 s 0 5448 800 5568 6 io_out[29]
port 98 nsew signal tristate
rlabel metal3 s 49200 35368 50000 35488 6 io_out[2]
port 99 nsew signal tristate
rlabel metal2 s 28354 51200 28410 52000 6 io_out[30]
port 100 nsew signal tristate
rlabel metal3 s 49200 46248 50000 46368 6 io_out[31]
port 101 nsew signal tristate
rlabel metal2 s 42522 0 42578 800 6 io_out[32]
port 102 nsew signal tristate
rlabel metal3 s 49200 10888 50000 11008 6 io_out[33]
port 103 nsew signal tristate
rlabel metal3 s 0 51008 800 51128 6 io_out[34]
port 104 nsew signal tristate
rlabel metal2 s 13542 0 13598 800 6 io_out[35]
port 105 nsew signal tristate
rlabel metal2 s 27066 51200 27122 52000 6 io_out[36]
port 106 nsew signal tristate
rlabel metal2 s 48318 51200 48374 52000 6 io_out[37]
port 107 nsew signal tristate
rlabel metal2 s 45742 51200 45798 52000 6 io_out[3]
port 108 nsew signal tristate
rlabel metal2 s 39946 51200 40002 52000 6 io_out[4]
port 109 nsew signal tristate
rlabel metal2 s 10322 51200 10378 52000 6 io_out[5]
port 110 nsew signal tristate
rlabel metal2 s 7102 51200 7158 52000 6 io_out[6]
port 111 nsew signal tristate
rlabel metal3 s 49200 34008 50000 34128 6 io_out[7]
port 112 nsew signal tristate
rlabel metal2 s 2594 0 2650 800 6 io_out[8]
port 113 nsew signal tristate
rlabel metal2 s 8390 51200 8446 52000 6 io_out[9]
port 114 nsew signal tristate
rlabel metal3 s 0 8168 800 8288 6 rambus_wb_ack_i
port 115 nsew signal input
rlabel metal3 s 49200 40128 50000 40248 6 rambus_wb_adr_o[0]
port 116 nsew signal tristate
rlabel metal3 s 0 46928 800 47048 6 rambus_wb_adr_o[1]
port 117 nsew signal tristate
rlabel metal2 s 10966 51200 11022 52000 6 rambus_wb_adr_o[2]
port 118 nsew signal tristate
rlabel metal3 s 49200 6128 50000 6248 6 rambus_wb_adr_o[3]
port 119 nsew signal tristate
rlabel metal3 s 49200 51008 50000 51128 6 rambus_wb_adr_o[4]
port 120 nsew signal tristate
rlabel metal3 s 49200 17688 50000 17808 6 rambus_wb_adr_o[5]
port 121 nsew signal tristate
rlabel metal3 s 49200 6808 50000 6928 6 rambus_wb_adr_o[6]
port 122 nsew signal tristate
rlabel metal3 s 49200 29248 50000 29368 6 rambus_wb_adr_o[7]
port 123 nsew signal tristate
rlabel metal2 s 9034 0 9090 800 6 rambus_wb_adr_o[8]
port 124 nsew signal tristate
rlabel metal3 s 0 2048 800 2168 6 rambus_wb_adr_o[9]
port 125 nsew signal tristate
rlabel metal3 s 0 18368 800 18488 6 rambus_wb_clk_o
port 126 nsew signal tristate
rlabel metal2 s 5170 51200 5226 52000 6 rambus_wb_cyc_o
port 127 nsew signal tristate
rlabel metal2 s 13542 51200 13598 52000 6 rambus_wb_dat_i[0]
port 128 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 rambus_wb_dat_i[10]
port 129 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 rambus_wb_dat_i[11]
port 130 nsew signal input
rlabel metal3 s 49200 688 50000 808 6 rambus_wb_dat_i[12]
port 131 nsew signal input
rlabel metal3 s 49200 13608 50000 13728 6 rambus_wb_dat_i[13]
port 132 nsew signal input
rlabel metal2 s 21914 51200 21970 52000 6 rambus_wb_dat_i[14]
port 133 nsew signal input
rlabel metal2 s 12898 51200 12954 52000 6 rambus_wb_dat_i[15]
port 134 nsew signal input
rlabel metal2 s 18050 51200 18106 52000 6 rambus_wb_dat_i[16]
port 135 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 rambus_wb_dat_i[17]
port 136 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 rambus_wb_dat_i[18]
port 137 nsew signal input
rlabel metal3 s 0 34688 800 34808 6 rambus_wb_dat_i[19]
port 138 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 rambus_wb_dat_i[1]
port 139 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 rambus_wb_dat_i[20]
port 140 nsew signal input
rlabel metal2 s 16118 51200 16174 52000 6 rambus_wb_dat_i[21]
port 141 nsew signal input
rlabel metal3 s 49200 8168 50000 8288 6 rambus_wb_dat_i[22]
port 142 nsew signal input
rlabel metal3 s 49200 31288 50000 31408 6 rambus_wb_dat_i[23]
port 143 nsew signal input
rlabel metal3 s 49200 33328 50000 33448 6 rambus_wb_dat_i[24]
port 144 nsew signal input
rlabel metal3 s 49200 38768 50000 38888 6 rambus_wb_dat_i[25]
port 145 nsew signal input
rlabel metal2 s 23846 51200 23902 52000 6 rambus_wb_dat_i[26]
port 146 nsew signal input
rlabel metal3 s 0 36728 800 36848 6 rambus_wb_dat_i[27]
port 147 nsew signal input
rlabel metal2 s 18 51200 74 52000 6 rambus_wb_dat_i[28]
port 148 nsew signal input
rlabel metal3 s 49200 42168 50000 42288 6 rambus_wb_dat_i[29]
port 149 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 rambus_wb_dat_i[2]
port 150 nsew signal input
rlabel metal3 s 49200 10208 50000 10328 6 rambus_wb_dat_i[30]
port 151 nsew signal input
rlabel metal2 s 14186 51200 14242 52000 6 rambus_wb_dat_i[31]
port 152 nsew signal input
rlabel metal3 s 49200 29928 50000 30048 6 rambus_wb_dat_i[3]
port 153 nsew signal input
rlabel metal3 s 49200 23808 50000 23928 6 rambus_wb_dat_i[4]
port 154 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 rambus_wb_dat_i[5]
port 155 nsew signal input
rlabel metal2 s 4526 51200 4582 52000 6 rambus_wb_dat_i[6]
port 156 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 rambus_wb_dat_i[7]
port 157 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 rambus_wb_dat_i[8]
port 158 nsew signal input
rlabel metal2 s 40590 51200 40646 52000 6 rambus_wb_dat_i[9]
port 159 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 rambus_wb_dat_o[0]
port 160 nsew signal tristate
rlabel metal2 s 30286 0 30342 800 6 rambus_wb_dat_o[10]
port 161 nsew signal tristate
rlabel metal2 s 20626 0 20682 800 6 rambus_wb_dat_o[11]
port 162 nsew signal tristate
rlabel metal2 s 41878 0 41934 800 6 rambus_wb_dat_o[12]
port 163 nsew signal tristate
rlabel metal3 s 49200 34688 50000 34808 6 rambus_wb_dat_o[13]
port 164 nsew signal tristate
rlabel metal3 s 0 50328 800 50448 6 rambus_wb_dat_o[14]
port 165 nsew signal tristate
rlabel metal2 s 42522 51200 42578 52000 6 rambus_wb_dat_o[15]
port 166 nsew signal tristate
rlabel metal2 s 1306 0 1362 800 6 rambus_wb_dat_o[16]
port 167 nsew signal tristate
rlabel metal3 s 0 29928 800 30048 6 rambus_wb_dat_o[17]
port 168 nsew signal tristate
rlabel metal2 s 18050 0 18106 800 6 rambus_wb_dat_o[18]
port 169 nsew signal tristate
rlabel metal2 s 20626 51200 20682 52000 6 rambus_wb_dat_o[19]
port 170 nsew signal tristate
rlabel metal3 s 0 10208 800 10328 6 rambus_wb_dat_o[1]
port 171 nsew signal tristate
rlabel metal2 s 15474 0 15530 800 6 rambus_wb_dat_o[20]
port 172 nsew signal tristate
rlabel metal2 s 30930 0 30986 800 6 rambus_wb_dat_o[21]
port 173 nsew signal tristate
rlabel metal3 s 0 31968 800 32088 6 rambus_wb_dat_o[22]
port 174 nsew signal tristate
rlabel metal3 s 49200 19728 50000 19848 6 rambus_wb_dat_o[23]
port 175 nsew signal tristate
rlabel metal2 s 30930 51200 30986 52000 6 rambus_wb_dat_o[24]
port 176 nsew signal tristate
rlabel metal3 s 0 16328 800 16448 6 rambus_wb_dat_o[25]
port 177 nsew signal tristate
rlabel metal2 s 23202 51200 23258 52000 6 rambus_wb_dat_o[26]
port 178 nsew signal tristate
rlabel metal3 s 0 28568 800 28688 6 rambus_wb_dat_o[27]
port 179 nsew signal tristate
rlabel metal3 s 49200 50328 50000 50448 6 rambus_wb_dat_o[28]
port 180 nsew signal tristate
rlabel metal3 s 0 48968 800 49088 6 rambus_wb_dat_o[29]
port 181 nsew signal tristate
rlabel metal2 s 31574 0 31630 800 6 rambus_wb_dat_o[2]
port 182 nsew signal tristate
rlabel metal3 s 49200 41488 50000 41608 6 rambus_wb_dat_o[30]
port 183 nsew signal tristate
rlabel metal2 s 46386 0 46442 800 6 rambus_wb_dat_o[31]
port 184 nsew signal tristate
rlabel metal2 s 17406 51200 17462 52000 6 rambus_wb_dat_o[3]
port 185 nsew signal tristate
rlabel metal3 s 0 32648 800 32768 6 rambus_wb_dat_o[4]
port 186 nsew signal tristate
rlabel metal2 s 32218 51200 32274 52000 6 rambus_wb_dat_o[5]
port 187 nsew signal tristate
rlabel metal2 s 5170 0 5226 800 6 rambus_wb_dat_o[6]
port 188 nsew signal tristate
rlabel metal3 s 49200 14288 50000 14408 6 rambus_wb_dat_o[7]
port 189 nsew signal tristate
rlabel metal2 s 23846 0 23902 800 6 rambus_wb_dat_o[8]
port 190 nsew signal tristate
rlabel metal2 s 12254 51200 12310 52000 6 rambus_wb_dat_o[9]
port 191 nsew signal tristate
rlabel metal3 s 0 8848 800 8968 6 rambus_wb_rst_o
port 192 nsew signal tristate
rlabel metal2 s 41234 0 41290 800 6 rambus_wb_sel_o[0]
port 193 nsew signal tristate
rlabel metal2 s 32862 51200 32918 52000 6 rambus_wb_sel_o[1]
port 194 nsew signal tristate
rlabel metal2 s 9678 51200 9734 52000 6 rambus_wb_sel_o[2]
port 195 nsew signal tristate
rlabel metal3 s 0 33328 800 33448 6 rambus_wb_sel_o[3]
port 196 nsew signal tristate
rlabel metal2 s 29642 51200 29698 52000 6 rambus_wb_stb_o
port 197 nsew signal tristate
rlabel metal3 s 0 4768 800 4888 6 rambus_wb_we_o
port 198 nsew signal tristate
rlabel metal4 s 4208 2128 4528 49552 6 vccd1
port 199 nsew power input
rlabel metal4 s 34928 2128 35248 49552 6 vccd1
port 199 nsew power input
rlabel metal4 s 19568 2128 19888 49552 6 vssd1
port 200 nsew ground input
rlabel metal3 s 49200 1368 50000 1488 6 wb_clk_i
port 201 nsew signal input
rlabel metal2 s 26422 51200 26478 52000 6 wb_rst_i
port 202 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 wbs_ack_o
port 203 nsew signal tristate
rlabel metal3 s 0 31288 800 31408 6 wbs_adr_i[0]
port 204 nsew signal input
rlabel metal2 s 38014 51200 38070 52000 6 wbs_adr_i[10]
port 205 nsew signal input
rlabel metal2 s 19982 51200 20038 52000 6 wbs_adr_i[11]
port 206 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 wbs_adr_i[12]
port 207 nsew signal input
rlabel metal2 s 6458 51200 6514 52000 6 wbs_adr_i[13]
port 208 nsew signal input
rlabel metal3 s 49200 27888 50000 28008 6 wbs_adr_i[14]
port 209 nsew signal input
rlabel metal3 s 0 688 800 808 6 wbs_adr_i[15]
port 210 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 wbs_adr_i[16]
port 211 nsew signal input
rlabel metal3 s 0 44208 800 44328 6 wbs_adr_i[17]
port 212 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 wbs_adr_i[18]
port 213 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 wbs_adr_i[19]
port 214 nsew signal input
rlabel metal2 s 44454 51200 44510 52000 6 wbs_adr_i[1]
port 215 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 wbs_adr_i[20]
port 216 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 wbs_adr_i[21]
port 217 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wbs_adr_i[22]
port 218 nsew signal input
rlabel metal3 s 49200 5448 50000 5568 6 wbs_adr_i[23]
port 219 nsew signal input
rlabel metal2 s 19338 51200 19394 52000 6 wbs_adr_i[24]
port 220 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_adr_i[25]
port 221 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_adr_i[26]
port 222 nsew signal input
rlabel metal2 s 28998 51200 29054 52000 6 wbs_adr_i[27]
port 223 nsew signal input
rlabel metal3 s 49200 22448 50000 22568 6 wbs_adr_i[28]
port 224 nsew signal input
rlabel metal3 s 49200 40808 50000 40928 6 wbs_adr_i[29]
port 225 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_adr_i[2]
port 226 nsew signal input
rlabel metal2 s 48962 51200 49018 52000 6 wbs_adr_i[30]
port 227 nsew signal input
rlabel metal3 s 49200 14968 50000 15088 6 wbs_adr_i[31]
port 228 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 wbs_adr_i[3]
port 229 nsew signal input
rlabel metal2 s 47674 51200 47730 52000 6 wbs_adr_i[4]
port 230 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 wbs_adr_i[5]
port 231 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 wbs_adr_i[6]
port 232 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 wbs_adr_i[7]
port 233 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 wbs_adr_i[8]
port 234 nsew signal input
rlabel metal3 s 49200 8848 50000 8968 6 wbs_adr_i[9]
port 235 nsew signal input
rlabel metal2 s 25778 51200 25834 52000 6 wbs_cyc_i
port 236 nsew signal input
rlabel metal3 s 49200 38088 50000 38208 6 wbs_dat_i[0]
port 237 nsew signal input
rlabel metal2 s 662 51200 718 52000 6 wbs_dat_i[10]
port 238 nsew signal input
rlabel metal2 s 3238 51200 3294 52000 6 wbs_dat_i[11]
port 239 nsew signal input
rlabel metal2 s 1950 51200 2006 52000 6 wbs_dat_i[12]
port 240 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wbs_dat_i[13]
port 241 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 wbs_dat_i[14]
port 242 nsew signal input
rlabel metal3 s 49200 21768 50000 21888 6 wbs_dat_i[15]
port 243 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 wbs_dat_i[16]
port 244 nsew signal input
rlabel metal2 s 41878 51200 41934 52000 6 wbs_dat_i[17]
port 245 nsew signal input
rlabel metal3 s 49200 48968 50000 49088 6 wbs_dat_i[18]
port 246 nsew signal input
rlabel metal2 s 11610 51200 11666 52000 6 wbs_dat_i[19]
port 247 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_dat_i[1]
port 248 nsew signal input
rlabel metal3 s 49200 25848 50000 25968 6 wbs_dat_i[20]
port 249 nsew signal input
rlabel metal3 s 49200 48288 50000 48408 6 wbs_dat_i[21]
port 250 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 wbs_dat_i[22]
port 251 nsew signal input
rlabel metal3 s 49200 36048 50000 36168 6 wbs_dat_i[23]
port 252 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 wbs_dat_i[24]
port 253 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 wbs_dat_i[25]
port 254 nsew signal input
rlabel metal2 s 47030 51200 47086 52000 6 wbs_dat_i[26]
port 255 nsew signal input
rlabel metal2 s 18694 51200 18750 52000 6 wbs_dat_i[27]
port 256 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_i[28]
port 257 nsew signal input
rlabel metal3 s 49200 27208 50000 27328 6 wbs_dat_i[29]
port 258 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 wbs_dat_i[2]
port 259 nsew signal input
rlabel metal3 s 49200 11568 50000 11688 6 wbs_dat_i[30]
port 260 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 wbs_dat_i[31]
port 261 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 wbs_dat_i[3]
port 262 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_dat_i[4]
port 263 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 wbs_dat_i[5]
port 264 nsew signal input
rlabel metal3 s 49200 19048 50000 19168 6 wbs_dat_i[6]
port 265 nsew signal input
rlabel metal2 s 43810 51200 43866 52000 6 wbs_dat_i[7]
port 266 nsew signal input
rlabel metal3 s 49200 42848 50000 42968 6 wbs_dat_i[8]
port 267 nsew signal input
rlabel metal3 s 49200 8 50000 128 6 wbs_dat_i[9]
port 268 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_o[0]
port 269 nsew signal tristate
rlabel metal3 s 49200 26528 50000 26648 6 wbs_dat_o[10]
port 270 nsew signal tristate
rlabel metal2 s 662 0 718 800 6 wbs_dat_o[11]
port 271 nsew signal tristate
rlabel metal3 s 49200 44888 50000 45008 6 wbs_dat_o[12]
port 272 nsew signal tristate
rlabel metal2 s 41234 51200 41290 52000 6 wbs_dat_o[13]
port 273 nsew signal tristate
rlabel metal3 s 49200 4088 50000 4208 6 wbs_dat_o[14]
port 274 nsew signal tristate
rlabel metal2 s 39302 51200 39358 52000 6 wbs_dat_o[15]
port 275 nsew signal tristate
rlabel metal3 s 0 19728 800 19848 6 wbs_dat_o[16]
port 276 nsew signal tristate
rlabel metal3 s 0 21768 800 21888 6 wbs_dat_o[17]
port 277 nsew signal tristate
rlabel metal2 s 32218 0 32274 800 6 wbs_dat_o[18]
port 278 nsew signal tristate
rlabel metal2 s 18 0 74 800 6 wbs_dat_o[19]
port 279 nsew signal tristate
rlabel metal2 s 38014 0 38070 800 6 wbs_dat_o[1]
port 280 nsew signal tristate
rlabel metal3 s 0 29248 800 29368 6 wbs_dat_o[20]
port 281 nsew signal tristate
rlabel metal3 s 0 4088 800 4208 6 wbs_dat_o[21]
port 282 nsew signal tristate
rlabel metal3 s 0 12928 800 13048 6 wbs_dat_o[22]
port 283 nsew signal tristate
rlabel metal3 s 0 21088 800 21208 6 wbs_dat_o[23]
port 284 nsew signal tristate
rlabel metal2 s 10322 0 10378 800 6 wbs_dat_o[24]
port 285 nsew signal tristate
rlabel metal2 s 3238 0 3294 800 6 wbs_dat_o[25]
port 286 nsew signal tristate
rlabel metal2 s 27710 51200 27766 52000 6 wbs_dat_o[26]
port 287 nsew signal tristate
rlabel metal2 s 16762 51200 16818 52000 6 wbs_dat_o[27]
port 288 nsew signal tristate
rlabel metal2 s 26422 0 26478 800 6 wbs_dat_o[28]
port 289 nsew signal tristate
rlabel metal2 s 36726 51200 36782 52000 6 wbs_dat_o[29]
port 290 nsew signal tristate
rlabel metal3 s 49200 12928 50000 13048 6 wbs_dat_o[2]
port 291 nsew signal tristate
rlabel metal3 s 0 36048 800 36168 6 wbs_dat_o[30]
port 292 nsew signal tristate
rlabel metal3 s 49200 39448 50000 39568 6 wbs_dat_o[31]
port 293 nsew signal tristate
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_o[3]
port 294 nsew signal tristate
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_o[4]
port 295 nsew signal tristate
rlabel metal3 s 0 6128 800 6248 6 wbs_dat_o[5]
port 296 nsew signal tristate
rlabel metal3 s 49200 37408 50000 37528 6 wbs_dat_o[6]
port 297 nsew signal tristate
rlabel metal2 s 29642 0 29698 800 6 wbs_dat_o[7]
port 298 nsew signal tristate
rlabel metal2 s 34150 51200 34206 52000 6 wbs_dat_o[8]
port 299 nsew signal tristate
rlabel metal2 s 33506 51200 33562 52000 6 wbs_dat_o[9]
port 300 nsew signal tristate
rlabel metal3 s 0 49648 800 49768 6 wbs_sel_i[0]
port 301 nsew signal input
rlabel metal2 s 5814 51200 5870 52000 6 wbs_sel_i[1]
port 302 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 wbs_sel_i[2]
port 303 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 wbs_sel_i[3]
port 304 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 wbs_stb_i
port 305 nsew signal input
rlabel metal3 s 49200 25168 50000 25288 6 wbs_we_i
port 306 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 50000 52000
<< end >>
