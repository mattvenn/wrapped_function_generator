magic
tech sky130A
magscale 1 2
timestamp 1651661543
<< viali >>
rect 3801 49249 3835 49283
rect 4261 49249 4295 49283
rect 10517 49249 10551 49283
rect 12725 49249 12759 49283
rect 14105 49249 14139 49283
rect 17877 49249 17911 49283
rect 18153 49249 18187 49283
rect 22569 49249 22603 49283
rect 24869 49249 24903 49283
rect 27629 49249 27663 49283
rect 29745 49249 29779 49283
rect 30941 49249 30975 49283
rect 40693 49249 40727 49283
rect 44465 49249 44499 49283
rect 46857 49249 46891 49283
rect 1869 49181 1903 49215
rect 2881 49181 2915 49215
rect 6837 49181 6871 49215
rect 7849 49181 7883 49215
rect 9873 49181 9907 49215
rect 11989 49181 12023 49215
rect 13001 49181 13035 49215
rect 14381 49181 14415 49215
rect 16129 49181 16163 49215
rect 16865 49181 16899 49215
rect 19349 49181 19383 49215
rect 20085 49181 20119 49215
rect 21281 49181 21315 49215
rect 22017 49181 22051 49215
rect 24409 49181 24443 49215
rect 26985 49181 27019 49215
rect 32965 49181 32999 49215
rect 35909 49181 35943 49215
rect 38117 49181 38151 49215
rect 39037 49181 39071 49215
rect 39865 49181 39899 49215
rect 42625 49181 42659 49215
rect 45201 49181 45235 49215
rect 47777 49181 47811 49215
rect 3985 49113 4019 49147
rect 12173 49113 12207 49147
rect 22201 49113 22235 49147
rect 24593 49113 24627 49147
rect 27169 49113 27203 49147
rect 29929 49113 29963 49147
rect 40049 49113 40083 49147
rect 42809 49113 42843 49147
rect 45385 49113 45419 49147
rect 1961 49045 1995 49079
rect 3157 49045 3191 49079
rect 6929 49045 6963 49079
rect 9045 49045 9079 49079
rect 19533 49045 19567 49079
rect 20269 49045 20303 49079
rect 21097 49045 21131 49079
rect 32137 49045 32171 49079
rect 38301 49045 38335 49079
rect 39221 49045 39255 49079
rect 48053 49045 48087 49079
rect 3341 48773 3375 48807
rect 25973 48773 26007 48807
rect 27445 48773 27479 48807
rect 28549 48773 28583 48807
rect 39221 48773 39255 48807
rect 40877 48773 40911 48807
rect 41521 48773 41555 48807
rect 47777 48773 47811 48807
rect 6653 48705 6687 48739
rect 8953 48705 8987 48739
rect 14013 48705 14047 48739
rect 15301 48705 15335 48739
rect 16681 48705 16715 48739
rect 21281 48705 21315 48739
rect 32137 48705 32171 48739
rect 34897 48705 34931 48739
rect 1501 48637 1535 48671
rect 1685 48637 1719 48671
rect 3801 48637 3835 48671
rect 3985 48637 4019 48671
rect 4721 48637 4755 48671
rect 6837 48637 6871 48671
rect 7849 48637 7883 48671
rect 9137 48637 9171 48671
rect 9689 48637 9723 48671
rect 11529 48637 11563 48671
rect 11713 48637 11747 48671
rect 12449 48637 12483 48671
rect 14289 48637 14323 48671
rect 15577 48637 15611 48671
rect 16865 48637 16899 48671
rect 17141 48637 17175 48671
rect 22293 48637 22327 48671
rect 22753 48637 22787 48671
rect 22937 48637 22971 48671
rect 23765 48637 23799 48671
rect 29193 48637 29227 48671
rect 29377 48637 29411 48671
rect 29653 48637 29687 48671
rect 32321 48637 32355 48671
rect 32873 48637 32907 48671
rect 35081 48637 35115 48671
rect 36093 48637 36127 48671
rect 38577 48637 38611 48671
rect 39037 48637 39071 48671
rect 42625 48637 42659 48671
rect 42809 48637 42843 48671
rect 43177 48637 43211 48671
rect 44925 48637 44959 48671
rect 45109 48637 45143 48671
rect 45753 48637 45787 48671
rect 27629 48569 27663 48603
rect 20269 48501 20303 48535
rect 25421 48501 25455 48535
rect 26065 48501 26099 48535
rect 28641 48501 28675 48535
rect 37473 48501 37507 48535
rect 41613 48501 41647 48535
rect 48053 48501 48087 48535
rect 9137 48297 9171 48331
rect 12081 48297 12115 48331
rect 30205 48297 30239 48331
rect 38761 48297 38795 48331
rect 7757 48229 7791 48263
rect 23673 48229 23707 48263
rect 28917 48229 28951 48263
rect 30849 48229 30883 48263
rect 39957 48229 39991 48263
rect 1869 48161 1903 48195
rect 5825 48161 5859 48195
rect 9689 48161 9723 48195
rect 10333 48161 10367 48195
rect 14933 48161 14967 48195
rect 16773 48161 16807 48195
rect 17417 48161 17451 48195
rect 19993 48161 20027 48195
rect 20729 48161 20763 48195
rect 25789 48161 25823 48195
rect 25973 48161 26007 48195
rect 27629 48161 27663 48195
rect 31401 48161 31435 48195
rect 32229 48161 32263 48195
rect 36369 48161 36403 48195
rect 37565 48161 37599 48195
rect 42533 48161 42567 48195
rect 48145 48161 48179 48195
rect 1409 48093 1443 48127
rect 4261 48093 4295 48127
rect 5365 48093 5399 48127
rect 7665 48093 7699 48127
rect 9045 48093 9079 48127
rect 11989 48093 12023 48127
rect 14473 48093 14507 48127
rect 22293 48093 22327 48127
rect 22569 48093 22603 48127
rect 23581 48093 23615 48127
rect 28273 48093 28307 48127
rect 28825 48093 28859 48127
rect 30113 48093 30147 48127
rect 30757 48093 30791 48127
rect 34069 48093 34103 48127
rect 35725 48093 35759 48127
rect 38669 48093 38703 48127
rect 39865 48093 39899 48127
rect 41061 48093 41095 48127
rect 43913 48093 43947 48127
rect 45017 48093 45051 48127
rect 46305 48093 46339 48127
rect 1593 48025 1627 48059
rect 4445 48025 4479 48059
rect 5549 48025 5583 48059
rect 9873 48025 9907 48059
rect 14657 48025 14691 48059
rect 16957 48025 16991 48059
rect 20177 48025 20211 48059
rect 24961 48025 24995 48059
rect 31585 48025 31619 48059
rect 35817 48025 35851 48059
rect 36553 48025 36587 48059
rect 41245 48025 41279 48059
rect 46489 48025 46523 48059
rect 25237 47957 25271 47991
rect 44097 47957 44131 47991
rect 45201 47957 45235 47991
rect 1501 47753 1535 47787
rect 3065 47753 3099 47787
rect 5457 47753 5491 47787
rect 9965 47753 9999 47787
rect 16773 47753 16807 47787
rect 17417 47753 17451 47787
rect 19717 47753 19751 47787
rect 21189 47753 21223 47787
rect 24225 47753 24259 47787
rect 32229 47753 32263 47787
rect 36185 47753 36219 47787
rect 40417 47753 40451 47787
rect 42717 47753 42751 47787
rect 43637 47753 43671 47787
rect 2145 47685 2179 47719
rect 33241 47685 33275 47719
rect 33977 47685 34011 47719
rect 46673 47685 46707 47719
rect 47777 47685 47811 47719
rect 1409 47617 1443 47651
rect 2973 47617 3007 47651
rect 3985 47617 4019 47651
rect 4629 47617 4663 47651
rect 5365 47617 5399 47651
rect 9873 47617 9907 47651
rect 11805 47617 11839 47651
rect 14657 47617 14691 47651
rect 16681 47617 16715 47651
rect 17325 47617 17359 47651
rect 19625 47617 19659 47651
rect 21097 47617 21131 47651
rect 21833 47617 21867 47651
rect 24133 47617 24167 47651
rect 25237 47617 25271 47651
rect 26985 47617 27019 47651
rect 27077 47617 27111 47651
rect 28089 47617 28123 47651
rect 30573 47617 30607 47651
rect 32137 47617 32171 47651
rect 33149 47617 33183 47651
rect 33793 47617 33827 47651
rect 36093 47617 36127 47651
rect 39773 47617 39807 47651
rect 40325 47617 40359 47651
rect 41245 47617 41279 47651
rect 41889 47617 41923 47651
rect 42625 47617 42659 47651
rect 43545 47617 43579 47651
rect 7481 47549 7515 47583
rect 7665 47549 7699 47583
rect 9229 47549 9263 47583
rect 22017 47549 22051 47583
rect 22293 47549 22327 47583
rect 25513 47549 25547 47583
rect 28273 47549 28307 47583
rect 28641 47549 28675 47583
rect 34805 47549 34839 47583
rect 44189 47549 44223 47583
rect 44373 47549 44407 47583
rect 45017 47549 45051 47583
rect 2237 47413 2271 47447
rect 4813 47413 4847 47447
rect 46949 47413 46983 47447
rect 47869 47413 47903 47447
rect 3985 47209 4019 47243
rect 5549 47209 5583 47243
rect 9045 47209 9079 47243
rect 14381 47209 14415 47243
rect 24593 47209 24627 47243
rect 26341 47209 26375 47243
rect 42993 47209 43027 47243
rect 43821 47209 43855 47243
rect 44373 47209 44407 47243
rect 45293 47209 45327 47243
rect 4629 47141 4663 47175
rect 1409 47073 1443 47107
rect 1869 47073 1903 47107
rect 5457 47005 5491 47039
rect 8953 47005 8987 47039
rect 14289 47005 14323 47039
rect 21833 47005 21867 47039
rect 25053 47005 25087 47039
rect 27353 47005 27387 47039
rect 27721 47005 27755 47039
rect 28457 47005 28491 47039
rect 28549 47005 28583 47039
rect 44281 47005 44315 47039
rect 45201 47005 45235 47039
rect 46305 47005 46339 47039
rect 48145 47005 48179 47039
rect 1593 46937 1627 46971
rect 46489 46937 46523 46971
rect 21925 46869 21959 46903
rect 2237 46665 2271 46699
rect 44649 46665 44683 46699
rect 47685 46665 47719 46699
rect 21281 46597 21315 46631
rect 24685 46597 24719 46631
rect 47041 46597 47075 46631
rect 1409 46529 1443 46563
rect 2145 46529 2179 46563
rect 2789 46529 2823 46563
rect 3617 46529 3651 46563
rect 4261 46529 4295 46563
rect 28273 46529 28307 46563
rect 44097 46529 44131 46563
rect 44557 46529 44591 46563
rect 47593 46529 47627 46563
rect 19441 46461 19475 46495
rect 19625 46461 19659 46495
rect 45201 46461 45235 46495
rect 45385 46461 45419 46495
rect 1593 46325 1627 46359
rect 2881 46325 2915 46359
rect 8125 46325 8159 46359
rect 26157 46325 26191 46359
rect 19717 46121 19751 46155
rect 44373 46121 44407 46155
rect 45201 46121 45235 46155
rect 1593 45985 1627 46019
rect 2973 45985 3007 46019
rect 25421 45985 25455 46019
rect 48145 45985 48179 46019
rect 1409 45917 1443 45951
rect 19625 45917 19659 45951
rect 25237 45917 25271 45951
rect 45661 45917 45695 45951
rect 46305 45917 46339 45951
rect 45753 45849 45787 45883
rect 46489 45849 46523 45883
rect 1869 45509 1903 45543
rect 46305 45509 46339 45543
rect 46949 45509 46983 45543
rect 2881 45441 2915 45475
rect 7941 45441 7975 45475
rect 23765 45441 23799 45475
rect 45109 45441 45143 45475
rect 45753 45441 45787 45475
rect 46213 45441 46247 45475
rect 46857 45441 46891 45475
rect 47593 45441 47627 45475
rect 8125 45373 8159 45407
rect 8401 45373 8435 45407
rect 24777 45373 24811 45407
rect 1961 45237 1995 45271
rect 47685 45237 47719 45271
rect 9045 45033 9079 45067
rect 45845 45033 45879 45067
rect 23213 44897 23247 44931
rect 46489 44897 46523 44931
rect 48145 44897 48179 44931
rect 2329 44829 2363 44863
rect 2973 44829 3007 44863
rect 8953 44829 8987 44863
rect 23029 44829 23063 44863
rect 46305 44829 46339 44863
rect 24777 44761 24811 44795
rect 3065 44693 3099 44727
rect 26065 44693 26099 44727
rect 2237 44421 2271 44455
rect 2053 44353 2087 44387
rect 23765 44353 23799 44387
rect 47777 44353 47811 44387
rect 2789 44285 2823 44319
rect 24777 44285 24811 44319
rect 47041 44149 47075 44183
rect 20269 43809 20303 43843
rect 25053 43809 25087 43843
rect 46305 43809 46339 43843
rect 1869 43741 1903 43775
rect 20085 43741 20119 43775
rect 23857 43741 23891 43775
rect 24501 43741 24535 43775
rect 2237 43673 2271 43707
rect 23489 43673 23523 43707
rect 46489 43673 46523 43707
rect 48145 43673 48179 43707
rect 27353 43401 27387 43435
rect 46949 43401 46983 43435
rect 1869 43333 1903 43367
rect 20545 43333 20579 43367
rect 20177 43265 20211 43299
rect 21925 43265 21959 43299
rect 22109 43265 22143 43299
rect 24685 43265 24719 43299
rect 24777 43265 24811 43299
rect 24869 43265 24903 43299
rect 25053 43265 25087 43299
rect 27169 43265 27203 43299
rect 27445 43265 27479 43299
rect 46857 43265 46891 43299
rect 47869 43265 47903 43299
rect 2145 43061 2179 43095
rect 22293 43061 22327 43095
rect 24409 43061 24443 43095
rect 26985 43061 27019 43095
rect 48053 43061 48087 43095
rect 19809 42653 19843 42687
rect 21373 42653 21407 42687
rect 24685 42653 24719 42687
rect 24952 42653 24986 42687
rect 26755 42653 26789 42687
rect 26893 42653 26927 42687
rect 26985 42653 27019 42687
rect 27169 42653 27203 42687
rect 28641 42653 28675 42687
rect 28825 42653 28859 42687
rect 28917 42653 28951 42687
rect 29561 42653 29595 42687
rect 20085 42585 20119 42619
rect 21640 42585 21674 42619
rect 23489 42585 23523 42619
rect 23673 42585 23707 42619
rect 23857 42585 23891 42619
rect 29806 42585 29840 42619
rect 47961 42585 47995 42619
rect 22753 42517 22787 42551
rect 26065 42517 26099 42551
rect 26525 42517 26559 42551
rect 28457 42517 28491 42551
rect 30941 42517 30975 42551
rect 48053 42517 48087 42551
rect 21833 42313 21867 42347
rect 25697 42313 25731 42347
rect 29837 42313 29871 42347
rect 30665 42313 30699 42347
rect 23489 42245 23523 42279
rect 23673 42245 23707 42279
rect 24562 42245 24596 42279
rect 27353 42245 27387 42279
rect 28702 42245 28736 42279
rect 15577 42177 15611 42211
rect 22109 42177 22143 42211
rect 22201 42177 22235 42211
rect 22293 42177 22327 42211
rect 22477 42177 22511 42211
rect 24317 42177 24351 42211
rect 27629 42177 27663 42211
rect 27721 42177 27755 42211
rect 27813 42177 27847 42211
rect 27997 42177 28031 42211
rect 30481 42177 30515 42211
rect 30757 42177 30791 42211
rect 28457 42109 28491 42143
rect 2053 41973 2087 42007
rect 15669 41973 15703 42007
rect 23857 41973 23891 42007
rect 30297 41973 30331 42007
rect 47777 41973 47811 42007
rect 24409 41769 24443 41803
rect 27353 41769 27387 41803
rect 27905 41769 27939 41803
rect 1409 41633 1443 41667
rect 1869 41633 1903 41667
rect 15761 41633 15795 41667
rect 16589 41633 16623 41667
rect 25973 41633 26007 41667
rect 29561 41633 29595 41667
rect 46305 41633 46339 41667
rect 15577 41565 15611 41599
rect 20545 41565 20579 41599
rect 22477 41565 22511 41599
rect 24685 41565 24719 41599
rect 24777 41565 24811 41599
rect 24869 41565 24903 41599
rect 25053 41565 25087 41599
rect 26240 41565 26274 41599
rect 28181 41565 28215 41599
rect 28273 41565 28307 41599
rect 28365 41565 28399 41599
rect 28549 41565 28583 41599
rect 48145 41565 48179 41599
rect 1593 41497 1627 41531
rect 20812 41497 20846 41531
rect 22744 41497 22778 41531
rect 29806 41497 29840 41531
rect 46489 41497 46523 41531
rect 21925 41429 21959 41463
rect 23857 41429 23891 41463
rect 30941 41429 30975 41463
rect 2605 41225 2639 41259
rect 22661 41225 22695 41259
rect 27721 41225 27755 41259
rect 29193 41225 29227 41259
rect 46765 41225 46799 41259
rect 22201 41157 22235 41191
rect 24133 41157 24167 41191
rect 28825 41157 28859 41191
rect 1869 41089 1903 41123
rect 2513 41089 2547 41123
rect 14749 41089 14783 41123
rect 15016 41089 15050 41123
rect 20821 41089 20855 41123
rect 20913 41089 20947 41123
rect 21005 41089 21039 41123
rect 21189 41089 21223 41123
rect 21833 41089 21867 41123
rect 22017 41089 22051 41123
rect 22891 41089 22925 41123
rect 23026 41092 23060 41126
rect 23126 41089 23160 41123
rect 23305 41089 23339 41123
rect 23765 41089 23799 41123
rect 23949 41089 23983 41123
rect 27997 41089 28031 41123
rect 28089 41089 28123 41123
rect 28181 41089 28215 41123
rect 28365 41089 28399 41123
rect 29009 41089 29043 41123
rect 29285 41089 29319 41123
rect 32577 41089 32611 41123
rect 46673 41089 46707 41123
rect 47961 41089 47995 41123
rect 32321 41021 32355 41055
rect 20545 40953 20579 40987
rect 1961 40885 1995 40919
rect 16129 40885 16163 40919
rect 33701 40885 33735 40919
rect 48053 40885 48087 40919
rect 23397 40681 23431 40715
rect 32873 40681 32907 40715
rect 29009 40613 29043 40647
rect 32321 40545 32355 40579
rect 33425 40545 33459 40579
rect 28825 40477 28859 40511
rect 31125 40477 31159 40511
rect 32137 40477 32171 40511
rect 33333 40477 33367 40511
rect 45845 40477 45879 40511
rect 46305 40477 46339 40511
rect 1869 40409 1903 40443
rect 23305 40409 23339 40443
rect 29745 40409 29779 40443
rect 29929 40409 29963 40443
rect 46489 40409 46523 40443
rect 48145 40409 48179 40443
rect 1961 40341 1995 40375
rect 30113 40341 30147 40375
rect 31125 40341 31159 40375
rect 31677 40341 31711 40375
rect 32045 40341 32079 40375
rect 33241 40341 33275 40375
rect 24777 40137 24811 40171
rect 29837 40137 29871 40171
rect 34345 40137 34379 40171
rect 46765 40137 46799 40171
rect 20361 40069 20395 40103
rect 20545 40069 20579 40103
rect 30205 40069 30239 40103
rect 31217 40069 31251 40103
rect 32321 40069 32355 40103
rect 23653 40001 23687 40035
rect 25651 40001 25685 40035
rect 25789 40001 25823 40035
rect 25881 40001 25915 40035
rect 26065 40001 26099 40035
rect 31401 40001 31435 40035
rect 32137 40001 32171 40035
rect 33232 40001 33266 40035
rect 46673 40001 46707 40035
rect 23397 39933 23431 39967
rect 30297 39933 30331 39967
rect 30389 39933 30423 39967
rect 32965 39933 32999 39967
rect 31585 39865 31619 39899
rect 2237 39797 2271 39831
rect 20729 39797 20763 39831
rect 25421 39797 25455 39831
rect 32505 39797 32539 39831
rect 47777 39797 47811 39831
rect 23213 39593 23247 39627
rect 32137 39593 32171 39627
rect 21281 39525 21315 39559
rect 24869 39457 24903 39491
rect 30297 39457 30331 39491
rect 33241 39457 33275 39491
rect 46305 39457 46339 39491
rect 48145 39457 48179 39491
rect 2881 39389 2915 39423
rect 19901 39389 19935 39423
rect 22109 39389 22143 39423
rect 23489 39389 23523 39423
rect 23581 39389 23615 39423
rect 23673 39389 23707 39423
rect 23857 39389 23891 39423
rect 25881 39389 25915 39423
rect 26137 39389 26171 39423
rect 27905 39389 27939 39423
rect 28181 39389 28215 39423
rect 32413 39389 32447 39423
rect 32502 39386 32536 39420
rect 32597 39389 32631 39423
rect 32781 39389 32815 39423
rect 33497 39389 33531 39423
rect 33609 39389 33643 39423
rect 33701 39389 33735 39423
rect 33885 39389 33919 39423
rect 34713 39389 34747 39423
rect 36553 39389 36587 39423
rect 20146 39321 20180 39355
rect 22293 39321 22327 39355
rect 24501 39321 24535 39355
rect 24685 39321 24719 39355
rect 27721 39321 27755 39355
rect 28089 39321 28123 39355
rect 30542 39321 30576 39355
rect 34958 39321 34992 39355
rect 36798 39321 36832 39355
rect 46489 39321 46523 39355
rect 2973 39253 3007 39287
rect 22477 39253 22511 39287
rect 27261 39253 27295 39287
rect 31677 39253 31711 39287
rect 36093 39253 36127 39287
rect 37933 39253 37967 39287
rect 19901 39049 19935 39083
rect 24225 39049 24259 39083
rect 26433 39049 26467 39083
rect 26985 39049 27019 39083
rect 27353 39049 27387 39083
rect 29193 39049 29227 39083
rect 29653 39049 29687 39083
rect 30389 39049 30423 39083
rect 36001 39049 36035 39083
rect 37657 39049 37691 39083
rect 46765 39049 46799 39083
rect 2237 38981 2271 39015
rect 33609 38981 33643 39015
rect 34253 38981 34287 39015
rect 37473 38981 37507 39015
rect 2053 38913 2087 38947
rect 20177 38913 20211 38947
rect 20269 38913 20303 38947
rect 20361 38913 20395 38947
rect 20545 38913 20579 38947
rect 22100 38913 22134 38947
rect 24133 38913 24167 38947
rect 25053 38913 25087 38947
rect 25320 38913 25354 38947
rect 27169 38913 27203 38947
rect 27445 38913 27479 38947
rect 29561 38913 29595 38947
rect 30665 38913 30699 38947
rect 30757 38913 30791 38947
rect 30849 38913 30883 38947
rect 31033 38913 31067 38947
rect 33425 38913 33459 38947
rect 34483 38913 34517 38947
rect 34618 38916 34652 38950
rect 34713 38913 34747 38947
rect 34897 38913 34931 38947
rect 36277 38913 36311 38947
rect 36366 38916 36400 38950
rect 36482 38916 36516 38950
rect 36645 38913 36679 38947
rect 37289 38913 37323 38947
rect 46673 38913 46707 38947
rect 48145 38913 48179 38947
rect 2789 38845 2823 38879
rect 21833 38845 21867 38879
rect 29837 38845 29871 38879
rect 33793 38777 33827 38811
rect 23213 38709 23247 38743
rect 47961 38709 47995 38743
rect 21741 38505 21775 38539
rect 24639 38505 24673 38539
rect 25697 38505 25731 38539
rect 23121 38437 23155 38471
rect 19257 38301 19291 38335
rect 22017 38301 22051 38335
rect 22109 38301 22143 38335
rect 22201 38301 22235 38335
rect 22385 38301 22419 38335
rect 24409 38301 24443 38335
rect 25973 38301 26007 38335
rect 26065 38301 26099 38335
rect 26157 38301 26191 38335
rect 26341 38301 26375 38335
rect 28641 38301 28675 38335
rect 28733 38301 28767 38335
rect 28825 38301 28859 38335
rect 29009 38301 29043 38335
rect 29561 38301 29595 38335
rect 32689 38301 32723 38335
rect 32781 38301 32815 38335
rect 32873 38301 32907 38335
rect 33057 38301 33091 38335
rect 35633 38301 35667 38335
rect 36277 38301 36311 38335
rect 47869 38301 47903 38335
rect 19502 38233 19536 38267
rect 22937 38233 22971 38267
rect 28365 38233 28399 38267
rect 29806 38233 29840 38267
rect 35449 38233 35483 38267
rect 36522 38233 36556 38267
rect 20637 38165 20671 38199
rect 30941 38165 30975 38199
rect 32413 38165 32447 38199
rect 35817 38165 35851 38199
rect 37657 38165 37691 38199
rect 48053 38165 48087 38199
rect 18613 37961 18647 37995
rect 22017 37961 22051 37995
rect 25697 37961 25731 37995
rect 27537 37961 27571 37995
rect 29193 37961 29227 37995
rect 36093 37961 36127 37995
rect 19901 37893 19935 37927
rect 23213 37893 23247 37927
rect 1869 37825 1903 37859
rect 18889 37825 18923 37859
rect 18981 37825 19015 37859
rect 19073 37825 19107 37859
rect 19257 37825 19291 37859
rect 19717 37825 19751 37859
rect 20637 37825 20671 37859
rect 21833 37825 21867 37859
rect 23029 37825 23063 37859
rect 23673 37825 23707 37859
rect 25605 37825 25639 37859
rect 27445 37825 27479 37859
rect 28825 37825 28859 37859
rect 29009 37825 29043 37859
rect 32413 37825 32447 37859
rect 32669 37825 32703 37859
rect 36349 37825 36383 37859
rect 36474 37825 36508 37859
rect 36574 37825 36608 37859
rect 36737 37825 36771 37859
rect 20085 37757 20119 37791
rect 23949 37757 23983 37791
rect 27721 37757 27755 37791
rect 2053 37689 2087 37723
rect 20821 37621 20855 37655
rect 27077 37621 27111 37655
rect 33793 37621 33827 37655
rect 32229 37417 32263 37451
rect 21557 37349 21591 37383
rect 28825 37349 28859 37383
rect 2053 37281 2087 37315
rect 30941 37281 30975 37315
rect 19533 37213 19567 37247
rect 19622 37213 19656 37247
rect 19717 37213 19751 37247
rect 19901 37213 19935 37247
rect 20729 37213 20763 37247
rect 24409 37213 24443 37247
rect 26709 37213 26743 37247
rect 28641 37213 28675 37247
rect 29561 37213 29595 37247
rect 32413 37213 32447 37247
rect 32689 37213 32723 37247
rect 33425 37213 33459 37247
rect 33517 37213 33551 37247
rect 33609 37213 33643 37247
rect 33793 37213 33827 37247
rect 36093 37213 36127 37247
rect 36185 37213 36219 37247
rect 36277 37207 36311 37241
rect 36461 37213 36495 37247
rect 1869 37145 1903 37179
rect 20545 37145 20579 37179
rect 21373 37145 21407 37179
rect 22661 37145 22695 37179
rect 22845 37145 22879 37179
rect 24593 37145 24627 37179
rect 25881 37145 25915 37179
rect 26065 37145 26099 37179
rect 26976 37145 27010 37179
rect 29745 37145 29779 37179
rect 30849 37145 30883 37179
rect 19257 37077 19291 37111
rect 23029 37077 23063 37111
rect 24777 37077 24811 37111
rect 26249 37077 26283 37111
rect 28089 37077 28123 37111
rect 29929 37077 29963 37111
rect 30389 37077 30423 37111
rect 30757 37077 30791 37111
rect 32597 37077 32631 37111
rect 33149 37077 33183 37111
rect 35817 37077 35851 37111
rect 25237 36873 25271 36907
rect 28273 36873 28307 36907
rect 28917 36873 28951 36907
rect 32873 36873 32907 36907
rect 36001 36873 36035 36907
rect 18880 36805 18914 36839
rect 20453 36805 20487 36839
rect 26985 36805 27019 36839
rect 28181 36805 28215 36839
rect 30266 36805 30300 36839
rect 34038 36805 34072 36839
rect 35817 36805 35851 36839
rect 18613 36737 18647 36771
rect 20637 36737 20671 36771
rect 22192 36737 22226 36771
rect 23857 36737 23891 36771
rect 24124 36737 24158 36771
rect 27261 36737 27295 36771
rect 27353 36737 27387 36771
rect 27445 36737 27479 36771
rect 27629 36737 27663 36771
rect 29193 36737 29227 36771
rect 29285 36737 29319 36771
rect 29382 36737 29416 36771
rect 29561 36737 29595 36771
rect 30021 36737 30055 36771
rect 32229 36737 32263 36771
rect 33057 36737 33091 36771
rect 33241 36737 33275 36771
rect 33333 36737 33367 36771
rect 35633 36737 35667 36771
rect 20821 36669 20855 36703
rect 21925 36669 21959 36703
rect 33793 36669 33827 36703
rect 19993 36601 20027 36635
rect 32413 36601 32447 36635
rect 23305 36533 23339 36567
rect 31401 36533 31435 36567
rect 35173 36533 35207 36567
rect 47777 36533 47811 36567
rect 21097 36329 21131 36363
rect 22477 36329 22511 36363
rect 24409 36329 24443 36363
rect 30849 36329 30883 36363
rect 37013 36329 37047 36363
rect 28365 36261 28399 36295
rect 31677 36261 31711 36295
rect 27261 36193 27295 36227
rect 27445 36193 27479 36227
rect 35633 36193 35667 36227
rect 46305 36193 46339 36227
rect 48145 36193 48179 36227
rect 2237 36125 2271 36159
rect 2881 36125 2915 36159
rect 19533 36125 19567 36159
rect 19625 36125 19659 36159
rect 19717 36125 19751 36159
rect 19901 36125 19935 36159
rect 20913 36125 20947 36159
rect 22753 36125 22787 36159
rect 22845 36125 22879 36159
rect 22937 36125 22971 36159
rect 23121 36125 23155 36159
rect 24685 36125 24719 36159
rect 24777 36125 24811 36159
rect 24869 36125 24903 36159
rect 25053 36125 25087 36159
rect 25973 36125 26007 36159
rect 26065 36125 26099 36159
rect 26157 36125 26191 36159
rect 26341 36125 26375 36159
rect 27169 36125 27203 36159
rect 29817 36125 29851 36159
rect 29926 36119 29960 36153
rect 30026 36125 30060 36159
rect 30205 36125 30239 36159
rect 31493 36125 31527 36159
rect 35889 36125 35923 36159
rect 21741 36057 21775 36091
rect 27997 36057 28031 36091
rect 28181 36057 28215 36091
rect 30757 36057 30791 36091
rect 46489 36057 46523 36091
rect 2973 35989 3007 36023
rect 19257 35989 19291 36023
rect 21833 35989 21867 36023
rect 25697 35989 25731 36023
rect 26801 35989 26835 36023
rect 29561 35989 29595 36023
rect 19993 35785 20027 35819
rect 20821 35785 20855 35819
rect 28365 35785 28399 35819
rect 29837 35785 29871 35819
rect 30205 35785 30239 35819
rect 2237 35717 2271 35751
rect 18880 35717 18914 35751
rect 20637 35717 20671 35751
rect 24685 35717 24719 35751
rect 26249 35717 26283 35751
rect 27230 35717 27264 35751
rect 29009 35717 29043 35751
rect 29377 35717 29411 35751
rect 31125 35717 31159 35751
rect 31309 35717 31343 35751
rect 2053 35649 2087 35683
rect 20453 35649 20487 35683
rect 21833 35649 21867 35683
rect 22569 35649 22603 35683
rect 24501 35649 24535 35683
rect 26985 35649 27019 35683
rect 29193 35649 29227 35683
rect 32367 35649 32401 35683
rect 32505 35649 32539 35683
rect 32618 35649 32652 35683
rect 32781 35649 32815 35683
rect 47869 35649 47903 35683
rect 2789 35581 2823 35615
rect 18613 35581 18647 35615
rect 26433 35581 26467 35615
rect 30297 35581 30331 35615
rect 30481 35581 30515 35615
rect 22753 35513 22787 35547
rect 22017 35445 22051 35479
rect 32137 35445 32171 35479
rect 46397 35445 46431 35479
rect 47041 35445 47075 35479
rect 48053 35445 48087 35479
rect 28457 35241 28491 35275
rect 31953 35241 31987 35275
rect 1685 35105 1719 35139
rect 21465 35105 21499 35139
rect 26893 35105 26927 35139
rect 32413 35105 32447 35139
rect 46305 35105 46339 35139
rect 48145 35105 48179 35139
rect 1409 35037 1443 35071
rect 17969 35037 18003 35071
rect 19257 35037 19291 35071
rect 21741 35037 21775 35071
rect 23489 35037 23523 35071
rect 26617 35037 26651 35071
rect 28273 35037 28307 35071
rect 29561 35037 29595 35071
rect 32669 35037 32703 35071
rect 45661 35037 45695 35071
rect 17785 34969 17819 35003
rect 19524 34969 19558 35003
rect 23305 34969 23339 35003
rect 24869 34969 24903 35003
rect 25053 34969 25087 35003
rect 29828 34969 29862 35003
rect 31585 34969 31619 35003
rect 31769 34969 31803 35003
rect 45753 34969 45787 35003
rect 46489 34969 46523 35003
rect 20637 34901 20671 34935
rect 30941 34901 30975 34935
rect 33793 34901 33827 34935
rect 18705 34697 18739 34731
rect 32781 34697 32815 34731
rect 47685 34697 47719 34731
rect 15853 34629 15887 34663
rect 19993 34629 20027 34663
rect 21097 34629 21131 34663
rect 26433 34629 26467 34663
rect 28733 34629 28767 34663
rect 33149 34629 33183 34663
rect 2053 34561 2087 34595
rect 14197 34561 14231 34595
rect 16957 34561 16991 34595
rect 17601 34561 17635 34595
rect 17785 34561 17819 34595
rect 18981 34561 19015 34595
rect 19073 34561 19107 34595
rect 19165 34561 19199 34595
rect 19349 34561 19383 34595
rect 19809 34561 19843 34595
rect 20913 34561 20947 34595
rect 22100 34561 22134 34595
rect 23949 34561 23983 34595
rect 24216 34561 24250 34595
rect 26249 34561 26283 34595
rect 28549 34561 28583 34595
rect 30573 34561 30607 34595
rect 46121 34561 46155 34595
rect 46765 34561 46799 34595
rect 47593 34561 47627 34595
rect 2697 34493 2731 34527
rect 14473 34493 14507 34527
rect 16773 34493 16807 34527
rect 20177 34493 20211 34527
rect 21833 34493 21867 34527
rect 26985 34493 27019 34527
rect 27261 34493 27295 34527
rect 29193 34493 29227 34527
rect 29469 34493 29503 34527
rect 33241 34493 33275 34527
rect 33425 34493 33459 34527
rect 46857 34493 46891 34527
rect 17693 34425 17727 34459
rect 23213 34425 23247 34459
rect 1593 34357 1627 34391
rect 2145 34357 2179 34391
rect 17141 34357 17175 34391
rect 21281 34357 21315 34391
rect 25329 34357 25363 34391
rect 30665 34357 30699 34391
rect 46213 34357 46247 34391
rect 17693 34153 17727 34187
rect 21465 34153 21499 34187
rect 22753 34153 22787 34187
rect 24409 34153 24443 34187
rect 19993 34085 20027 34119
rect 1409 34017 1443 34051
rect 1593 34017 1627 34051
rect 2789 34017 2823 34051
rect 11713 34017 11747 34051
rect 13093 34017 13127 34051
rect 15577 34017 15611 34051
rect 23857 34017 23891 34051
rect 28365 34017 28399 34051
rect 32689 34017 32723 34051
rect 32781 34017 32815 34051
rect 33977 34017 34011 34051
rect 46305 34017 46339 34051
rect 46489 34017 46523 34051
rect 48145 34017 48179 34051
rect 17417 33949 17451 33983
rect 18613 33949 18647 33983
rect 21741 33949 21775 33983
rect 21833 33949 21867 33983
rect 21925 33949 21959 33983
rect 22109 33949 22143 33983
rect 22569 33949 22603 33983
rect 23489 33949 23523 33983
rect 24685 33949 24719 33983
rect 24777 33949 24811 33983
rect 24869 33949 24903 33983
rect 25053 33949 25087 33983
rect 27169 33949 27203 33983
rect 27258 33949 27292 33983
rect 27353 33949 27387 33983
rect 27537 33949 27571 33983
rect 28181 33949 28215 33983
rect 31401 33949 31435 33983
rect 31493 33949 31527 33983
rect 31585 33949 31619 33983
rect 31769 33949 31803 33983
rect 32597 33949 32631 33983
rect 11897 33881 11931 33915
rect 15844 33881 15878 33915
rect 18429 33881 18463 33915
rect 19809 33881 19843 33915
rect 23673 33881 23707 33915
rect 27997 33881 28031 33915
rect 29653 33881 29687 33915
rect 29837 33881 29871 33915
rect 31125 33881 31159 33915
rect 33885 33881 33919 33915
rect 16957 33813 16991 33847
rect 17877 33813 17911 33847
rect 26893 33813 26927 33847
rect 30021 33813 30055 33847
rect 32229 33813 32263 33847
rect 33425 33813 33459 33847
rect 33793 33813 33827 33847
rect 11897 33609 11931 33643
rect 14749 33609 14783 33643
rect 15301 33609 15335 33643
rect 15485 33609 15519 33643
rect 27445 33609 27479 33643
rect 27905 33609 27939 33643
rect 29929 33609 29963 33643
rect 30389 33609 30423 33643
rect 32505 33609 32539 33643
rect 36277 33609 36311 33643
rect 16865 33541 16899 33575
rect 23305 33541 23339 33575
rect 24041 33541 24075 33575
rect 26249 33541 26283 33575
rect 28917 33541 28951 33575
rect 32137 33541 32171 33575
rect 1777 33473 1811 33507
rect 11805 33473 11839 33507
rect 14657 33473 14691 33507
rect 14841 33473 14875 33507
rect 15482 33473 15516 33507
rect 15853 33473 15887 33507
rect 16681 33473 16715 33507
rect 16957 33473 16991 33507
rect 19349 33473 19383 33507
rect 23123 33473 23157 33507
rect 24225 33473 24259 33507
rect 27813 33473 27847 33507
rect 28733 33473 28767 33507
rect 30297 33473 30331 33507
rect 32321 33473 32355 33507
rect 33057 33473 33091 33507
rect 33324 33473 33358 33507
rect 34897 33473 34931 33507
rect 35153 33473 35187 33507
rect 46489 33473 46523 33507
rect 1961 33405 1995 33439
rect 2789 33405 2823 33439
rect 15945 33405 15979 33439
rect 17509 33405 17543 33439
rect 17785 33405 17819 33439
rect 19073 33405 19107 33439
rect 28089 33405 28123 33439
rect 30481 33405 30515 33439
rect 46213 33405 46247 33439
rect 16681 33337 16715 33371
rect 26433 33337 26467 33371
rect 34437 33337 34471 33371
rect 24409 33269 24443 33303
rect 47777 33269 47811 33303
rect 2237 33065 2271 33099
rect 23765 33065 23799 33099
rect 31401 33065 31435 33099
rect 31953 33065 31987 33099
rect 15945 32997 15979 33031
rect 18061 32997 18095 33031
rect 19257 32929 19291 32963
rect 33425 32929 33459 32963
rect 46305 32929 46339 32963
rect 48053 32929 48087 32963
rect 2145 32861 2179 32895
rect 2973 32861 3007 32895
rect 15761 32861 15795 32895
rect 18337 32861 18371 32895
rect 18426 32855 18460 32889
rect 18526 32861 18560 32895
rect 18705 32861 18739 32895
rect 24409 32861 24443 32895
rect 27077 32861 27111 32895
rect 27333 32861 27367 32895
rect 30021 32861 30055 32895
rect 32229 32861 32263 32895
rect 32321 32861 32355 32895
rect 32413 32861 32447 32895
rect 32597 32861 32631 32895
rect 33057 32861 33091 32895
rect 19502 32793 19536 32827
rect 23673 32793 23707 32827
rect 24654 32793 24688 32827
rect 30266 32793 30300 32827
rect 33241 32793 33275 32827
rect 46489 32793 46523 32827
rect 20637 32725 20671 32759
rect 25789 32725 25823 32759
rect 28457 32725 28491 32759
rect 15669 32521 15703 32555
rect 16773 32521 16807 32555
rect 20269 32521 20303 32555
rect 23857 32521 23891 32555
rect 28825 32521 28859 32555
rect 29377 32521 29411 32555
rect 20085 32453 20119 32487
rect 20821 32453 20855 32487
rect 30573 32453 30607 32487
rect 2053 32385 2087 32419
rect 13369 32385 13403 32419
rect 13636 32385 13670 32419
rect 15393 32385 15427 32419
rect 16681 32385 16715 32419
rect 16865 32385 16899 32419
rect 19027 32385 19061 32419
rect 19165 32385 19199 32419
rect 19257 32385 19291 32419
rect 19441 32385 19475 32419
rect 19901 32385 19935 32419
rect 22293 32385 22327 32419
rect 23029 32385 23063 32419
rect 23213 32385 23247 32419
rect 24113 32385 24147 32419
rect 24206 32388 24240 32422
rect 24317 32385 24351 32419
rect 24501 32385 24535 32419
rect 26249 32385 26283 32419
rect 27353 32385 27387 32419
rect 27442 32385 27476 32419
rect 27558 32385 27592 32419
rect 27721 32385 27755 32419
rect 28733 32385 28767 32419
rect 29607 32385 29641 32419
rect 29758 32391 29792 32425
rect 29858 32388 29892 32422
rect 30021 32385 30055 32419
rect 47685 32385 47719 32419
rect 2237 32317 2271 32351
rect 3065 32317 3099 32351
rect 15669 32317 15703 32351
rect 22477 32317 22511 32351
rect 47869 32317 47903 32351
rect 14749 32181 14783 32215
rect 15485 32181 15519 32215
rect 18797 32181 18831 32215
rect 20913 32181 20947 32215
rect 23397 32181 23431 32215
rect 26341 32181 26375 32215
rect 27077 32181 27111 32215
rect 30665 32181 30699 32215
rect 1593 31977 1627 32011
rect 2973 31977 3007 32011
rect 14105 31977 14139 32011
rect 17417 31977 17451 32011
rect 18705 31977 18739 32011
rect 20637 31977 20671 32011
rect 22109 31977 22143 32011
rect 25789 31977 25823 32011
rect 27629 31909 27663 31943
rect 31033 31909 31067 31943
rect 31769 31909 31803 31943
rect 19257 31841 19291 31875
rect 23213 31841 23247 31875
rect 24409 31841 24443 31875
rect 28089 31841 28123 31875
rect 28273 31841 28307 31875
rect 47593 31841 47627 31875
rect 1409 31773 1443 31807
rect 2329 31773 2363 31807
rect 2881 31773 2915 31807
rect 14289 31773 14323 31807
rect 14473 31773 14507 31807
rect 14565 31773 14599 31807
rect 15393 31773 15427 31807
rect 17233 31773 17267 31807
rect 18521 31773 18555 31807
rect 19513 31773 19547 31807
rect 21465 31773 21499 31807
rect 22365 31773 22399 31807
rect 22458 31770 22492 31804
rect 22569 31767 22603 31801
rect 22753 31773 22787 31807
rect 23489 31773 23523 31807
rect 23581 31773 23615 31807
rect 23673 31773 23707 31807
rect 23857 31773 23891 31807
rect 24665 31773 24699 31807
rect 29791 31773 29825 31807
rect 29929 31773 29963 31807
rect 30026 31773 30060 31807
rect 30205 31773 30239 31807
rect 31585 31773 31619 31807
rect 32597 31773 32631 31807
rect 32689 31773 32723 31807
rect 32781 31773 32815 31807
rect 32965 31773 32999 31807
rect 47317 31773 47351 31807
rect 12265 31705 12299 31739
rect 12438 31705 12472 31739
rect 15660 31705 15694 31739
rect 18337 31705 18371 31739
rect 26801 31705 26835 31739
rect 26985 31705 27019 31739
rect 30665 31705 30699 31739
rect 30849 31705 30883 31739
rect 12633 31637 12667 31671
rect 16773 31637 16807 31671
rect 21557 31637 21591 31671
rect 27169 31637 27203 31671
rect 27997 31637 28031 31671
rect 29561 31637 29595 31671
rect 32321 31637 32355 31671
rect 13185 31433 13219 31467
rect 16037 31433 16071 31467
rect 17049 31433 17083 31467
rect 18705 31433 18739 31467
rect 20637 31433 20671 31467
rect 23213 31433 23247 31467
rect 29009 31433 29043 31467
rect 30297 31433 30331 31467
rect 30757 31433 30791 31467
rect 32597 31433 32631 31467
rect 14933 31365 14967 31399
rect 15853 31365 15887 31399
rect 23940 31365 23974 31399
rect 33324 31365 33358 31399
rect 1961 31297 1995 31331
rect 9772 31297 9806 31331
rect 11805 31297 11839 31331
rect 12061 31297 12095 31331
rect 15117 31297 15151 31331
rect 16129 31297 16163 31331
rect 16681 31297 16715 31331
rect 18889 31297 18923 31331
rect 19349 31297 19383 31331
rect 20913 31297 20947 31331
rect 21005 31297 21039 31331
rect 21097 31297 21131 31331
rect 21281 31297 21315 31331
rect 22089 31297 22123 31331
rect 26019 31297 26053 31331
rect 26157 31297 26191 31331
rect 26249 31297 26283 31331
rect 26433 31297 26467 31331
rect 28917 31297 28951 31331
rect 30665 31297 30699 31331
rect 32229 31297 32263 31331
rect 32413 31297 32447 31331
rect 33057 31297 33091 31331
rect 2145 31229 2179 31263
rect 3065 31229 3099 31263
rect 9505 31229 9539 31263
rect 15393 31229 15427 31263
rect 16773 31229 16807 31263
rect 19625 31229 19659 31263
rect 21833 31229 21867 31263
rect 23673 31229 23707 31263
rect 27261 31229 27295 31263
rect 27537 31229 27571 31263
rect 29101 31229 29135 31263
rect 30849 31229 30883 31263
rect 15853 31161 15887 31195
rect 25053 31161 25087 31195
rect 10885 31093 10919 31127
rect 15301 31093 15335 31127
rect 16681 31093 16715 31127
rect 25789 31093 25823 31127
rect 28549 31093 28583 31127
rect 34437 31093 34471 31127
rect 2881 30889 2915 30923
rect 10425 30889 10459 30923
rect 11805 30889 11839 30923
rect 16405 30889 16439 30923
rect 21741 30889 21775 30923
rect 22569 30889 22603 30923
rect 28549 30889 28583 30923
rect 32873 30889 32907 30923
rect 9965 30753 9999 30787
rect 20729 30753 20763 30787
rect 23029 30753 23063 30787
rect 33425 30753 33459 30787
rect 2053 30685 2087 30719
rect 2789 30685 2823 30719
rect 10655 30685 10689 30719
rect 10793 30685 10827 30719
rect 10885 30685 10919 30719
rect 11069 30685 11103 30719
rect 12081 30685 12115 30719
rect 12173 30685 12207 30719
rect 12265 30685 12299 30719
rect 12449 30685 12483 30719
rect 13277 30685 13311 30719
rect 14105 30685 14139 30719
rect 16681 30685 16715 30719
rect 19533 30685 19567 30719
rect 19625 30685 19659 30719
rect 19717 30685 19751 30719
rect 19901 30685 19935 30719
rect 20361 30685 20395 30719
rect 21373 30685 21407 30719
rect 22201 30685 22235 30719
rect 23305 30685 23339 30719
rect 26341 30685 26375 30719
rect 28181 30685 28215 30719
rect 28365 30685 28399 30719
rect 29745 30685 29779 30719
rect 30001 30685 30035 30719
rect 32229 30685 32263 30719
rect 33333 30685 33367 30719
rect 9597 30617 9631 30651
rect 9781 30617 9815 30651
rect 13369 30617 13403 30651
rect 14289 30617 14323 30651
rect 15945 30617 15979 30651
rect 16405 30617 16439 30651
rect 20545 30617 20579 30651
rect 21557 30617 21591 30651
rect 22385 30617 22419 30651
rect 26586 30617 26620 30651
rect 32045 30617 32079 30651
rect 32413 30617 32447 30651
rect 16589 30549 16623 30583
rect 19257 30549 19291 30583
rect 27721 30549 27755 30583
rect 31125 30549 31159 30583
rect 33241 30549 33275 30583
rect 29561 30345 29595 30379
rect 10425 30277 10459 30311
rect 17877 30277 17911 30311
rect 18429 30277 18463 30311
rect 19340 30277 19374 30311
rect 23397 30277 23431 30311
rect 29469 30277 29503 30311
rect 32505 30277 32539 30311
rect 33854 30277 33888 30311
rect 1777 30209 1811 30243
rect 4813 30209 4847 30243
rect 8760 30209 8794 30243
rect 10609 30209 10643 30243
rect 17695 30209 17729 30243
rect 21005 30209 21039 30243
rect 21833 30209 21867 30243
rect 23213 30209 23247 30243
rect 27793 30209 27827 30243
rect 32781 30209 32815 30243
rect 32873 30209 32907 30243
rect 32965 30209 32999 30243
rect 33149 30209 33183 30243
rect 47961 30209 47995 30243
rect 1961 30141 1995 30175
rect 2789 30141 2823 30175
rect 8493 30141 8527 30175
rect 19073 30141 19107 30175
rect 22109 30141 22143 30175
rect 27537 30141 27571 30175
rect 33609 30141 33643 30175
rect 4629 30073 4663 30107
rect 18613 30073 18647 30107
rect 20453 30073 20487 30107
rect 9873 30005 9907 30039
rect 10793 30005 10827 30039
rect 21189 30005 21223 30039
rect 28917 30005 28951 30039
rect 34989 30005 35023 30039
rect 48053 30005 48087 30039
rect 2145 29801 2179 29835
rect 10241 29801 10275 29835
rect 12265 29801 12299 29835
rect 33425 29801 33459 29835
rect 12449 29665 12483 29699
rect 16313 29665 16347 29699
rect 23029 29665 23063 29699
rect 27537 29665 27571 29699
rect 33885 29665 33919 29699
rect 33977 29665 34011 29699
rect 38025 29665 38059 29699
rect 1593 29597 1627 29631
rect 2053 29597 2087 29631
rect 2697 29597 2731 29631
rect 9137 29597 9171 29631
rect 10517 29597 10551 29631
rect 10609 29597 10643 29631
rect 10701 29597 10735 29631
rect 10885 29597 10919 29631
rect 12541 29597 12575 29631
rect 14381 29597 14415 29631
rect 14657 29597 14691 29631
rect 15853 29597 15887 29631
rect 16589 29597 16623 29631
rect 20085 29597 20119 29631
rect 20729 29597 20763 29631
rect 20913 29597 20947 29631
rect 23305 29597 23339 29631
rect 24685 29597 24719 29631
rect 24777 29597 24811 29631
rect 24869 29597 24903 29631
rect 25053 29597 25087 29631
rect 25605 29597 25639 29631
rect 27813 29597 27847 29631
rect 31401 29597 31435 29631
rect 32781 29597 32815 29631
rect 36185 29597 36219 29631
rect 12265 29529 12299 29563
rect 17969 29529 18003 29563
rect 18153 29529 18187 29563
rect 31217 29529 31251 29563
rect 32597 29529 32631 29563
rect 36369 29529 36403 29563
rect 2789 29461 2823 29495
rect 8953 29461 8987 29495
rect 12725 29461 12759 29495
rect 14197 29461 14231 29495
rect 14565 29461 14599 29495
rect 15669 29461 15703 29495
rect 18337 29461 18371 29495
rect 20177 29461 20211 29495
rect 21097 29461 21131 29495
rect 24409 29461 24443 29495
rect 25697 29461 25731 29495
rect 31585 29461 31619 29495
rect 32965 29461 32999 29495
rect 33793 29461 33827 29495
rect 9229 29257 9263 29291
rect 13737 29257 13771 29291
rect 18061 29257 18095 29291
rect 19901 29257 19935 29291
rect 24041 29257 24075 29291
rect 25881 29257 25915 29291
rect 36461 29257 36495 29291
rect 1961 29189 1995 29223
rect 8116 29189 8150 29223
rect 9689 29189 9723 29223
rect 9889 29189 9923 29223
rect 15485 29189 15519 29223
rect 24746 29189 24780 29223
rect 27537 29189 27571 29223
rect 32505 29189 32539 29223
rect 1777 29121 1811 29155
rect 11529 29121 11563 29155
rect 11785 29121 11819 29155
rect 13461 29121 13495 29155
rect 13645 29121 13679 29155
rect 14381 29121 14415 29155
rect 15761 29121 15795 29155
rect 15853 29121 15887 29155
rect 15945 29121 15979 29155
rect 16129 29121 16163 29155
rect 16681 29121 16715 29155
rect 16948 29121 16982 29155
rect 18521 29121 18555 29155
rect 18777 29121 18811 29155
rect 20591 29121 20625 29155
rect 20729 29121 20763 29155
rect 20821 29121 20855 29155
rect 21005 29121 21039 29155
rect 22063 29121 22097 29155
rect 22198 29124 22232 29158
rect 22298 29121 22332 29155
rect 22477 29121 22511 29155
rect 23673 29121 23707 29155
rect 23857 29121 23891 29155
rect 27353 29121 27387 29155
rect 27997 29121 28031 29155
rect 28179 29121 28213 29155
rect 31033 29121 31067 29155
rect 31125 29121 31159 29155
rect 31217 29121 31251 29155
rect 31401 29121 31435 29155
rect 32735 29121 32769 29155
rect 32873 29121 32907 29155
rect 32965 29124 32999 29158
rect 33143 29121 33177 29155
rect 33701 29121 33735 29155
rect 33957 29121 33991 29155
rect 36369 29121 36403 29155
rect 47593 29121 47627 29155
rect 3341 29053 3375 29087
rect 7849 29053 7883 29087
rect 24501 29053 24535 29087
rect 29469 29053 29503 29087
rect 29745 29053 29779 29087
rect 10057 28985 10091 29019
rect 21833 28985 21867 29019
rect 28365 28985 28399 29019
rect 35081 28985 35115 29019
rect 4261 28917 4295 28951
rect 9873 28917 9907 28951
rect 12909 28917 12943 28951
rect 14473 28917 14507 28951
rect 20361 28917 20395 28951
rect 30757 28917 30791 28951
rect 47685 28917 47719 28951
rect 8217 28713 8251 28747
rect 8401 28713 8435 28747
rect 11345 28713 11379 28747
rect 15669 28713 15703 28747
rect 17417 28713 17451 28747
rect 21373 28713 21407 28747
rect 28273 28713 28307 28747
rect 31493 28713 31527 28747
rect 33425 28713 33459 28747
rect 7849 28645 7883 28679
rect 1409 28577 1443 28611
rect 2789 28577 2823 28611
rect 9597 28577 9631 28611
rect 9781 28577 9815 28611
rect 12173 28577 12207 28611
rect 13277 28577 13311 28611
rect 13553 28577 13587 28611
rect 16129 28577 16163 28611
rect 21833 28577 21867 28611
rect 24685 28577 24719 28611
rect 28733 28577 28767 28611
rect 28917 28577 28951 28611
rect 30481 28577 30515 28611
rect 31953 28577 31987 28611
rect 32137 28577 32171 28611
rect 32965 28577 32999 28611
rect 33977 28577 34011 28611
rect 46489 28577 46523 28611
rect 48145 28577 48179 28611
rect 9689 28509 9723 28543
rect 9873 28509 9907 28543
rect 11529 28509 11563 28543
rect 12265 28509 12299 28543
rect 12357 28509 12391 28543
rect 12449 28509 12483 28543
rect 13185 28509 13219 28543
rect 14289 28509 14323 28543
rect 16405 28509 16439 28543
rect 17673 28509 17707 28543
rect 17782 28509 17816 28543
rect 17882 28509 17916 28543
rect 18061 28509 18095 28543
rect 19993 28509 20027 28543
rect 22100 28509 22134 28543
rect 27353 28509 27387 28543
rect 30297 28509 30331 28543
rect 31861 28509 31895 28543
rect 33885 28509 33919 28543
rect 46305 28509 46339 28543
rect 1593 28441 1627 28475
rect 8217 28441 8251 28475
rect 14556 28441 14590 28475
rect 20260 28441 20294 28475
rect 24930 28441 24964 28475
rect 32781 28441 32815 28475
rect 9413 28373 9447 28407
rect 11989 28373 12023 28407
rect 23213 28373 23247 28407
rect 26065 28373 26099 28407
rect 27445 28373 27479 28407
rect 28641 28373 28675 28407
rect 29837 28373 29871 28407
rect 30205 28373 30239 28407
rect 33793 28373 33827 28407
rect 2329 28169 2363 28203
rect 12173 28169 12207 28203
rect 13001 28169 13035 28203
rect 13093 28169 13127 28203
rect 14657 28169 14691 28203
rect 17049 28169 17083 28203
rect 23305 28169 23339 28203
rect 24501 28169 24535 28203
rect 33885 28169 33919 28203
rect 8401 28101 8435 28135
rect 11989 28101 12023 28135
rect 16681 28101 16715 28135
rect 16865 28101 16899 28135
rect 2237 28033 2271 28067
rect 7941 28033 7975 28067
rect 8585 28033 8619 28067
rect 9505 28033 9539 28067
rect 10517 28033 10551 28067
rect 10701 28033 10735 28067
rect 12909 28033 12943 28067
rect 13829 28033 13863 28067
rect 14013 28033 14047 28067
rect 14197 28033 14231 28067
rect 14841 28033 14875 28067
rect 22063 28033 22097 28067
rect 22201 28033 22235 28067
rect 22293 28033 22327 28067
rect 22477 28033 22511 28067
rect 22937 28033 22971 28067
rect 23121 28033 23155 28067
rect 24731 28033 24765 28067
rect 24869 28033 24903 28067
rect 24961 28033 24995 28067
rect 25145 28033 25179 28067
rect 27977 28033 28011 28067
rect 30205 28033 30239 28067
rect 30472 28033 30506 28067
rect 32761 28033 32795 28067
rect 47961 28033 47995 28067
rect 9229 27965 9263 27999
rect 11621 27965 11655 27999
rect 13277 27965 13311 27999
rect 27721 27965 27755 27999
rect 32505 27965 32539 27999
rect 12725 27897 12759 27931
rect 7757 27829 7791 27863
rect 8769 27829 8803 27863
rect 10609 27829 10643 27863
rect 11989 27829 12023 27863
rect 21833 27829 21867 27863
rect 29101 27829 29135 27863
rect 31585 27829 31619 27863
rect 48053 27829 48087 27863
rect 9873 27625 9907 27659
rect 12725 27625 12759 27659
rect 24961 27625 24995 27659
rect 12909 27557 12943 27591
rect 27261 27557 27295 27591
rect 30205 27557 30239 27591
rect 30941 27557 30975 27591
rect 47685 27557 47719 27591
rect 12541 27489 12575 27523
rect 22017 27489 22051 27523
rect 1593 27421 1627 27455
rect 2053 27421 2087 27455
rect 2881 27421 2915 27455
rect 7021 27421 7055 27455
rect 9597 27421 9631 27455
rect 9689 27421 9723 27455
rect 10333 27421 10367 27455
rect 12725 27421 12759 27455
rect 17969 27421 18003 27455
rect 20269 27421 20303 27455
rect 27537 27421 27571 27455
rect 27626 27421 27660 27455
rect 27742 27421 27776 27455
rect 27905 27421 27939 27455
rect 29837 27421 29871 27455
rect 31171 27421 31205 27455
rect 31309 27421 31343 27455
rect 31401 27421 31435 27455
rect 31585 27421 31619 27455
rect 32137 27421 32171 27455
rect 7288 27353 7322 27387
rect 10517 27353 10551 27387
rect 12449 27353 12483 27387
rect 18153 27353 18187 27387
rect 20821 27353 20855 27387
rect 22262 27353 22296 27387
rect 24593 27353 24627 27387
rect 24777 27353 24811 27387
rect 30021 27353 30055 27387
rect 2145 27285 2179 27319
rect 8401 27285 8435 27319
rect 10701 27285 10735 27319
rect 18337 27285 18371 27319
rect 23397 27285 23431 27319
rect 32229 27285 32263 27319
rect 8519 27081 8553 27115
rect 12081 27081 12115 27115
rect 23397 27081 23431 27115
rect 1961 27013 1995 27047
rect 8309 27013 8343 27047
rect 9505 27013 9539 27047
rect 11989 27013 12023 27047
rect 19073 27013 19107 27047
rect 23029 27013 23063 27047
rect 26433 27013 26467 27047
rect 28641 27013 28675 27047
rect 34897 27013 34931 27047
rect 1777 26945 1811 26979
rect 9137 26945 9171 26979
rect 10425 26945 10459 26979
rect 14013 26945 14047 26979
rect 14102 26945 14136 26979
rect 14197 26945 14231 26979
rect 14381 26945 14415 26979
rect 15577 26945 15611 26979
rect 16911 26945 16945 26979
rect 17046 26945 17080 26979
rect 17162 26945 17196 26979
rect 17325 26945 17359 26979
rect 18061 26945 18095 26979
rect 18153 26945 18187 26979
rect 18245 26945 18279 26979
rect 18429 26945 18463 26979
rect 18889 26945 18923 26979
rect 20269 26945 20303 26979
rect 23213 26945 23247 26979
rect 24961 26945 24995 26979
rect 25053 26945 25087 26979
rect 25166 26951 25200 26985
rect 25329 26945 25363 26979
rect 26065 26945 26099 26979
rect 26249 26945 26283 26979
rect 27629 26945 27663 26979
rect 27718 26951 27752 26985
rect 27813 26945 27847 26979
rect 27997 26945 28031 26979
rect 28457 26945 28491 26979
rect 31217 26945 31251 26979
rect 32873 26945 32907 26979
rect 32965 26945 32999 26979
rect 33057 26945 33091 26979
rect 33241 26945 33275 26979
rect 35081 26945 35115 26979
rect 2789 26877 2823 26911
rect 10149 26877 10183 26911
rect 15301 26877 15335 26911
rect 20545 26877 20579 26911
rect 28825 26877 28859 26911
rect 8677 26809 8711 26843
rect 8493 26741 8527 26775
rect 9505 26741 9539 26775
rect 9689 26741 9723 26775
rect 13737 26741 13771 26775
rect 16681 26741 16715 26775
rect 17785 26741 17819 26775
rect 19257 26741 19291 26775
rect 24685 26741 24719 26775
rect 27353 26741 27387 26775
rect 31309 26741 31343 26775
rect 32597 26741 32631 26775
rect 35265 26741 35299 26775
rect 11437 26537 11471 26571
rect 13461 26537 13495 26571
rect 26709 26537 26743 26571
rect 29561 26537 29595 26571
rect 31769 26537 31803 26571
rect 10333 26469 10367 26503
rect 11621 26469 11655 26503
rect 20637 26469 20671 26503
rect 34161 26469 34195 26503
rect 1409 26401 1443 26435
rect 2789 26401 2823 26435
rect 16773 26401 16807 26435
rect 24869 26401 24903 26435
rect 27169 26401 27203 26435
rect 27353 26401 27387 26435
rect 30021 26401 30055 26435
rect 30113 26401 30147 26435
rect 37013 26401 37047 26435
rect 8953 26333 8987 26367
rect 12173 26333 12207 26367
rect 13369 26333 13403 26367
rect 13553 26333 13587 26367
rect 14197 26333 14231 26367
rect 14464 26333 14498 26367
rect 17029 26333 17063 26367
rect 19257 26333 19291 26367
rect 25125 26333 25159 26367
rect 30941 26333 30975 26367
rect 31585 26333 31619 26367
rect 32781 26333 32815 26367
rect 33037 26333 33071 26367
rect 34989 26333 35023 26367
rect 35081 26333 35115 26367
rect 35173 26333 35207 26367
rect 35357 26333 35391 26367
rect 1593 26265 1627 26299
rect 9220 26265 9254 26299
rect 11253 26265 11287 26299
rect 11469 26265 11503 26299
rect 12357 26265 12391 26299
rect 19502 26265 19536 26299
rect 31125 26265 31159 26299
rect 37197 26265 37231 26299
rect 38853 26265 38887 26299
rect 47961 26265 47995 26299
rect 48145 26265 48179 26299
rect 12541 26197 12575 26231
rect 15577 26197 15611 26231
rect 18153 26197 18187 26231
rect 26249 26197 26283 26231
rect 27077 26197 27111 26231
rect 29929 26197 29963 26231
rect 34713 26197 34747 26231
rect 2237 25993 2271 26027
rect 9137 25993 9171 26027
rect 10333 25993 10367 26027
rect 15301 25993 15335 26027
rect 17601 25993 17635 26027
rect 19533 25993 19567 26027
rect 20269 25993 20303 26027
rect 27353 25993 27387 26027
rect 29285 25993 29319 26027
rect 34345 25993 34379 26027
rect 37381 25993 37415 26027
rect 12081 25925 12115 25959
rect 33977 25925 34011 25959
rect 35418 25925 35452 25959
rect 1409 25857 1443 25891
rect 2145 25857 2179 25891
rect 7113 25857 7147 25891
rect 9321 25857 9355 25891
rect 9965 25857 9999 25891
rect 12817 25857 12851 25891
rect 14933 25857 14967 25891
rect 15761 25857 15795 25891
rect 17233 25857 17267 25891
rect 17417 25857 17451 25891
rect 18409 25857 18443 25891
rect 20085 25857 20119 25891
rect 20821 25857 20855 25891
rect 22477 25857 22511 25891
rect 23489 25857 23523 25891
rect 23756 25857 23790 25891
rect 25605 25857 25639 25891
rect 25697 25857 25731 25891
rect 25789 25857 25823 25891
rect 25973 25857 26007 25891
rect 27169 25857 27203 25891
rect 28161 25857 28195 25891
rect 30757 25857 30791 25891
rect 32137 25857 32171 25891
rect 33057 25857 33091 25891
rect 34161 25857 34195 25891
rect 37289 25857 37323 25891
rect 15025 25789 15059 25823
rect 18153 25789 18187 25823
rect 25329 25789 25363 25823
rect 27905 25789 27939 25823
rect 30941 25789 30975 25823
rect 35173 25789 35207 25823
rect 11713 25721 11747 25755
rect 36553 25721 36587 25755
rect 1593 25653 1627 25687
rect 7205 25653 7239 25687
rect 10333 25653 10367 25687
rect 10517 25653 10551 25687
rect 12081 25653 12115 25687
rect 12265 25653 12299 25687
rect 13001 25653 13035 25687
rect 15853 25653 15887 25687
rect 20913 25653 20947 25687
rect 22569 25653 22603 25687
rect 24869 25653 24903 25687
rect 11069 25449 11103 25483
rect 12725 25449 12759 25483
rect 24777 25449 24811 25483
rect 27537 25449 27571 25483
rect 6561 25313 6595 25347
rect 6745 25313 6779 25347
rect 8125 25313 8159 25347
rect 17877 25313 17911 25347
rect 20177 25313 20211 25347
rect 20361 25313 20395 25347
rect 21557 25313 21591 25347
rect 30573 25313 30607 25347
rect 31769 25313 31803 25347
rect 37381 25313 37415 25347
rect 9137 25245 9171 25279
rect 10885 25245 10919 25279
rect 11621 25245 11655 25279
rect 11713 25245 11747 25279
rect 12725 25245 12759 25279
rect 13001 25245 13035 25279
rect 14105 25245 14139 25279
rect 14289 25245 14323 25279
rect 18107 25245 18141 25279
rect 18245 25245 18279 25279
rect 18337 25245 18371 25279
rect 18521 25245 18555 25279
rect 24409 25245 24443 25279
rect 27353 25245 27387 25279
rect 28621 25245 28655 25279
rect 28733 25245 28767 25279
rect 28825 25245 28859 25279
rect 29009 25245 29043 25279
rect 29929 25245 29963 25279
rect 30389 25245 30423 25279
rect 32689 25245 32723 25279
rect 34989 25245 35023 25279
rect 35081 25245 35115 25279
rect 35173 25245 35207 25279
rect 35357 25245 35391 25279
rect 36737 25245 36771 25279
rect 47869 25245 47903 25279
rect 10701 25177 10735 25211
rect 24593 25177 24627 25211
rect 29561 25177 29595 25211
rect 29745 25177 29779 25211
rect 32956 25177 32990 25211
rect 36829 25177 36863 25211
rect 37565 25177 37599 25211
rect 39221 25177 39255 25211
rect 8953 25109 8987 25143
rect 11897 25109 11931 25143
rect 12909 25109 12943 25143
rect 14473 25109 14507 25143
rect 28365 25109 28399 25143
rect 34069 25109 34103 25143
rect 34713 25109 34747 25143
rect 48053 25109 48087 25143
rect 30757 24905 30791 24939
rect 31401 24905 31435 24939
rect 14841 24837 14875 24871
rect 22100 24837 22134 24871
rect 27813 24837 27847 24871
rect 28013 24837 28047 24871
rect 32505 24837 32539 24871
rect 35624 24837 35658 24871
rect 7757 24769 7791 24803
rect 8024 24769 8058 24803
rect 10149 24769 10183 24803
rect 10333 24769 10367 24803
rect 14933 24769 14967 24803
rect 26065 24769 26099 24803
rect 26985 24769 27019 24803
rect 27169 24769 27203 24803
rect 27353 24769 27387 24803
rect 28733 24769 28767 24803
rect 28917 24769 28951 24803
rect 29633 24769 29667 24803
rect 31217 24769 31251 24803
rect 37473 24769 37507 24803
rect 38117 24769 38151 24803
rect 47593 24769 47627 24803
rect 14473 24701 14507 24735
rect 21833 24701 21867 24735
rect 29377 24701 29411 24735
rect 34253 24701 34287 24735
rect 35357 24701 35391 24735
rect 23213 24633 23247 24667
rect 9137 24565 9171 24599
rect 10241 24565 10275 24599
rect 14657 24565 14691 24599
rect 26065 24565 26099 24599
rect 27997 24565 28031 24599
rect 28181 24565 28215 24599
rect 36737 24565 36771 24599
rect 37565 24565 37599 24599
rect 38209 24565 38243 24599
rect 47041 24565 47075 24599
rect 47685 24565 47719 24599
rect 9873 24361 9907 24395
rect 12725 24361 12759 24395
rect 23397 24361 23431 24395
rect 30113 24361 30147 24395
rect 32413 24361 32447 24395
rect 33333 24361 33367 24395
rect 35909 24361 35943 24395
rect 9321 24293 9355 24327
rect 9413 24293 9447 24327
rect 11161 24293 11195 24327
rect 10241 24225 10275 24259
rect 11805 24225 11839 24259
rect 13093 24225 13127 24259
rect 13185 24225 13219 24259
rect 14473 24225 14507 24259
rect 37657 24225 37691 24259
rect 46305 24225 46339 24259
rect 46489 24225 46523 24259
rect 48145 24225 48179 24259
rect 10057 24157 10091 24191
rect 10149 24157 10183 24191
rect 10333 24157 10367 24191
rect 11897 24157 11931 24191
rect 12909 24157 12943 24191
rect 13001 24157 13035 24191
rect 14105 24157 14139 24191
rect 14289 24157 14323 24191
rect 14381 24157 14415 24191
rect 14657 24157 14691 24191
rect 15301 24157 15335 24191
rect 15485 24157 15519 24191
rect 16037 24157 16071 24191
rect 17785 24157 17819 24191
rect 18337 24157 18371 24191
rect 18429 24157 18463 24191
rect 18521 24157 18555 24191
rect 18705 24157 18739 24191
rect 24409 24157 24443 24191
rect 26065 24157 26099 24191
rect 26249 24157 26283 24191
rect 26709 24157 26743 24191
rect 28549 24157 28583 24191
rect 28733 24157 28767 24191
rect 33609 24157 33643 24191
rect 33701 24157 33735 24191
rect 33793 24157 33827 24191
rect 33977 24157 34011 24191
rect 35081 24157 35115 24191
rect 35541 24157 35575 24191
rect 37473 24157 37507 24191
rect 1869 24089 1903 24123
rect 2053 24089 2087 24123
rect 8953 24089 8987 24123
rect 10977 24089 11011 24123
rect 16304 24089 16338 24123
rect 20453 24089 20487 24123
rect 20637 24089 20671 24123
rect 22109 24089 22143 24123
rect 26976 24089 27010 24123
rect 30021 24089 30055 24123
rect 31125 24089 31159 24123
rect 34713 24089 34747 24123
rect 34897 24089 34931 24123
rect 35725 24089 35759 24123
rect 39313 24089 39347 24123
rect 12265 24021 12299 24055
rect 14841 24021 14875 24055
rect 15485 24021 15519 24055
rect 17417 24021 17451 24055
rect 18061 24021 18095 24055
rect 20821 24021 20855 24055
rect 24501 24021 24535 24055
rect 26157 24021 26191 24055
rect 28089 24021 28123 24055
rect 28641 24021 28675 24055
rect 8861 23817 8895 23851
rect 10977 23817 11011 23851
rect 14013 23817 14047 23851
rect 15777 23817 15811 23851
rect 16681 23817 16715 23851
rect 27813 23817 27847 23851
rect 29653 23817 29687 23851
rect 48053 23817 48087 23851
rect 14933 23749 14967 23783
rect 15577 23749 15611 23783
rect 18490 23749 18524 23783
rect 24317 23749 24351 23783
rect 25421 23749 25455 23783
rect 47961 23749 47995 23783
rect 8401 23681 8435 23715
rect 9321 23681 9355 23715
rect 10241 23681 10275 23715
rect 10425 23681 10459 23715
rect 10609 23681 10643 23715
rect 10793 23681 10827 23715
rect 11529 23681 11563 23715
rect 11713 23681 11747 23715
rect 11805 23681 11839 23715
rect 11902 23671 11936 23705
rect 12633 23681 12667 23715
rect 13829 23681 13863 23715
rect 14105 23681 14139 23715
rect 14749 23681 14783 23715
rect 16957 23681 16991 23715
rect 17049 23681 17083 23715
rect 17141 23681 17175 23715
rect 17325 23681 17359 23715
rect 20913 23681 20947 23715
rect 21005 23681 21039 23715
rect 21102 23684 21136 23718
rect 21281 23681 21315 23715
rect 22477 23681 22511 23715
rect 22744 23681 22778 23715
rect 24593 23681 24627 23715
rect 24682 23681 24716 23715
rect 24777 23681 24811 23715
rect 24961 23681 24995 23715
rect 25605 23681 25639 23715
rect 27445 23681 27479 23715
rect 27629 23681 27663 23715
rect 29837 23681 29871 23715
rect 30113 23681 30147 23715
rect 31033 23681 31067 23715
rect 31309 23681 31343 23715
rect 32137 23681 32171 23715
rect 33333 23681 33367 23715
rect 34713 23681 34747 23715
rect 34818 23681 34852 23715
rect 34918 23687 34952 23721
rect 35081 23681 35115 23715
rect 35541 23681 35575 23715
rect 35733 23681 35767 23715
rect 37381 23681 37415 23715
rect 10517 23613 10551 23647
rect 18245 23613 18279 23647
rect 30757 23613 30791 23647
rect 31217 23613 31251 23647
rect 37565 23613 37599 23647
rect 39221 23613 39255 23647
rect 11529 23545 11563 23579
rect 23857 23545 23891 23579
rect 31493 23545 31527 23579
rect 35909 23545 35943 23579
rect 2053 23477 2087 23511
rect 8677 23477 8711 23511
rect 9413 23477 9447 23511
rect 9781 23477 9815 23511
rect 12449 23477 12483 23511
rect 13645 23477 13679 23511
rect 15117 23477 15151 23511
rect 15761 23477 15795 23511
rect 15945 23477 15979 23511
rect 19625 23477 19659 23511
rect 20637 23477 20671 23511
rect 25789 23477 25823 23511
rect 30297 23477 30331 23511
rect 31033 23477 31067 23511
rect 34437 23477 34471 23511
rect 25789 23273 25823 23307
rect 27445 23273 27479 23307
rect 29929 23273 29963 23307
rect 10609 23205 10643 23239
rect 13369 23205 13403 23239
rect 16865 23205 16899 23239
rect 19625 23205 19659 23239
rect 1409 23137 1443 23171
rect 2789 23137 2823 23171
rect 10333 23137 10367 23171
rect 10425 23137 10459 23171
rect 14105 23137 14139 23171
rect 15669 23137 15703 23171
rect 24409 23137 24443 23171
rect 29745 23137 29779 23171
rect 34713 23137 34747 23171
rect 9965 23069 9999 23103
rect 11989 23069 12023 23103
rect 14381 23069 14415 23103
rect 15577 23069 15611 23103
rect 16681 23069 16715 23103
rect 17325 23069 17359 23103
rect 17581 23069 17615 23103
rect 20453 23069 20487 23103
rect 22293 23069 22327 23103
rect 26801 23069 26835 23103
rect 26985 23069 27019 23103
rect 27629 23069 27663 23103
rect 28549 23069 28583 23103
rect 29929 23069 29963 23103
rect 30665 23069 30699 23103
rect 31769 23069 31803 23103
rect 33333 23069 33367 23103
rect 48145 23069 48179 23103
rect 1593 23001 1627 23035
rect 12256 23001 12290 23035
rect 16497 23001 16531 23035
rect 19257 23001 19291 23035
rect 19441 23001 19475 23035
rect 20720 23001 20754 23035
rect 22538 23001 22572 23035
rect 24676 23001 24710 23035
rect 28181 23001 28215 23035
rect 29653 23001 29687 23035
rect 31033 23001 31067 23035
rect 34958 23001 34992 23035
rect 15945 22933 15979 22967
rect 18705 22933 18739 22967
rect 21833 22933 21867 22967
rect 23673 22933 23707 22967
rect 30113 22933 30147 22967
rect 36093 22933 36127 22967
rect 47961 22933 47995 22967
rect 2605 22729 2639 22763
rect 10977 22729 11011 22763
rect 14473 22729 14507 22763
rect 17877 22729 17911 22763
rect 24041 22729 24075 22763
rect 2053 22661 2087 22695
rect 13277 22661 13311 22695
rect 13493 22661 13527 22695
rect 14381 22661 14415 22695
rect 14590 22661 14624 22695
rect 20637 22661 20671 22695
rect 25145 22661 25179 22695
rect 25789 22661 25823 22695
rect 31033 22661 31067 22695
rect 1869 22593 1903 22627
rect 2513 22593 2547 22627
rect 9873 22593 9907 22627
rect 10701 22593 10735 22627
rect 17601 22593 17635 22627
rect 18107 22593 18141 22627
rect 18245 22593 18279 22627
rect 18337 22593 18371 22627
rect 18521 22593 18555 22627
rect 20913 22593 20947 22627
rect 21005 22593 21039 22627
rect 21102 22593 21136 22627
rect 21281 22593 21315 22627
rect 24225 22593 24259 22627
rect 24409 22593 24443 22627
rect 24501 22593 24535 22627
rect 24961 22593 24995 22627
rect 25237 22593 25271 22627
rect 25697 22593 25731 22627
rect 25881 22593 25915 22627
rect 29469 22593 29503 22627
rect 29745 22593 29779 22627
rect 31349 22593 31383 22627
rect 32229 22593 32263 22627
rect 32781 22593 32815 22627
rect 35725 22593 35759 22627
rect 35909 22593 35943 22627
rect 47593 22593 47627 22627
rect 47777 22593 47811 22627
rect 9965 22525 9999 22559
rect 10241 22525 10275 22559
rect 10977 22525 11011 22559
rect 14112 22525 14146 22559
rect 29561 22525 29595 22559
rect 31217 22525 31251 22559
rect 33425 22525 33459 22559
rect 33609 22525 33643 22559
rect 35265 22525 35299 22559
rect 10793 22457 10827 22491
rect 13645 22457 13679 22491
rect 24961 22457 24995 22491
rect 31493 22457 31527 22491
rect 13461 22389 13495 22423
rect 14749 22389 14783 22423
rect 29469 22389 29503 22423
rect 29929 22389 29963 22423
rect 31033 22389 31067 22423
rect 36093 22389 36127 22423
rect 47685 22389 47719 22423
rect 18153 22185 18187 22219
rect 20913 22185 20947 22219
rect 28825 22185 28859 22219
rect 29745 22185 29779 22219
rect 30205 22185 30239 22219
rect 30849 22185 30883 22219
rect 31309 22185 31343 22219
rect 47869 22185 47903 22219
rect 10057 22117 10091 22151
rect 14289 22117 14323 22151
rect 20085 22117 20119 22151
rect 36369 22117 36403 22151
rect 14473 22049 14507 22083
rect 25605 22049 25639 22083
rect 28641 22049 28675 22083
rect 29837 22049 29871 22083
rect 30941 22049 30975 22083
rect 47409 22049 47443 22083
rect 6837 21981 6871 22015
rect 9965 21981 9999 22015
rect 14197 21981 14231 22015
rect 17785 21981 17819 22015
rect 17969 21981 18003 22015
rect 19901 21981 19935 22015
rect 25145 21981 25179 22015
rect 25513 21981 25547 22015
rect 26249 21981 26283 22015
rect 26433 21981 26467 22015
rect 26893 21981 26927 22015
rect 28825 21981 28859 22015
rect 30021 21981 30055 22015
rect 31125 21981 31159 22015
rect 31953 21981 31987 22015
rect 33793 21981 33827 22015
rect 33885 21981 33919 22015
rect 33977 21981 34011 22015
rect 34161 21981 34195 22015
rect 34989 21981 35023 22015
rect 36921 21981 36955 22015
rect 47501 21981 47535 22015
rect 47869 21981 47903 22015
rect 7104 21913 7138 21947
rect 10241 21913 10275 21947
rect 14473 21913 14507 21947
rect 20545 21913 20579 21947
rect 20729 21913 20763 21947
rect 28549 21913 28583 21947
rect 29561 21913 29595 21947
rect 30849 21913 30883 21947
rect 32597 21913 32631 21947
rect 33517 21913 33551 21947
rect 35234 21913 35268 21947
rect 37105 21913 37139 21947
rect 38761 21913 38795 21947
rect 8217 21845 8251 21879
rect 9965 21845 9999 21879
rect 25237 21845 25271 21879
rect 26433 21845 26467 21879
rect 26985 21845 27019 21879
rect 29009 21845 29043 21879
rect 30573 21845 30607 21879
rect 48053 21845 48087 21879
rect 14657 21641 14691 21675
rect 15761 21641 15795 21675
rect 19533 21641 19567 21675
rect 25053 21641 25087 21675
rect 25973 21641 26007 21675
rect 29837 21641 29871 21675
rect 31585 21641 31619 21675
rect 32597 21641 32631 21675
rect 33149 21641 33183 21675
rect 36369 21641 36403 21675
rect 37381 21641 37415 21675
rect 22928 21573 22962 21607
rect 26341 21573 26375 21607
rect 26985 21573 27019 21607
rect 47961 21573 47995 21607
rect 7297 21505 7331 21539
rect 14197 21505 14231 21539
rect 14473 21505 14507 21539
rect 15393 21505 15427 21539
rect 19717 21505 19751 21539
rect 20177 21505 20211 21539
rect 21099 21505 21133 21539
rect 21833 21505 21867 21539
rect 22017 21505 22051 21539
rect 22661 21505 22695 21539
rect 24961 21505 24995 21539
rect 26065 21505 26099 21539
rect 26157 21505 26191 21539
rect 27261 21505 27295 21539
rect 28273 21505 28307 21539
rect 28549 21505 28583 21539
rect 29377 21505 29411 21539
rect 29653 21505 29687 21539
rect 31125 21505 31159 21539
rect 31401 21505 31435 21539
rect 32137 21505 32171 21539
rect 32413 21505 32447 21539
rect 33057 21505 33091 21539
rect 36277 21505 36311 21539
rect 37289 21505 37323 21539
rect 7481 21437 7515 21471
rect 7757 21437 7791 21471
rect 11529 21437 11563 21471
rect 11713 21437 11747 21471
rect 13093 21437 13127 21471
rect 14381 21437 14415 21471
rect 15301 21437 15335 21471
rect 25789 21437 25823 21471
rect 27169 21437 27203 21471
rect 28365 21437 28399 21471
rect 29561 21437 29595 21471
rect 31217 21437 31251 21471
rect 32321 21437 32355 21471
rect 33701 21437 33735 21471
rect 33885 21437 33919 21471
rect 35541 21437 35575 21471
rect 29101 21369 29135 21403
rect 14473 21301 14507 21335
rect 20361 21301 20395 21335
rect 21189 21301 21223 21335
rect 22201 21301 22235 21335
rect 24041 21301 24075 21335
rect 27261 21301 27295 21335
rect 27445 21301 27479 21335
rect 28273 21301 28307 21335
rect 28733 21301 28767 21335
rect 29377 21301 29411 21335
rect 30757 21301 30791 21335
rect 31401 21301 31435 21335
rect 32137 21301 32171 21335
rect 48053 21301 48087 21335
rect 7573 21097 7607 21131
rect 12173 21097 12207 21131
rect 22477 21097 22511 21131
rect 27445 21097 27479 21131
rect 28365 21097 28399 21131
rect 28825 21097 28859 21131
rect 29837 21097 29871 21131
rect 31217 21097 31251 21131
rect 14473 20961 14507 20995
rect 16865 20961 16899 20995
rect 25605 20961 25639 20995
rect 26801 20961 26835 20995
rect 26893 20961 26927 20995
rect 27629 20961 27663 20995
rect 28457 20961 28491 20995
rect 29653 20961 29687 20995
rect 36093 20961 36127 20995
rect 36277 20961 36311 20995
rect 7481 20893 7515 20927
rect 12081 20893 12115 20927
rect 13165 20893 13199 20927
rect 13274 20893 13308 20927
rect 13390 20893 13424 20927
rect 13547 20893 13581 20927
rect 19717 20893 19751 20927
rect 21005 20893 21039 20927
rect 21281 20893 21315 20927
rect 22753 20893 22787 20927
rect 22845 20893 22879 20927
rect 22937 20893 22971 20927
rect 23121 20893 23155 20927
rect 25513 20893 25547 20927
rect 25697 20893 25731 20927
rect 26433 20893 26467 20927
rect 27445 20893 27479 20927
rect 27721 20893 27755 20927
rect 28365 20893 28399 20927
rect 28641 20893 28675 20927
rect 29837 20893 29871 20927
rect 31401 20893 31435 20927
rect 31493 20893 31527 20927
rect 33425 20893 33459 20927
rect 38393 20893 38427 20927
rect 14105 20825 14139 20859
rect 14289 20825 14323 20859
rect 17132 20825 17166 20859
rect 26341 20825 26375 20859
rect 29561 20825 29595 20859
rect 31217 20825 31251 20859
rect 37933 20825 37967 20859
rect 12909 20757 12943 20791
rect 18245 20757 18279 20791
rect 19809 20757 19843 20791
rect 27905 20757 27939 20791
rect 30021 20757 30055 20791
rect 31677 20757 31711 20791
rect 33517 20757 33551 20791
rect 38485 20757 38519 20791
rect 17509 20553 17543 20587
rect 13338 20485 13372 20519
rect 22661 20485 22695 20519
rect 27445 20485 27479 20519
rect 30573 20485 30607 20519
rect 30849 20485 30883 20519
rect 33701 20485 33735 20519
rect 37473 20485 37507 20519
rect 39129 20485 39163 20519
rect 4813 20417 4847 20451
rect 11529 20417 11563 20451
rect 11713 20417 11747 20451
rect 13093 20417 13127 20451
rect 15761 20417 15795 20451
rect 15853 20417 15887 20451
rect 15945 20417 15979 20451
rect 16129 20417 16163 20451
rect 17765 20417 17799 20451
rect 17874 20423 17908 20457
rect 17969 20417 18003 20451
rect 18153 20417 18187 20451
rect 18889 20417 18923 20451
rect 19800 20417 19834 20451
rect 21833 20417 21867 20451
rect 22017 20417 22051 20451
rect 22109 20417 22143 20451
rect 23857 20417 23891 20451
rect 28641 20417 28675 20451
rect 28917 20417 28951 20451
rect 29561 20417 29595 20451
rect 29745 20417 29779 20451
rect 29837 20417 29871 20451
rect 31125 20417 31159 20451
rect 32873 20417 32907 20451
rect 47593 20417 47627 20451
rect 8769 20349 8803 20383
rect 8953 20349 8987 20383
rect 10425 20349 10459 20383
rect 17233 20349 17267 20383
rect 19533 20349 19567 20383
rect 24041 20349 24075 20383
rect 28825 20349 28859 20383
rect 31033 20349 31067 20383
rect 33517 20349 33551 20383
rect 34069 20349 34103 20383
rect 37289 20349 37323 20383
rect 21833 20281 21867 20315
rect 29101 20281 29135 20315
rect 31309 20281 31343 20315
rect 4905 20213 4939 20247
rect 11897 20213 11931 20247
rect 14473 20213 14507 20247
rect 15485 20213 15519 20247
rect 18981 20213 19015 20247
rect 20913 20213 20947 20247
rect 22753 20213 22787 20247
rect 27721 20213 27755 20247
rect 28641 20213 28675 20247
rect 29561 20213 29595 20247
rect 30021 20213 30055 20247
rect 30849 20213 30883 20247
rect 32965 20213 32999 20247
rect 47685 20213 47719 20247
rect 8309 20009 8343 20043
rect 11713 20009 11747 20043
rect 14749 20009 14783 20043
rect 16957 20009 16991 20043
rect 17693 20009 17727 20043
rect 19717 20009 19751 20043
rect 28457 20009 28491 20043
rect 28917 20009 28951 20043
rect 30389 20009 30423 20043
rect 30573 20009 30607 20043
rect 33885 20009 33919 20043
rect 20913 19941 20947 19975
rect 4721 19873 4755 19907
rect 4905 19873 4939 19907
rect 5549 19873 5583 19907
rect 10333 19873 10367 19907
rect 12633 19873 12667 19907
rect 21833 19873 21867 19907
rect 28549 19873 28583 19907
rect 30205 19873 30239 19907
rect 46489 19873 46523 19907
rect 2053 19805 2087 19839
rect 8217 19805 8251 19839
rect 9459 19805 9493 19839
rect 9597 19805 9631 19839
rect 9689 19805 9723 19839
rect 9873 19805 9907 19839
rect 12081 19805 12115 19839
rect 12357 19805 12391 19839
rect 15209 19805 15243 19839
rect 18245 19805 18279 19839
rect 19901 19805 19935 19839
rect 20177 19805 20211 19839
rect 20729 19805 20763 19839
rect 21649 19805 21683 19839
rect 22385 19805 22419 19839
rect 27261 19805 27295 19839
rect 27353 19805 27387 19839
rect 28457 19805 28491 19839
rect 28733 19805 28767 19839
rect 30113 19805 30147 19839
rect 30389 19805 30423 19839
rect 33793 19805 33827 19839
rect 46305 19805 46339 19839
rect 10600 19737 10634 19771
rect 14381 19737 14415 19771
rect 14565 19737 14599 19771
rect 15476 19737 15510 19771
rect 16865 19737 16899 19771
rect 17325 19737 17359 19771
rect 17509 19737 17543 19771
rect 18613 19737 18647 19771
rect 31585 19737 31619 19771
rect 48145 19737 48179 19771
rect 9229 19669 9263 19703
rect 16589 19669 16623 19703
rect 20085 19669 20119 19703
rect 22477 19669 22511 19703
rect 27261 19669 27295 19703
rect 32873 19669 32907 19703
rect 9413 19465 9447 19499
rect 10241 19465 10275 19499
rect 11529 19465 11563 19499
rect 21281 19465 21315 19499
rect 24777 19465 24811 19499
rect 8300 19397 8334 19431
rect 10057 19397 10091 19431
rect 12725 19397 12759 19431
rect 17233 19397 17267 19431
rect 18797 19397 18831 19431
rect 20453 19397 20487 19431
rect 25881 19397 25915 19431
rect 26985 19397 27019 19431
rect 27169 19397 27203 19431
rect 33333 19397 33367 19431
rect 1777 19329 1811 19363
rect 8033 19329 8067 19363
rect 9873 19329 9907 19363
rect 11805 19329 11839 19363
rect 11897 19329 11931 19363
rect 11989 19329 12023 19363
rect 12173 19329 12207 19363
rect 13645 19329 13679 19363
rect 14289 19329 14323 19363
rect 14473 19329 14507 19363
rect 15117 19329 15151 19363
rect 19717 19329 19751 19363
rect 20353 19329 20387 19363
rect 21097 19329 21131 19363
rect 21281 19329 21315 19363
rect 21833 19329 21867 19363
rect 22845 19329 22879 19363
rect 23101 19329 23135 19363
rect 24685 19329 24719 19363
rect 25697 19329 25731 19363
rect 32137 19329 32171 19363
rect 36461 19329 36495 19363
rect 37289 19329 37323 19363
rect 47869 19329 47903 19363
rect 1961 19261 1995 19295
rect 2237 19261 2271 19295
rect 12909 19261 12943 19295
rect 13829 19261 13863 19295
rect 14657 19261 14691 19295
rect 15393 19261 15427 19295
rect 25513 19261 25547 19295
rect 33149 19261 33183 19295
rect 34161 19261 34195 19295
rect 19073 19193 19107 19227
rect 27353 19193 27387 19227
rect 32321 19193 32355 19227
rect 17325 19125 17359 19159
rect 19809 19125 19843 19159
rect 22017 19125 22051 19159
rect 24225 19125 24259 19159
rect 36553 19125 36587 19159
rect 37381 19125 37415 19159
rect 48053 19125 48087 19159
rect 2237 18921 2271 18955
rect 22385 18921 22419 18955
rect 33333 18921 33367 18955
rect 47685 18921 47719 18955
rect 23857 18853 23891 18887
rect 24409 18853 24443 18887
rect 14473 18785 14507 18819
rect 21097 18785 21131 18819
rect 23581 18785 23615 18819
rect 25053 18785 25087 18819
rect 36553 18785 36587 18819
rect 2145 18717 2179 18751
rect 9321 18717 9355 18751
rect 9413 18717 9447 18751
rect 9505 18717 9539 18751
rect 9689 18717 9723 18751
rect 11621 18717 11655 18751
rect 11710 18717 11744 18751
rect 11805 18717 11839 18751
rect 11989 18717 12023 18751
rect 13185 18717 13219 18751
rect 13274 18717 13308 18751
rect 13374 18717 13408 18751
rect 13553 18717 13587 18751
rect 14289 18717 14323 18751
rect 16129 18717 16163 18751
rect 17141 18717 17175 18751
rect 19901 18717 19935 18751
rect 19993 18717 20027 18751
rect 20085 18717 20119 18751
rect 20269 18717 20303 18751
rect 21557 18717 21591 18751
rect 21741 18717 21775 18751
rect 22569 18717 22603 18751
rect 22845 18717 22879 18751
rect 23489 18717 23523 18751
rect 25605 18717 25639 18751
rect 25881 18717 25915 18751
rect 26801 18717 26835 18751
rect 27445 18717 27479 18751
rect 27629 18717 27663 18751
rect 29745 18717 29779 18751
rect 31953 18717 31987 18751
rect 34897 18717 34931 18751
rect 36369 18717 36403 18751
rect 14105 18649 14139 18683
rect 17386 18649 17420 18683
rect 20729 18649 20763 18683
rect 20913 18649 20947 18683
rect 24869 18649 24903 18683
rect 27813 18649 27847 18683
rect 32220 18649 32254 18683
rect 34713 18649 34747 18683
rect 38209 18649 38243 18683
rect 9045 18581 9079 18615
rect 11345 18581 11379 18615
rect 12909 18581 12943 18615
rect 16221 18581 16255 18615
rect 18521 18581 18555 18615
rect 19625 18581 19659 18615
rect 21649 18581 21683 18615
rect 22753 18581 22787 18615
rect 24777 18581 24811 18615
rect 25697 18581 25731 18615
rect 26893 18581 26927 18615
rect 29561 18581 29595 18615
rect 35081 18581 35115 18615
rect 10885 18377 10919 18411
rect 11897 18377 11931 18411
rect 14381 18377 14415 18411
rect 15945 18377 15979 18411
rect 16865 18377 16899 18411
rect 24133 18377 24167 18411
rect 26065 18377 26099 18411
rect 27261 18377 27295 18411
rect 28181 18377 28215 18411
rect 32137 18377 32171 18411
rect 35633 18377 35667 18411
rect 11529 18309 11563 18343
rect 13246 18309 13280 18343
rect 29622 18309 29656 18343
rect 33609 18309 33643 18343
rect 37473 18309 37507 18343
rect 39129 18309 39163 18343
rect 2053 18241 2087 18275
rect 6837 18241 6871 18275
rect 7481 18241 7515 18275
rect 7748 18241 7782 18275
rect 9669 18241 9703 18275
rect 9781 18241 9815 18275
rect 9873 18241 9907 18275
rect 10057 18241 10091 18275
rect 10517 18241 10551 18275
rect 10701 18241 10735 18275
rect 11713 18241 11747 18275
rect 13001 18241 13035 18275
rect 15853 18241 15887 18275
rect 17095 18241 17129 18275
rect 17230 18244 17264 18278
rect 17325 18244 17359 18278
rect 17509 18241 17543 18275
rect 19901 18241 19935 18275
rect 20168 18241 20202 18275
rect 23581 18241 23615 18275
rect 23765 18241 23799 18275
rect 23857 18241 23891 18275
rect 23949 18241 23983 18275
rect 24777 18241 24811 18275
rect 25053 18241 25087 18275
rect 27258 18241 27292 18275
rect 28549 18241 28583 18275
rect 32413 18241 32447 18275
rect 32518 18241 32552 18275
rect 32618 18241 32652 18275
rect 32781 18241 32815 18275
rect 33241 18241 33275 18275
rect 33425 18241 33459 18275
rect 34520 18241 34554 18275
rect 36093 18241 36127 18275
rect 36277 18241 36311 18275
rect 37289 18241 37323 18275
rect 24961 18173 24995 18207
rect 26157 18173 26191 18207
rect 26341 18173 26375 18207
rect 27721 18173 27755 18207
rect 28641 18173 28675 18207
rect 28733 18173 28767 18207
rect 29377 18173 29411 18207
rect 34253 18173 34287 18207
rect 25237 18105 25271 18139
rect 25697 18105 25731 18139
rect 27077 18105 27111 18139
rect 30757 18105 30791 18139
rect 2145 18037 2179 18071
rect 2881 18037 2915 18071
rect 6929 18037 6963 18071
rect 8861 18037 8895 18071
rect 9413 18037 9447 18071
rect 21281 18037 21315 18071
rect 25053 18037 25087 18071
rect 27629 18037 27663 18071
rect 36461 18037 36495 18071
rect 24777 17833 24811 17867
rect 25605 17833 25639 17867
rect 26249 17833 26283 17867
rect 33149 17833 33183 17867
rect 36185 17833 36219 17867
rect 18153 17765 18187 17799
rect 26617 17765 26651 17799
rect 28733 17765 28767 17799
rect 1409 17697 1443 17731
rect 1593 17697 1627 17731
rect 2789 17697 2823 17731
rect 6745 17697 6779 17731
rect 7021 17697 7055 17731
rect 8953 17697 8987 17731
rect 15761 17697 15795 17731
rect 16037 17697 16071 17731
rect 24593 17697 24627 17731
rect 25789 17697 25823 17731
rect 26525 17697 26559 17731
rect 27261 17697 27295 17731
rect 32137 17697 32171 17731
rect 37289 17697 37323 17731
rect 39129 17697 39163 17731
rect 10793 17629 10827 17663
rect 14933 17629 14967 17663
rect 15577 17629 15611 17663
rect 20361 17629 20395 17663
rect 24777 17629 24811 17663
rect 25513 17629 25547 17663
rect 26433 17629 26467 17663
rect 26709 17629 26743 17663
rect 27537 17629 27571 17663
rect 28549 17629 28583 17663
rect 29561 17629 29595 17663
rect 31861 17629 31895 17663
rect 33425 17629 33459 17663
rect 33517 17629 33551 17663
rect 33609 17629 33643 17663
rect 33793 17629 33827 17663
rect 34805 17629 34839 17663
rect 36645 17629 36679 17663
rect 47685 17629 47719 17663
rect 6837 17561 6871 17595
rect 9220 17561 9254 17595
rect 11060 17561 11094 17595
rect 14749 17561 14783 17595
rect 17969 17561 18003 17595
rect 19533 17561 19567 17595
rect 19717 17561 19751 17595
rect 20606 17561 20640 17595
rect 24501 17561 24535 17595
rect 25789 17561 25823 17595
rect 29806 17561 29840 17595
rect 35050 17561 35084 17595
rect 36737 17561 36771 17595
rect 37473 17561 37507 17595
rect 10333 17493 10367 17527
rect 12173 17493 12207 17527
rect 15117 17493 15151 17527
rect 19901 17493 19935 17527
rect 21741 17493 21775 17527
rect 24961 17493 24995 17527
rect 30941 17493 30975 17527
rect 1961 17289 1995 17323
rect 24777 17289 24811 17323
rect 25881 17289 25915 17323
rect 27261 17289 27295 17323
rect 27721 17289 27755 17323
rect 28181 17289 28215 17323
rect 29653 17289 29687 17323
rect 33885 17289 33919 17323
rect 9413 17221 9447 17255
rect 9781 17221 9815 17255
rect 20821 17221 20855 17255
rect 21005 17221 21039 17255
rect 23489 17221 23523 17255
rect 24685 17221 24719 17255
rect 36461 17221 36495 17255
rect 1869 17153 1903 17187
rect 9597 17153 9631 17187
rect 14565 17153 14599 17187
rect 14821 17153 14855 17187
rect 17305 17153 17339 17187
rect 19993 17153 20027 17187
rect 20085 17153 20119 17187
rect 20177 17153 20211 17187
rect 20361 17153 20395 17187
rect 23213 17153 23247 17187
rect 23361 17153 23395 17187
rect 23581 17153 23615 17187
rect 23678 17153 23712 17187
rect 25513 17153 25547 17187
rect 25651 17153 25685 17187
rect 25973 17153 26007 17187
rect 26985 17153 27019 17187
rect 27077 17153 27111 17187
rect 28089 17153 28123 17187
rect 28917 17153 28951 17187
rect 29101 17151 29135 17185
rect 29469 17153 29503 17187
rect 32321 17153 32355 17187
rect 34141 17153 34175 17187
rect 34250 17156 34284 17190
rect 34345 17153 34379 17187
rect 34529 17153 34563 17187
rect 35265 17153 35299 17187
rect 35357 17153 35391 17187
rect 35470 17156 35504 17190
rect 35633 17153 35667 17187
rect 36093 17153 36127 17187
rect 36277 17153 36311 17187
rect 37289 17153 37323 17187
rect 46765 17153 46799 17187
rect 17049 17085 17083 17119
rect 21189 17085 21223 17119
rect 24961 17085 24995 17119
rect 27261 17085 27295 17119
rect 28365 17085 28399 17119
rect 29187 17085 29221 17119
rect 29285 17085 29319 17119
rect 15945 17017 15979 17051
rect 19717 17017 19751 17051
rect 25789 17017 25823 17051
rect 18429 16949 18463 16983
rect 23857 16949 23891 16983
rect 24317 16949 24351 16983
rect 32137 16949 32171 16983
rect 34989 16949 35023 16983
rect 37381 16949 37415 16983
rect 46857 16949 46891 16983
rect 47777 16949 47811 16983
rect 14565 16745 14599 16779
rect 16865 16745 16899 16779
rect 18613 16745 18647 16779
rect 20637 16745 20671 16779
rect 23857 16745 23891 16779
rect 24409 16745 24443 16779
rect 26709 16745 26743 16779
rect 36093 16745 36127 16779
rect 9965 16609 9999 16643
rect 13553 16609 13587 16643
rect 19257 16609 19291 16643
rect 22477 16609 22511 16643
rect 34713 16609 34747 16643
rect 36921 16609 36955 16643
rect 38577 16609 38611 16643
rect 46305 16609 46339 16643
rect 46489 16609 46523 16643
rect 48145 16609 48179 16643
rect 2237 16541 2271 16575
rect 2881 16541 2915 16575
rect 11805 16541 11839 16575
rect 13369 16541 13403 16575
rect 14841 16541 14875 16575
rect 14930 16541 14964 16575
rect 15025 16541 15059 16575
rect 15209 16541 15243 16575
rect 15899 16541 15933 16575
rect 16037 16541 16071 16575
rect 16129 16541 16163 16575
rect 16313 16541 16347 16575
rect 17141 16541 17175 16575
rect 17233 16541 17267 16575
rect 17325 16541 17359 16575
rect 17509 16541 17543 16575
rect 22744 16541 22778 16575
rect 24685 16541 24719 16575
rect 26893 16541 26927 16575
rect 27169 16541 27203 16575
rect 27721 16541 27755 16575
rect 32229 16541 32263 16575
rect 32321 16541 32355 16575
rect 32413 16541 32447 16575
rect 32597 16541 32631 16575
rect 33241 16541 33275 16575
rect 34969 16541 35003 16575
rect 10149 16473 10183 16507
rect 13185 16473 13219 16507
rect 18521 16473 18555 16507
rect 19524 16473 19558 16507
rect 24409 16473 24443 16507
rect 24593 16473 24627 16507
rect 33057 16473 33091 16507
rect 37105 16473 37139 16507
rect 2973 16405 3007 16439
rect 15669 16405 15703 16439
rect 27077 16405 27111 16439
rect 27905 16405 27939 16439
rect 31953 16405 31987 16439
rect 33425 16405 33459 16439
rect 10149 16201 10183 16235
rect 13737 16201 13771 16235
rect 17233 16201 17267 16235
rect 17877 16201 17911 16235
rect 18981 16201 19015 16235
rect 20913 16201 20947 16235
rect 24777 16201 24811 16235
rect 2237 16133 2271 16167
rect 12624 16133 12658 16167
rect 17049 16133 17083 16167
rect 24317 16133 24351 16167
rect 28549 16133 28583 16167
rect 30297 16133 30331 16167
rect 32382 16133 32416 16167
rect 2053 16065 2087 16099
rect 10057 16065 10091 16099
rect 12357 16065 12391 16099
rect 14473 16065 14507 16099
rect 16865 16065 16899 16099
rect 17693 16065 17727 16099
rect 19257 16065 19291 16099
rect 19349 16065 19383 16099
rect 19441 16065 19475 16099
rect 19625 16065 19659 16099
rect 20729 16065 20763 16099
rect 24593 16065 24627 16099
rect 27261 16065 27295 16099
rect 28365 16065 28399 16099
rect 29009 16065 29043 16099
rect 29193 16065 29227 16099
rect 29561 16065 29595 16099
rect 32137 16065 32171 16099
rect 47593 16065 47627 16099
rect 2789 15997 2823 16031
rect 14197 15997 14231 16031
rect 24501 15997 24535 16031
rect 27537 15997 27571 16031
rect 29285 15997 29319 16031
rect 29377 15997 29411 16031
rect 24593 15861 24627 15895
rect 27353 15861 27387 15895
rect 27445 15861 27479 15895
rect 29745 15861 29779 15895
rect 30389 15861 30423 15895
rect 33517 15861 33551 15895
rect 47041 15861 47075 15895
rect 47685 15861 47719 15895
rect 15209 15657 15243 15691
rect 24777 15657 24811 15691
rect 26249 15657 26283 15691
rect 28273 15657 28307 15691
rect 27123 15589 27157 15623
rect 9229 15521 9263 15555
rect 10977 15521 11011 15555
rect 11529 15521 11563 15555
rect 17693 15521 17727 15555
rect 19257 15521 19291 15555
rect 26433 15521 26467 15555
rect 28825 15521 28859 15555
rect 46305 15521 46339 15555
rect 46489 15521 46523 15555
rect 48145 15521 48179 15555
rect 14335 15453 14369 15487
rect 14470 15447 14504 15481
rect 14565 15453 14599 15487
rect 14749 15453 14783 15487
rect 15393 15453 15427 15487
rect 16497 15453 16531 15487
rect 16586 15453 16620 15487
rect 16702 15453 16736 15487
rect 16865 15453 16899 15487
rect 18429 15453 18463 15487
rect 19533 15453 19567 15487
rect 20821 15453 20855 15487
rect 20910 15447 20944 15481
rect 21005 15453 21039 15487
rect 21189 15453 21223 15487
rect 21649 15453 21683 15487
rect 24685 15453 24719 15487
rect 24869 15453 24903 15487
rect 24961 15453 24995 15487
rect 25145 15453 25179 15487
rect 26157 15453 26191 15487
rect 26893 15453 26927 15487
rect 29837 15453 29871 15487
rect 30093 15453 30127 15487
rect 32505 15453 32539 15487
rect 34989 15453 35023 15487
rect 9413 15385 9447 15419
rect 11713 15385 11747 15419
rect 13369 15385 13403 15419
rect 17325 15385 17359 15419
rect 17509 15385 17543 15419
rect 18245 15385 18279 15419
rect 21833 15385 21867 15419
rect 28641 15385 28675 15419
rect 31769 15385 31803 15419
rect 32689 15385 32723 15419
rect 35173 15385 35207 15419
rect 14105 15317 14139 15351
rect 16221 15317 16255 15351
rect 20545 15317 20579 15351
rect 22017 15317 22051 15351
rect 24409 15317 24443 15351
rect 26433 15317 26467 15351
rect 28733 15317 28767 15351
rect 31217 15317 31251 15351
rect 31861 15317 31895 15351
rect 35357 15317 35391 15351
rect 9597 15113 9631 15147
rect 10609 15113 10643 15147
rect 14565 15113 14599 15147
rect 18061 15113 18095 15147
rect 22201 15113 22235 15147
rect 25881 15113 25915 15147
rect 27537 15113 27571 15147
rect 27905 15113 27939 15147
rect 30941 15113 30975 15147
rect 48053 15113 48087 15147
rect 14381 15045 14415 15079
rect 16948 15045 16982 15079
rect 30481 15045 30515 15079
rect 9505 14977 9539 15011
rect 10517 14977 10551 15011
rect 12357 14977 12391 15011
rect 12624 14977 12658 15011
rect 14197 14977 14231 15011
rect 16681 14977 16715 15011
rect 18521 14977 18555 15011
rect 19901 14977 19935 15011
rect 20157 14977 20191 15011
rect 21833 14977 21867 15011
rect 22017 14977 22051 15011
rect 22661 14977 22695 15011
rect 26065 14977 26099 15011
rect 26157 14977 26191 15011
rect 27997 14977 28031 15011
rect 29285 14977 29319 15011
rect 29469 14977 29503 15011
rect 29837 14977 29871 15011
rect 30757 14977 30791 15011
rect 32689 14977 32723 15011
rect 32794 14977 32828 15011
rect 32894 14977 32928 15011
rect 33057 14977 33091 15011
rect 35440 14977 35474 15011
rect 46857 14977 46891 15011
rect 47961 14977 47995 15011
rect 26249 14909 26283 14943
rect 26341 14909 26375 14943
rect 28181 14909 28215 14943
rect 29561 14909 29595 14943
rect 29653 14909 29687 14943
rect 30573 14909 30607 14943
rect 35173 14909 35207 14943
rect 21281 14841 21315 14875
rect 22845 14841 22879 14875
rect 13737 14773 13771 14807
rect 18613 14773 18647 14807
rect 30021 14773 30055 14807
rect 30481 14773 30515 14807
rect 32413 14773 32447 14807
rect 36553 14773 36587 14807
rect 46949 14773 46983 14807
rect 27721 14569 27755 14603
rect 31401 14569 31435 14603
rect 35173 14569 35207 14603
rect 19717 14501 19751 14535
rect 22201 14501 22235 14535
rect 26341 14501 26375 14535
rect 20821 14433 20855 14467
rect 33977 14433 34011 14467
rect 46305 14433 46339 14467
rect 46489 14433 46523 14467
rect 12449 14365 12483 14399
rect 14749 14365 14783 14399
rect 14933 14365 14967 14399
rect 18521 14365 18555 14399
rect 19993 14365 20027 14399
rect 20085 14365 20119 14399
rect 20177 14365 20211 14399
rect 20361 14365 20395 14399
rect 21077 14365 21111 14399
rect 22753 14365 22787 14399
rect 24961 14365 24995 14399
rect 27261 14365 27295 14399
rect 27905 14365 27939 14399
rect 28181 14365 28215 14399
rect 30021 14365 30055 14399
rect 30277 14365 30311 14399
rect 32781 14365 32815 14399
rect 32873 14365 32907 14399
rect 32965 14365 32999 14399
rect 33149 14365 33183 14399
rect 33793 14365 33827 14399
rect 35403 14365 35437 14399
rect 35541 14365 35575 14399
rect 35633 14365 35667 14399
rect 35817 14365 35851 14399
rect 36553 14365 36587 14399
rect 36642 14365 36676 14399
rect 36737 14365 36771 14399
rect 36921 14365 36955 14399
rect 18705 14297 18739 14331
rect 25228 14297 25262 14331
rect 26985 14297 27019 14331
rect 28641 14297 28675 14331
rect 28825 14297 28859 14331
rect 33609 14297 33643 14331
rect 48145 14297 48179 14331
rect 12541 14229 12575 14263
rect 14841 14229 14875 14263
rect 22845 14229 22879 14263
rect 27083 14229 27117 14263
rect 27169 14229 27203 14263
rect 28089 14229 28123 14263
rect 29009 14229 29043 14263
rect 32505 14229 32539 14263
rect 36277 14229 36311 14263
rect 16865 14025 16899 14059
rect 20545 14025 20579 14059
rect 22385 14025 22419 14059
rect 25513 14025 25547 14059
rect 26157 14025 26191 14059
rect 30297 14025 30331 14059
rect 31585 14025 31619 14059
rect 33977 14025 34011 14059
rect 48053 14025 48087 14059
rect 12633 13957 12667 13991
rect 15669 13957 15703 13991
rect 16773 13957 16807 13991
rect 22293 13957 22327 13991
rect 30205 13957 30239 13991
rect 31217 13957 31251 13991
rect 35348 13957 35382 13991
rect 2053 13889 2087 13923
rect 8125 13889 8159 13923
rect 12449 13889 12483 13923
rect 14841 13889 14875 13923
rect 14933 13889 14967 13923
rect 15577 13889 15611 13923
rect 17785 13889 17819 13923
rect 20361 13889 20395 13923
rect 23397 13889 23431 13923
rect 23664 13889 23698 13923
rect 25881 13889 25915 13923
rect 27537 13889 27571 13923
rect 27813 13889 27847 13923
rect 29285 13889 29319 13923
rect 29377 13889 29411 13923
rect 31401 13889 31435 13923
rect 32597 13889 32631 13923
rect 32853 13889 32887 13923
rect 35081 13889 35115 13923
rect 47869 13889 47903 13923
rect 8309 13821 8343 13855
rect 8585 13821 8619 13855
rect 12909 13821 12943 13855
rect 15117 13821 15151 13855
rect 17969 13821 18003 13855
rect 19441 13821 19475 13855
rect 25973 13821 26007 13855
rect 27721 13821 27755 13855
rect 29469 13821 29503 13855
rect 28917 13753 28951 13787
rect 2145 13685 2179 13719
rect 2881 13685 2915 13719
rect 15025 13685 15059 13719
rect 24777 13685 24811 13719
rect 27537 13685 27571 13719
rect 27997 13685 28031 13719
rect 36461 13685 36495 13719
rect 8309 13481 8343 13515
rect 16037 13481 16071 13515
rect 26893 13481 26927 13515
rect 28825 13481 28859 13515
rect 33793 13481 33827 13515
rect 36553 13481 36587 13515
rect 30849 13413 30883 13447
rect 1409 13345 1443 13379
rect 1593 13345 1627 13379
rect 2789 13345 2823 13379
rect 14657 13345 14691 13379
rect 19901 13345 19935 13379
rect 26157 13345 26191 13379
rect 26985 13345 27019 13379
rect 29837 13345 29871 13379
rect 32413 13345 32447 13379
rect 8217 13277 8251 13311
rect 18153 13277 18187 13311
rect 18245 13277 18279 13311
rect 18337 13277 18371 13311
rect 18521 13277 18555 13311
rect 19717 13277 19751 13311
rect 20361 13277 20395 13311
rect 22477 13277 22511 13311
rect 25237 13277 25271 13311
rect 25973 13277 26007 13311
rect 26709 13277 26743 13311
rect 26801 13277 26835 13311
rect 27997 13277 28031 13311
rect 29561 13277 29595 13311
rect 29745 13277 29779 13311
rect 29929 13277 29963 13311
rect 30113 13277 30147 13311
rect 30757 13277 30791 13311
rect 30941 13277 30975 13311
rect 31769 13277 31803 13311
rect 32669 13277 32703 13311
rect 35357 13277 35391 13311
rect 35446 13277 35480 13311
rect 35541 13277 35575 13311
rect 35725 13277 35759 13311
rect 36369 13277 36403 13311
rect 14924 13209 14958 13243
rect 17233 13209 17267 13243
rect 17417 13209 17451 13243
rect 22744 13209 22778 13243
rect 28733 13209 28767 13243
rect 36185 13209 36219 13243
rect 17877 13141 17911 13175
rect 20453 13141 20487 13175
rect 23857 13141 23891 13175
rect 25329 13141 25363 13175
rect 28089 13141 28123 13175
rect 30297 13141 30331 13175
rect 31861 13141 31895 13175
rect 35081 13141 35115 13175
rect 19993 12937 20027 12971
rect 23673 12937 23707 12971
rect 29285 12937 29319 12971
rect 16948 12869 16982 12903
rect 19901 12869 19935 12903
rect 20729 12869 20763 12903
rect 35234 12869 35268 12903
rect 1685 12801 1719 12835
rect 14105 12801 14139 12835
rect 16681 12801 16715 12835
rect 18521 12801 18555 12835
rect 24501 12801 24535 12835
rect 24685 12801 24719 12835
rect 24777 12801 24811 12835
rect 25053 12801 25087 12835
rect 25237 12801 25271 12835
rect 27813 12801 27847 12835
rect 29377 12801 29411 12835
rect 32413 12801 32447 12835
rect 34989 12801 35023 12835
rect 1409 12733 1443 12767
rect 14289 12733 14323 12767
rect 14565 12733 14599 12767
rect 18797 12733 18831 12767
rect 23765 12733 23799 12767
rect 23949 12733 23983 12767
rect 24869 12733 24903 12767
rect 29469 12733 29503 12767
rect 32137 12733 32171 12767
rect 18061 12597 18095 12631
rect 20821 12597 20855 12631
rect 23305 12597 23339 12631
rect 27905 12597 27939 12631
rect 28917 12597 28951 12631
rect 36369 12597 36403 12631
rect 14289 12393 14323 12427
rect 18705 12393 18739 12427
rect 23581 12393 23615 12427
rect 26893 12393 26927 12427
rect 31309 12393 31343 12427
rect 35357 12393 35391 12427
rect 16037 12257 16071 12291
rect 20269 12257 20303 12291
rect 27721 12257 27755 12291
rect 29929 12257 29963 12291
rect 14197 12189 14231 12223
rect 15393 12189 15427 12223
rect 18521 12189 18555 12223
rect 19441 12189 19475 12223
rect 20085 12189 20119 12223
rect 23489 12189 23523 12223
rect 23673 12189 23707 12223
rect 26709 12189 26743 12223
rect 27445 12189 27479 12223
rect 29009 12189 29043 12223
rect 30196 12189 30230 12223
rect 34989 12189 35023 12223
rect 35173 12189 35207 12223
rect 15485 12121 15519 12155
rect 16221 12121 16255 12155
rect 17877 12121 17911 12155
rect 18337 12121 18371 12155
rect 19257 12121 19291 12155
rect 21925 12121 21959 12155
rect 28825 12121 28859 12155
rect 19625 12053 19659 12087
rect 19901 11849 19935 11883
rect 27077 11781 27111 11815
rect 17785 11713 17819 11747
rect 18788 11713 18822 11747
rect 20545 11713 20579 11747
rect 21833 11713 21867 11747
rect 25789 11713 25823 11747
rect 25973 11713 26007 11747
rect 26065 11713 26099 11747
rect 27721 11713 27755 11747
rect 28457 11713 28491 11747
rect 28641 11713 28675 11747
rect 29469 11713 29503 11747
rect 18521 11645 18555 11679
rect 20361 11645 20395 11679
rect 22109 11645 22143 11679
rect 29561 11645 29595 11679
rect 29653 11645 29687 11679
rect 28549 11577 28583 11611
rect 17969 11509 18003 11543
rect 20729 11509 20763 11543
rect 25605 11509 25639 11543
rect 27169 11509 27203 11543
rect 27905 11509 27939 11543
rect 29101 11509 29135 11543
rect 18429 11305 18463 11339
rect 19257 11305 19291 11339
rect 26617 11305 26651 11339
rect 27537 11305 27571 11339
rect 31861 11305 31895 11339
rect 28273 11237 28307 11271
rect 29837 11237 29871 11271
rect 2053 11169 2087 11203
rect 24501 11169 24535 11203
rect 28825 11169 28859 11203
rect 2513 11101 2547 11135
rect 18337 11101 18371 11135
rect 19533 11101 19567 11135
rect 19622 11101 19656 11135
rect 19717 11101 19751 11135
rect 19901 11101 19935 11135
rect 20637 11101 20671 11135
rect 20729 11101 20763 11135
rect 20913 11101 20947 11135
rect 21005 11101 21039 11135
rect 21833 11101 21867 11135
rect 23213 11101 23247 11135
rect 23361 11101 23395 11135
rect 23489 11101 23523 11135
rect 23719 11101 23753 11135
rect 24409 11101 24443 11135
rect 24593 11101 24627 11135
rect 25237 11101 25271 11135
rect 25504 11101 25538 11135
rect 27813 11101 27847 11135
rect 30021 11101 30055 11135
rect 30481 11101 30515 11135
rect 30737 11101 30771 11135
rect 32689 11101 32723 11135
rect 33517 11101 33551 11135
rect 47225 11101 47259 11135
rect 48053 11101 48087 11135
rect 1869 11033 1903 11067
rect 2605 11033 2639 11067
rect 22017 11033 22051 11067
rect 23581 11033 23615 11067
rect 27537 11033 27571 11067
rect 28641 11033 28675 11067
rect 32873 11033 32907 11067
rect 20453 10965 20487 10999
rect 22201 10965 22235 10999
rect 23857 10965 23891 10999
rect 27721 10965 27755 10999
rect 28733 10965 28767 10999
rect 33057 10965 33091 10999
rect 33609 10965 33643 10999
rect 47317 10965 47351 10999
rect 26433 10761 26467 10795
rect 27997 10761 28031 10795
rect 19892 10693 19926 10727
rect 29009 10693 29043 10727
rect 2145 10625 2179 10659
rect 18613 10625 18647 10659
rect 18705 10625 18739 10659
rect 18797 10625 18831 10659
rect 18981 10625 19015 10659
rect 19625 10625 19659 10659
rect 22109 10625 22143 10659
rect 22201 10625 22235 10659
rect 22293 10625 22327 10659
rect 22477 10625 22511 10659
rect 23029 10625 23063 10659
rect 23296 10625 23330 10659
rect 24869 10625 24903 10659
rect 25053 10625 25087 10659
rect 25697 10625 25731 10659
rect 25881 10625 25915 10659
rect 26065 10625 26099 10659
rect 26249 10625 26283 10659
rect 26985 10625 27019 10659
rect 27169 10625 27203 10659
rect 27629 10625 27663 10659
rect 32393 10625 32427 10659
rect 32502 10625 32536 10659
rect 32597 10631 32631 10665
rect 32781 10625 32815 10659
rect 33609 10625 33643 10659
rect 35449 10625 35483 10659
rect 47777 10625 47811 10659
rect 25237 10557 25271 10591
rect 25973 10557 26007 10591
rect 27721 10557 27755 10591
rect 33793 10557 33827 10591
rect 21005 10489 21039 10523
rect 27077 10489 27111 10523
rect 29193 10489 29227 10523
rect 47961 10489 47995 10523
rect 1685 10421 1719 10455
rect 2237 10421 2271 10455
rect 2973 10421 3007 10455
rect 18337 10421 18371 10455
rect 21833 10421 21867 10455
rect 24409 10421 24443 10455
rect 27813 10421 27847 10455
rect 32137 10421 32171 10455
rect 19625 10217 19659 10251
rect 22385 10217 22419 10251
rect 26065 10217 26099 10251
rect 27813 10217 27847 10251
rect 28917 10217 28951 10251
rect 33793 10217 33827 10251
rect 1409 10081 1443 10115
rect 1593 10081 1627 10115
rect 2789 10081 2823 10115
rect 17049 10081 17083 10115
rect 21005 10081 21039 10115
rect 23581 10081 23615 10115
rect 23765 10081 23799 10115
rect 25237 10081 25271 10115
rect 28273 10081 28307 10115
rect 28641 10081 28675 10115
rect 30113 10081 30147 10115
rect 46305 10081 46339 10115
rect 46489 10081 46523 10115
rect 48145 10081 48179 10115
rect 17316 10013 17350 10047
rect 20361 10013 20395 10047
rect 21272 10013 21306 10047
rect 25053 10013 25087 10047
rect 25973 10013 26007 10047
rect 27445 10013 27479 10047
rect 28733 10013 28767 10047
rect 29929 10013 29963 10047
rect 32413 10013 32447 10047
rect 32669 10013 32703 10047
rect 19257 9945 19291 9979
rect 19441 9945 19475 9979
rect 20545 9945 20579 9979
rect 23489 9945 23523 9979
rect 26801 9945 26835 9979
rect 26985 9945 27019 9979
rect 27629 9945 27663 9979
rect 18429 9877 18463 9911
rect 23121 9877 23155 9911
rect 24685 9877 24719 9911
rect 25145 9877 25179 9911
rect 29561 9877 29595 9911
rect 30021 9877 30055 9911
rect 24869 9673 24903 9707
rect 24225 9605 24259 9639
rect 25329 9605 25363 9639
rect 31493 9605 31527 9639
rect 32781 9605 32815 9639
rect 1777 9537 1811 9571
rect 17601 9537 17635 9571
rect 23213 9537 23247 9571
rect 24501 9537 24535 9571
rect 24685 9537 24719 9571
rect 25605 9537 25639 9571
rect 27813 9537 27847 9571
rect 27997 9537 28031 9571
rect 28089 9537 28123 9571
rect 29101 9537 29135 9571
rect 29193 9537 29227 9571
rect 29929 9537 29963 9571
rect 30113 9537 30147 9571
rect 30297 9537 30331 9571
rect 30481 9537 30515 9571
rect 31401 9537 31435 9571
rect 1961 9469 1995 9503
rect 2789 9469 2823 9503
rect 17785 9469 17819 9503
rect 18245 9469 18279 9503
rect 23305 9469 23339 9503
rect 23581 9469 23615 9503
rect 25421 9469 25455 9503
rect 29377 9469 29411 9503
rect 30205 9469 30239 9503
rect 32597 9469 32631 9503
rect 33149 9469 33183 9503
rect 24409 9333 24443 9367
rect 25329 9333 25363 9367
rect 25789 9333 25823 9367
rect 27813 9333 27847 9367
rect 28733 9333 28767 9367
rect 30665 9333 30699 9367
rect 18061 9129 18095 9163
rect 23857 9129 23891 9163
rect 27905 9129 27939 9163
rect 28089 9129 28123 9163
rect 31401 9129 31435 9163
rect 27077 9061 27111 9095
rect 48145 9061 48179 9095
rect 24869 8993 24903 9027
rect 27813 8993 27847 9027
rect 17969 8925 18003 8959
rect 24593 8925 24627 8959
rect 24777 8925 24811 8959
rect 26985 8925 27019 8959
rect 27169 8925 27203 8959
rect 27629 8925 27663 8959
rect 27905 8925 27939 8959
rect 28549 8925 28583 8959
rect 30021 8925 30055 8959
rect 30288 8925 30322 8959
rect 32459 8925 32493 8959
rect 32597 8925 32631 8959
rect 32694 8925 32728 8959
rect 32873 8925 32907 8959
rect 33333 8925 33367 8959
rect 33425 8925 33459 8959
rect 46765 8925 46799 8959
rect 23489 8857 23523 8891
rect 23673 8857 23707 8891
rect 28733 8857 28767 8891
rect 47961 8857 47995 8891
rect 24409 8789 24443 8823
rect 28917 8789 28951 8823
rect 32229 8789 32263 8823
rect 46857 8789 46891 8823
rect 23581 8585 23615 8619
rect 28549 8585 28583 8619
rect 29561 8585 29595 8619
rect 18245 8517 18279 8551
rect 19594 8517 19628 8551
rect 23397 8517 23431 8551
rect 29101 8517 29135 8551
rect 32658 8517 32692 8551
rect 1869 8449 1903 8483
rect 18521 8449 18555 8483
rect 18610 8452 18644 8486
rect 18705 8449 18739 8483
rect 18889 8449 18923 8483
rect 19349 8449 19383 8483
rect 23673 8449 23707 8483
rect 24133 8449 24167 8483
rect 24317 8449 24351 8483
rect 27445 8449 27479 8483
rect 28181 8449 28215 8483
rect 29377 8449 29411 8483
rect 32413 8449 32447 8483
rect 47869 8449 47903 8483
rect 27721 8381 27755 8415
rect 28273 8381 28307 8415
rect 29285 8381 29319 8415
rect 2145 8313 2179 8347
rect 20729 8313 20763 8347
rect 23397 8313 23431 8347
rect 27261 8313 27295 8347
rect 48053 8313 48087 8347
rect 24225 8245 24259 8279
rect 27629 8245 27663 8279
rect 28181 8245 28215 8279
rect 29101 8245 29135 8279
rect 33793 8245 33827 8279
rect 47041 8245 47075 8279
rect 19625 8041 19659 8075
rect 28089 8041 28123 8075
rect 33425 8041 33459 8075
rect 2145 7905 2179 7939
rect 17601 7905 17635 7939
rect 20821 7905 20855 7939
rect 23581 7905 23615 7939
rect 23765 7905 23799 7939
rect 24685 7905 24719 7939
rect 25697 7905 25731 7939
rect 28273 7905 28307 7939
rect 31217 7905 31251 7939
rect 46305 7905 46339 7939
rect 17233 7837 17267 7871
rect 18337 7837 18371 7871
rect 18442 7831 18476 7865
rect 18542 7834 18576 7868
rect 18705 7837 18739 7871
rect 19257 7837 19291 7871
rect 19441 7837 19475 7871
rect 24409 7837 24443 7871
rect 24593 7837 24627 7871
rect 24777 7837 24811 7871
rect 24961 7837 24995 7871
rect 27997 7837 28031 7871
rect 33241 7837 33275 7871
rect 1869 7769 1903 7803
rect 17417 7769 17451 7803
rect 21005 7769 21039 7803
rect 22661 7769 22695 7803
rect 23489 7769 23523 7803
rect 25881 7769 25915 7803
rect 27537 7769 27571 7803
rect 31462 7769 31496 7803
rect 33057 7769 33091 7803
rect 46489 7769 46523 7803
rect 48145 7769 48179 7803
rect 18061 7701 18095 7735
rect 23121 7701 23155 7735
rect 25145 7701 25179 7735
rect 28549 7701 28583 7735
rect 32597 7701 32631 7735
rect 18521 7497 18555 7531
rect 21005 7497 21039 7531
rect 24869 7497 24903 7531
rect 28181 7497 28215 7531
rect 30941 7497 30975 7531
rect 20269 7429 20303 7463
rect 23756 7429 23790 7463
rect 33057 7429 33091 7463
rect 17141 7361 17175 7395
rect 17408 7361 17442 7395
rect 20085 7361 20119 7395
rect 20913 7361 20947 7395
rect 23489 7361 23523 7395
rect 26065 7361 26099 7395
rect 27353 7361 27387 7395
rect 28549 7361 28583 7395
rect 28641 7361 28675 7395
rect 29377 7361 29411 7395
rect 29561 7361 29595 7395
rect 29745 7361 29779 7395
rect 29929 7361 29963 7395
rect 31197 7361 31231 7395
rect 31309 7361 31343 7395
rect 31401 7361 31435 7395
rect 31585 7361 31619 7395
rect 32137 7361 32171 7395
rect 26157 7293 26191 7327
rect 27445 7293 27479 7327
rect 27537 7293 27571 7327
rect 28733 7293 28767 7327
rect 29653 7293 29687 7327
rect 32873 7293 32907 7327
rect 33333 7293 33367 7327
rect 26433 7225 26467 7259
rect 2053 7157 2087 7191
rect 20453 7157 20487 7191
rect 26985 7157 27019 7191
rect 30113 7157 30147 7191
rect 32229 7157 32263 7191
rect 1409 6817 1443 6851
rect 2789 6817 2823 6851
rect 20269 6817 20303 6851
rect 27261 6817 27295 6851
rect 31861 6817 31895 6851
rect 32137 6817 32171 6851
rect 18337 6749 18371 6783
rect 26249 6749 26283 6783
rect 26433 6749 26467 6783
rect 26893 6749 26927 6783
rect 27077 6749 27111 6783
rect 27169 6749 27203 6783
rect 27445 6749 27479 6783
rect 29561 6749 29595 6783
rect 29828 6749 29862 6783
rect 31677 6749 31711 6783
rect 1593 6681 1627 6715
rect 20536 6681 20570 6715
rect 22661 6681 22695 6715
rect 22845 6681 22879 6715
rect 26065 6681 26099 6715
rect 18429 6613 18463 6647
rect 21649 6613 21683 6647
rect 23029 6613 23063 6647
rect 27629 6613 27663 6647
rect 30941 6613 30975 6647
rect 2237 6409 2271 6443
rect 28825 6409 28859 6443
rect 18337 6341 18371 6375
rect 22201 6341 22235 6375
rect 32137 6341 32171 6375
rect 32505 6341 32539 6375
rect 2145 6273 2179 6307
rect 18153 6273 18187 6307
rect 20729 6273 20763 6307
rect 20821 6273 20855 6307
rect 20913 6273 20947 6307
rect 21097 6273 21131 6307
rect 21833 6273 21867 6307
rect 22017 6273 22051 6307
rect 23029 6273 23063 6307
rect 23121 6273 23155 6307
rect 23213 6273 23247 6307
rect 23397 6273 23431 6307
rect 27445 6273 27479 6307
rect 27712 6273 27746 6307
rect 32321 6273 32355 6307
rect 19533 6205 19567 6239
rect 20453 6069 20487 6103
rect 22753 6069 22787 6103
rect 21649 5797 21683 5831
rect 20269 5729 20303 5763
rect 2145 5661 2179 5695
rect 2973 5661 3007 5695
rect 3801 5661 3835 5695
rect 19257 5661 19291 5695
rect 20536 5661 20570 5695
rect 22477 5661 22511 5695
rect 47869 5661 47903 5695
rect 22722 5593 22756 5627
rect 2237 5525 2271 5559
rect 3893 5525 3927 5559
rect 19349 5525 19383 5559
rect 23857 5525 23891 5559
rect 48053 5525 48087 5559
rect 20637 5321 20671 5355
rect 22109 5321 22143 5355
rect 24777 5321 24811 5355
rect 2329 5253 2363 5287
rect 18521 5253 18555 5287
rect 20177 5253 20211 5287
rect 2145 5185 2179 5219
rect 20913 5185 20947 5219
rect 21005 5185 21039 5219
rect 21097 5185 21131 5219
rect 21281 5185 21315 5219
rect 22339 5185 22373 5219
rect 22477 5185 22511 5219
rect 22569 5185 22603 5219
rect 22753 5185 22787 5219
rect 23397 5185 23431 5219
rect 23664 5185 23698 5219
rect 47593 5185 47627 5219
rect 2789 5117 2823 5151
rect 18337 5117 18371 5151
rect 1685 4981 1719 5015
rect 47041 4981 47075 5015
rect 47685 4981 47719 5015
rect 22293 4777 22327 4811
rect 1409 4641 1443 4675
rect 1593 4641 1627 4675
rect 2789 4641 2823 4675
rect 46305 4641 46339 4675
rect 46489 4641 46523 4675
rect 48145 4641 48179 4675
rect 4629 4573 4663 4607
rect 11713 4573 11747 4607
rect 12357 4573 12391 4607
rect 18521 4573 18555 4607
rect 21925 4573 21959 4607
rect 22109 4573 22143 4607
rect 31493 4573 31527 4607
rect 39865 4573 39899 4607
rect 11805 4437 11839 4471
rect 12449 4437 12483 4471
rect 18613 4437 18647 4471
rect 39957 4437 39991 4471
rect 40509 4437 40543 4471
rect 11713 4165 11747 4199
rect 47961 4165 47995 4199
rect 4169 4097 4203 4131
rect 4813 4097 4847 4131
rect 11529 4097 11563 4131
rect 13829 4097 13863 4131
rect 15209 4097 15243 4131
rect 19993 4097 20027 4131
rect 23305 4097 23339 4131
rect 26065 4097 26099 4131
rect 30941 4097 30975 4131
rect 32137 4097 32171 4131
rect 36185 4097 36219 4131
rect 37841 4097 37875 4131
rect 37933 4097 37967 4131
rect 40509 4097 40543 4131
rect 41337 4097 41371 4131
rect 46857 4097 46891 4131
rect 9137 4029 9171 4063
rect 9321 4029 9355 4063
rect 9597 4029 9631 4063
rect 12541 4029 12575 4063
rect 38669 4029 38703 4063
rect 38853 4029 38887 4063
rect 48145 3961 48179 3995
rect 2053 3893 2087 3927
rect 3617 3893 3651 3927
rect 4261 3893 4295 3927
rect 4905 3893 4939 3927
rect 6653 3893 6687 3927
rect 13921 3893 13955 3927
rect 15301 3893 15335 3927
rect 18245 3893 18279 3927
rect 20085 3893 20119 3927
rect 20913 3893 20947 3927
rect 23397 3893 23431 3927
rect 26157 3893 26191 3927
rect 30021 3893 30055 3927
rect 31033 3893 31067 3927
rect 32229 3893 32263 3927
rect 32965 3893 32999 3927
rect 36277 3893 36311 3927
rect 41429 3893 41463 3927
rect 42625 3893 42659 3927
rect 44281 3893 44315 3927
rect 44925 3893 44959 3927
rect 46949 3893 46983 3927
rect 9321 3689 9355 3723
rect 38853 3689 38887 3723
rect 1409 3553 1443 3587
rect 1869 3553 1903 3587
rect 3801 3553 3835 3587
rect 3985 3553 4019 3587
rect 4261 3553 4295 3587
rect 11805 3553 11839 3587
rect 12541 3553 12575 3587
rect 15117 3553 15151 3587
rect 15485 3553 15519 3587
rect 20269 3553 20303 3587
rect 20637 3553 20671 3587
rect 25973 3553 26007 3587
rect 26433 3553 26467 3587
rect 31677 3553 31711 3587
rect 36461 3553 36495 3587
rect 36737 3553 36771 3587
rect 41613 3553 41647 3587
rect 41889 3553 41923 3587
rect 46489 3553 46523 3587
rect 6101 3485 6135 3519
rect 6929 3485 6963 3519
rect 7481 3485 7515 3519
rect 9229 3485 9263 3519
rect 11161 3485 11195 3519
rect 11621 3485 11655 3519
rect 14105 3485 14139 3519
rect 14933 3485 14967 3519
rect 20085 3485 20119 3519
rect 23673 3485 23707 3519
rect 25789 3485 25823 3519
rect 29009 3485 29043 3519
rect 29553 3485 29587 3519
rect 30205 3485 30239 3519
rect 31217 3485 31251 3519
rect 36277 3485 36311 3519
rect 39865 3485 39899 3519
rect 40969 3485 41003 3519
rect 41429 3485 41463 3519
rect 43913 3485 43947 3519
rect 45017 3485 45051 3519
rect 45845 3485 45879 3519
rect 46305 3485 46339 3519
rect 1593 3417 1627 3451
rect 29653 3417 29687 3451
rect 31401 3417 31435 3451
rect 48145 3417 48179 3451
rect 6193 3349 6227 3383
rect 7573 3349 7607 3383
rect 14197 3349 14231 3383
rect 30297 3349 30331 3383
rect 39957 3349 39991 3383
rect 44005 3349 44039 3383
rect 45109 3349 45143 3383
rect 2145 3145 2179 3179
rect 22845 3145 22879 3179
rect 26985 3145 27019 3179
rect 46489 3145 46523 3179
rect 48053 3145 48087 3179
rect 4169 3077 4203 3111
rect 6561 3077 6595 3111
rect 10241 3077 10275 3111
rect 18153 3077 18187 3111
rect 23581 3077 23615 3111
rect 29929 3077 29963 3111
rect 32413 3077 32447 3111
rect 40233 3077 40267 3111
rect 44189 3077 44223 3111
rect 2053 3009 2087 3043
rect 6377 3009 6411 3043
rect 8953 3009 8987 3043
rect 10057 3009 10091 3043
rect 12265 3009 12299 3043
rect 14565 3009 14599 3043
rect 15485 3009 15519 3043
rect 17969 3009 18003 3043
rect 20453 3009 20487 3043
rect 20913 3009 20947 3043
rect 22753 3009 22787 3043
rect 23397 3009 23431 3043
rect 26065 3009 26099 3043
rect 27169 3009 27203 3043
rect 29745 3009 29779 3043
rect 36553 3009 36587 3043
rect 42441 3009 42475 3043
rect 43269 3009 43303 3043
rect 44005 3009 44039 3043
rect 46305 3009 46339 3043
rect 47869 3009 47903 3043
rect 3985 2941 4019 2975
rect 5181 2941 5215 2975
rect 6837 2941 6871 2975
rect 8677 2941 8711 2975
rect 12449 2941 12483 2975
rect 12909 2941 12943 2975
rect 18429 2941 18463 2975
rect 23857 2941 23891 2975
rect 30297 2941 30331 2975
rect 32229 2941 32263 2975
rect 33425 2941 33459 2975
rect 40049 2941 40083 2975
rect 41245 2941 41279 2975
rect 44465 2941 44499 2975
rect 14749 2873 14783 2907
rect 43453 2873 43487 2907
rect 21005 2805 21039 2839
rect 39589 2805 39623 2839
rect 42533 2805 42567 2839
rect 12449 2601 12483 2635
rect 2973 2533 3007 2567
rect 4813 2533 4847 2567
rect 10425 2533 10459 2567
rect 20361 2533 20395 2567
rect 27353 2533 27387 2567
rect 28181 2533 28215 2567
rect 34161 2533 34195 2567
rect 6469 2465 6503 2499
rect 6653 2465 6687 2499
rect 7021 2465 7055 2499
rect 8953 2465 8987 2499
rect 14565 2465 14599 2499
rect 21833 2465 21867 2499
rect 22017 2465 22051 2499
rect 22293 2465 22327 2499
rect 26249 2465 26283 2499
rect 29561 2465 29595 2499
rect 29745 2465 29779 2499
rect 30941 2465 30975 2499
rect 35357 2465 35391 2499
rect 39865 2465 39899 2499
rect 40049 2465 40083 2499
rect 40325 2465 40359 2499
rect 42441 2465 42475 2499
rect 42625 2465 42659 2499
rect 42901 2465 42935 2499
rect 45017 2465 45051 2499
rect 45201 2465 45235 2499
rect 45569 2465 45603 2499
rect 2789 2397 2823 2431
rect 4629 2397 4663 2431
rect 10241 2397 10275 2431
rect 13093 2397 13127 2431
rect 14105 2397 14139 2431
rect 17509 2397 17543 2431
rect 25513 2397 25547 2431
rect 27169 2397 27203 2431
rect 32965 2397 32999 2431
rect 36461 2397 36495 2431
rect 38485 2397 38519 2431
rect 38761 2397 38795 2431
rect 1869 2329 1903 2363
rect 2237 2329 2271 2363
rect 14289 2329 14323 2363
rect 20177 2329 20211 2363
rect 25329 2329 25363 2363
rect 26065 2329 26099 2363
rect 27997 2329 28031 2363
rect 33977 2329 34011 2363
rect 35173 2329 35207 2363
rect 36277 2329 36311 2363
rect 47777 2329 47811 2363
rect 9183 2261 9217 2295
rect 17693 2261 17727 2295
rect 33149 2261 33183 2295
rect 47869 2261 47903 2295
<< metal1 >>
rect 41414 50192 41420 50244
rect 41472 50232 41478 50244
rect 46842 50232 46848 50244
rect 41472 50204 46848 50232
rect 41472 50192 41478 50204
rect 46842 50192 46848 50204
rect 46900 50192 46906 50244
rect 3418 49716 3424 49768
rect 3476 49756 3482 49768
rect 9214 49756 9220 49768
rect 3476 49728 9220 49756
rect 3476 49716 3482 49728
rect 9214 49716 9220 49728
rect 9272 49716 9278 49768
rect 21266 49716 21272 49768
rect 21324 49756 21330 49768
rect 46750 49756 46756 49768
rect 21324 49728 46756 49756
rect 21324 49716 21330 49728
rect 46750 49716 46756 49728
rect 46808 49716 46814 49768
rect 1104 49530 48852 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 48852 49530
rect 1104 49456 48852 49478
rect 23842 49348 23848 49360
rect 21284 49320 23848 49348
rect 3789 49283 3847 49289
rect 3789 49249 3801 49283
rect 3835 49280 3847 49283
rect 3970 49280 3976 49292
rect 3835 49252 3976 49280
rect 3835 49249 3847 49252
rect 3789 49243 3847 49249
rect 3970 49240 3976 49252
rect 4028 49240 4034 49292
rect 4062 49240 4068 49292
rect 4120 49280 4126 49292
rect 4249 49283 4307 49289
rect 4249 49280 4261 49283
rect 4120 49252 4261 49280
rect 4120 49240 4126 49252
rect 4249 49249 4261 49252
rect 4295 49249 4307 49283
rect 4249 49243 4307 49249
rect 8662 49240 8668 49292
rect 8720 49280 8726 49292
rect 10505 49283 10563 49289
rect 10505 49280 10517 49283
rect 8720 49252 10517 49280
rect 8720 49240 8726 49252
rect 10505 49249 10517 49252
rect 10551 49249 10563 49283
rect 12710 49280 12716 49292
rect 12671 49252 12716 49280
rect 10505 49243 10563 49249
rect 12710 49240 12716 49252
rect 12768 49240 12774 49292
rect 13814 49240 13820 49292
rect 13872 49280 13878 49292
rect 14093 49283 14151 49289
rect 14093 49280 14105 49283
rect 13872 49252 14105 49280
rect 13872 49240 13878 49252
rect 14093 49249 14105 49252
rect 14139 49249 14151 49283
rect 14093 49243 14151 49249
rect 17865 49283 17923 49289
rect 17865 49249 17877 49283
rect 17911 49280 17923 49283
rect 18046 49280 18052 49292
rect 17911 49252 18052 49280
rect 17911 49249 17923 49252
rect 17865 49243 17923 49249
rect 18046 49240 18052 49252
rect 18104 49240 18110 49292
rect 18141 49283 18199 49289
rect 18141 49249 18153 49283
rect 18187 49280 18199 49283
rect 20438 49280 20444 49292
rect 18187 49252 20444 49280
rect 18187 49249 18199 49252
rect 18141 49243 18199 49249
rect 20438 49240 20444 49252
rect 20496 49240 20502 49292
rect 658 49172 664 49224
rect 716 49212 722 49224
rect 1857 49215 1915 49221
rect 1857 49212 1869 49215
rect 716 49184 1869 49212
rect 716 49172 722 49184
rect 1857 49181 1869 49184
rect 1903 49181 1915 49215
rect 1857 49175 1915 49181
rect 2869 49215 2927 49221
rect 2869 49181 2881 49215
rect 2915 49212 2927 49215
rect 3234 49212 3240 49224
rect 2915 49184 3240 49212
rect 2915 49181 2927 49184
rect 2869 49175 2927 49181
rect 3234 49172 3240 49184
rect 3292 49172 3298 49224
rect 6454 49172 6460 49224
rect 6512 49212 6518 49224
rect 6825 49215 6883 49221
rect 6825 49212 6837 49215
rect 6512 49184 6837 49212
rect 6512 49172 6518 49184
rect 6825 49181 6837 49184
rect 6871 49181 6883 49215
rect 6825 49175 6883 49181
rect 7837 49215 7895 49221
rect 7837 49181 7849 49215
rect 7883 49181 7895 49215
rect 9858 49212 9864 49224
rect 9819 49184 9864 49212
rect 7837 49175 7895 49181
rect 3973 49147 4031 49153
rect 3973 49113 3985 49147
rect 4019 49144 4031 49147
rect 5442 49144 5448 49156
rect 4019 49116 5448 49144
rect 4019 49113 4031 49116
rect 3973 49107 4031 49113
rect 5442 49104 5448 49116
rect 5500 49104 5506 49156
rect 6638 49104 6644 49156
rect 6696 49144 6702 49156
rect 7852 49144 7880 49175
rect 9858 49172 9864 49184
rect 9916 49172 9922 49224
rect 11606 49172 11612 49224
rect 11664 49212 11670 49224
rect 11977 49215 12035 49221
rect 11977 49212 11989 49215
rect 11664 49184 11989 49212
rect 11664 49172 11670 49184
rect 11977 49181 11989 49184
rect 12023 49181 12035 49215
rect 12986 49212 12992 49224
rect 12947 49184 12992 49212
rect 11977 49175 12035 49181
rect 12986 49172 12992 49184
rect 13044 49172 13050 49224
rect 14366 49212 14372 49224
rect 14327 49184 14372 49212
rect 14366 49172 14372 49184
rect 14424 49172 14430 49224
rect 16117 49215 16175 49221
rect 16117 49181 16129 49215
rect 16163 49212 16175 49215
rect 16574 49212 16580 49224
rect 16163 49184 16580 49212
rect 16163 49181 16175 49184
rect 16117 49175 16175 49181
rect 16574 49172 16580 49184
rect 16632 49172 16638 49224
rect 16666 49172 16672 49224
rect 16724 49212 16730 49224
rect 16853 49215 16911 49221
rect 16853 49212 16865 49215
rect 16724 49184 16865 49212
rect 16724 49172 16730 49184
rect 16853 49181 16865 49184
rect 16899 49181 16911 49215
rect 19334 49212 19340 49224
rect 19295 49184 19340 49212
rect 16853 49175 16911 49181
rect 19334 49172 19340 49184
rect 19392 49172 19398 49224
rect 19978 49172 19984 49224
rect 20036 49212 20042 49224
rect 21284 49221 21312 49320
rect 23842 49308 23848 49320
rect 23900 49308 23906 49360
rect 40034 49308 40040 49360
rect 40092 49348 40098 49360
rect 40092 49320 40724 49348
rect 40092 49308 40098 49320
rect 22554 49280 22560 49292
rect 22515 49252 22560 49280
rect 22554 49240 22560 49252
rect 22612 49240 22618 49292
rect 24762 49240 24768 49292
rect 24820 49280 24826 49292
rect 24857 49283 24915 49289
rect 24857 49280 24869 49283
rect 24820 49252 24869 49280
rect 24820 49240 24826 49252
rect 24857 49249 24869 49252
rect 24903 49249 24915 49283
rect 27614 49280 27620 49292
rect 27575 49252 27620 49280
rect 24857 49243 24915 49249
rect 27614 49240 27620 49252
rect 27672 49240 27678 49292
rect 29733 49283 29791 49289
rect 29733 49249 29745 49283
rect 29779 49280 29791 49283
rect 30558 49280 30564 49292
rect 29779 49252 30564 49280
rect 29779 49249 29791 49252
rect 29733 49243 29791 49249
rect 30558 49240 30564 49252
rect 30616 49240 30622 49292
rect 30926 49280 30932 49292
rect 30887 49252 30932 49280
rect 30926 49240 30932 49252
rect 30984 49240 30990 49292
rect 40586 49280 40592 49292
rect 39040 49252 40592 49280
rect 20073 49215 20131 49221
rect 20073 49212 20085 49215
rect 20036 49184 20085 49212
rect 20036 49172 20042 49184
rect 20073 49181 20085 49184
rect 20119 49181 20131 49215
rect 20073 49175 20131 49181
rect 21269 49215 21327 49221
rect 21269 49181 21281 49215
rect 21315 49181 21327 49215
rect 22002 49212 22008 49224
rect 21963 49184 22008 49212
rect 21269 49175 21327 49181
rect 22002 49172 22008 49184
rect 22060 49172 22066 49224
rect 24394 49212 24400 49224
rect 24355 49184 24400 49212
rect 24394 49172 24400 49184
rect 24452 49172 24458 49224
rect 26970 49212 26976 49224
rect 26931 49184 26976 49212
rect 26970 49172 26976 49184
rect 27028 49172 27034 49224
rect 31938 49172 31944 49224
rect 31996 49212 32002 49224
rect 32953 49215 33011 49221
rect 32953 49212 32965 49215
rect 31996 49184 32965 49212
rect 31996 49172 32002 49184
rect 32953 49181 32965 49184
rect 32999 49181 33011 49215
rect 32953 49175 33011 49181
rect 34882 49172 34888 49224
rect 34940 49212 34946 49224
rect 35897 49215 35955 49221
rect 35897 49212 35909 49215
rect 34940 49184 35909 49212
rect 34940 49172 34946 49184
rect 35897 49181 35909 49184
rect 35943 49181 35955 49215
rect 38102 49212 38108 49224
rect 38063 49184 38108 49212
rect 35897 49175 35955 49181
rect 38102 49172 38108 49184
rect 38160 49172 38166 49224
rect 39040 49221 39068 49252
rect 40586 49240 40592 49252
rect 40644 49240 40650 49292
rect 40696 49289 40724 49320
rect 40681 49283 40739 49289
rect 40681 49249 40693 49283
rect 40727 49249 40739 49283
rect 40681 49243 40739 49249
rect 44453 49283 44511 49289
rect 44453 49249 44465 49283
rect 44499 49280 44511 49283
rect 46658 49280 46664 49292
rect 44499 49252 46664 49280
rect 44499 49249 44511 49252
rect 44453 49243 44511 49249
rect 46658 49240 46664 49252
rect 46716 49240 46722 49292
rect 46842 49280 46848 49292
rect 46803 49252 46848 49280
rect 46842 49240 46848 49252
rect 46900 49240 46906 49292
rect 39025 49215 39083 49221
rect 39025 49181 39037 49215
rect 39071 49181 39083 49215
rect 39025 49175 39083 49181
rect 39758 49172 39764 49224
rect 39816 49212 39822 49224
rect 39853 49215 39911 49221
rect 39853 49212 39865 49215
rect 39816 49184 39865 49212
rect 39816 49172 39822 49184
rect 39853 49181 39865 49184
rect 39899 49181 39911 49215
rect 39853 49175 39911 49181
rect 41966 49172 41972 49224
rect 42024 49212 42030 49224
rect 42613 49215 42671 49221
rect 42613 49212 42625 49215
rect 42024 49184 42625 49212
rect 42024 49172 42030 49184
rect 42613 49181 42625 49184
rect 42659 49181 42671 49215
rect 42613 49175 42671 49181
rect 44082 49172 44088 49224
rect 44140 49212 44146 49224
rect 45189 49215 45247 49221
rect 45189 49212 45201 49215
rect 44140 49184 45201 49212
rect 44140 49172 44146 49184
rect 45189 49181 45201 49184
rect 45235 49181 45247 49215
rect 45189 49175 45247 49181
rect 47765 49215 47823 49221
rect 47765 49181 47777 49215
rect 47811 49212 47823 49215
rect 48958 49212 48964 49224
rect 47811 49184 48964 49212
rect 47811 49181 47823 49184
rect 47765 49175 47823 49181
rect 48958 49172 48964 49184
rect 49016 49172 49022 49224
rect 12158 49144 12164 49156
rect 6696 49116 7880 49144
rect 12119 49116 12164 49144
rect 6696 49104 6702 49116
rect 12158 49104 12164 49116
rect 12216 49104 12222 49156
rect 22186 49144 22192 49156
rect 22147 49116 22192 49144
rect 22186 49104 22192 49116
rect 22244 49104 22250 49156
rect 24578 49144 24584 49156
rect 24539 49116 24584 49144
rect 24578 49104 24584 49116
rect 24636 49104 24642 49156
rect 27154 49144 27160 49156
rect 27115 49116 27160 49144
rect 27154 49104 27160 49116
rect 27212 49104 27218 49156
rect 29914 49144 29920 49156
rect 29875 49116 29920 49144
rect 29914 49104 29920 49116
rect 29972 49104 29978 49156
rect 40034 49144 40040 49156
rect 39995 49116 40040 49144
rect 40034 49104 40040 49116
rect 40092 49104 40098 49156
rect 42797 49147 42855 49153
rect 42797 49113 42809 49147
rect 42843 49144 42855 49147
rect 43714 49144 43720 49156
rect 42843 49116 43720 49144
rect 42843 49113 42855 49116
rect 42797 49107 42855 49113
rect 43714 49104 43720 49116
rect 43772 49104 43778 49156
rect 45370 49144 45376 49156
rect 45331 49116 45376 49144
rect 45370 49104 45376 49116
rect 45428 49104 45434 49156
rect 1670 49036 1676 49088
rect 1728 49076 1734 49088
rect 1949 49079 2007 49085
rect 1949 49076 1961 49079
rect 1728 49048 1961 49076
rect 1728 49036 1734 49048
rect 1949 49045 1961 49048
rect 1995 49045 2007 49079
rect 3142 49076 3148 49088
rect 3103 49048 3148 49076
rect 1949 49039 2007 49045
rect 3142 49036 3148 49048
rect 3200 49036 3206 49088
rect 6914 49036 6920 49088
rect 6972 49076 6978 49088
rect 6972 49048 7017 49076
rect 6972 49036 6978 49048
rect 8938 49036 8944 49088
rect 8996 49076 9002 49088
rect 9033 49079 9091 49085
rect 9033 49076 9045 49079
rect 8996 49048 9045 49076
rect 8996 49036 9002 49048
rect 9033 49045 9045 49048
rect 9079 49045 9091 49079
rect 9033 49039 9091 49045
rect 19521 49079 19579 49085
rect 19521 49045 19533 49079
rect 19567 49076 19579 49079
rect 20162 49076 20168 49088
rect 19567 49048 20168 49076
rect 19567 49045 19579 49048
rect 19521 49039 19579 49045
rect 20162 49036 20168 49048
rect 20220 49036 20226 49088
rect 20257 49079 20315 49085
rect 20257 49045 20269 49079
rect 20303 49076 20315 49079
rect 20346 49076 20352 49088
rect 20303 49048 20352 49076
rect 20303 49045 20315 49048
rect 20257 49039 20315 49045
rect 20346 49036 20352 49048
rect 20404 49036 20410 49088
rect 21085 49079 21143 49085
rect 21085 49045 21097 49079
rect 21131 49076 21143 49079
rect 23474 49076 23480 49088
rect 21131 49048 23480 49076
rect 21131 49045 21143 49048
rect 21085 49039 21143 49045
rect 23474 49036 23480 49048
rect 23532 49036 23538 49088
rect 32122 49076 32128 49088
rect 32083 49048 32128 49076
rect 32122 49036 32128 49048
rect 32180 49036 32186 49088
rect 38286 49076 38292 49088
rect 38247 49048 38292 49076
rect 38286 49036 38292 49048
rect 38344 49036 38350 49088
rect 39206 49076 39212 49088
rect 39167 49048 39212 49076
rect 39206 49036 39212 49048
rect 39264 49036 39270 49088
rect 47946 49036 47952 49088
rect 48004 49076 48010 49088
rect 48041 49079 48099 49085
rect 48041 49076 48053 49079
rect 48004 49048 48053 49076
rect 48004 49036 48010 49048
rect 48041 49045 48053 49048
rect 48087 49045 48099 49079
rect 48041 49039 48099 49045
rect 1104 48986 48852 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 48852 48986
rect 1104 48912 48852 48934
rect 20162 48832 20168 48884
rect 20220 48872 20226 48884
rect 26786 48872 26792 48884
rect 20220 48844 26792 48872
rect 20220 48832 20226 48844
rect 26786 48832 26792 48844
rect 26844 48832 26850 48884
rect 2866 48764 2872 48816
rect 2924 48804 2930 48816
rect 3329 48807 3387 48813
rect 3329 48804 3341 48807
rect 2924 48776 3341 48804
rect 2924 48764 2930 48776
rect 3329 48773 3341 48776
rect 3375 48773 3387 48807
rect 3329 48767 3387 48773
rect 14366 48764 14372 48816
rect 14424 48804 14430 48816
rect 22922 48804 22928 48816
rect 14424 48776 22928 48804
rect 14424 48764 14430 48776
rect 22922 48764 22928 48776
rect 22980 48764 22986 48816
rect 25774 48764 25780 48816
rect 25832 48804 25838 48816
rect 25961 48807 26019 48813
rect 25961 48804 25973 48807
rect 25832 48776 25973 48804
rect 25832 48764 25838 48776
rect 25961 48773 25973 48776
rect 26007 48773 26019 48807
rect 25961 48767 26019 48773
rect 26418 48764 26424 48816
rect 26476 48804 26482 48816
rect 27433 48807 27491 48813
rect 27433 48804 27445 48807
rect 26476 48776 27445 48804
rect 26476 48764 26482 48776
rect 27433 48773 27445 48776
rect 27479 48773 27491 48807
rect 27433 48767 27491 48773
rect 28537 48807 28595 48813
rect 28537 48773 28549 48807
rect 28583 48804 28595 48807
rect 28994 48804 29000 48816
rect 28583 48776 29000 48804
rect 28583 48773 28595 48776
rect 28537 48767 28595 48773
rect 28994 48764 29000 48776
rect 29052 48764 29058 48816
rect 38746 48764 38752 48816
rect 38804 48804 38810 48816
rect 39209 48807 39267 48813
rect 39209 48804 39221 48807
rect 38804 48776 39221 48804
rect 38804 48764 38810 48776
rect 39209 48773 39221 48776
rect 39255 48773 39267 48807
rect 39209 48767 39267 48773
rect 40865 48807 40923 48813
rect 40865 48773 40877 48807
rect 40911 48804 40923 48807
rect 41414 48804 41420 48816
rect 40911 48776 41420 48804
rect 40911 48773 40923 48776
rect 40865 48767 40923 48773
rect 41414 48764 41420 48776
rect 41472 48764 41478 48816
rect 41509 48807 41567 48813
rect 41509 48773 41521 48807
rect 41555 48804 41567 48807
rect 41874 48804 41880 48816
rect 41555 48776 41880 48804
rect 41555 48773 41567 48776
rect 41509 48767 41567 48773
rect 41874 48764 41880 48776
rect 41932 48764 41938 48816
rect 47762 48804 47768 48816
rect 47723 48776 47768 48804
rect 47762 48764 47768 48776
rect 47820 48764 47826 48816
rect 6638 48736 6644 48748
rect 6599 48708 6644 48736
rect 6638 48696 6644 48708
rect 6696 48696 6702 48748
rect 8938 48736 8944 48748
rect 8899 48708 8944 48736
rect 8938 48696 8944 48708
rect 8996 48696 9002 48748
rect 13998 48736 14004 48748
rect 13959 48708 14004 48736
rect 13998 48696 14004 48708
rect 14056 48696 14062 48748
rect 15289 48739 15347 48745
rect 15289 48705 15301 48739
rect 15335 48736 15347 48739
rect 16114 48736 16120 48748
rect 15335 48708 16120 48736
rect 15335 48705 15347 48708
rect 15289 48699 15347 48705
rect 16114 48696 16120 48708
rect 16172 48696 16178 48748
rect 16666 48736 16672 48748
rect 16627 48708 16672 48736
rect 16666 48696 16672 48708
rect 16724 48696 16730 48748
rect 21269 48739 21327 48745
rect 21269 48705 21281 48739
rect 21315 48736 21327 48739
rect 22002 48736 22008 48748
rect 21315 48708 22008 48736
rect 21315 48705 21327 48708
rect 21269 48699 21327 48705
rect 22002 48696 22008 48708
rect 22060 48696 22066 48748
rect 32122 48736 32128 48748
rect 32083 48708 32128 48736
rect 32122 48696 32128 48708
rect 32180 48696 32186 48748
rect 34882 48736 34888 48748
rect 34843 48708 34888 48736
rect 34882 48696 34888 48708
rect 34940 48696 34946 48748
rect 1489 48671 1547 48677
rect 1489 48637 1501 48671
rect 1535 48637 1547 48671
rect 1489 48631 1547 48637
rect 1673 48671 1731 48677
rect 1673 48637 1685 48671
rect 1719 48668 1731 48671
rect 3050 48668 3056 48680
rect 1719 48640 3056 48668
rect 1719 48637 1731 48640
rect 1673 48631 1731 48637
rect 1504 48600 1532 48631
rect 3050 48628 3056 48640
rect 3108 48628 3114 48680
rect 3786 48668 3792 48680
rect 3747 48640 3792 48668
rect 3786 48628 3792 48640
rect 3844 48628 3850 48680
rect 3973 48671 4031 48677
rect 3973 48637 3985 48671
rect 4019 48668 4031 48671
rect 4062 48668 4068 48680
rect 4019 48640 4068 48668
rect 4019 48637 4031 48640
rect 3973 48631 4031 48637
rect 4062 48628 4068 48640
rect 4120 48628 4126 48680
rect 4706 48668 4712 48680
rect 4667 48640 4712 48668
rect 4706 48628 4712 48640
rect 4764 48628 4770 48680
rect 6825 48671 6883 48677
rect 6825 48637 6837 48671
rect 6871 48668 6883 48671
rect 7742 48668 7748 48680
rect 6871 48640 7748 48668
rect 6871 48637 6883 48640
rect 6825 48631 6883 48637
rect 7742 48628 7748 48640
rect 7800 48628 7806 48680
rect 7837 48671 7895 48677
rect 7837 48637 7849 48671
rect 7883 48637 7895 48671
rect 9122 48668 9128 48680
rect 9083 48640 9128 48668
rect 7837 48631 7895 48637
rect 3878 48600 3884 48612
rect 1504 48572 3884 48600
rect 3878 48560 3884 48572
rect 3936 48560 3942 48612
rect 7098 48560 7104 48612
rect 7156 48600 7162 48612
rect 7852 48600 7880 48631
rect 9122 48628 9128 48640
rect 9180 48628 9186 48680
rect 9674 48668 9680 48680
rect 9635 48640 9680 48668
rect 9674 48628 9680 48640
rect 9732 48628 9738 48680
rect 11514 48668 11520 48680
rect 11475 48640 11520 48668
rect 11514 48628 11520 48640
rect 11572 48628 11578 48680
rect 11698 48668 11704 48680
rect 11659 48640 11704 48668
rect 11698 48628 11704 48640
rect 11756 48628 11762 48680
rect 12434 48628 12440 48680
rect 12492 48668 12498 48680
rect 14277 48671 14335 48677
rect 12492 48640 12537 48668
rect 12492 48628 12498 48640
rect 14277 48637 14289 48671
rect 14323 48637 14335 48671
rect 14277 48631 14335 48637
rect 15565 48671 15623 48677
rect 15565 48637 15577 48671
rect 15611 48637 15623 48671
rect 16850 48668 16856 48680
rect 16811 48640 16856 48668
rect 15565 48631 15623 48637
rect 7156 48572 7880 48600
rect 7156 48560 7162 48572
rect 14292 48532 14320 48631
rect 15580 48600 15608 48631
rect 16850 48628 16856 48640
rect 16908 48628 16914 48680
rect 16942 48628 16948 48680
rect 17000 48668 17006 48680
rect 17129 48671 17187 48677
rect 17129 48668 17141 48671
rect 17000 48640 17141 48668
rect 17000 48628 17006 48640
rect 17129 48637 17141 48640
rect 17175 48637 17187 48671
rect 17129 48631 17187 48637
rect 22281 48671 22339 48677
rect 22281 48637 22293 48671
rect 22327 48668 22339 48671
rect 22741 48671 22799 48677
rect 22741 48668 22753 48671
rect 22327 48640 22753 48668
rect 22327 48637 22339 48640
rect 22281 48631 22339 48637
rect 22741 48637 22753 48640
rect 22787 48637 22799 48671
rect 22741 48631 22799 48637
rect 22925 48671 22983 48677
rect 22925 48637 22937 48671
rect 22971 48668 22983 48671
rect 23658 48668 23664 48680
rect 22971 48640 23664 48668
rect 22971 48637 22983 48640
rect 22925 48631 22983 48637
rect 23658 48628 23664 48640
rect 23716 48628 23722 48680
rect 23753 48671 23811 48677
rect 23753 48637 23765 48671
rect 23799 48637 23811 48671
rect 23753 48631 23811 48637
rect 29181 48671 29239 48677
rect 29181 48637 29193 48671
rect 29227 48668 29239 48671
rect 29227 48640 29316 48668
rect 29227 48637 29239 48640
rect 29181 48631 29239 48637
rect 18598 48600 18604 48612
rect 15580 48572 18604 48600
rect 18598 48560 18604 48572
rect 18656 48560 18662 48612
rect 20806 48600 20812 48612
rect 20088 48572 20812 48600
rect 20088 48532 20116 48572
rect 20806 48560 20812 48572
rect 20864 48560 20870 48612
rect 23198 48560 23204 48612
rect 23256 48600 23262 48612
rect 23768 48600 23796 48631
rect 29288 48612 29316 48640
rect 29362 48628 29368 48680
rect 29420 48668 29426 48680
rect 29638 48668 29644 48680
rect 29420 48640 29465 48668
rect 29599 48640 29644 48668
rect 29420 48628 29426 48640
rect 29638 48628 29644 48640
rect 29696 48628 29702 48680
rect 32306 48668 32312 48680
rect 32267 48640 32312 48668
rect 32306 48628 32312 48640
rect 32364 48628 32370 48680
rect 32858 48668 32864 48680
rect 32819 48640 32864 48668
rect 32858 48628 32864 48640
rect 32916 48628 32922 48680
rect 35069 48671 35127 48677
rect 35069 48637 35081 48671
rect 35115 48668 35127 48671
rect 36078 48668 36084 48680
rect 35115 48640 35894 48668
rect 36039 48640 36084 48668
rect 35115 48637 35127 48640
rect 35069 48631 35127 48637
rect 27614 48600 27620 48612
rect 23256 48572 23796 48600
rect 27575 48572 27620 48600
rect 23256 48560 23262 48572
rect 27614 48560 27620 48572
rect 27672 48560 27678 48612
rect 29270 48560 29276 48612
rect 29328 48560 29334 48612
rect 35866 48600 35894 48640
rect 36078 48628 36084 48640
rect 36136 48628 36142 48680
rect 38565 48671 38623 48677
rect 38565 48637 38577 48671
rect 38611 48668 38623 48671
rect 39025 48671 39083 48677
rect 39025 48668 39037 48671
rect 38611 48640 39037 48668
rect 38611 48637 38623 48640
rect 38565 48631 38623 48637
rect 39025 48637 39037 48640
rect 39071 48637 39083 48671
rect 39025 48631 39083 48637
rect 42613 48671 42671 48677
rect 42613 48637 42625 48671
rect 42659 48637 42671 48671
rect 42794 48668 42800 48680
rect 42755 48640 42800 48668
rect 42613 48631 42671 48637
rect 36170 48600 36176 48612
rect 35866 48572 36176 48600
rect 36170 48560 36176 48572
rect 36228 48560 36234 48612
rect 42628 48600 42656 48631
rect 42794 48628 42800 48640
rect 42852 48628 42858 48680
rect 43162 48668 43168 48680
rect 43123 48640 43168 48668
rect 43162 48628 43168 48640
rect 43220 48628 43226 48680
rect 44910 48668 44916 48680
rect 44871 48640 44916 48668
rect 44910 48628 44916 48640
rect 44968 48628 44974 48680
rect 45094 48668 45100 48680
rect 45055 48640 45100 48668
rect 45094 48628 45100 48640
rect 45152 48628 45158 48680
rect 45738 48668 45744 48680
rect 45699 48640 45744 48668
rect 45738 48628 45744 48640
rect 45796 48628 45802 48680
rect 42978 48600 42984 48612
rect 42628 48572 42984 48600
rect 42978 48560 42984 48572
rect 43036 48560 43042 48612
rect 20254 48532 20260 48544
rect 14292 48504 20116 48532
rect 20215 48504 20260 48532
rect 20254 48492 20260 48504
rect 20312 48492 20318 48544
rect 25406 48532 25412 48544
rect 25367 48504 25412 48532
rect 25406 48492 25412 48504
rect 25464 48492 25470 48544
rect 25498 48492 25504 48544
rect 25556 48532 25562 48544
rect 26053 48535 26111 48541
rect 26053 48532 26065 48535
rect 25556 48504 26065 48532
rect 25556 48492 25562 48504
rect 26053 48501 26065 48504
rect 26099 48501 26111 48535
rect 26053 48495 26111 48501
rect 28442 48492 28448 48544
rect 28500 48532 28506 48544
rect 28629 48535 28687 48541
rect 28629 48532 28641 48535
rect 28500 48504 28641 48532
rect 28500 48492 28506 48504
rect 28629 48501 28641 48504
rect 28675 48501 28687 48535
rect 28629 48495 28687 48501
rect 33778 48492 33784 48544
rect 33836 48532 33842 48544
rect 34146 48532 34152 48544
rect 33836 48504 34152 48532
rect 33836 48492 33842 48504
rect 34146 48492 34152 48504
rect 34204 48492 34210 48544
rect 37458 48532 37464 48544
rect 37419 48504 37464 48532
rect 37458 48492 37464 48504
rect 37516 48492 37522 48544
rect 41598 48532 41604 48544
rect 41559 48504 41604 48532
rect 41598 48492 41604 48504
rect 41656 48492 41662 48544
rect 48041 48535 48099 48541
rect 48041 48501 48053 48535
rect 48087 48532 48099 48535
rect 48222 48532 48228 48544
rect 48087 48504 48228 48532
rect 48087 48501 48099 48504
rect 48041 48495 48099 48501
rect 48222 48492 48228 48504
rect 48280 48492 48286 48544
rect 1104 48442 48852 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 48852 48442
rect 1104 48368 48852 48390
rect 9122 48328 9128 48340
rect 9083 48300 9128 48328
rect 9122 48288 9128 48300
rect 9180 48288 9186 48340
rect 11698 48288 11704 48340
rect 11756 48328 11762 48340
rect 12069 48331 12127 48337
rect 12069 48328 12081 48331
rect 11756 48300 12081 48328
rect 11756 48288 11762 48300
rect 12069 48297 12081 48300
rect 12115 48297 12127 48331
rect 12069 48291 12127 48297
rect 29914 48288 29920 48340
rect 29972 48328 29978 48340
rect 30193 48331 30251 48337
rect 30193 48328 30205 48331
rect 29972 48300 30205 48328
rect 29972 48288 29978 48300
rect 30193 48297 30205 48300
rect 30239 48297 30251 48331
rect 38746 48328 38752 48340
rect 38707 48300 38752 48328
rect 30193 48291 30251 48297
rect 38746 48288 38752 48300
rect 38804 48288 38810 48340
rect 14 48220 20 48272
rect 72 48260 78 48272
rect 7742 48260 7748 48272
rect 72 48232 4292 48260
rect 7703 48232 7748 48260
rect 72 48220 78 48232
rect 1302 48152 1308 48204
rect 1360 48192 1366 48204
rect 1857 48195 1915 48201
rect 1857 48192 1869 48195
rect 1360 48164 1869 48192
rect 1360 48152 1366 48164
rect 1857 48161 1869 48164
rect 1903 48161 1915 48195
rect 1857 48155 1915 48161
rect 4264 48133 4292 48232
rect 7742 48220 7748 48232
rect 7800 48220 7806 48272
rect 17126 48220 17132 48272
rect 17184 48260 17190 48272
rect 23658 48260 23664 48272
rect 17184 48232 23520 48260
rect 23619 48232 23664 48260
rect 17184 48220 17190 48232
rect 5166 48152 5172 48204
rect 5224 48192 5230 48204
rect 5813 48195 5871 48201
rect 5813 48192 5825 48195
rect 5224 48164 5825 48192
rect 5224 48152 5230 48164
rect 5813 48161 5825 48164
rect 5859 48161 5871 48195
rect 5813 48155 5871 48161
rect 9677 48195 9735 48201
rect 9677 48161 9689 48195
rect 9723 48192 9735 48195
rect 9858 48192 9864 48204
rect 9723 48164 9864 48192
rect 9723 48161 9735 48164
rect 9677 48155 9735 48161
rect 9858 48152 9864 48164
rect 9916 48152 9922 48204
rect 10318 48192 10324 48204
rect 10279 48164 10324 48192
rect 10318 48152 10324 48164
rect 10376 48152 10382 48204
rect 14918 48192 14924 48204
rect 14879 48164 14924 48192
rect 14918 48152 14924 48164
rect 14976 48152 14982 48204
rect 16574 48152 16580 48204
rect 16632 48192 16638 48204
rect 16761 48195 16819 48201
rect 16761 48192 16773 48195
rect 16632 48164 16773 48192
rect 16632 48152 16638 48164
rect 16761 48161 16773 48164
rect 16807 48161 16819 48195
rect 17402 48192 17408 48204
rect 17363 48164 17408 48192
rect 16761 48155 16819 48161
rect 17402 48152 17408 48164
rect 17460 48152 17466 48204
rect 19981 48195 20039 48201
rect 19981 48161 19993 48195
rect 20027 48192 20039 48195
rect 20254 48192 20260 48204
rect 20027 48164 20260 48192
rect 20027 48161 20039 48164
rect 19981 48155 20039 48161
rect 20254 48152 20260 48164
rect 20312 48152 20318 48204
rect 20622 48152 20628 48204
rect 20680 48192 20686 48204
rect 20717 48195 20775 48201
rect 20717 48192 20729 48195
rect 20680 48164 20729 48192
rect 20680 48152 20686 48164
rect 20717 48161 20729 48164
rect 20763 48161 20775 48195
rect 20717 48155 20775 48161
rect 21376 48164 23428 48192
rect 1397 48127 1455 48133
rect 1397 48093 1409 48127
rect 1443 48093 1455 48127
rect 1397 48087 1455 48093
rect 4249 48127 4307 48133
rect 4249 48093 4261 48127
rect 4295 48093 4307 48127
rect 5350 48124 5356 48136
rect 5311 48096 5356 48124
rect 4249 48087 4307 48093
rect 1412 47988 1440 48087
rect 5350 48084 5356 48096
rect 5408 48084 5414 48136
rect 7098 48084 7104 48136
rect 7156 48124 7162 48136
rect 7653 48127 7711 48133
rect 7653 48124 7665 48127
rect 7156 48096 7665 48124
rect 7156 48084 7162 48096
rect 7653 48093 7665 48096
rect 7699 48124 7711 48127
rect 8938 48124 8944 48136
rect 7699 48096 8944 48124
rect 7699 48093 7711 48096
rect 7653 48087 7711 48093
rect 8938 48084 8944 48096
rect 8996 48084 9002 48136
rect 9033 48127 9091 48133
rect 9033 48093 9045 48127
rect 9079 48124 9091 48127
rect 9122 48124 9128 48136
rect 9079 48096 9128 48124
rect 9079 48093 9091 48096
rect 9033 48087 9091 48093
rect 9122 48084 9128 48096
rect 9180 48084 9186 48136
rect 11974 48124 11980 48136
rect 11935 48096 11980 48124
rect 11974 48084 11980 48096
rect 12032 48084 12038 48136
rect 14458 48124 14464 48136
rect 14419 48096 14464 48124
rect 14458 48084 14464 48096
rect 14516 48084 14522 48136
rect 1578 48056 1584 48068
rect 1539 48028 1584 48056
rect 1578 48016 1584 48028
rect 1636 48016 1642 48068
rect 4430 48056 4436 48068
rect 4391 48028 4436 48056
rect 4430 48016 4436 48028
rect 4488 48016 4494 48068
rect 5534 48056 5540 48068
rect 5495 48028 5540 48056
rect 5534 48016 5540 48028
rect 5592 48016 5598 48068
rect 9861 48059 9919 48065
rect 9861 48025 9873 48059
rect 9907 48056 9919 48059
rect 9950 48056 9956 48068
rect 9907 48028 9956 48056
rect 9907 48025 9919 48028
rect 9861 48019 9919 48025
rect 9950 48016 9956 48028
rect 10008 48016 10014 48068
rect 14366 48016 14372 48068
rect 14424 48056 14430 48068
rect 14645 48059 14703 48065
rect 14645 48056 14657 48059
rect 14424 48028 14657 48056
rect 14424 48016 14430 48028
rect 14645 48025 14657 48028
rect 14691 48025 14703 48059
rect 14645 48019 14703 48025
rect 16945 48059 17003 48065
rect 16945 48025 16957 48059
rect 16991 48056 17003 48059
rect 17402 48056 17408 48068
rect 16991 48028 17408 48056
rect 16991 48025 17003 48028
rect 16945 48019 17003 48025
rect 17402 48016 17408 48028
rect 17460 48016 17466 48068
rect 20162 48056 20168 48068
rect 20123 48028 20168 48056
rect 20162 48016 20168 48028
rect 20220 48016 20226 48068
rect 4706 47988 4712 48000
rect 1412 47960 4712 47988
rect 4706 47948 4712 47960
rect 4764 47948 4770 48000
rect 7374 47948 7380 48000
rect 7432 47988 7438 48000
rect 21376 47988 21404 48164
rect 21910 48084 21916 48136
rect 21968 48124 21974 48136
rect 22281 48127 22339 48133
rect 22281 48124 22293 48127
rect 21968 48096 22293 48124
rect 21968 48084 21974 48096
rect 22281 48093 22293 48096
rect 22327 48093 22339 48127
rect 22281 48087 22339 48093
rect 22557 48127 22615 48133
rect 22557 48093 22569 48127
rect 22603 48093 22615 48127
rect 22557 48087 22615 48093
rect 7432 47960 21404 47988
rect 7432 47948 7438 47960
rect 21634 47948 21640 48000
rect 21692 47988 21698 48000
rect 22572 47988 22600 48087
rect 23400 48056 23428 48164
rect 23492 48124 23520 48232
rect 23658 48220 23664 48232
rect 23716 48220 23722 48272
rect 25314 48220 25320 48272
rect 25372 48260 25378 48272
rect 28905 48263 28963 48269
rect 25372 48232 26004 48260
rect 25372 48220 25378 48232
rect 25406 48152 25412 48204
rect 25464 48192 25470 48204
rect 25976 48201 26004 48232
rect 28905 48229 28917 48263
rect 28951 48260 28963 48263
rect 29362 48260 29368 48272
rect 28951 48232 29368 48260
rect 28951 48229 28963 48232
rect 28905 48223 28963 48229
rect 29362 48220 29368 48232
rect 29420 48220 29426 48272
rect 30837 48263 30895 48269
rect 30837 48229 30849 48263
rect 30883 48260 30895 48263
rect 32306 48260 32312 48272
rect 30883 48232 32312 48260
rect 30883 48229 30895 48232
rect 30837 48223 30895 48229
rect 32306 48220 32312 48232
rect 32364 48220 32370 48272
rect 36722 48220 36728 48272
rect 36780 48260 36786 48272
rect 39945 48263 40003 48269
rect 36780 48232 37596 48260
rect 36780 48220 36786 48232
rect 25777 48195 25835 48201
rect 25777 48192 25789 48195
rect 25464 48164 25789 48192
rect 25464 48152 25470 48164
rect 25777 48161 25789 48164
rect 25823 48161 25835 48195
rect 25777 48155 25835 48161
rect 25961 48195 26019 48201
rect 25961 48161 25973 48195
rect 26007 48161 26019 48195
rect 25961 48155 26019 48161
rect 27617 48195 27675 48201
rect 27617 48161 27629 48195
rect 27663 48192 27675 48195
rect 27706 48192 27712 48204
rect 27663 48164 27712 48192
rect 27663 48161 27675 48164
rect 27617 48155 27675 48161
rect 27706 48152 27712 48164
rect 27764 48152 27770 48204
rect 31389 48195 31447 48201
rect 31389 48161 31401 48195
rect 31435 48192 31447 48195
rect 31938 48192 31944 48204
rect 31435 48164 31944 48192
rect 31435 48161 31447 48164
rect 31389 48155 31447 48161
rect 31938 48152 31944 48164
rect 31996 48152 32002 48204
rect 32214 48192 32220 48204
rect 32175 48164 32220 48192
rect 32214 48152 32220 48164
rect 32272 48152 32278 48204
rect 36357 48195 36415 48201
rect 36357 48161 36369 48195
rect 36403 48192 36415 48195
rect 37458 48192 37464 48204
rect 36403 48164 37464 48192
rect 36403 48161 36415 48164
rect 36357 48155 36415 48161
rect 37458 48152 37464 48164
rect 37516 48152 37522 48204
rect 37568 48201 37596 48232
rect 39945 48229 39957 48263
rect 39991 48260 40003 48263
rect 40034 48260 40040 48272
rect 39991 48232 40040 48260
rect 39991 48229 40003 48232
rect 39945 48223 40003 48229
rect 40034 48220 40040 48232
rect 40092 48220 40098 48272
rect 47026 48220 47032 48272
rect 47084 48260 47090 48272
rect 49602 48260 49608 48272
rect 47084 48232 49608 48260
rect 47084 48220 47090 48232
rect 49602 48220 49608 48232
rect 49660 48220 49666 48272
rect 37553 48195 37611 48201
rect 37553 48161 37565 48195
rect 37599 48161 37611 48195
rect 42518 48192 42524 48204
rect 42479 48164 42524 48192
rect 37553 48155 37611 48161
rect 42518 48152 42524 48164
rect 42576 48152 42582 48204
rect 48133 48195 48191 48201
rect 48133 48161 48145 48195
rect 48179 48192 48191 48195
rect 48314 48192 48320 48204
rect 48179 48164 48320 48192
rect 48179 48161 48191 48164
rect 48133 48155 48191 48161
rect 48314 48152 48320 48164
rect 48372 48152 48378 48204
rect 23569 48127 23627 48133
rect 23569 48124 23581 48127
rect 23492 48096 23581 48124
rect 23569 48093 23581 48096
rect 23615 48124 23627 48127
rect 23842 48124 23848 48136
rect 23615 48096 23848 48124
rect 23615 48093 23627 48096
rect 23569 48087 23627 48093
rect 23842 48084 23848 48096
rect 23900 48084 23906 48136
rect 23952 48096 25452 48124
rect 23952 48056 23980 48096
rect 24946 48056 24952 48068
rect 23400 48028 23980 48056
rect 24907 48028 24952 48056
rect 24946 48016 24952 48028
rect 25004 48016 25010 48068
rect 25222 47988 25228 48000
rect 21692 47960 22600 47988
rect 25183 47960 25228 47988
rect 21692 47948 21698 47960
rect 25222 47948 25228 47960
rect 25280 47948 25286 48000
rect 25424 47988 25452 48096
rect 28074 48084 28080 48136
rect 28132 48124 28138 48136
rect 28261 48127 28319 48133
rect 28261 48124 28273 48127
rect 28132 48096 28273 48124
rect 28132 48084 28138 48096
rect 28261 48093 28273 48096
rect 28307 48093 28319 48127
rect 28261 48087 28319 48093
rect 28813 48127 28871 48133
rect 28813 48093 28825 48127
rect 28859 48093 28871 48127
rect 30098 48124 30104 48136
rect 30059 48096 30104 48124
rect 28813 48087 28871 48093
rect 28166 48016 28172 48068
rect 28224 48056 28230 48068
rect 28828 48056 28856 48087
rect 30098 48084 30104 48096
rect 30156 48084 30162 48136
rect 30742 48124 30748 48136
rect 30703 48096 30748 48124
rect 30742 48084 30748 48096
rect 30800 48084 30806 48136
rect 33778 48084 33784 48136
rect 33836 48124 33842 48136
rect 34057 48127 34115 48133
rect 34057 48124 34069 48127
rect 33836 48096 34069 48124
rect 33836 48084 33842 48096
rect 34057 48093 34069 48096
rect 34103 48093 34115 48127
rect 35710 48124 35716 48136
rect 35671 48096 35716 48124
rect 34057 48087 34115 48093
rect 35710 48084 35716 48096
rect 35768 48084 35774 48136
rect 38654 48124 38660 48136
rect 38615 48096 38660 48124
rect 38654 48084 38660 48096
rect 38712 48084 38718 48136
rect 39850 48124 39856 48136
rect 39811 48096 39856 48124
rect 39850 48084 39856 48096
rect 39908 48084 39914 48136
rect 41046 48124 41052 48136
rect 41007 48096 41052 48124
rect 41046 48084 41052 48096
rect 41104 48084 41110 48136
rect 43898 48124 43904 48136
rect 43859 48096 43904 48124
rect 43898 48084 43904 48096
rect 43956 48084 43962 48136
rect 44450 48084 44456 48136
rect 44508 48124 44514 48136
rect 45005 48127 45063 48133
rect 45005 48124 45017 48127
rect 44508 48096 45017 48124
rect 44508 48084 44514 48096
rect 45005 48093 45017 48096
rect 45051 48093 45063 48127
rect 46293 48127 46351 48133
rect 46293 48124 46305 48127
rect 45005 48087 45063 48093
rect 45526 48096 46305 48124
rect 28224 48028 28856 48056
rect 31573 48059 31631 48065
rect 28224 48016 28230 48028
rect 31573 48025 31585 48059
rect 31619 48056 31631 48059
rect 32214 48056 32220 48068
rect 31619 48028 32220 48056
rect 31619 48025 31631 48028
rect 31573 48019 31631 48025
rect 32214 48016 32220 48028
rect 32272 48016 32278 48068
rect 35805 48059 35863 48065
rect 35805 48025 35817 48059
rect 35851 48056 35863 48059
rect 36541 48059 36599 48065
rect 36541 48056 36553 48059
rect 35851 48028 36553 48056
rect 35851 48025 35863 48028
rect 35805 48019 35863 48025
rect 36541 48025 36553 48028
rect 36587 48025 36599 48059
rect 36541 48019 36599 48025
rect 40402 48016 40408 48068
rect 40460 48056 40466 48068
rect 41233 48059 41291 48065
rect 41233 48056 41245 48059
rect 40460 48028 41245 48056
rect 40460 48016 40466 48028
rect 41233 48025 41245 48028
rect 41279 48025 41291 48059
rect 41233 48019 41291 48025
rect 43806 48016 43812 48068
rect 43864 48056 43870 48068
rect 45526 48056 45554 48096
rect 46293 48093 46305 48096
rect 46339 48093 46351 48127
rect 46293 48087 46351 48093
rect 43864 48028 45554 48056
rect 46477 48059 46535 48065
rect 43864 48016 43870 48028
rect 46477 48025 46489 48059
rect 46523 48056 46535 48059
rect 47670 48056 47676 48068
rect 46523 48028 47676 48056
rect 46523 48025 46535 48028
rect 46477 48019 46535 48025
rect 47670 48016 47676 48028
rect 47728 48016 47734 48068
rect 32122 47988 32128 48000
rect 25424 47960 32128 47988
rect 32122 47948 32128 47960
rect 32180 47948 32186 48000
rect 43990 47948 43996 48000
rect 44048 47988 44054 48000
rect 44085 47991 44143 47997
rect 44085 47988 44097 47991
rect 44048 47960 44097 47988
rect 44048 47948 44054 47960
rect 44085 47957 44097 47960
rect 44131 47957 44143 47991
rect 45186 47988 45192 48000
rect 45147 47960 45192 47988
rect 44085 47951 44143 47957
rect 45186 47948 45192 47960
rect 45244 47948 45250 48000
rect 1104 47898 48852 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 48852 47898
rect 1104 47824 48852 47846
rect 1489 47787 1547 47793
rect 1489 47753 1501 47787
rect 1535 47784 1547 47787
rect 1578 47784 1584 47796
rect 1535 47756 1584 47784
rect 1535 47753 1547 47756
rect 1489 47747 1547 47753
rect 1578 47744 1584 47756
rect 1636 47744 1642 47796
rect 3050 47784 3056 47796
rect 3011 47756 3056 47784
rect 3050 47744 3056 47756
rect 3108 47744 3114 47796
rect 5442 47784 5448 47796
rect 5403 47756 5448 47784
rect 5442 47744 5448 47756
rect 5500 47744 5506 47796
rect 7466 47744 7472 47796
rect 7524 47784 7530 47796
rect 8662 47784 8668 47796
rect 7524 47756 8668 47784
rect 7524 47744 7530 47756
rect 8662 47744 8668 47756
rect 8720 47744 8726 47796
rect 9950 47784 9956 47796
rect 9911 47756 9956 47784
rect 9950 47744 9956 47756
rect 10008 47744 10014 47796
rect 16761 47787 16819 47793
rect 16761 47753 16773 47787
rect 16807 47784 16819 47787
rect 16850 47784 16856 47796
rect 16807 47756 16856 47784
rect 16807 47753 16819 47756
rect 16761 47747 16819 47753
rect 16850 47744 16856 47756
rect 16908 47744 16914 47796
rect 17402 47784 17408 47796
rect 17363 47756 17408 47784
rect 17402 47744 17408 47756
rect 17460 47744 17466 47796
rect 19705 47787 19763 47793
rect 19705 47753 19717 47787
rect 19751 47784 19763 47787
rect 20162 47784 20168 47796
rect 19751 47756 20168 47784
rect 19751 47753 19763 47756
rect 19705 47747 19763 47753
rect 20162 47744 20168 47756
rect 20220 47744 20226 47796
rect 21177 47787 21235 47793
rect 21177 47753 21189 47787
rect 21223 47784 21235 47787
rect 22186 47784 22192 47796
rect 21223 47756 22192 47784
rect 21223 47753 21235 47756
rect 21177 47747 21235 47753
rect 22186 47744 22192 47756
rect 22244 47744 22250 47796
rect 24213 47787 24271 47793
rect 24213 47753 24225 47787
rect 24259 47784 24271 47787
rect 24578 47784 24584 47796
rect 24259 47756 24584 47784
rect 24259 47753 24271 47756
rect 24213 47747 24271 47753
rect 24578 47744 24584 47756
rect 24636 47744 24642 47796
rect 24762 47744 24768 47796
rect 24820 47784 24826 47796
rect 30742 47784 30748 47796
rect 24820 47756 30748 47784
rect 24820 47744 24826 47756
rect 30742 47744 30748 47756
rect 30800 47744 30806 47796
rect 32214 47784 32220 47796
rect 32175 47756 32220 47784
rect 32214 47744 32220 47756
rect 32272 47744 32278 47796
rect 36170 47784 36176 47796
rect 32324 47756 35894 47784
rect 36131 47756 36176 47784
rect 2130 47716 2136 47728
rect 2091 47688 2136 47716
rect 2130 47676 2136 47688
rect 2188 47676 2194 47728
rect 3326 47676 3332 47728
rect 3384 47716 3390 47728
rect 24946 47716 24952 47728
rect 3384 47688 21680 47716
rect 3384 47676 3390 47688
rect 1397 47651 1455 47657
rect 1397 47617 1409 47651
rect 1443 47617 1455 47651
rect 1397 47611 1455 47617
rect 2961 47651 3019 47657
rect 2961 47617 2973 47651
rect 3007 47648 3019 47651
rect 3510 47648 3516 47660
rect 3007 47620 3516 47648
rect 3007 47617 3019 47620
rect 2961 47611 3019 47617
rect 1412 47580 1440 47611
rect 3510 47608 3516 47620
rect 3568 47608 3574 47660
rect 3786 47608 3792 47660
rect 3844 47648 3850 47660
rect 3973 47651 4031 47657
rect 3973 47648 3985 47651
rect 3844 47620 3985 47648
rect 3844 47608 3850 47620
rect 3973 47617 3985 47620
rect 4019 47617 4031 47651
rect 4614 47648 4620 47660
rect 4575 47620 4620 47648
rect 3973 47611 4031 47617
rect 4614 47608 4620 47620
rect 4672 47608 4678 47660
rect 5353 47651 5411 47657
rect 5353 47617 5365 47651
rect 5399 47648 5411 47651
rect 7374 47648 7380 47660
rect 5399 47620 7380 47648
rect 5399 47617 5411 47620
rect 5353 47611 5411 47617
rect 7374 47608 7380 47620
rect 7432 47608 7438 47660
rect 8938 47608 8944 47660
rect 8996 47648 9002 47660
rect 9861 47651 9919 47657
rect 9861 47648 9873 47651
rect 8996 47620 9873 47648
rect 8996 47608 9002 47620
rect 9861 47617 9873 47620
rect 9907 47617 9919 47651
rect 9861 47611 9919 47617
rect 11514 47608 11520 47660
rect 11572 47648 11578 47660
rect 11793 47651 11851 47657
rect 11793 47648 11805 47651
rect 11572 47620 11805 47648
rect 11572 47608 11578 47620
rect 11793 47617 11805 47620
rect 11839 47617 11851 47651
rect 11793 47611 11851 47617
rect 14458 47608 14464 47660
rect 14516 47648 14522 47660
rect 14645 47651 14703 47657
rect 14645 47648 14657 47651
rect 14516 47620 14657 47648
rect 14516 47608 14522 47620
rect 14645 47617 14657 47620
rect 14691 47617 14703 47651
rect 16666 47648 16672 47660
rect 16627 47620 16672 47648
rect 14645 47611 14703 47617
rect 16666 47608 16672 47620
rect 16724 47608 16730 47660
rect 17310 47648 17316 47660
rect 17271 47620 17316 47648
rect 17310 47608 17316 47620
rect 17368 47608 17374 47660
rect 19613 47651 19671 47657
rect 19613 47617 19625 47651
rect 19659 47648 19671 47651
rect 20070 47648 20076 47660
rect 19659 47620 20076 47648
rect 19659 47617 19671 47620
rect 19613 47611 19671 47617
rect 20070 47608 20076 47620
rect 20128 47608 20134 47660
rect 21085 47651 21143 47657
rect 21085 47617 21097 47651
rect 21131 47617 21143 47651
rect 21085 47611 21143 47617
rect 2498 47580 2504 47592
rect 1412 47552 2504 47580
rect 2498 47540 2504 47552
rect 2556 47580 2562 47592
rect 7466 47580 7472 47592
rect 2556 47552 6914 47580
rect 7427 47552 7472 47580
rect 2556 47540 2562 47552
rect 4430 47472 4436 47524
rect 4488 47512 4494 47524
rect 5442 47512 5448 47524
rect 4488 47484 5448 47512
rect 4488 47472 4494 47484
rect 5442 47472 5448 47484
rect 5500 47472 5506 47524
rect 6886 47512 6914 47552
rect 7466 47540 7472 47552
rect 7524 47540 7530 47592
rect 7653 47583 7711 47589
rect 7653 47549 7665 47583
rect 7699 47580 7711 47583
rect 9030 47580 9036 47592
rect 7699 47552 9036 47580
rect 7699 47549 7711 47552
rect 7653 47543 7711 47549
rect 9030 47540 9036 47552
rect 9088 47540 9094 47592
rect 9214 47580 9220 47592
rect 9175 47552 9220 47580
rect 9214 47540 9220 47552
rect 9272 47540 9278 47592
rect 11974 47540 11980 47592
rect 12032 47580 12038 47592
rect 17126 47580 17132 47592
rect 12032 47552 17132 47580
rect 12032 47540 12038 47552
rect 17126 47540 17132 47552
rect 17184 47540 17190 47592
rect 17218 47512 17224 47524
rect 6886 47484 17224 47512
rect 17218 47472 17224 47484
rect 17276 47472 17282 47524
rect 21100 47512 21128 47611
rect 21652 47512 21680 47688
rect 21836 47688 24952 47716
rect 21836 47657 21864 47688
rect 24946 47676 24952 47688
rect 25004 47676 25010 47728
rect 25056 47688 26832 47716
rect 21821 47651 21879 47657
rect 21821 47617 21833 47651
rect 21867 47617 21879 47651
rect 21821 47611 21879 47617
rect 24121 47651 24179 47657
rect 24121 47617 24133 47651
rect 24167 47648 24179 47651
rect 24210 47648 24216 47660
rect 24167 47620 24216 47648
rect 24167 47617 24179 47620
rect 24121 47611 24179 47617
rect 24210 47608 24216 47620
rect 24268 47648 24274 47660
rect 25056 47648 25084 47688
rect 25222 47648 25228 47660
rect 24268 47620 25084 47648
rect 25183 47620 25228 47648
rect 24268 47608 24274 47620
rect 25222 47608 25228 47620
rect 25280 47608 25286 47660
rect 22002 47580 22008 47592
rect 21963 47552 22008 47580
rect 22002 47540 22008 47552
rect 22060 47540 22066 47592
rect 22281 47583 22339 47589
rect 22281 47549 22293 47583
rect 22327 47549 22339 47583
rect 22281 47543 22339 47549
rect 22296 47512 22324 47543
rect 25130 47540 25136 47592
rect 25188 47580 25194 47592
rect 25501 47583 25559 47589
rect 25501 47580 25513 47583
rect 25188 47552 25513 47580
rect 25188 47540 25194 47552
rect 25501 47549 25513 47552
rect 25547 47580 25559 47583
rect 26694 47580 26700 47592
rect 25547 47552 26700 47580
rect 25547 47549 25559 47552
rect 25501 47543 25559 47549
rect 26694 47540 26700 47552
rect 26752 47540 26758 47592
rect 26804 47580 26832 47688
rect 26988 47688 30052 47716
rect 26878 47608 26884 47660
rect 26936 47648 26942 47660
rect 26988 47657 27016 47688
rect 26973 47651 27031 47657
rect 26973 47648 26985 47651
rect 26936 47620 26985 47648
rect 26936 47608 26942 47620
rect 26973 47617 26985 47620
rect 27019 47617 27031 47651
rect 26973 47611 27031 47617
rect 27065 47651 27123 47657
rect 27065 47617 27077 47651
rect 27111 47648 27123 47651
rect 27154 47648 27160 47660
rect 27111 47620 27160 47648
rect 27111 47617 27123 47620
rect 27065 47611 27123 47617
rect 27154 47608 27160 47620
rect 27212 47608 27218 47660
rect 28074 47648 28080 47660
rect 28035 47620 28080 47648
rect 28074 47608 28080 47620
rect 28132 47608 28138 47660
rect 27522 47580 27528 47592
rect 26804 47552 27528 47580
rect 27522 47540 27528 47552
rect 27580 47540 27586 47592
rect 28261 47583 28319 47589
rect 28261 47549 28273 47583
rect 28307 47580 28319 47583
rect 28534 47580 28540 47592
rect 28307 47552 28540 47580
rect 28307 47549 28319 47552
rect 28261 47543 28319 47549
rect 28534 47540 28540 47552
rect 28592 47540 28598 47592
rect 28629 47583 28687 47589
rect 28629 47549 28641 47583
rect 28675 47549 28687 47583
rect 29546 47580 29552 47592
rect 28629 47543 28687 47549
rect 28736 47552 29552 47580
rect 25406 47512 25412 47524
rect 21100 47484 21588 47512
rect 21652 47484 22324 47512
rect 24228 47484 25412 47512
rect 1946 47404 1952 47456
rect 2004 47444 2010 47456
rect 2225 47447 2283 47453
rect 2225 47444 2237 47447
rect 2004 47416 2237 47444
rect 2004 47404 2010 47416
rect 2225 47413 2237 47416
rect 2271 47413 2283 47447
rect 4798 47444 4804 47456
rect 4759 47416 4804 47444
rect 2225 47407 2283 47413
rect 4798 47404 4804 47416
rect 4856 47404 4862 47456
rect 21560 47444 21588 47484
rect 24228 47444 24256 47484
rect 25406 47472 25412 47484
rect 25464 47472 25470 47524
rect 28350 47472 28356 47524
rect 28408 47512 28414 47524
rect 28644 47512 28672 47543
rect 28408 47484 28672 47512
rect 28408 47472 28414 47484
rect 21560 47416 24256 47444
rect 24302 47404 24308 47456
rect 24360 47444 24366 47456
rect 28736 47444 28764 47552
rect 29546 47540 29552 47552
rect 29604 47540 29610 47592
rect 30024 47512 30052 47688
rect 30098 47676 30104 47728
rect 30156 47716 30162 47728
rect 32324 47716 32352 47756
rect 30156 47688 32352 47716
rect 33229 47719 33287 47725
rect 30156 47676 30162 47688
rect 33229 47685 33241 47719
rect 33275 47716 33287 47719
rect 33965 47719 34023 47725
rect 33965 47716 33977 47719
rect 33275 47688 33977 47716
rect 33275 47685 33287 47688
rect 33229 47679 33287 47685
rect 33965 47685 33977 47688
rect 34011 47685 34023 47719
rect 35866 47716 35894 47756
rect 36170 47744 36176 47756
rect 36228 47744 36234 47796
rect 40402 47784 40408 47796
rect 40363 47756 40408 47784
rect 40402 47744 40408 47756
rect 40460 47744 40466 47796
rect 42705 47787 42763 47793
rect 42705 47753 42717 47787
rect 42751 47784 42763 47787
rect 42794 47784 42800 47796
rect 42751 47756 42800 47784
rect 42751 47753 42763 47756
rect 42705 47747 42763 47753
rect 42794 47744 42800 47756
rect 42852 47744 42858 47796
rect 43625 47787 43683 47793
rect 43625 47753 43637 47787
rect 43671 47784 43683 47787
rect 45370 47784 45376 47796
rect 43671 47756 45376 47784
rect 43671 47753 43683 47756
rect 43625 47747 43683 47753
rect 45370 47744 45376 47756
rect 45428 47744 45434 47796
rect 46658 47716 46664 47728
rect 35866 47688 43576 47716
rect 46619 47688 46664 47716
rect 33965 47679 34023 47685
rect 43548 47660 43576 47688
rect 46658 47676 46664 47688
rect 46716 47676 46722 47728
rect 47765 47719 47823 47725
rect 47765 47685 47777 47719
rect 47811 47716 47823 47719
rect 47854 47716 47860 47728
rect 47811 47688 47860 47716
rect 47811 47685 47823 47688
rect 47765 47679 47823 47685
rect 47854 47676 47860 47688
rect 47912 47676 47918 47728
rect 30558 47648 30564 47660
rect 30519 47620 30564 47648
rect 30558 47608 30564 47620
rect 30616 47608 30622 47660
rect 31846 47608 31852 47660
rect 31904 47648 31910 47660
rect 32122 47648 32128 47660
rect 31904 47620 32128 47648
rect 31904 47608 31910 47620
rect 32122 47608 32128 47620
rect 32180 47608 32186 47660
rect 33134 47648 33140 47660
rect 33095 47620 33140 47648
rect 33134 47608 33140 47620
rect 33192 47608 33198 47660
rect 33778 47648 33784 47660
rect 33739 47620 33784 47648
rect 33778 47608 33784 47620
rect 33836 47608 33842 47660
rect 36078 47648 36084 47660
rect 36039 47620 36084 47648
rect 36078 47608 36084 47620
rect 36136 47608 36142 47660
rect 39758 47648 39764 47660
rect 39719 47620 39764 47648
rect 39758 47608 39764 47620
rect 39816 47608 39822 47660
rect 40310 47648 40316 47660
rect 40271 47620 40316 47648
rect 40310 47608 40316 47620
rect 40368 47608 40374 47660
rect 41046 47608 41052 47660
rect 41104 47648 41110 47660
rect 41233 47651 41291 47657
rect 41233 47648 41245 47651
rect 41104 47620 41245 47648
rect 41104 47608 41110 47620
rect 41233 47617 41245 47620
rect 41279 47617 41291 47651
rect 41233 47611 41291 47617
rect 41877 47651 41935 47657
rect 41877 47617 41889 47651
rect 41923 47648 41935 47651
rect 41966 47648 41972 47660
rect 41923 47620 41972 47648
rect 41923 47617 41935 47620
rect 41877 47611 41935 47617
rect 41966 47608 41972 47620
rect 42024 47608 42030 47660
rect 42613 47651 42671 47657
rect 42613 47617 42625 47651
rect 42659 47617 42671 47651
rect 43530 47648 43536 47660
rect 43443 47620 43536 47648
rect 42613 47611 42671 47617
rect 34790 47580 34796 47592
rect 34751 47552 34796 47580
rect 34790 47540 34796 47552
rect 34848 47540 34854 47592
rect 42628 47580 42656 47611
rect 43530 47608 43536 47620
rect 43588 47608 43594 47660
rect 44174 47580 44180 47592
rect 38626 47552 42656 47580
rect 44135 47552 44180 47580
rect 38626 47512 38654 47552
rect 30024 47484 38654 47512
rect 24360 47416 28764 47444
rect 42628 47444 42656 47552
rect 44174 47540 44180 47552
rect 44232 47540 44238 47592
rect 44358 47580 44364 47592
rect 44319 47552 44364 47580
rect 44358 47540 44364 47552
rect 44416 47540 44422 47592
rect 45002 47580 45008 47592
rect 44963 47552 45008 47580
rect 45002 47540 45008 47552
rect 45060 47540 45066 47592
rect 47578 47512 47584 47524
rect 45526 47484 47584 47512
rect 45526 47444 45554 47484
rect 47578 47472 47584 47484
rect 47636 47472 47642 47524
rect 42628 47416 45554 47444
rect 46937 47447 46995 47453
rect 24360 47404 24366 47416
rect 46937 47413 46949 47447
rect 46983 47444 46995 47447
rect 47118 47444 47124 47456
rect 46983 47416 47124 47444
rect 46983 47413 46995 47416
rect 46937 47407 46995 47413
rect 47118 47404 47124 47416
rect 47176 47404 47182 47456
rect 47762 47404 47768 47456
rect 47820 47444 47826 47456
rect 47857 47447 47915 47453
rect 47857 47444 47869 47447
rect 47820 47416 47869 47444
rect 47820 47404 47826 47416
rect 47857 47413 47869 47416
rect 47903 47413 47915 47447
rect 47857 47407 47915 47413
rect 1104 47354 48852 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 48852 47354
rect 1104 47280 48852 47302
rect 3970 47240 3976 47252
rect 3931 47212 3976 47240
rect 3970 47200 3976 47212
rect 4028 47200 4034 47252
rect 5534 47240 5540 47252
rect 5495 47212 5540 47240
rect 5534 47200 5540 47212
rect 5592 47200 5598 47252
rect 9030 47240 9036 47252
rect 8991 47212 9036 47240
rect 9030 47200 9036 47212
rect 9088 47200 9094 47252
rect 14366 47240 14372 47252
rect 14327 47212 14372 47240
rect 14366 47200 14372 47212
rect 14424 47200 14430 47252
rect 16666 47200 16672 47252
rect 16724 47240 16730 47252
rect 24302 47240 24308 47252
rect 16724 47212 24308 47240
rect 16724 47200 16730 47212
rect 24302 47200 24308 47212
rect 24360 47200 24366 47252
rect 24394 47200 24400 47252
rect 24452 47240 24458 47252
rect 24581 47243 24639 47249
rect 24581 47240 24593 47243
rect 24452 47212 24593 47240
rect 24452 47200 24458 47212
rect 24581 47209 24593 47212
rect 24627 47209 24639 47243
rect 24581 47203 24639 47209
rect 24854 47200 24860 47252
rect 24912 47240 24918 47252
rect 26142 47240 26148 47252
rect 24912 47212 26148 47240
rect 24912 47200 24918 47212
rect 26142 47200 26148 47212
rect 26200 47240 26206 47252
rect 26329 47243 26387 47249
rect 26329 47240 26341 47243
rect 26200 47212 26341 47240
rect 26200 47200 26206 47212
rect 26329 47209 26341 47212
rect 26375 47209 26387 47243
rect 26329 47203 26387 47209
rect 26694 47200 26700 47252
rect 26752 47240 26758 47252
rect 36078 47240 36084 47252
rect 26752 47212 36084 47240
rect 26752 47200 26758 47212
rect 36078 47200 36084 47212
rect 36136 47240 36142 47252
rect 37182 47240 37188 47252
rect 36136 47212 37188 47240
rect 36136 47200 36142 47212
rect 37182 47200 37188 47212
rect 37240 47200 37246 47252
rect 42978 47240 42984 47252
rect 42939 47212 42984 47240
rect 42978 47200 42984 47212
rect 43036 47200 43042 47252
rect 43806 47240 43812 47252
rect 43767 47212 43812 47240
rect 43806 47200 43812 47212
rect 43864 47200 43870 47252
rect 44358 47240 44364 47252
rect 44319 47212 44364 47240
rect 44358 47200 44364 47212
rect 44416 47200 44422 47252
rect 45094 47200 45100 47252
rect 45152 47240 45158 47252
rect 45281 47243 45339 47249
rect 45281 47240 45293 47243
rect 45152 47212 45293 47240
rect 45152 47200 45158 47212
rect 45281 47209 45293 47212
rect 45327 47209 45339 47243
rect 45281 47203 45339 47209
rect 3602 47172 3608 47184
rect 1412 47144 3608 47172
rect 1412 47113 1440 47144
rect 3602 47132 3608 47144
rect 3660 47132 3666 47184
rect 3878 47132 3884 47184
rect 3936 47172 3942 47184
rect 4617 47175 4675 47181
rect 4617 47172 4629 47175
rect 3936 47144 4629 47172
rect 3936 47132 3942 47144
rect 4617 47141 4629 47144
rect 4663 47141 4675 47175
rect 4617 47135 4675 47141
rect 17310 47132 17316 47184
rect 17368 47172 17374 47184
rect 17368 47144 35894 47172
rect 17368 47132 17374 47144
rect 1397 47107 1455 47113
rect 1397 47073 1409 47107
rect 1443 47073 1455 47107
rect 1854 47104 1860 47116
rect 1815 47076 1860 47104
rect 1397 47067 1455 47073
rect 1854 47064 1860 47076
rect 1912 47064 1918 47116
rect 9122 47064 9128 47116
rect 9180 47104 9186 47116
rect 24762 47104 24768 47116
rect 9180 47076 24768 47104
rect 9180 47064 9186 47076
rect 24762 47064 24768 47076
rect 24820 47064 24826 47116
rect 33134 47104 33140 47116
rect 24964 47076 33140 47104
rect 4890 46996 4896 47048
rect 4948 47036 4954 47048
rect 5445 47039 5503 47045
rect 5445 47036 5457 47039
rect 4948 47008 5457 47036
rect 4948 46996 4954 47008
rect 5445 47005 5457 47008
rect 5491 47005 5503 47039
rect 5445 46999 5503 47005
rect 8941 47039 8999 47045
rect 8941 47005 8953 47039
rect 8987 47036 8999 47039
rect 9398 47036 9404 47048
rect 8987 47008 9404 47036
rect 8987 47005 8999 47008
rect 8941 46999 8999 47005
rect 9398 46996 9404 47008
rect 9456 46996 9462 47048
rect 14274 47036 14280 47048
rect 14235 47008 14280 47036
rect 14274 46996 14280 47008
rect 14332 46996 14338 47048
rect 21726 46996 21732 47048
rect 21784 47036 21790 47048
rect 21821 47039 21879 47045
rect 21821 47036 21833 47039
rect 21784 47008 21833 47036
rect 21784 46996 21790 47008
rect 21821 47005 21833 47008
rect 21867 47005 21879 47039
rect 24854 47036 24860 47048
rect 21821 46999 21879 47005
rect 21928 47008 24860 47036
rect 1578 46968 1584 46980
rect 1539 46940 1584 46968
rect 1578 46928 1584 46940
rect 1636 46928 1642 46980
rect 15470 46928 15476 46980
rect 15528 46968 15534 46980
rect 16574 46968 16580 46980
rect 15528 46940 16580 46968
rect 15528 46928 15534 46940
rect 16574 46928 16580 46940
rect 16632 46928 16638 46980
rect 17218 46928 17224 46980
rect 17276 46968 17282 46980
rect 21928 46968 21956 47008
rect 24854 46996 24860 47008
rect 24912 46996 24918 47048
rect 17276 46940 21956 46968
rect 17276 46928 17282 46940
rect 22002 46928 22008 46980
rect 22060 46968 22066 46980
rect 24964 46968 24992 47076
rect 33134 47064 33140 47076
rect 33192 47104 33198 47116
rect 33686 47104 33692 47116
rect 33192 47076 33692 47104
rect 33192 47064 33198 47076
rect 33686 47064 33692 47076
rect 33744 47064 33750 47116
rect 35866 47104 35894 47144
rect 35866 47076 45232 47104
rect 25041 47039 25099 47045
rect 25041 47005 25053 47039
rect 25087 47036 25099 47039
rect 25222 47036 25228 47048
rect 25087 47008 25228 47036
rect 25087 47005 25099 47008
rect 25041 46999 25099 47005
rect 25222 46996 25228 47008
rect 25280 47036 25286 47048
rect 27341 47039 27399 47045
rect 27341 47036 27353 47039
rect 25280 47008 27353 47036
rect 25280 46996 25286 47008
rect 27341 47005 27353 47008
rect 27387 47005 27399 47039
rect 27341 46999 27399 47005
rect 27522 46996 27528 47048
rect 27580 47036 27586 47048
rect 27709 47039 27767 47045
rect 27709 47036 27721 47039
rect 27580 47008 27721 47036
rect 27580 46996 27586 47008
rect 27709 47005 27721 47008
rect 27755 47005 27767 47039
rect 27709 46999 27767 47005
rect 22060 46940 24992 46968
rect 22060 46928 22066 46940
rect 21910 46900 21916 46912
rect 21871 46872 21916 46900
rect 21910 46860 21916 46872
rect 21968 46860 21974 46912
rect 27724 46900 27752 46999
rect 28258 46996 28264 47048
rect 28316 47036 28322 47048
rect 28445 47039 28503 47045
rect 28445 47036 28457 47039
rect 28316 47008 28457 47036
rect 28316 46996 28322 47008
rect 28445 47005 28457 47008
rect 28491 47005 28503 47039
rect 28445 46999 28503 47005
rect 28534 46996 28540 47048
rect 28592 47036 28598 47048
rect 45204 47045 45232 47076
rect 44269 47039 44327 47045
rect 28592 47008 28637 47036
rect 28592 46996 28598 47008
rect 44269 47005 44281 47039
rect 44315 47005 44327 47039
rect 44269 46999 44327 47005
rect 45189 47039 45247 47045
rect 45189 47005 45201 47039
rect 45235 47036 45247 47039
rect 45554 47036 45560 47048
rect 45235 47008 45560 47036
rect 45235 47005 45247 47008
rect 45189 46999 45247 47005
rect 44284 46968 44312 46999
rect 45554 46996 45560 47008
rect 45612 46996 45618 47048
rect 46290 47036 46296 47048
rect 46251 47008 46296 47036
rect 46290 46996 46296 47008
rect 46348 46996 46354 47048
rect 48130 47036 48136 47048
rect 48091 47008 48136 47036
rect 48130 46996 48136 47008
rect 48188 46996 48194 47048
rect 44542 46968 44548 46980
rect 28736 46940 44548 46968
rect 28736 46900 28764 46940
rect 44542 46928 44548 46940
rect 44600 46928 44606 46980
rect 46474 46968 46480 46980
rect 46435 46940 46480 46968
rect 46474 46928 46480 46940
rect 46532 46928 46538 46980
rect 27724 46872 28764 46900
rect 1104 46810 48852 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 48852 46810
rect 1104 46736 48852 46758
rect 1578 46656 1584 46708
rect 1636 46696 1642 46708
rect 2225 46699 2283 46705
rect 2225 46696 2237 46699
rect 1636 46668 2237 46696
rect 1636 46656 1642 46668
rect 2225 46665 2237 46668
rect 2271 46665 2283 46699
rect 2225 46659 2283 46665
rect 43714 46656 43720 46708
rect 43772 46696 43778 46708
rect 44637 46699 44695 46705
rect 44637 46696 44649 46699
rect 43772 46668 44649 46696
rect 43772 46656 43778 46668
rect 44637 46665 44649 46668
rect 44683 46665 44695 46699
rect 47670 46696 47676 46708
rect 47631 46668 47676 46696
rect 44637 46659 44695 46665
rect 47670 46656 47676 46668
rect 47728 46656 47734 46708
rect 21266 46628 21272 46640
rect 21227 46600 21272 46628
rect 21266 46588 21272 46600
rect 21324 46588 21330 46640
rect 24673 46631 24731 46637
rect 24673 46597 24685 46631
rect 24719 46628 24731 46631
rect 25222 46628 25228 46640
rect 24719 46600 25228 46628
rect 24719 46597 24731 46600
rect 24673 46591 24731 46597
rect 25222 46588 25228 46600
rect 25280 46588 25286 46640
rect 47026 46628 47032 46640
rect 46987 46600 47032 46628
rect 47026 46588 47032 46600
rect 47084 46588 47090 46640
rect 1394 46560 1400 46572
rect 1355 46532 1400 46560
rect 1394 46520 1400 46532
rect 1452 46520 1458 46572
rect 2130 46560 2136 46572
rect 2091 46532 2136 46560
rect 2130 46520 2136 46532
rect 2188 46520 2194 46572
rect 2777 46563 2835 46569
rect 2777 46529 2789 46563
rect 2823 46529 2835 46563
rect 3602 46560 3608 46572
rect 3563 46532 3608 46560
rect 2777 46523 2835 46529
rect 2792 46492 2820 46523
rect 3602 46520 3608 46532
rect 3660 46520 3666 46572
rect 4249 46563 4307 46569
rect 4249 46529 4261 46563
rect 4295 46560 4307 46563
rect 4706 46560 4712 46572
rect 4295 46532 4712 46560
rect 4295 46529 4307 46532
rect 4249 46523 4307 46529
rect 4706 46520 4712 46532
rect 4764 46520 4770 46572
rect 26970 46520 26976 46572
rect 27028 46560 27034 46572
rect 28261 46563 28319 46569
rect 28261 46560 28273 46563
rect 27028 46532 28273 46560
rect 27028 46520 27034 46532
rect 28261 46529 28273 46532
rect 28307 46529 28319 46563
rect 44082 46560 44088 46572
rect 44043 46532 44088 46560
rect 28261 46523 28319 46529
rect 44082 46520 44088 46532
rect 44140 46520 44146 46572
rect 44542 46560 44548 46572
rect 44503 46532 44548 46560
rect 44542 46520 44548 46532
rect 44600 46520 44606 46572
rect 47578 46560 47584 46572
rect 47539 46532 47584 46560
rect 47578 46520 47584 46532
rect 47636 46520 47642 46572
rect 3050 46492 3056 46504
rect 2792 46464 3056 46492
rect 3050 46452 3056 46464
rect 3108 46492 3114 46504
rect 14274 46492 14280 46504
rect 3108 46464 14280 46492
rect 3108 46452 3114 46464
rect 14274 46452 14280 46464
rect 14332 46452 14338 46504
rect 19334 46452 19340 46504
rect 19392 46492 19398 46504
rect 19429 46495 19487 46501
rect 19429 46492 19441 46495
rect 19392 46464 19441 46492
rect 19392 46452 19398 46464
rect 19429 46461 19441 46464
rect 19475 46461 19487 46495
rect 19429 46455 19487 46461
rect 19613 46495 19671 46501
rect 19613 46461 19625 46495
rect 19659 46492 19671 46495
rect 19702 46492 19708 46504
rect 19659 46464 19708 46492
rect 19659 46461 19671 46464
rect 19613 46455 19671 46461
rect 19702 46452 19708 46464
rect 19760 46452 19766 46504
rect 45186 46492 45192 46504
rect 45147 46464 45192 46492
rect 45186 46452 45192 46464
rect 45244 46452 45250 46504
rect 45373 46495 45431 46501
rect 45373 46461 45385 46495
rect 45419 46492 45431 46495
rect 46106 46492 46112 46504
rect 45419 46464 46112 46492
rect 45419 46461 45431 46464
rect 45373 46455 45431 46461
rect 46106 46452 46112 46464
rect 46164 46452 46170 46504
rect 4890 46384 4896 46436
rect 4948 46424 4954 46436
rect 4948 46396 22094 46424
rect 4948 46384 4954 46396
rect 1578 46356 1584 46368
rect 1539 46328 1584 46356
rect 1578 46316 1584 46328
rect 1636 46316 1642 46368
rect 2866 46356 2872 46368
rect 2827 46328 2872 46356
rect 2866 46316 2872 46328
rect 2924 46316 2930 46368
rect 7926 46316 7932 46368
rect 7984 46356 7990 46368
rect 8113 46359 8171 46365
rect 8113 46356 8125 46359
rect 7984 46328 8125 46356
rect 7984 46316 7990 46328
rect 8113 46325 8125 46328
rect 8159 46325 8171 46359
rect 22066 46356 22094 46396
rect 26145 46359 26203 46365
rect 26145 46356 26157 46359
rect 22066 46328 26157 46356
rect 8113 46319 8171 46325
rect 26145 46325 26157 46328
rect 26191 46356 26203 46359
rect 28074 46356 28080 46368
rect 26191 46328 28080 46356
rect 26191 46325 26203 46328
rect 26145 46319 26203 46325
rect 28074 46316 28080 46328
rect 28132 46316 28138 46368
rect 1104 46266 48852 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 48852 46266
rect 1104 46192 48852 46214
rect 19702 46152 19708 46164
rect 19663 46124 19708 46152
rect 19702 46112 19708 46124
rect 19760 46112 19766 46164
rect 44174 46112 44180 46164
rect 44232 46152 44238 46164
rect 44361 46155 44419 46161
rect 44361 46152 44373 46155
rect 44232 46124 44373 46152
rect 44232 46112 44238 46124
rect 44361 46121 44373 46124
rect 44407 46121 44419 46155
rect 44361 46115 44419 46121
rect 44910 46112 44916 46164
rect 44968 46152 44974 46164
rect 45189 46155 45247 46161
rect 45189 46152 45201 46155
rect 44968 46124 45201 46152
rect 44968 46112 44974 46124
rect 45189 46121 45201 46124
rect 45235 46121 45247 46155
rect 45189 46115 45247 46121
rect 1581 46019 1639 46025
rect 1581 45985 1593 46019
rect 1627 46016 1639 46019
rect 2866 46016 2872 46028
rect 1627 45988 2872 46016
rect 1627 45985 1639 45988
rect 1581 45979 1639 45985
rect 2866 45976 2872 45988
rect 2924 45976 2930 46028
rect 2958 45976 2964 46028
rect 3016 46016 3022 46028
rect 25406 46016 25412 46028
rect 3016 45988 3061 46016
rect 25367 45988 25412 46016
rect 3016 45976 3022 45988
rect 25406 45976 25412 45988
rect 25464 45976 25470 46028
rect 48130 46016 48136 46028
rect 48091 45988 48136 46016
rect 48130 45976 48136 45988
rect 48188 45976 48194 46028
rect 1397 45951 1455 45957
rect 1397 45917 1409 45951
rect 1443 45917 1455 45951
rect 1397 45911 1455 45917
rect 19613 45951 19671 45957
rect 19613 45917 19625 45951
rect 19659 45948 19671 45951
rect 20070 45948 20076 45960
rect 19659 45920 20076 45948
rect 19659 45917 19671 45920
rect 19613 45911 19671 45917
rect 1412 45880 1440 45911
rect 20070 45908 20076 45920
rect 20128 45908 20134 45960
rect 25222 45948 25228 45960
rect 25183 45920 25228 45948
rect 25222 45908 25228 45920
rect 25280 45908 25286 45960
rect 45646 45948 45652 45960
rect 45607 45920 45652 45948
rect 45646 45908 45652 45920
rect 45704 45908 45710 45960
rect 45830 45908 45836 45960
rect 45888 45948 45894 45960
rect 46293 45951 46351 45957
rect 46293 45948 46305 45951
rect 45888 45920 46305 45948
rect 45888 45908 45894 45920
rect 46293 45917 46305 45920
rect 46339 45917 46351 45951
rect 46293 45911 46351 45917
rect 2866 45880 2872 45892
rect 1412 45852 2872 45880
rect 2866 45840 2872 45852
rect 2924 45840 2930 45892
rect 45741 45883 45799 45889
rect 45741 45849 45753 45883
rect 45787 45880 45799 45883
rect 46477 45883 46535 45889
rect 46477 45880 46489 45883
rect 45787 45852 46489 45880
rect 45787 45849 45799 45852
rect 45741 45843 45799 45849
rect 46477 45849 46489 45852
rect 46523 45849 46535 45883
rect 46477 45843 46535 45849
rect 1104 45722 48852 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 48852 45722
rect 1104 45648 48852 45670
rect 1854 45540 1860 45552
rect 1815 45512 1860 45540
rect 1854 45500 1860 45512
rect 1912 45500 1918 45552
rect 38626 45512 45968 45540
rect 2866 45472 2872 45484
rect 2827 45444 2872 45472
rect 2866 45432 2872 45444
rect 2924 45432 2930 45484
rect 7926 45472 7932 45484
rect 7887 45444 7932 45472
rect 7926 45432 7932 45444
rect 7984 45432 7990 45484
rect 23750 45472 23756 45484
rect 23711 45444 23756 45472
rect 23750 45432 23756 45444
rect 23808 45432 23814 45484
rect 26142 45432 26148 45484
rect 26200 45472 26206 45484
rect 38626 45472 38654 45512
rect 26200 45444 38654 45472
rect 45097 45475 45155 45481
rect 26200 45432 26206 45444
rect 45097 45441 45109 45475
rect 45143 45472 45155 45475
rect 45186 45472 45192 45484
rect 45143 45444 45192 45472
rect 45143 45441 45155 45444
rect 45097 45435 45155 45441
rect 45186 45432 45192 45444
rect 45244 45432 45250 45484
rect 45741 45475 45799 45481
rect 45741 45441 45753 45475
rect 45787 45472 45799 45475
rect 45830 45472 45836 45484
rect 45787 45444 45836 45472
rect 45787 45441 45799 45444
rect 45741 45435 45799 45441
rect 45830 45432 45836 45444
rect 45888 45432 45894 45484
rect 45940 45472 45968 45512
rect 46106 45500 46112 45552
rect 46164 45540 46170 45552
rect 46293 45543 46351 45549
rect 46293 45540 46305 45543
rect 46164 45512 46305 45540
rect 46164 45500 46170 45512
rect 46293 45509 46305 45512
rect 46339 45509 46351 45543
rect 46293 45503 46351 45509
rect 46474 45500 46480 45552
rect 46532 45540 46538 45552
rect 46937 45543 46995 45549
rect 46937 45540 46949 45543
rect 46532 45512 46949 45540
rect 46532 45500 46538 45512
rect 46937 45509 46949 45512
rect 46983 45509 46995 45543
rect 46937 45503 46995 45509
rect 46198 45472 46204 45484
rect 45940 45444 46204 45472
rect 46198 45432 46204 45444
rect 46256 45432 46262 45484
rect 46845 45475 46903 45481
rect 46845 45441 46857 45475
rect 46891 45441 46903 45475
rect 47578 45472 47584 45484
rect 47539 45444 47584 45472
rect 46845 45435 46903 45441
rect 8110 45404 8116 45416
rect 8071 45376 8116 45404
rect 8110 45364 8116 45376
rect 8168 45364 8174 45416
rect 8386 45404 8392 45416
rect 8347 45376 8392 45404
rect 8386 45364 8392 45376
rect 8444 45364 8450 45416
rect 24118 45364 24124 45416
rect 24176 45404 24182 45416
rect 24765 45407 24823 45413
rect 24765 45404 24777 45407
rect 24176 45376 24777 45404
rect 24176 45364 24182 45376
rect 24765 45373 24777 45376
rect 24811 45404 24823 45407
rect 46860 45404 46888 45435
rect 47578 45432 47584 45444
rect 47636 45432 47642 45484
rect 24811 45376 38654 45404
rect 24811 45373 24823 45376
rect 24765 45367 24823 45373
rect 38626 45336 38654 45376
rect 45756 45376 46888 45404
rect 45756 45348 45784 45376
rect 45738 45336 45744 45348
rect 38626 45308 45744 45336
rect 45738 45296 45744 45308
rect 45796 45296 45802 45348
rect 1486 45228 1492 45280
rect 1544 45268 1550 45280
rect 1949 45271 2007 45277
rect 1949 45268 1961 45271
rect 1544 45240 1961 45268
rect 1544 45228 1550 45240
rect 1949 45237 1961 45240
rect 1995 45237 2007 45271
rect 1949 45231 2007 45237
rect 46474 45228 46480 45280
rect 46532 45268 46538 45280
rect 47673 45271 47731 45277
rect 47673 45268 47685 45271
rect 46532 45240 47685 45268
rect 46532 45228 46538 45240
rect 47673 45237 47685 45240
rect 47719 45237 47731 45271
rect 47673 45231 47731 45237
rect 1104 45178 48852 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 48852 45178
rect 1104 45104 48852 45126
rect 8110 45024 8116 45076
rect 8168 45064 8174 45076
rect 9033 45067 9091 45073
rect 9033 45064 9045 45067
rect 8168 45036 9045 45064
rect 8168 45024 8174 45036
rect 9033 45033 9045 45036
rect 9079 45033 9091 45067
rect 9033 45027 9091 45033
rect 45833 45067 45891 45073
rect 45833 45033 45845 45067
rect 45879 45064 45891 45067
rect 46290 45064 46296 45076
rect 45879 45036 46296 45064
rect 45879 45033 45891 45036
rect 45833 45027 45891 45033
rect 46290 45024 46296 45036
rect 46348 45024 46354 45076
rect 15102 44928 15108 44940
rect 6886 44900 15108 44928
rect 2038 44820 2044 44872
rect 2096 44860 2102 44872
rect 2317 44863 2375 44869
rect 2317 44860 2329 44863
rect 2096 44832 2329 44860
rect 2096 44820 2102 44832
rect 2317 44829 2329 44832
rect 2363 44829 2375 44863
rect 2317 44823 2375 44829
rect 2961 44863 3019 44869
rect 2961 44829 2973 44863
rect 3007 44860 3019 44863
rect 6886 44860 6914 44900
rect 15102 44888 15108 44900
rect 15160 44888 15166 44940
rect 22370 44888 22376 44940
rect 22428 44928 22434 44940
rect 23201 44931 23259 44937
rect 23201 44928 23213 44931
rect 22428 44900 23213 44928
rect 22428 44888 22434 44900
rect 23201 44897 23213 44900
rect 23247 44928 23259 44931
rect 30098 44928 30104 44940
rect 23247 44900 30104 44928
rect 23247 44897 23259 44900
rect 23201 44891 23259 44897
rect 30098 44888 30104 44900
rect 30156 44888 30162 44940
rect 46474 44928 46480 44940
rect 46435 44900 46480 44928
rect 46474 44888 46480 44900
rect 46532 44888 46538 44940
rect 48130 44928 48136 44940
rect 48091 44900 48136 44928
rect 48130 44888 48136 44900
rect 48188 44888 48194 44940
rect 8938 44860 8944 44872
rect 3007 44832 6914 44860
rect 8899 44832 8944 44860
rect 3007 44829 3019 44832
rect 2961 44823 3019 44829
rect 8938 44820 8944 44832
rect 8996 44820 9002 44872
rect 23017 44863 23075 44869
rect 23017 44829 23029 44863
rect 23063 44860 23075 44863
rect 46290 44860 46296 44872
rect 23063 44832 23796 44860
rect 46251 44832 46296 44860
rect 23063 44829 23075 44832
rect 23017 44823 23075 44829
rect 23768 44804 23796 44832
rect 46290 44820 46296 44832
rect 46348 44820 46354 44872
rect 6886 44764 12434 44792
rect 2222 44684 2228 44736
rect 2280 44724 2286 44736
rect 3053 44727 3111 44733
rect 3053 44724 3065 44727
rect 2280 44696 3065 44724
rect 2280 44684 2286 44696
rect 3053 44693 3065 44696
rect 3099 44693 3111 44727
rect 3053 44687 3111 44693
rect 3510 44684 3516 44736
rect 3568 44724 3574 44736
rect 6886 44724 6914 44764
rect 3568 44696 6914 44724
rect 12406 44724 12434 44764
rect 23750 44752 23756 44804
rect 23808 44792 23814 44804
rect 24765 44795 24823 44801
rect 24765 44792 24777 44795
rect 23808 44764 24777 44792
rect 23808 44752 23814 44764
rect 24765 44761 24777 44764
rect 24811 44761 24823 44795
rect 24765 44755 24823 44761
rect 25590 44724 25596 44736
rect 12406 44696 25596 44724
rect 3568 44684 3574 44696
rect 25590 44684 25596 44696
rect 25648 44724 25654 44736
rect 26053 44727 26111 44733
rect 26053 44724 26065 44727
rect 25648 44696 26065 44724
rect 25648 44684 25654 44696
rect 26053 44693 26065 44696
rect 26099 44724 26111 44727
rect 38654 44724 38660 44736
rect 26099 44696 38660 44724
rect 26099 44693 26111 44696
rect 26053 44687 26111 44693
rect 38654 44684 38660 44696
rect 38712 44724 38718 44736
rect 38712 44696 38759 44724
rect 38712 44684 38718 44696
rect 1104 44634 48852 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 48852 44634
rect 1104 44560 48852 44582
rect 2222 44452 2228 44464
rect 2183 44424 2228 44452
rect 2222 44412 2228 44424
rect 2280 44412 2286 44464
rect 2038 44384 2044 44396
rect 1999 44356 2044 44384
rect 2038 44344 2044 44356
rect 2096 44344 2102 44396
rect 23750 44384 23756 44396
rect 23711 44356 23756 44384
rect 23750 44344 23756 44356
rect 23808 44344 23814 44396
rect 46290 44344 46296 44396
rect 46348 44384 46354 44396
rect 47765 44387 47823 44393
rect 47765 44384 47777 44387
rect 46348 44356 47777 44384
rect 46348 44344 46354 44356
rect 47765 44353 47777 44356
rect 47811 44353 47823 44387
rect 47765 44347 47823 44353
rect 2774 44316 2780 44328
rect 2735 44288 2780 44316
rect 2774 44276 2780 44288
rect 2832 44276 2838 44328
rect 23842 44276 23848 44328
rect 23900 44316 23906 44328
rect 24762 44316 24768 44328
rect 23900 44288 24768 44316
rect 23900 44276 23906 44288
rect 24762 44276 24768 44288
rect 24820 44276 24826 44328
rect 47026 44180 47032 44192
rect 46987 44152 47032 44180
rect 47026 44140 47032 44152
rect 47084 44140 47090 44192
rect 1104 44090 48852 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 48852 44090
rect 1104 44016 48852 44038
rect 8938 43868 8944 43920
rect 8996 43908 9002 43920
rect 8996 43880 25084 43908
rect 8996 43868 9002 43880
rect 15102 43800 15108 43852
rect 15160 43840 15166 43852
rect 25056 43849 25084 43880
rect 20257 43843 20315 43849
rect 20257 43840 20269 43843
rect 15160 43812 20269 43840
rect 15160 43800 15166 43812
rect 20257 43809 20269 43812
rect 20303 43840 20315 43843
rect 25041 43843 25099 43849
rect 20303 43812 24992 43840
rect 20303 43809 20315 43812
rect 20257 43803 20315 43809
rect 1854 43772 1860 43784
rect 1815 43744 1860 43772
rect 1854 43732 1860 43744
rect 1912 43732 1918 43784
rect 20073 43775 20131 43781
rect 20073 43741 20085 43775
rect 20119 43772 20131 43775
rect 20162 43772 20168 43784
rect 20119 43744 20168 43772
rect 20119 43741 20131 43744
rect 20073 43735 20131 43741
rect 20162 43732 20168 43744
rect 20220 43732 20226 43784
rect 23750 43732 23756 43784
rect 23808 43772 23814 43784
rect 23845 43775 23903 43781
rect 23845 43772 23857 43775
rect 23808 43744 23857 43772
rect 23808 43732 23814 43744
rect 23845 43741 23857 43744
rect 23891 43772 23903 43775
rect 24489 43775 24547 43781
rect 24489 43772 24501 43775
rect 23891 43744 24501 43772
rect 23891 43741 23903 43744
rect 23845 43735 23903 43741
rect 24489 43741 24501 43744
rect 24535 43741 24547 43775
rect 24964 43772 24992 43812
rect 25041 43809 25053 43843
rect 25087 43840 25099 43843
rect 46293 43843 46351 43849
rect 25087 43812 35894 43840
rect 25087 43809 25099 43812
rect 25041 43803 25099 43809
rect 26878 43772 26884 43784
rect 24964 43744 26884 43772
rect 24489 43735 24547 43741
rect 26878 43732 26884 43744
rect 26936 43732 26942 43784
rect 2225 43707 2283 43713
rect 2225 43673 2237 43707
rect 2271 43704 2283 43707
rect 2314 43704 2320 43716
rect 2271 43676 2320 43704
rect 2271 43673 2283 43676
rect 2225 43667 2283 43673
rect 2314 43664 2320 43676
rect 2372 43664 2378 43716
rect 23477 43707 23535 43713
rect 23477 43673 23489 43707
rect 23523 43704 23535 43707
rect 23566 43704 23572 43716
rect 23523 43676 23572 43704
rect 23523 43673 23535 43676
rect 23477 43667 23535 43673
rect 23566 43664 23572 43676
rect 23624 43704 23630 43716
rect 24946 43704 24952 43716
rect 23624 43676 24952 43704
rect 23624 43664 23630 43676
rect 24946 43664 24952 43676
rect 25004 43664 25010 43716
rect 35866 43704 35894 43812
rect 46293 43809 46305 43843
rect 46339 43840 46351 43843
rect 47026 43840 47032 43852
rect 46339 43812 47032 43840
rect 46339 43809 46351 43812
rect 46293 43803 46351 43809
rect 47026 43800 47032 43812
rect 47084 43800 47090 43852
rect 45830 43704 45836 43716
rect 35866 43676 45836 43704
rect 45830 43664 45836 43676
rect 45888 43664 45894 43716
rect 46477 43707 46535 43713
rect 46477 43673 46489 43707
rect 46523 43704 46535 43707
rect 46934 43704 46940 43716
rect 46523 43676 46940 43704
rect 46523 43673 46535 43676
rect 46477 43667 46535 43673
rect 46934 43664 46940 43676
rect 46992 43664 46998 43716
rect 48130 43704 48136 43716
rect 48091 43676 48136 43704
rect 48130 43664 48136 43676
rect 48188 43664 48194 43716
rect 1104 43546 48852 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 48852 43546
rect 1104 43472 48852 43494
rect 27341 43435 27399 43441
rect 27341 43401 27353 43435
rect 27387 43432 27399 43435
rect 28810 43432 28816 43444
rect 27387 43404 28816 43432
rect 27387 43401 27399 43404
rect 27341 43395 27399 43401
rect 28810 43392 28816 43404
rect 28868 43392 28874 43444
rect 46934 43432 46940 43444
rect 46895 43404 46940 43432
rect 46934 43392 46940 43404
rect 46992 43392 46998 43444
rect 1854 43364 1860 43376
rect 1815 43336 1860 43364
rect 1854 43324 1860 43336
rect 1912 43324 1918 43376
rect 20530 43364 20536 43376
rect 6886 43336 20536 43364
rect 2130 43188 2136 43240
rect 2188 43228 2194 43240
rect 6886 43228 6914 43336
rect 20530 43324 20536 43336
rect 20588 43364 20594 43376
rect 20588 43336 31754 43364
rect 20588 43324 20594 43336
rect 20162 43296 20168 43308
rect 20123 43268 20168 43296
rect 20162 43256 20168 43268
rect 20220 43256 20226 43308
rect 21913 43299 21971 43305
rect 21913 43265 21925 43299
rect 21959 43296 21971 43299
rect 22002 43296 22008 43308
rect 21959 43268 22008 43296
rect 21959 43265 21971 43268
rect 21913 43259 21971 43265
rect 22002 43256 22008 43268
rect 22060 43256 22066 43308
rect 22097 43299 22155 43305
rect 22097 43265 22109 43299
rect 22143 43296 22155 43299
rect 22738 43296 22744 43308
rect 22143 43268 22744 43296
rect 22143 43265 22155 43268
rect 22097 43259 22155 43265
rect 22738 43256 22744 43268
rect 22796 43256 22802 43308
rect 24670 43296 24676 43308
rect 24631 43268 24676 43296
rect 24670 43256 24676 43268
rect 24728 43256 24734 43308
rect 24765 43299 24823 43305
rect 24765 43265 24777 43299
rect 24811 43265 24823 43299
rect 24765 43259 24823 43265
rect 2188 43200 6914 43228
rect 2188 43188 2194 43200
rect 24578 43188 24584 43240
rect 24636 43228 24642 43240
rect 24780 43228 24808 43259
rect 24854 43256 24860 43308
rect 24912 43296 24918 43308
rect 24912 43268 24957 43296
rect 24912 43256 24918 43268
rect 25038 43256 25044 43308
rect 25096 43296 25102 43308
rect 27154 43296 27160 43308
rect 25096 43268 25141 43296
rect 27115 43268 27160 43296
rect 25096 43256 25102 43268
rect 27154 43256 27160 43268
rect 27212 43256 27218 43308
rect 27430 43256 27436 43308
rect 27488 43296 27494 43308
rect 27488 43268 27533 43296
rect 27488 43256 27494 43268
rect 24636 43200 24808 43228
rect 31726 43228 31754 43336
rect 45830 43256 45836 43308
rect 45888 43296 45894 43308
rect 46845 43299 46903 43305
rect 46845 43296 46857 43299
rect 45888 43268 46857 43296
rect 45888 43256 45894 43268
rect 46845 43265 46857 43268
rect 46891 43265 46903 43299
rect 47854 43296 47860 43308
rect 47815 43268 47860 43296
rect 46845 43259 46903 43265
rect 47854 43256 47860 43268
rect 47912 43256 47918 43308
rect 40310 43228 40316 43240
rect 31726 43200 40316 43228
rect 24636 43188 24642 43200
rect 40310 43188 40316 43200
rect 40368 43188 40374 43240
rect 2133 43095 2191 43101
rect 2133 43061 2145 43095
rect 2179 43092 2191 43095
rect 2406 43092 2412 43104
rect 2179 43064 2412 43092
rect 2179 43061 2191 43064
rect 2133 43055 2191 43061
rect 2406 43052 2412 43064
rect 2464 43052 2470 43104
rect 22278 43092 22284 43104
rect 22239 43064 22284 43092
rect 22278 43052 22284 43064
rect 22336 43052 22342 43104
rect 24397 43095 24455 43101
rect 24397 43061 24409 43095
rect 24443 43092 24455 43095
rect 24946 43092 24952 43104
rect 24443 43064 24952 43092
rect 24443 43061 24455 43064
rect 24397 43055 24455 43061
rect 24946 43052 24952 43064
rect 25004 43052 25010 43104
rect 26970 43092 26976 43104
rect 26931 43064 26976 43092
rect 26970 43052 26976 43064
rect 27028 43052 27034 43104
rect 47210 43052 47216 43104
rect 47268 43092 47274 43104
rect 48041 43095 48099 43101
rect 48041 43092 48053 43095
rect 47268 43064 48053 43092
rect 47268 43052 47274 43064
rect 48041 43061 48053 43064
rect 48087 43061 48099 43095
rect 48041 43055 48099 43061
rect 1104 43002 48852 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 48852 43002
rect 1104 42928 48852 42950
rect 29086 42752 29092 42764
rect 28644 42724 29092 42752
rect 19797 42687 19855 42693
rect 19797 42653 19809 42687
rect 19843 42684 19855 42687
rect 20162 42684 20168 42696
rect 19843 42656 20168 42684
rect 19843 42653 19855 42656
rect 19797 42647 19855 42653
rect 20162 42644 20168 42656
rect 20220 42644 20226 42696
rect 21358 42684 21364 42696
rect 21319 42656 21364 42684
rect 21358 42644 21364 42656
rect 21416 42644 21422 42696
rect 24026 42644 24032 42696
rect 24084 42684 24090 42696
rect 24946 42693 24952 42696
rect 24673 42687 24731 42693
rect 24673 42684 24685 42687
rect 24084 42656 24685 42684
rect 24084 42644 24090 42656
rect 24673 42653 24685 42656
rect 24719 42653 24731 42687
rect 24940 42684 24952 42693
rect 24907 42656 24952 42684
rect 24673 42647 24731 42653
rect 24940 42647 24952 42656
rect 24946 42644 24952 42647
rect 25004 42644 25010 42696
rect 25682 42644 25688 42696
rect 25740 42684 25746 42696
rect 26743 42687 26801 42693
rect 26743 42684 26755 42687
rect 25740 42656 26755 42684
rect 25740 42644 25746 42656
rect 26743 42653 26755 42656
rect 26789 42653 26801 42687
rect 26878 42684 26884 42696
rect 26839 42656 26884 42684
rect 26743 42647 26801 42653
rect 26878 42644 26884 42656
rect 26936 42644 26942 42696
rect 26970 42644 26976 42696
rect 27028 42684 27034 42696
rect 27157 42687 27215 42693
rect 27028 42656 27073 42684
rect 27028 42644 27034 42656
rect 27157 42653 27169 42687
rect 27203 42684 27215 42687
rect 27522 42684 27528 42696
rect 27203 42656 27528 42684
rect 27203 42653 27215 42656
rect 27157 42647 27215 42653
rect 27522 42644 27528 42656
rect 27580 42684 27586 42696
rect 27982 42684 27988 42696
rect 27580 42656 27988 42684
rect 27580 42644 27586 42656
rect 27982 42644 27988 42656
rect 28040 42644 28046 42696
rect 28644 42693 28672 42724
rect 29086 42712 29092 42724
rect 29144 42712 29150 42764
rect 28629 42687 28687 42693
rect 28629 42653 28641 42687
rect 28675 42653 28687 42687
rect 28810 42684 28816 42696
rect 28771 42656 28816 42684
rect 28629 42647 28687 42653
rect 28810 42644 28816 42656
rect 28868 42644 28874 42696
rect 28905 42687 28963 42693
rect 28905 42653 28917 42687
rect 28951 42684 28963 42687
rect 29362 42684 29368 42696
rect 28951 42656 29368 42684
rect 28951 42653 28963 42656
rect 28905 42647 28963 42653
rect 29362 42644 29368 42656
rect 29420 42644 29426 42696
rect 29546 42684 29552 42696
rect 29507 42656 29552 42684
rect 29546 42644 29552 42656
rect 29604 42644 29610 42696
rect 20070 42616 20076 42628
rect 20031 42588 20076 42616
rect 20070 42576 20076 42588
rect 20128 42576 20134 42628
rect 21628 42619 21686 42625
rect 21628 42585 21640 42619
rect 21674 42616 21686 42619
rect 21818 42616 21824 42628
rect 21674 42588 21824 42616
rect 21674 42585 21686 42588
rect 21628 42579 21686 42585
rect 21818 42576 21824 42588
rect 21876 42576 21882 42628
rect 23382 42576 23388 42628
rect 23440 42616 23446 42628
rect 23477 42619 23535 42625
rect 23477 42616 23489 42619
rect 23440 42588 23489 42616
rect 23440 42576 23446 42588
rect 23477 42585 23489 42588
rect 23523 42585 23535 42619
rect 23477 42579 23535 42585
rect 23661 42619 23719 42625
rect 23661 42585 23673 42619
rect 23707 42585 23719 42619
rect 23661 42579 23719 42585
rect 23845 42619 23903 42625
rect 23845 42585 23857 42619
rect 23891 42616 23903 42619
rect 24854 42616 24860 42628
rect 23891 42588 24860 42616
rect 23891 42585 23903 42588
rect 23845 42579 23903 42585
rect 22738 42548 22744 42560
rect 22699 42520 22744 42548
rect 22738 42508 22744 42520
rect 22796 42508 22802 42560
rect 23676 42548 23704 42579
rect 24854 42576 24860 42588
rect 24912 42576 24918 42628
rect 27890 42576 27896 42628
rect 27948 42616 27954 42628
rect 29794 42619 29852 42625
rect 29794 42616 29806 42619
rect 27948 42588 29806 42616
rect 27948 42576 27954 42588
rect 29794 42585 29806 42588
rect 29840 42585 29852 42619
rect 47946 42616 47952 42628
rect 47907 42588 47952 42616
rect 29794 42579 29852 42585
rect 47946 42576 47952 42588
rect 48004 42576 48010 42628
rect 26053 42551 26111 42557
rect 26053 42548 26065 42551
rect 23676 42520 26065 42548
rect 26053 42517 26065 42520
rect 26099 42548 26111 42551
rect 26142 42548 26148 42560
rect 26099 42520 26148 42548
rect 26099 42517 26111 42520
rect 26053 42511 26111 42517
rect 26142 42508 26148 42520
rect 26200 42508 26206 42560
rect 26510 42548 26516 42560
rect 26471 42520 26516 42548
rect 26510 42508 26516 42520
rect 26568 42508 26574 42560
rect 27798 42508 27804 42560
rect 27856 42548 27862 42560
rect 28445 42551 28503 42557
rect 28445 42548 28457 42551
rect 27856 42520 28457 42548
rect 27856 42508 27862 42520
rect 28445 42517 28457 42520
rect 28491 42517 28503 42551
rect 28445 42511 28503 42517
rect 30190 42508 30196 42560
rect 30248 42548 30254 42560
rect 30929 42551 30987 42557
rect 30929 42548 30941 42551
rect 30248 42520 30941 42548
rect 30248 42508 30254 42520
rect 30929 42517 30941 42520
rect 30975 42517 30987 42551
rect 48038 42548 48044 42560
rect 47999 42520 48044 42548
rect 30929 42511 30987 42517
rect 48038 42508 48044 42520
rect 48096 42508 48102 42560
rect 1104 42458 48852 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 48852 42458
rect 1104 42384 48852 42406
rect 5442 42304 5448 42356
rect 5500 42344 5506 42356
rect 21818 42344 21824 42356
rect 5500 42316 6914 42344
rect 21779 42316 21824 42344
rect 5500 42304 5506 42316
rect 6886 42276 6914 42316
rect 21818 42304 21824 42316
rect 21876 42304 21882 42356
rect 22094 42304 22100 42356
rect 22152 42344 22158 42356
rect 23382 42344 23388 42356
rect 22152 42316 23388 42344
rect 22152 42304 22158 42316
rect 23382 42304 23388 42316
rect 23440 42344 23446 42356
rect 25682 42344 25688 42356
rect 23440 42316 23520 42344
rect 23440 42304 23446 42316
rect 23492 42285 23520 42316
rect 23676 42316 25688 42344
rect 23676 42285 23704 42316
rect 25682 42304 25688 42316
rect 25740 42304 25746 42356
rect 29178 42344 29184 42356
rect 27264 42316 29184 42344
rect 23477 42279 23535 42285
rect 6886 42248 22140 42276
rect 15565 42211 15623 42217
rect 15565 42177 15577 42211
rect 15611 42208 15623 42211
rect 21726 42208 21732 42220
rect 15611 42180 21732 42208
rect 15611 42177 15623 42180
rect 15565 42171 15623 42177
rect 21726 42168 21732 42180
rect 21784 42168 21790 42220
rect 22112 42217 22140 42248
rect 23477 42245 23489 42279
rect 23523 42245 23535 42279
rect 23477 42239 23535 42245
rect 23661 42279 23719 42285
rect 23661 42245 23673 42279
rect 23707 42245 23719 42279
rect 23661 42239 23719 42245
rect 23842 42236 23848 42288
rect 23900 42276 23906 42288
rect 24550 42279 24608 42285
rect 24550 42276 24562 42279
rect 23900 42248 24562 42276
rect 23900 42236 23906 42248
rect 24550 42245 24562 42248
rect 24596 42245 24608 42279
rect 24550 42239 24608 42245
rect 24670 42236 24676 42288
rect 24728 42276 24734 42288
rect 27264 42276 27292 42316
rect 29178 42304 29184 42316
rect 29236 42304 29242 42356
rect 29362 42304 29368 42356
rect 29420 42344 29426 42356
rect 29638 42344 29644 42356
rect 29420 42316 29644 42344
rect 29420 42304 29426 42316
rect 29638 42304 29644 42316
rect 29696 42344 29702 42356
rect 29825 42347 29883 42353
rect 29825 42344 29837 42347
rect 29696 42316 29837 42344
rect 29696 42304 29702 42316
rect 29825 42313 29837 42316
rect 29871 42313 29883 42347
rect 29825 42307 29883 42313
rect 29914 42304 29920 42356
rect 29972 42344 29978 42356
rect 30653 42347 30711 42353
rect 30653 42344 30665 42347
rect 29972 42316 30665 42344
rect 29972 42304 29978 42316
rect 30653 42313 30665 42316
rect 30699 42313 30711 42347
rect 30653 42307 30711 42313
rect 30834 42304 30840 42356
rect 30892 42344 30898 42356
rect 48038 42344 48044 42356
rect 30892 42316 48044 42344
rect 30892 42304 30898 42316
rect 48038 42304 48044 42316
rect 48096 42304 48102 42356
rect 24728 42248 27292 42276
rect 27341 42279 27399 42285
rect 24728 42236 24734 42248
rect 27341 42245 27353 42279
rect 27387 42276 27399 42279
rect 28690 42279 28748 42285
rect 28690 42276 28702 42279
rect 27387 42248 28702 42276
rect 27387 42245 27399 42248
rect 27341 42239 27399 42245
rect 28690 42245 28702 42248
rect 28736 42245 28748 42279
rect 28690 42239 28748 42245
rect 28810 42236 28816 42288
rect 28868 42236 28874 42288
rect 22097 42211 22155 42217
rect 22097 42177 22109 42211
rect 22143 42177 22155 42211
rect 22097 42171 22155 42177
rect 22189 42211 22247 42217
rect 22189 42177 22201 42211
rect 22235 42177 22247 42211
rect 22189 42171 22247 42177
rect 21450 42100 21456 42152
rect 21508 42140 21514 42152
rect 22204 42140 22232 42171
rect 22278 42168 22284 42220
rect 22336 42208 22342 42220
rect 22465 42211 22523 42217
rect 22336 42180 22381 42208
rect 22336 42168 22342 42180
rect 22465 42177 22477 42211
rect 22511 42208 22523 42211
rect 23934 42208 23940 42220
rect 22511 42180 23940 42208
rect 22511 42177 22523 42180
rect 22465 42171 22523 42177
rect 23934 42168 23940 42180
rect 23992 42168 23998 42220
rect 24026 42168 24032 42220
rect 24084 42208 24090 42220
rect 24305 42211 24363 42217
rect 24305 42208 24317 42211
rect 24084 42180 24317 42208
rect 24084 42168 24090 42180
rect 24305 42177 24317 42180
rect 24351 42177 24363 42211
rect 27617 42211 27675 42217
rect 27617 42208 27629 42211
rect 24305 42171 24363 42177
rect 24412 42180 27629 42208
rect 23658 42140 23664 42152
rect 21508 42112 23664 42140
rect 21508 42100 21514 42112
rect 23658 42100 23664 42112
rect 23716 42100 23722 42152
rect 24412 42140 24440 42180
rect 27617 42177 27629 42180
rect 27663 42177 27675 42211
rect 27617 42171 27675 42177
rect 27709 42211 27767 42217
rect 27709 42177 27721 42211
rect 27755 42177 27767 42211
rect 27709 42171 27767 42177
rect 24320 42112 24440 42140
rect 22738 42032 22744 42084
rect 22796 42072 22802 42084
rect 24320 42072 24348 42112
rect 27724 42084 27752 42171
rect 27798 42168 27804 42220
rect 27856 42208 27862 42220
rect 27856 42180 27901 42208
rect 27856 42168 27862 42180
rect 27982 42168 27988 42220
rect 28040 42208 28046 42220
rect 28828 42208 28856 42236
rect 29914 42208 29920 42220
rect 28040 42180 28085 42208
rect 28828 42180 29920 42208
rect 28040 42168 28046 42180
rect 29914 42168 29920 42180
rect 29972 42168 29978 42220
rect 30469 42211 30527 42217
rect 30469 42208 30481 42211
rect 30024 42180 30481 42208
rect 28445 42143 28503 42149
rect 28445 42109 28457 42143
rect 28491 42109 28503 42143
rect 28445 42103 28503 42109
rect 22796 42044 24348 42072
rect 22796 42032 22802 42044
rect 27706 42032 27712 42084
rect 27764 42032 27770 42084
rect 1394 41964 1400 42016
rect 1452 42004 1458 42016
rect 2041 42007 2099 42013
rect 2041 42004 2053 42007
rect 1452 41976 2053 42004
rect 1452 41964 1458 41976
rect 2041 41973 2053 41976
rect 2087 41973 2099 42007
rect 2041 41967 2099 41973
rect 15657 42007 15715 42013
rect 15657 41973 15669 42007
rect 15703 42004 15715 42007
rect 15746 42004 15752 42016
rect 15703 41976 15752 42004
rect 15703 41973 15715 41976
rect 15657 41967 15715 41973
rect 15746 41964 15752 41976
rect 15804 41964 15810 42016
rect 23845 42007 23903 42013
rect 23845 41973 23857 42007
rect 23891 42004 23903 42007
rect 24946 42004 24952 42016
rect 23891 41976 24952 42004
rect 23891 41973 23903 41976
rect 23845 41967 23903 41973
rect 24946 41964 24952 41976
rect 25004 41964 25010 42016
rect 25958 41964 25964 42016
rect 26016 42004 26022 42016
rect 28460 42004 28488 42103
rect 26016 41976 28488 42004
rect 26016 41964 26022 41976
rect 29086 41964 29092 42016
rect 29144 42004 29150 42016
rect 30024 42004 30052 42180
rect 30469 42177 30481 42180
rect 30515 42177 30527 42211
rect 30469 42171 30527 42177
rect 30745 42211 30803 42217
rect 30745 42177 30757 42211
rect 30791 42177 30803 42211
rect 30745 42171 30803 42177
rect 30190 42100 30196 42152
rect 30248 42140 30254 42152
rect 30760 42140 30788 42171
rect 30248 42112 30788 42140
rect 30248 42100 30254 42112
rect 30282 42004 30288 42016
rect 29144 41976 30052 42004
rect 30243 41976 30288 42004
rect 29144 41964 29150 41976
rect 30282 41964 30288 41976
rect 30340 41964 30346 42016
rect 46290 41964 46296 42016
rect 46348 42004 46354 42016
rect 47765 42007 47823 42013
rect 47765 42004 47777 42007
rect 46348 41976 47777 42004
rect 46348 41964 46354 41976
rect 47765 41973 47777 41976
rect 47811 41973 47823 42007
rect 47765 41967 47823 41973
rect 1104 41914 48852 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 48852 41914
rect 1104 41840 48852 41862
rect 23842 41760 23848 41812
rect 23900 41800 23906 41812
rect 24397 41803 24455 41809
rect 24397 41800 24409 41803
rect 23900 41772 24409 41800
rect 23900 41760 23906 41772
rect 24397 41769 24409 41772
rect 24443 41769 24455 41803
rect 24397 41763 24455 41769
rect 26142 41760 26148 41812
rect 26200 41800 26206 41812
rect 27341 41803 27399 41809
rect 26200 41772 27016 41800
rect 26200 41760 26206 41772
rect 24026 41692 24032 41744
rect 24084 41732 24090 41744
rect 24762 41732 24768 41744
rect 24084 41704 24768 41732
rect 24084 41692 24090 41704
rect 24762 41692 24768 41704
rect 24820 41692 24826 41744
rect 1394 41664 1400 41676
rect 1355 41636 1400 41664
rect 1394 41624 1400 41636
rect 1452 41624 1458 41676
rect 1854 41664 1860 41676
rect 1815 41636 1860 41664
rect 1854 41624 1860 41636
rect 1912 41624 1918 41676
rect 15746 41664 15752 41676
rect 15707 41636 15752 41664
rect 15746 41624 15752 41636
rect 15804 41624 15810 41676
rect 16574 41664 16580 41676
rect 16535 41636 16580 41664
rect 16574 41624 16580 41636
rect 16632 41624 16638 41676
rect 24780 41664 24808 41692
rect 25958 41664 25964 41676
rect 24780 41636 25964 41664
rect 25958 41624 25964 41636
rect 26016 41624 26022 41676
rect 15562 41596 15568 41608
rect 15523 41568 15568 41596
rect 15562 41556 15568 41568
rect 15620 41556 15626 41608
rect 20533 41599 20591 41605
rect 20533 41565 20545 41599
rect 20579 41596 20591 41599
rect 20622 41596 20628 41608
rect 20579 41568 20628 41596
rect 20579 41565 20591 41568
rect 20533 41559 20591 41565
rect 20622 41556 20628 41568
rect 20680 41596 20686 41608
rect 21358 41596 21364 41608
rect 20680 41568 21364 41596
rect 20680 41556 20686 41568
rect 21358 41556 21364 41568
rect 21416 41596 21422 41608
rect 22465 41599 22523 41605
rect 22465 41596 22477 41599
rect 21416 41568 22477 41596
rect 21416 41556 21422 41568
rect 22465 41565 22477 41568
rect 22511 41565 22523 41599
rect 22465 41559 22523 41565
rect 24026 41556 24032 41608
rect 24084 41596 24090 41608
rect 24673 41599 24731 41605
rect 24673 41596 24685 41599
rect 24084 41568 24685 41596
rect 24084 41556 24090 41568
rect 24673 41565 24685 41568
rect 24719 41565 24731 41599
rect 24673 41559 24731 41565
rect 24765 41599 24823 41605
rect 24765 41565 24777 41599
rect 24811 41565 24823 41599
rect 24765 41559 24823 41565
rect 24857 41599 24915 41605
rect 24857 41565 24869 41599
rect 24903 41596 24915 41599
rect 24946 41596 24952 41608
rect 24903 41568 24952 41596
rect 24903 41565 24915 41568
rect 24857 41559 24915 41565
rect 1581 41531 1639 41537
rect 1581 41497 1593 41531
rect 1627 41528 1639 41531
rect 2590 41528 2596 41540
rect 1627 41500 2596 41528
rect 1627 41497 1639 41500
rect 1581 41491 1639 41497
rect 2590 41488 2596 41500
rect 2648 41488 2654 41540
rect 20800 41531 20858 41537
rect 20800 41497 20812 41531
rect 20846 41528 20858 41531
rect 20898 41528 20904 41540
rect 20846 41500 20904 41528
rect 20846 41497 20858 41500
rect 20800 41491 20858 41497
rect 20898 41488 20904 41500
rect 20956 41488 20962 41540
rect 22738 41537 22744 41540
rect 22732 41491 22744 41537
rect 22796 41528 22802 41540
rect 22796 41500 22832 41528
rect 22738 41488 22744 41491
rect 22796 41488 22802 41500
rect 23658 41488 23664 41540
rect 23716 41528 23722 41540
rect 24578 41528 24584 41540
rect 23716 41500 24584 41528
rect 23716 41488 23722 41500
rect 24578 41488 24584 41500
rect 24636 41528 24642 41540
rect 24780 41528 24808 41559
rect 24946 41556 24952 41568
rect 25004 41556 25010 41608
rect 25038 41556 25044 41608
rect 25096 41596 25102 41608
rect 26228 41599 26286 41605
rect 25096 41568 25141 41596
rect 25096 41556 25102 41568
rect 26228 41565 26240 41599
rect 26274 41596 26286 41599
rect 26510 41596 26516 41608
rect 26274 41568 26516 41596
rect 26274 41565 26286 41568
rect 26228 41559 26286 41565
rect 26510 41556 26516 41568
rect 26568 41556 26574 41608
rect 26988 41596 27016 41772
rect 27341 41769 27353 41803
rect 27387 41800 27399 41803
rect 27430 41800 27436 41812
rect 27387 41772 27436 41800
rect 27387 41769 27399 41772
rect 27341 41763 27399 41769
rect 27430 41760 27436 41772
rect 27488 41760 27494 41812
rect 27890 41800 27896 41812
rect 27851 41772 27896 41800
rect 27890 41760 27896 41772
rect 27948 41760 27954 41812
rect 30282 41800 30288 41812
rect 28368 41772 30288 41800
rect 27706 41624 27712 41676
rect 27764 41664 27770 41676
rect 27764 41636 28304 41664
rect 27764 41624 27770 41636
rect 28276 41605 28304 41636
rect 28368 41605 28396 41772
rect 30282 41760 30288 41772
rect 30340 41760 30346 41812
rect 29546 41664 29552 41676
rect 29507 41636 29552 41664
rect 29546 41624 29552 41636
rect 29604 41624 29610 41676
rect 46290 41664 46296 41676
rect 46251 41636 46296 41664
rect 46290 41624 46296 41636
rect 46348 41624 46354 41676
rect 28169 41599 28227 41605
rect 28169 41596 28181 41599
rect 26988 41568 28181 41596
rect 28169 41565 28181 41568
rect 28215 41565 28227 41599
rect 28169 41559 28227 41565
rect 28261 41599 28319 41605
rect 28261 41565 28273 41599
rect 28307 41565 28319 41599
rect 28261 41559 28319 41565
rect 28353 41599 28411 41605
rect 28353 41565 28365 41599
rect 28399 41565 28411 41599
rect 28353 41559 28411 41565
rect 28537 41599 28595 41605
rect 28537 41565 28549 41599
rect 28583 41565 28595 41599
rect 48130 41596 48136 41608
rect 48091 41568 48136 41596
rect 28537 41559 28595 41565
rect 24636 41500 24808 41528
rect 24636 41488 24642 41500
rect 21913 41463 21971 41469
rect 21913 41429 21925 41463
rect 21959 41460 21971 41463
rect 22002 41460 22008 41472
rect 21959 41432 22008 41460
rect 21959 41429 21971 41432
rect 21913 41423 21971 41429
rect 22002 41420 22008 41432
rect 22060 41460 22066 41472
rect 23198 41460 23204 41472
rect 22060 41432 23204 41460
rect 22060 41420 22066 41432
rect 23198 41420 23204 41432
rect 23256 41420 23262 41472
rect 23842 41460 23848 41472
rect 23803 41432 23848 41460
rect 23842 41420 23848 41432
rect 23900 41420 23906 41472
rect 23934 41420 23940 41472
rect 23992 41460 23998 41472
rect 25056 41460 25084 41556
rect 27522 41488 27528 41540
rect 27580 41528 27586 41540
rect 28552 41528 28580 41559
rect 48130 41556 48136 41568
rect 48188 41556 48194 41608
rect 27580 41500 28580 41528
rect 27580 41488 27586 41500
rect 28994 41488 29000 41540
rect 29052 41528 29058 41540
rect 29794 41531 29852 41537
rect 29794 41528 29806 41531
rect 29052 41500 29806 41528
rect 29052 41488 29058 41500
rect 29794 41497 29806 41500
rect 29840 41497 29852 41531
rect 46474 41528 46480 41540
rect 46435 41500 46480 41528
rect 29794 41491 29852 41497
rect 46474 41488 46480 41500
rect 46532 41488 46538 41540
rect 23992 41432 25084 41460
rect 23992 41420 23998 41432
rect 26510 41420 26516 41472
rect 26568 41460 26574 41472
rect 27154 41460 27160 41472
rect 26568 41432 27160 41460
rect 26568 41420 26574 41432
rect 27154 41420 27160 41432
rect 27212 41460 27218 41472
rect 29086 41460 29092 41472
rect 27212 41432 29092 41460
rect 27212 41420 27218 41432
rect 29086 41420 29092 41432
rect 29144 41420 29150 41472
rect 30926 41460 30932 41472
rect 30839 41432 30932 41460
rect 30926 41420 30932 41432
rect 30984 41460 30990 41472
rect 33318 41460 33324 41472
rect 30984 41432 33324 41460
rect 30984 41420 30990 41432
rect 33318 41420 33324 41432
rect 33376 41420 33382 41472
rect 1104 41370 48852 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 48852 41370
rect 1104 41296 48852 41318
rect 2590 41256 2596 41268
rect 2551 41228 2596 41256
rect 2590 41216 2596 41228
rect 2648 41216 2654 41268
rect 22649 41259 22707 41265
rect 6886 41228 22600 41256
rect 1854 41120 1860 41132
rect 1815 41092 1860 41120
rect 1854 41080 1860 41092
rect 1912 41080 1918 41132
rect 2130 41080 2136 41132
rect 2188 41120 2194 41132
rect 2501 41123 2559 41129
rect 2501 41120 2513 41123
rect 2188 41092 2513 41120
rect 2188 41080 2194 41092
rect 2501 41089 2513 41092
rect 2547 41120 2559 41123
rect 6886 41120 6914 41228
rect 15194 41188 15200 41200
rect 14752 41160 15200 41188
rect 14752 41129 14780 41160
rect 15194 41148 15200 41160
rect 15252 41148 15258 41200
rect 22189 41191 22247 41197
rect 22189 41188 22201 41191
rect 21008 41160 22201 41188
rect 15010 41129 15016 41132
rect 2547 41092 6914 41120
rect 14737 41123 14795 41129
rect 2547 41089 2559 41092
rect 2501 41083 2559 41089
rect 14737 41089 14749 41123
rect 14783 41089 14795 41123
rect 14737 41083 14795 41089
rect 15004 41083 15016 41129
rect 15068 41120 15074 41132
rect 20806 41120 20812 41132
rect 15068 41092 15104 41120
rect 20767 41092 20812 41120
rect 15010 41080 15016 41083
rect 15068 41080 15074 41092
rect 20806 41080 20812 41092
rect 20864 41080 20870 41132
rect 21008 41129 21036 41160
rect 22189 41157 22201 41160
rect 22235 41157 22247 41191
rect 22572 41188 22600 41228
rect 22649 41225 22661 41259
rect 22695 41256 22707 41259
rect 22738 41256 22744 41268
rect 22695 41228 22744 41256
rect 22695 41225 22707 41228
rect 22649 41219 22707 41225
rect 22738 41216 22744 41228
rect 22796 41216 22802 41268
rect 24210 41256 24216 41268
rect 22848 41228 24216 41256
rect 22848 41188 22876 41228
rect 24210 41216 24216 41228
rect 24268 41216 24274 41268
rect 27709 41259 27767 41265
rect 27709 41225 27721 41259
rect 27755 41256 27767 41259
rect 28994 41256 29000 41268
rect 27755 41228 29000 41256
rect 27755 41225 27767 41228
rect 27709 41219 27767 41225
rect 28994 41216 29000 41228
rect 29052 41216 29058 41268
rect 29178 41256 29184 41268
rect 29139 41228 29184 41256
rect 29178 41216 29184 41228
rect 29236 41216 29242 41268
rect 46474 41216 46480 41268
rect 46532 41256 46538 41268
rect 46753 41259 46811 41265
rect 46753 41256 46765 41259
rect 46532 41228 46765 41256
rect 46532 41216 46538 41228
rect 46753 41225 46765 41228
rect 46799 41225 46811 41259
rect 46753 41219 46811 41225
rect 24121 41191 24179 41197
rect 24121 41188 24133 41191
rect 22572 41160 22876 41188
rect 23124 41160 24133 41188
rect 22189 41151 22247 41157
rect 20901 41123 20959 41129
rect 20901 41089 20913 41123
rect 20947 41089 20959 41123
rect 20901 41083 20959 41089
rect 20993 41123 21051 41129
rect 20993 41089 21005 41123
rect 21039 41089 21051 41123
rect 21174 41120 21180 41132
rect 21135 41092 21180 41120
rect 20993 41083 21051 41089
rect 20916 41052 20944 41083
rect 21174 41080 21180 41092
rect 21232 41080 21238 41132
rect 21821 41123 21879 41129
rect 21821 41089 21833 41123
rect 21867 41089 21879 41123
rect 22002 41120 22008 41132
rect 21963 41092 22008 41120
rect 21821 41083 21879 41089
rect 21450 41052 21456 41064
rect 20916 41024 21456 41052
rect 21450 41012 21456 41024
rect 21508 41012 21514 41064
rect 20533 40987 20591 40993
rect 20533 40953 20545 40987
rect 20579 40984 20591 40987
rect 20898 40984 20904 40996
rect 20579 40956 20904 40984
rect 20579 40953 20591 40956
rect 20533 40947 20591 40953
rect 20898 40944 20904 40956
rect 20956 40944 20962 40996
rect 1394 40876 1400 40928
rect 1452 40916 1458 40928
rect 1949 40919 2007 40925
rect 1949 40916 1961 40919
rect 1452 40888 1961 40916
rect 1452 40876 1458 40888
rect 1949 40885 1961 40888
rect 1995 40885 2007 40919
rect 1949 40879 2007 40885
rect 15654 40876 15660 40928
rect 15712 40916 15718 40928
rect 16117 40919 16175 40925
rect 16117 40916 16129 40919
rect 15712 40888 16129 40916
rect 15712 40876 15718 40888
rect 16117 40885 16129 40888
rect 16163 40885 16175 40919
rect 21836 40916 21864 41083
rect 22002 41080 22008 41092
rect 22060 41080 22066 41132
rect 22830 41080 22836 41132
rect 22888 41129 22894 41132
rect 22888 41123 22937 41129
rect 23011 41123 23017 41135
rect 22888 41089 22891 41123
rect 22925 41089 22937 41123
rect 22972 41095 23017 41123
rect 22888 41083 22937 41089
rect 23011 41083 23017 41095
rect 23069 41083 23075 41135
rect 23124 41129 23152 41160
rect 24121 41157 24133 41160
rect 24167 41157 24179 41191
rect 24121 41151 24179 41157
rect 25222 41148 25228 41200
rect 25280 41188 25286 41200
rect 26878 41188 26884 41200
rect 25280 41160 26884 41188
rect 25280 41148 25286 41160
rect 26878 41148 26884 41160
rect 26936 41188 26942 41200
rect 28813 41191 28871 41197
rect 28813 41188 28825 41191
rect 26936 41160 28120 41188
rect 26936 41148 26942 41160
rect 23114 41123 23172 41129
rect 23114 41089 23126 41123
rect 23160 41089 23172 41123
rect 23290 41120 23296 41132
rect 23251 41092 23296 41120
rect 23114 41083 23172 41089
rect 22888 41080 22894 41083
rect 23290 41080 23296 41092
rect 23348 41080 23354 41132
rect 23658 41080 23664 41132
rect 23716 41120 23722 41132
rect 23753 41123 23811 41129
rect 23753 41120 23765 41123
rect 23716 41092 23765 41120
rect 23716 41080 23722 41092
rect 23753 41089 23765 41092
rect 23799 41089 23811 41123
rect 23753 41083 23811 41089
rect 23842 41080 23848 41132
rect 23900 41120 23906 41132
rect 28092 41129 28120 41160
rect 28184 41160 28825 41188
rect 28184 41129 28212 41160
rect 28813 41157 28825 41160
rect 28859 41157 28871 41191
rect 28813 41151 28871 41157
rect 23937 41123 23995 41129
rect 23937 41120 23949 41123
rect 23900 41092 23949 41120
rect 23900 41080 23906 41092
rect 23937 41089 23949 41092
rect 23983 41089 23995 41123
rect 23937 41083 23995 41089
rect 27985 41123 28043 41129
rect 27985 41089 27997 41123
rect 28031 41089 28043 41123
rect 27985 41083 28043 41089
rect 28077 41123 28135 41129
rect 28077 41089 28089 41123
rect 28123 41089 28135 41123
rect 28077 41083 28135 41089
rect 28169 41123 28227 41129
rect 28169 41089 28181 41123
rect 28215 41089 28227 41123
rect 28169 41083 28227 41089
rect 28353 41123 28411 41129
rect 28353 41089 28365 41123
rect 28399 41089 28411 41123
rect 28353 41083 28411 41089
rect 28997 41123 29055 41129
rect 28997 41089 29009 41123
rect 29043 41120 29055 41123
rect 29086 41120 29092 41132
rect 29043 41092 29092 41120
rect 29043 41089 29055 41092
rect 28997 41083 29055 41089
rect 23198 41012 23204 41064
rect 23256 41052 23262 41064
rect 28000 41052 28028 41083
rect 23256 41024 28028 41052
rect 23256 41012 23262 41024
rect 23290 40944 23296 40996
rect 23348 40984 23354 40996
rect 27430 40984 27436 40996
rect 23348 40956 27436 40984
rect 23348 40944 23354 40956
rect 27430 40944 27436 40956
rect 27488 40984 27494 40996
rect 28368 40984 28396 41083
rect 29086 41080 29092 41092
rect 29144 41080 29150 41132
rect 29273 41123 29331 41129
rect 29273 41089 29285 41123
rect 29319 41120 29331 41123
rect 30926 41120 30932 41132
rect 29319 41092 30932 41120
rect 29319 41089 29331 41092
rect 29273 41083 29331 41089
rect 30926 41080 30932 41092
rect 30984 41080 30990 41132
rect 32122 41080 32128 41132
rect 32180 41120 32186 41132
rect 32565 41123 32623 41129
rect 32565 41120 32577 41123
rect 32180 41092 32577 41120
rect 32180 41080 32186 41092
rect 32565 41089 32577 41092
rect 32611 41089 32623 41123
rect 46658 41120 46664 41132
rect 46619 41092 46664 41120
rect 32565 41083 32623 41089
rect 46658 41080 46664 41092
rect 46716 41080 46722 41132
rect 47946 41120 47952 41132
rect 47907 41092 47952 41120
rect 47946 41080 47952 41092
rect 48004 41080 48010 41132
rect 29546 41012 29552 41064
rect 29604 41052 29610 41064
rect 30282 41052 30288 41064
rect 29604 41024 30288 41052
rect 29604 41012 29610 41024
rect 30282 41012 30288 41024
rect 30340 41052 30346 41064
rect 32306 41052 32312 41064
rect 30340 41024 32312 41052
rect 30340 41012 30346 41024
rect 32306 41012 32312 41024
rect 32364 41012 32370 41064
rect 27488 40956 28396 40984
rect 27488 40944 27494 40956
rect 22094 40916 22100 40928
rect 21836 40888 22100 40916
rect 16117 40879 16175 40885
rect 22094 40876 22100 40888
rect 22152 40916 22158 40928
rect 22462 40916 22468 40928
rect 22152 40888 22468 40916
rect 22152 40876 22158 40888
rect 22462 40876 22468 40888
rect 22520 40876 22526 40928
rect 23106 40876 23112 40928
rect 23164 40916 23170 40928
rect 25222 40916 25228 40928
rect 23164 40888 25228 40916
rect 23164 40876 23170 40888
rect 25222 40876 25228 40888
rect 25280 40876 25286 40928
rect 33689 40919 33747 40925
rect 33689 40885 33701 40919
rect 33735 40916 33747 40919
rect 33778 40916 33784 40928
rect 33735 40888 33784 40916
rect 33735 40885 33747 40888
rect 33689 40879 33747 40885
rect 33778 40876 33784 40888
rect 33836 40876 33842 40928
rect 47394 40876 47400 40928
rect 47452 40916 47458 40928
rect 48041 40919 48099 40925
rect 48041 40916 48053 40919
rect 47452 40888 48053 40916
rect 47452 40876 47458 40888
rect 48041 40885 48053 40888
rect 48087 40885 48099 40919
rect 48041 40879 48099 40885
rect 1104 40826 48852 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 48852 40826
rect 1104 40752 48852 40774
rect 23290 40672 23296 40724
rect 23348 40712 23354 40724
rect 23385 40715 23443 40721
rect 23385 40712 23397 40715
rect 23348 40684 23397 40712
rect 23348 40672 23354 40684
rect 23385 40681 23397 40684
rect 23431 40681 23443 40715
rect 23385 40675 23443 40681
rect 27338 40672 27344 40724
rect 27396 40712 27402 40724
rect 27396 40684 31708 40712
rect 27396 40672 27402 40684
rect 28810 40604 28816 40656
rect 28868 40644 28874 40656
rect 28997 40647 29055 40653
rect 28997 40644 29009 40647
rect 28868 40616 29009 40644
rect 28868 40604 28874 40616
rect 28997 40613 29009 40616
rect 29043 40613 29055 40647
rect 31680 40644 31708 40684
rect 32214 40672 32220 40724
rect 32272 40712 32278 40724
rect 32861 40715 32919 40721
rect 32861 40712 32873 40715
rect 32272 40684 32873 40712
rect 32272 40672 32278 40684
rect 32861 40681 32873 40684
rect 32907 40681 32919 40715
rect 32861 40675 32919 40681
rect 31680 40616 32076 40644
rect 28997 40607 29055 40613
rect 28813 40511 28871 40517
rect 28813 40477 28825 40511
rect 28859 40508 28871 40511
rect 29178 40508 29184 40520
rect 28859 40480 29184 40508
rect 28859 40477 28871 40480
rect 28813 40471 28871 40477
rect 29178 40468 29184 40480
rect 29236 40508 29242 40520
rect 31110 40508 31116 40520
rect 29236 40480 30972 40508
rect 31071 40480 31116 40508
rect 29236 40468 29242 40480
rect 1854 40440 1860 40452
rect 1815 40412 1860 40440
rect 1854 40400 1860 40412
rect 1912 40400 1918 40452
rect 23293 40443 23351 40449
rect 23293 40409 23305 40443
rect 23339 40440 23351 40443
rect 23382 40440 23388 40452
rect 23339 40412 23388 40440
rect 23339 40409 23351 40412
rect 23293 40403 23351 40409
rect 23382 40400 23388 40412
rect 23440 40400 23446 40452
rect 29733 40443 29791 40449
rect 29733 40409 29745 40443
rect 29779 40440 29791 40443
rect 29822 40440 29828 40452
rect 29779 40412 29828 40440
rect 29779 40409 29791 40412
rect 29733 40403 29791 40409
rect 29822 40400 29828 40412
rect 29880 40400 29886 40452
rect 29917 40443 29975 40449
rect 29917 40409 29929 40443
rect 29963 40440 29975 40443
rect 30742 40440 30748 40452
rect 29963 40412 30748 40440
rect 29963 40409 29975 40412
rect 29917 40403 29975 40409
rect 1949 40375 2007 40381
rect 1949 40341 1961 40375
rect 1995 40372 2007 40375
rect 17126 40372 17132 40384
rect 1995 40344 17132 40372
rect 1995 40341 2007 40344
rect 1949 40335 2007 40341
rect 17126 40332 17132 40344
rect 17184 40332 17190 40384
rect 23658 40332 23664 40384
rect 23716 40372 23722 40384
rect 29932 40372 29960 40403
rect 30742 40400 30748 40412
rect 30800 40400 30806 40452
rect 23716 40344 29960 40372
rect 30101 40375 30159 40381
rect 23716 40332 23722 40344
rect 30101 40341 30113 40375
rect 30147 40372 30159 40375
rect 30834 40372 30840 40384
rect 30147 40344 30840 40372
rect 30147 40341 30159 40344
rect 30101 40335 30159 40341
rect 30834 40332 30840 40344
rect 30892 40332 30898 40384
rect 30944 40372 30972 40480
rect 31110 40468 31116 40480
rect 31168 40468 31174 40520
rect 32048 40508 32076 40616
rect 32309 40579 32367 40585
rect 32309 40545 32321 40579
rect 32355 40576 32367 40579
rect 32398 40576 32404 40588
rect 32355 40548 32404 40576
rect 32355 40545 32367 40548
rect 32309 40539 32367 40545
rect 32398 40536 32404 40548
rect 32456 40576 32462 40588
rect 32950 40576 32956 40588
rect 32456 40548 32956 40576
rect 32456 40536 32462 40548
rect 32950 40536 32956 40548
rect 33008 40576 33014 40588
rect 33413 40579 33471 40585
rect 33413 40576 33425 40579
rect 33008 40548 33425 40576
rect 33008 40536 33014 40548
rect 33413 40545 33425 40548
rect 33459 40545 33471 40579
rect 33413 40539 33471 40545
rect 32125 40511 32183 40517
rect 32125 40508 32137 40511
rect 32048 40480 32137 40508
rect 32125 40477 32137 40480
rect 32171 40477 32183 40511
rect 33318 40508 33324 40520
rect 33279 40480 33324 40508
rect 32125 40471 32183 40477
rect 33318 40468 33324 40480
rect 33376 40468 33382 40520
rect 45833 40511 45891 40517
rect 45833 40477 45845 40511
rect 45879 40508 45891 40511
rect 46293 40511 46351 40517
rect 46293 40508 46305 40511
rect 45879 40480 46305 40508
rect 45879 40477 45891 40480
rect 45833 40471 45891 40477
rect 46293 40477 46305 40480
rect 46339 40477 46351 40511
rect 46293 40471 46351 40477
rect 31754 40440 31760 40452
rect 31312 40412 31760 40440
rect 31113 40375 31171 40381
rect 31113 40372 31125 40375
rect 30944 40344 31125 40372
rect 31113 40341 31125 40344
rect 31159 40372 31171 40375
rect 31312 40372 31340 40412
rect 31754 40400 31760 40412
rect 31812 40400 31818 40452
rect 33778 40440 33784 40452
rect 33152 40412 33784 40440
rect 31662 40372 31668 40384
rect 31159 40344 31340 40372
rect 31623 40344 31668 40372
rect 31159 40341 31171 40344
rect 31113 40335 31171 40341
rect 31662 40332 31668 40344
rect 31720 40332 31726 40384
rect 32033 40375 32091 40381
rect 32033 40341 32045 40375
rect 32079 40372 32091 40375
rect 33152 40372 33180 40412
rect 33778 40400 33784 40412
rect 33836 40400 33842 40452
rect 46474 40440 46480 40452
rect 46435 40412 46480 40440
rect 46474 40400 46480 40412
rect 46532 40400 46538 40452
rect 48130 40440 48136 40452
rect 48091 40412 48136 40440
rect 48130 40400 48136 40412
rect 48188 40400 48194 40452
rect 32079 40344 33180 40372
rect 33229 40375 33287 40381
rect 32079 40341 32091 40344
rect 32033 40335 32091 40341
rect 33229 40341 33241 40375
rect 33275 40372 33287 40375
rect 33410 40372 33416 40384
rect 33275 40344 33416 40372
rect 33275 40341 33287 40344
rect 33229 40335 33287 40341
rect 33410 40332 33416 40344
rect 33468 40332 33474 40384
rect 1104 40282 48852 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 48852 40282
rect 1104 40208 48852 40230
rect 24765 40171 24823 40177
rect 24765 40137 24777 40171
rect 24811 40137 24823 40171
rect 29822 40168 29828 40180
rect 29783 40140 29828 40168
rect 24765 40131 24823 40137
rect 20349 40103 20407 40109
rect 20349 40069 20361 40103
rect 20395 40100 20407 40103
rect 20533 40103 20591 40109
rect 20395 40072 20484 40100
rect 20395 40069 20407 40072
rect 20349 40063 20407 40069
rect 20456 40032 20484 40072
rect 20533 40069 20545 40103
rect 20579 40100 20591 40103
rect 21266 40100 21272 40112
rect 20579 40072 21272 40100
rect 20579 40069 20591 40072
rect 20533 40063 20591 40069
rect 21266 40060 21272 40072
rect 21324 40060 21330 40112
rect 23842 40060 23848 40112
rect 23900 40100 23906 40112
rect 24486 40100 24492 40112
rect 23900 40072 24492 40100
rect 23900 40060 23906 40072
rect 24486 40060 24492 40072
rect 24544 40060 24550 40112
rect 20456 40004 20576 40032
rect 20548 39976 20576 40004
rect 22002 39992 22008 40044
rect 22060 40032 22066 40044
rect 22060 39992 22094 40032
rect 23198 39992 23204 40044
rect 23256 40032 23262 40044
rect 23641 40035 23699 40041
rect 23641 40032 23653 40035
rect 23256 40004 23653 40032
rect 23256 39992 23262 40004
rect 23641 40001 23653 40004
rect 23687 40001 23699 40035
rect 24780 40032 24808 40131
rect 29822 40128 29828 40140
rect 29880 40128 29886 40180
rect 32214 40168 32220 40180
rect 31220 40140 32220 40168
rect 26970 40100 26976 40112
rect 25884 40072 26976 40100
rect 24854 40032 24860 40044
rect 24767 40004 24860 40032
rect 23641 39995 23699 40001
rect 24854 39992 24860 40004
rect 24912 40032 24918 40044
rect 25639 40035 25697 40041
rect 25639 40032 25651 40035
rect 24912 40004 25651 40032
rect 24912 39992 24918 40004
rect 25639 40001 25651 40004
rect 25685 40001 25697 40035
rect 25774 40032 25780 40044
rect 25735 40004 25780 40032
rect 25639 39995 25697 40001
rect 25774 39992 25780 40004
rect 25832 39992 25838 40044
rect 25884 40041 25912 40072
rect 26970 40060 26976 40072
rect 27028 40060 27034 40112
rect 30193 40103 30251 40109
rect 30193 40069 30205 40103
rect 30239 40100 30251 40103
rect 31018 40100 31024 40112
rect 30239 40072 31024 40100
rect 30239 40069 30251 40072
rect 30193 40063 30251 40069
rect 31018 40060 31024 40072
rect 31076 40060 31082 40112
rect 31220 40109 31248 40140
rect 32214 40128 32220 40140
rect 32272 40128 32278 40180
rect 33410 40128 33416 40180
rect 33468 40168 33474 40180
rect 34333 40171 34391 40177
rect 34333 40168 34345 40171
rect 33468 40140 34345 40168
rect 33468 40128 33474 40140
rect 34333 40137 34345 40140
rect 34379 40137 34391 40171
rect 34333 40131 34391 40137
rect 46474 40128 46480 40180
rect 46532 40168 46538 40180
rect 46753 40171 46811 40177
rect 46753 40168 46765 40171
rect 46532 40140 46765 40168
rect 46532 40128 46538 40140
rect 46753 40137 46765 40140
rect 46799 40137 46811 40171
rect 46753 40131 46811 40137
rect 31205 40103 31263 40109
rect 31205 40069 31217 40103
rect 31251 40069 31263 40103
rect 31205 40063 31263 40069
rect 31662 40060 31668 40112
rect 31720 40100 31726 40112
rect 32309 40103 32367 40109
rect 32309 40100 32321 40103
rect 31720 40072 31800 40100
rect 31720 40060 31726 40072
rect 25869 40035 25927 40041
rect 25869 40001 25881 40035
rect 25915 40001 25927 40035
rect 26050 40032 26056 40044
rect 26011 40004 26056 40032
rect 25869 39995 25927 40001
rect 26050 39992 26056 40004
rect 26108 39992 26114 40044
rect 29822 39992 29828 40044
rect 29880 40032 29886 40044
rect 29880 40004 30420 40032
rect 29880 39992 29886 40004
rect 20530 39924 20536 39976
rect 20588 39924 20594 39976
rect 22066 39964 22094 39992
rect 23290 39964 23296 39976
rect 22066 39936 23296 39964
rect 23290 39924 23296 39936
rect 23348 39924 23354 39976
rect 30392 39973 30420 40004
rect 30742 39992 30748 40044
rect 30800 40032 30806 40044
rect 31389 40035 31447 40041
rect 31389 40032 31401 40035
rect 30800 40004 31401 40032
rect 30800 39992 30806 40004
rect 31389 40001 31401 40004
rect 31435 40001 31447 40035
rect 31772 40032 31800 40072
rect 32232 40072 32321 40100
rect 32125 40035 32183 40041
rect 32125 40032 32137 40035
rect 31772 40004 32137 40032
rect 31389 39995 31447 40001
rect 32125 40001 32137 40004
rect 32171 40001 32183 40035
rect 32125 39995 32183 40001
rect 23385 39967 23443 39973
rect 23385 39933 23397 39967
rect 23431 39933 23443 39967
rect 23385 39927 23443 39933
rect 30285 39967 30343 39973
rect 30285 39933 30297 39967
rect 30331 39933 30343 39967
rect 30285 39927 30343 39933
rect 30377 39967 30435 39973
rect 30377 39933 30389 39967
rect 30423 39933 30435 39967
rect 31404 39964 31432 39995
rect 32232 39964 32260 40072
rect 32309 40069 32321 40072
rect 32355 40069 32367 40103
rect 32309 40063 32367 40069
rect 32968 40072 33456 40100
rect 31404 39936 32260 39964
rect 30377 39927 30435 39933
rect 2038 39788 2044 39840
rect 2096 39828 2102 39840
rect 2225 39831 2283 39837
rect 2225 39828 2237 39831
rect 2096 39800 2237 39828
rect 2096 39788 2102 39800
rect 2225 39797 2237 39800
rect 2271 39797 2283 39831
rect 2225 39791 2283 39797
rect 5534 39788 5540 39840
rect 5592 39828 5598 39840
rect 6086 39828 6092 39840
rect 5592 39800 6092 39828
rect 5592 39788 5598 39800
rect 6086 39788 6092 39800
rect 6144 39828 6150 39840
rect 17218 39828 17224 39840
rect 6144 39800 17224 39828
rect 6144 39788 6150 39800
rect 17218 39788 17224 39800
rect 17276 39788 17282 39840
rect 20346 39788 20352 39840
rect 20404 39828 20410 39840
rect 20717 39831 20775 39837
rect 20717 39828 20729 39831
rect 20404 39800 20729 39828
rect 20404 39788 20410 39800
rect 20717 39797 20729 39800
rect 20763 39797 20775 39831
rect 23400 39828 23428 39927
rect 24394 39856 24400 39908
rect 24452 39896 24458 39908
rect 24452 39868 26096 39896
rect 24452 39856 24458 39868
rect 24762 39828 24768 39840
rect 23400 39800 24768 39828
rect 20717 39791 20775 39797
rect 24762 39788 24768 39800
rect 24820 39788 24826 39840
rect 25409 39831 25467 39837
rect 25409 39797 25421 39831
rect 25455 39828 25467 39831
rect 25958 39828 25964 39840
rect 25455 39800 25964 39828
rect 25455 39797 25467 39800
rect 25409 39791 25467 39797
rect 25958 39788 25964 39800
rect 26016 39788 26022 39840
rect 26068 39828 26096 39868
rect 30190 39856 30196 39908
rect 30248 39896 30254 39908
rect 30300 39896 30328 39927
rect 32306 39924 32312 39976
rect 32364 39964 32370 39976
rect 32968 39973 32996 40072
rect 33226 40041 33232 40044
rect 33220 39995 33232 40041
rect 33284 40032 33290 40044
rect 33428 40032 33456 40072
rect 35894 40032 35900 40044
rect 33284 40004 33320 40032
rect 33428 40004 35900 40032
rect 33226 39992 33232 39995
rect 33284 39992 33290 40004
rect 35894 39992 35900 40004
rect 35952 39992 35958 40044
rect 37182 39992 37188 40044
rect 37240 40032 37246 40044
rect 46661 40035 46719 40041
rect 46661 40032 46673 40035
rect 37240 40004 46673 40032
rect 37240 39992 37246 40004
rect 46661 40001 46673 40004
rect 46707 40001 46719 40035
rect 46661 39995 46719 40001
rect 32953 39967 33011 39973
rect 32953 39964 32965 39967
rect 32364 39936 32965 39964
rect 32364 39924 32370 39936
rect 32953 39933 32965 39936
rect 32999 39933 33011 39967
rect 32953 39927 33011 39933
rect 30248 39868 30328 39896
rect 31573 39899 31631 39905
rect 30248 39856 30254 39868
rect 31573 39865 31585 39899
rect 31619 39896 31631 39899
rect 31619 39868 32720 39896
rect 31619 39865 31631 39868
rect 31573 39859 31631 39865
rect 32398 39828 32404 39840
rect 26068 39800 32404 39828
rect 32398 39788 32404 39800
rect 32456 39788 32462 39840
rect 32490 39788 32496 39840
rect 32548 39828 32554 39840
rect 32692 39828 32720 39868
rect 33962 39828 33968 39840
rect 32548 39800 32593 39828
rect 32692 39800 33968 39828
rect 32548 39788 32554 39800
rect 33962 39788 33968 39800
rect 34020 39788 34026 39840
rect 46290 39788 46296 39840
rect 46348 39828 46354 39840
rect 47765 39831 47823 39837
rect 47765 39828 47777 39831
rect 46348 39800 47777 39828
rect 46348 39788 46354 39800
rect 47765 39797 47777 39800
rect 47811 39797 47823 39831
rect 47765 39791 47823 39797
rect 1104 39738 48852 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 48852 39738
rect 1104 39664 48852 39686
rect 17218 39584 17224 39636
rect 17276 39624 17282 39636
rect 23198 39624 23204 39636
rect 17276 39596 22094 39624
rect 23159 39596 23204 39624
rect 17276 39584 17282 39596
rect 21266 39556 21272 39568
rect 21227 39528 21272 39556
rect 21266 39516 21272 39528
rect 21324 39516 21330 39568
rect 22066 39556 22094 39596
rect 23198 39584 23204 39596
rect 23256 39584 23262 39636
rect 23290 39584 23296 39636
rect 23348 39624 23354 39636
rect 31846 39624 31852 39636
rect 23348 39596 31852 39624
rect 23348 39584 23354 39596
rect 31846 39584 31852 39596
rect 31904 39584 31910 39636
rect 32122 39624 32128 39636
rect 32083 39596 32128 39624
rect 32122 39584 32128 39596
rect 32180 39584 32186 39636
rect 25130 39556 25136 39568
rect 22066 39528 25136 39556
rect 25130 39516 25136 39528
rect 25188 39516 25194 39568
rect 32490 39516 32496 39568
rect 32548 39556 32554 39568
rect 32548 39528 32628 39556
rect 32548 39516 32554 39528
rect 24857 39491 24915 39497
rect 24857 39488 24869 39491
rect 23676 39460 24869 39488
rect 2869 39423 2927 39429
rect 2869 39389 2881 39423
rect 2915 39420 2927 39423
rect 5534 39420 5540 39432
rect 2915 39392 5540 39420
rect 2915 39389 2927 39392
rect 2869 39383 2927 39389
rect 5534 39380 5540 39392
rect 5592 39380 5598 39432
rect 19889 39423 19947 39429
rect 19889 39389 19901 39423
rect 19935 39420 19947 39423
rect 20714 39420 20720 39432
rect 19935 39392 20720 39420
rect 19935 39389 19947 39392
rect 19889 39383 19947 39389
rect 20714 39380 20720 39392
rect 20772 39420 20778 39432
rect 21818 39420 21824 39432
rect 20772 39392 21824 39420
rect 20772 39380 20778 39392
rect 21818 39380 21824 39392
rect 21876 39380 21882 39432
rect 22097 39423 22155 39429
rect 22097 39389 22109 39423
rect 22143 39420 22155 39423
rect 22462 39420 22468 39432
rect 22143 39392 22468 39420
rect 22143 39389 22155 39392
rect 22097 39383 22155 39389
rect 22462 39380 22468 39392
rect 22520 39380 22526 39432
rect 23474 39420 23480 39432
rect 23435 39392 23480 39420
rect 23474 39380 23480 39392
rect 23532 39380 23538 39432
rect 23676 39429 23704 39460
rect 24857 39457 24869 39460
rect 24903 39457 24915 39491
rect 27246 39488 27252 39500
rect 24857 39451 24915 39457
rect 26988 39460 27252 39488
rect 23569 39423 23627 39429
rect 23569 39389 23581 39423
rect 23615 39389 23627 39423
rect 23569 39383 23627 39389
rect 23661 39423 23719 39429
rect 23661 39389 23673 39423
rect 23707 39389 23719 39423
rect 23661 39383 23719 39389
rect 23845 39423 23903 39429
rect 23845 39389 23857 39423
rect 23891 39420 23903 39423
rect 23934 39420 23940 39432
rect 23891 39392 23940 39420
rect 23891 39389 23903 39392
rect 23845 39383 23903 39389
rect 19978 39312 19984 39364
rect 20036 39352 20042 39364
rect 20134 39355 20192 39361
rect 20134 39352 20146 39355
rect 20036 39324 20146 39352
rect 20036 39312 20042 39324
rect 20134 39321 20146 39324
rect 20180 39321 20192 39355
rect 20134 39315 20192 39321
rect 22281 39355 22339 39361
rect 22281 39321 22293 39355
rect 22327 39352 22339 39355
rect 23584 39352 23612 39383
rect 23934 39380 23940 39392
rect 23992 39380 23998 39432
rect 24762 39380 24768 39432
rect 24820 39420 24826 39432
rect 25869 39423 25927 39429
rect 25869 39420 25881 39423
rect 24820 39392 25881 39420
rect 24820 39380 24826 39392
rect 25869 39389 25881 39392
rect 25915 39389 25927 39423
rect 25869 39383 25927 39389
rect 25958 39380 25964 39432
rect 26016 39420 26022 39432
rect 26125 39423 26183 39429
rect 26125 39420 26137 39423
rect 26016 39392 26137 39420
rect 26016 39380 26022 39392
rect 26125 39389 26137 39392
rect 26171 39389 26183 39423
rect 26125 39383 26183 39389
rect 26418 39380 26424 39432
rect 26476 39420 26482 39432
rect 26988 39420 27016 39460
rect 27246 39448 27252 39460
rect 27304 39488 27310 39500
rect 30282 39488 30288 39500
rect 27304 39460 28212 39488
rect 30243 39460 30288 39488
rect 27304 39448 27310 39460
rect 27893 39423 27951 39429
rect 26476 39392 27016 39420
rect 27080 39392 27844 39420
rect 26476 39380 26482 39392
rect 24394 39352 24400 39364
rect 22327 39324 23520 39352
rect 23584 39324 24400 39352
rect 22327 39321 22339 39324
rect 22281 39315 22339 39321
rect 23492 39296 23520 39324
rect 23676 39296 23704 39324
rect 24394 39312 24400 39324
rect 24452 39312 24458 39364
rect 24489 39355 24547 39361
rect 24489 39321 24501 39355
rect 24535 39321 24547 39355
rect 24489 39315 24547 39321
rect 24673 39355 24731 39361
rect 24673 39321 24685 39355
rect 24719 39352 24731 39355
rect 24854 39352 24860 39364
rect 24719 39324 24860 39352
rect 24719 39321 24731 39324
rect 24673 39315 24731 39321
rect 2222 39244 2228 39296
rect 2280 39284 2286 39296
rect 2961 39287 3019 39293
rect 2961 39284 2973 39287
rect 2280 39256 2973 39284
rect 2280 39244 2286 39256
rect 2961 39253 2973 39256
rect 3007 39253 3019 39287
rect 2961 39247 3019 39253
rect 22186 39244 22192 39296
rect 22244 39284 22250 39296
rect 22465 39287 22523 39293
rect 22465 39284 22477 39287
rect 22244 39256 22477 39284
rect 22244 39244 22250 39256
rect 22465 39253 22477 39256
rect 22511 39253 22523 39287
rect 22465 39247 22523 39253
rect 23474 39244 23480 39296
rect 23532 39244 23538 39296
rect 23658 39244 23664 39296
rect 23716 39244 23722 39296
rect 24504 39284 24532 39315
rect 24854 39312 24860 39324
rect 24912 39312 24918 39364
rect 24946 39312 24952 39364
rect 25004 39352 25010 39364
rect 27080 39352 27108 39392
rect 25004 39324 27108 39352
rect 25004 39312 25010 39324
rect 27154 39312 27160 39364
rect 27212 39352 27218 39364
rect 27709 39355 27767 39361
rect 27709 39352 27721 39355
rect 27212 39324 27721 39352
rect 27212 39312 27218 39324
rect 27709 39321 27721 39324
rect 27755 39321 27767 39355
rect 27709 39315 27767 39321
rect 24578 39284 24584 39296
rect 24504 39256 24584 39284
rect 24578 39244 24584 39256
rect 24636 39244 24642 39296
rect 27249 39287 27307 39293
rect 27249 39253 27261 39287
rect 27295 39284 27307 39287
rect 27430 39284 27436 39296
rect 27295 39256 27436 39284
rect 27295 39253 27307 39256
rect 27249 39247 27307 39253
rect 27430 39244 27436 39256
rect 27488 39244 27494 39296
rect 27816 39284 27844 39392
rect 27893 39389 27905 39423
rect 27939 39420 27951 39423
rect 27982 39420 27988 39432
rect 27939 39392 27988 39420
rect 27939 39389 27951 39392
rect 27893 39383 27951 39389
rect 27982 39380 27988 39392
rect 28040 39380 28046 39432
rect 28184 39429 28212 39460
rect 30282 39448 30288 39460
rect 30340 39448 30346 39500
rect 28169 39423 28227 39429
rect 28169 39389 28181 39423
rect 28215 39389 28227 39423
rect 28169 39383 28227 39389
rect 32306 39380 32312 39432
rect 32364 39420 32370 39432
rect 32600 39429 32628 39528
rect 33226 39488 33232 39500
rect 33187 39460 33232 39488
rect 33226 39448 33232 39460
rect 33284 39448 33290 39500
rect 33318 39448 33324 39500
rect 33376 39488 33382 39500
rect 46290 39488 46296 39500
rect 33376 39460 33640 39488
rect 46251 39460 46296 39488
rect 33376 39448 33382 39460
rect 32401 39423 32459 39429
rect 32401 39420 32413 39423
rect 32364 39392 32413 39420
rect 32364 39380 32370 39392
rect 32401 39389 32413 39392
rect 32447 39389 32459 39423
rect 32401 39383 32459 39389
rect 32490 39420 32548 39426
rect 32490 39386 32502 39420
rect 32536 39386 32548 39420
rect 32490 39380 32548 39386
rect 32585 39423 32643 39429
rect 32585 39389 32597 39423
rect 32631 39389 32643 39423
rect 32585 39383 32643 39389
rect 32766 39380 32772 39432
rect 32824 39420 32830 39432
rect 33502 39429 33508 39432
rect 33485 39423 33508 39429
rect 32824 39392 32869 39420
rect 32824 39380 32830 39392
rect 33485 39389 33497 39423
rect 33485 39383 33508 39389
rect 33502 39380 33508 39383
rect 33560 39380 33566 39432
rect 33612 39429 33640 39460
rect 46290 39448 46296 39460
rect 46348 39448 46354 39500
rect 48130 39488 48136 39500
rect 48091 39460 48136 39488
rect 48130 39448 48136 39460
rect 48188 39448 48194 39500
rect 33597 39423 33655 39429
rect 33597 39389 33609 39423
rect 33643 39389 33655 39423
rect 33597 39383 33655 39389
rect 33689 39423 33747 39429
rect 33689 39389 33701 39423
rect 33735 39389 33747 39423
rect 33870 39420 33876 39432
rect 33831 39392 33876 39420
rect 33689 39383 33747 39389
rect 28074 39352 28080 39364
rect 27987 39324 28080 39352
rect 28074 39312 28080 39324
rect 28132 39352 28138 39364
rect 28810 39352 28816 39364
rect 28132 39324 28816 39352
rect 28132 39312 28138 39324
rect 28810 39312 28816 39324
rect 28868 39312 28874 39364
rect 30374 39312 30380 39364
rect 30432 39352 30438 39364
rect 30530 39355 30588 39361
rect 30530 39352 30542 39355
rect 30432 39324 30542 39352
rect 30432 39312 30438 39324
rect 30530 39321 30542 39324
rect 30576 39321 30588 39355
rect 32508 39352 32536 39380
rect 33318 39352 33324 39364
rect 32508 39324 33324 39352
rect 30530 39315 30588 39321
rect 33318 39312 33324 39324
rect 33376 39312 33382 39364
rect 33704 39352 33732 39383
rect 33870 39380 33876 39392
rect 33928 39380 33934 39432
rect 34701 39423 34759 39429
rect 34701 39389 34713 39423
rect 34747 39420 34759 39423
rect 35894 39420 35900 39432
rect 34747 39392 35900 39420
rect 34747 39389 34759 39392
rect 34701 39383 34759 39389
rect 35894 39380 35900 39392
rect 35952 39420 35958 39432
rect 36541 39423 36599 39429
rect 36541 39420 36553 39423
rect 35952 39392 36553 39420
rect 35952 39380 35958 39392
rect 36541 39389 36553 39392
rect 36587 39389 36599 39423
rect 36541 39383 36599 39389
rect 33962 39352 33968 39364
rect 33704 39324 33968 39352
rect 33962 39312 33968 39324
rect 34020 39312 34026 39364
rect 34238 39312 34244 39364
rect 34296 39352 34302 39364
rect 34946 39355 35004 39361
rect 34946 39352 34958 39355
rect 34296 39324 34958 39352
rect 34296 39312 34302 39324
rect 34946 39321 34958 39324
rect 34992 39321 35004 39355
rect 34946 39315 35004 39321
rect 35986 39312 35992 39364
rect 36044 39352 36050 39364
rect 36786 39355 36844 39361
rect 36786 39352 36798 39355
rect 36044 39324 36798 39352
rect 36044 39312 36050 39324
rect 36786 39321 36798 39324
rect 36832 39321 36844 39355
rect 36786 39315 36844 39321
rect 46477 39355 46535 39361
rect 46477 39321 46489 39355
rect 46523 39352 46535 39355
rect 46750 39352 46756 39364
rect 46523 39324 46756 39352
rect 46523 39321 46535 39324
rect 46477 39315 46535 39321
rect 46750 39312 46756 39324
rect 46808 39312 46814 39364
rect 30926 39284 30932 39296
rect 27816 39256 30932 39284
rect 30926 39244 30932 39256
rect 30984 39244 30990 39296
rect 31018 39244 31024 39296
rect 31076 39284 31082 39296
rect 31662 39284 31668 39296
rect 31076 39256 31668 39284
rect 31076 39244 31082 39256
rect 31662 39244 31668 39256
rect 31720 39244 31726 39296
rect 33594 39244 33600 39296
rect 33652 39284 33658 39296
rect 36081 39287 36139 39293
rect 36081 39284 36093 39287
rect 33652 39256 36093 39284
rect 33652 39244 33658 39256
rect 36081 39253 36093 39256
rect 36127 39253 36139 39287
rect 36081 39247 36139 39253
rect 37458 39244 37464 39296
rect 37516 39284 37522 39296
rect 37921 39287 37979 39293
rect 37921 39284 37933 39287
rect 37516 39256 37933 39284
rect 37516 39244 37522 39256
rect 37921 39253 37933 39256
rect 37967 39253 37979 39287
rect 37921 39247 37979 39253
rect 1104 39194 48852 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 48852 39194
rect 1104 39120 48852 39142
rect 19889 39083 19947 39089
rect 19889 39049 19901 39083
rect 19935 39080 19947 39083
rect 19978 39080 19984 39092
rect 19935 39052 19984 39080
rect 19935 39049 19947 39052
rect 19889 39043 19947 39049
rect 19978 39040 19984 39052
rect 20036 39040 20042 39092
rect 24213 39083 24271 39089
rect 24213 39049 24225 39083
rect 24259 39080 24271 39083
rect 26050 39080 26056 39092
rect 24259 39052 26056 39080
rect 24259 39049 24271 39052
rect 24213 39043 24271 39049
rect 26050 39040 26056 39052
rect 26108 39040 26114 39092
rect 26418 39080 26424 39092
rect 26379 39052 26424 39080
rect 26418 39040 26424 39052
rect 26476 39040 26482 39092
rect 26970 39080 26976 39092
rect 26931 39052 26976 39080
rect 26970 39040 26976 39052
rect 27028 39040 27034 39092
rect 27341 39083 27399 39089
rect 27341 39049 27353 39083
rect 27387 39080 27399 39083
rect 28074 39080 28080 39092
rect 27387 39052 28080 39080
rect 27387 39049 27399 39052
rect 27341 39043 27399 39049
rect 28074 39040 28080 39052
rect 28132 39040 28138 39092
rect 29086 39040 29092 39092
rect 29144 39080 29150 39092
rect 29181 39083 29239 39089
rect 29181 39080 29193 39083
rect 29144 39052 29193 39080
rect 29144 39040 29150 39052
rect 29181 39049 29193 39052
rect 29227 39049 29239 39083
rect 29638 39080 29644 39092
rect 29599 39052 29644 39080
rect 29181 39043 29239 39049
rect 29638 39040 29644 39052
rect 29696 39040 29702 39092
rect 30374 39080 30380 39092
rect 30335 39052 30380 39080
rect 30374 39040 30380 39052
rect 30432 39040 30438 39092
rect 31846 39040 31852 39092
rect 31904 39080 31910 39092
rect 35986 39080 35992 39092
rect 31904 39052 34928 39080
rect 35947 39052 35992 39080
rect 31904 39040 31910 39052
rect 2222 39012 2228 39024
rect 2183 38984 2228 39012
rect 2222 38972 2228 38984
rect 2280 38972 2286 39024
rect 33318 39012 33324 39024
rect 23124 38984 30696 39012
rect 2038 38944 2044 38956
rect 1999 38916 2044 38944
rect 2038 38904 2044 38916
rect 2096 38904 2102 38956
rect 18598 38904 18604 38956
rect 18656 38944 18662 38956
rect 20165 38947 20223 38953
rect 20165 38944 20177 38947
rect 18656 38916 20177 38944
rect 18656 38904 18662 38916
rect 20165 38913 20177 38916
rect 20211 38913 20223 38947
rect 20165 38907 20223 38913
rect 20257 38947 20315 38953
rect 20257 38913 20269 38947
rect 20303 38913 20315 38947
rect 20257 38907 20315 38913
rect 2774 38876 2780 38888
rect 2735 38848 2780 38876
rect 2774 38836 2780 38848
rect 2832 38836 2838 38888
rect 20272 38876 20300 38907
rect 20346 38904 20352 38956
rect 20404 38944 20410 38956
rect 20533 38947 20591 38953
rect 20404 38916 20449 38944
rect 20404 38904 20410 38916
rect 20533 38913 20545 38947
rect 20579 38944 20591 38947
rect 21910 38944 21916 38956
rect 20579 38916 21916 38944
rect 20579 38913 20591 38916
rect 20533 38907 20591 38913
rect 21910 38904 21916 38916
rect 21968 38904 21974 38956
rect 22094 38953 22100 38956
rect 22088 38907 22100 38953
rect 22152 38944 22158 38956
rect 22152 38916 22188 38944
rect 22094 38904 22100 38907
rect 22152 38904 22158 38916
rect 20622 38876 20628 38888
rect 20272 38848 20628 38876
rect 20622 38836 20628 38848
rect 20680 38836 20686 38888
rect 21818 38876 21824 38888
rect 21779 38848 21824 38876
rect 21818 38836 21824 38848
rect 21876 38836 21882 38888
rect 21266 38700 21272 38752
rect 21324 38740 21330 38752
rect 23124 38740 23152 38984
rect 23382 38904 23388 38956
rect 23440 38944 23446 38956
rect 24121 38947 24179 38953
rect 24121 38944 24133 38947
rect 23440 38916 24133 38944
rect 23440 38904 23446 38916
rect 24121 38913 24133 38916
rect 24167 38913 24179 38947
rect 24121 38907 24179 38913
rect 24762 38904 24768 38956
rect 24820 38944 24826 38956
rect 25041 38947 25099 38953
rect 25041 38944 25053 38947
rect 24820 38916 25053 38944
rect 24820 38904 24826 38916
rect 25041 38913 25053 38916
rect 25087 38913 25099 38947
rect 25041 38907 25099 38913
rect 25308 38947 25366 38953
rect 25308 38913 25320 38947
rect 25354 38944 25366 38947
rect 25682 38944 25688 38956
rect 25354 38916 25688 38944
rect 25354 38913 25366 38916
rect 25308 38907 25366 38913
rect 25682 38904 25688 38916
rect 25740 38904 25746 38956
rect 25866 38904 25872 38956
rect 25924 38944 25930 38956
rect 27157 38947 27215 38953
rect 27157 38944 27169 38947
rect 25924 38916 27169 38944
rect 25924 38904 25930 38916
rect 27157 38913 27169 38916
rect 27203 38913 27215 38947
rect 27157 38907 27215 38913
rect 23750 38836 23756 38888
rect 23808 38876 23814 38888
rect 24670 38876 24676 38888
rect 23808 38848 24676 38876
rect 23808 38836 23814 38848
rect 24670 38836 24676 38848
rect 24728 38836 24734 38888
rect 27172 38876 27200 38907
rect 27430 38904 27436 38956
rect 27488 38944 27494 38956
rect 29549 38947 29607 38953
rect 27488 38916 27533 38944
rect 27488 38904 27494 38916
rect 29549 38913 29561 38947
rect 29595 38944 29607 38947
rect 30374 38944 30380 38956
rect 29595 38916 30380 38944
rect 29595 38913 29607 38916
rect 29549 38907 29607 38913
rect 30374 38904 30380 38916
rect 30432 38904 30438 38956
rect 30668 38953 30696 38984
rect 30760 38984 33324 39012
rect 30760 38953 30788 38984
rect 33318 38972 33324 38984
rect 33376 38972 33382 39024
rect 33594 39012 33600 39024
rect 33555 38984 33600 39012
rect 33594 38972 33600 38984
rect 33652 38972 33658 39024
rect 34238 39012 34244 39024
rect 34199 38984 34244 39012
rect 34238 38972 34244 38984
rect 34296 38972 34302 39024
rect 34330 38972 34336 39024
rect 34388 39012 34394 39024
rect 34900 39012 34928 39052
rect 35986 39040 35992 39052
rect 36044 39040 36050 39092
rect 36078 39040 36084 39092
rect 36136 39080 36142 39092
rect 37645 39083 37703 39089
rect 37645 39080 37657 39083
rect 36136 39052 36413 39080
rect 36136 39040 36142 39052
rect 36170 39012 36176 39024
rect 34388 38984 34652 39012
rect 34388 38972 34394 38984
rect 34624 38956 34652 38984
rect 34900 38984 36176 39012
rect 30653 38947 30711 38953
rect 30653 38913 30665 38947
rect 30699 38913 30711 38947
rect 30653 38907 30711 38913
rect 30745 38947 30803 38953
rect 30745 38913 30757 38947
rect 30791 38913 30803 38947
rect 30745 38907 30803 38913
rect 27982 38876 27988 38888
rect 27172 38848 27988 38876
rect 27982 38836 27988 38848
rect 28040 38876 28046 38888
rect 28902 38876 28908 38888
rect 28040 38848 28908 38876
rect 28040 38836 28046 38848
rect 28902 38836 28908 38848
rect 28960 38836 28966 38888
rect 29822 38876 29828 38888
rect 29783 38848 29828 38876
rect 29822 38836 29828 38848
rect 29880 38836 29886 38888
rect 25976 38780 29224 38808
rect 21324 38712 23152 38740
rect 23201 38743 23259 38749
rect 21324 38700 21330 38712
rect 23201 38709 23213 38743
rect 23247 38740 23259 38743
rect 23474 38740 23480 38752
rect 23247 38712 23480 38740
rect 23247 38709 23259 38712
rect 23201 38703 23259 38709
rect 23474 38700 23480 38712
rect 23532 38700 23538 38752
rect 24578 38700 24584 38752
rect 24636 38740 24642 38752
rect 25976 38740 26004 38780
rect 24636 38712 26004 38740
rect 29196 38740 29224 38780
rect 29270 38768 29276 38820
rect 29328 38808 29334 38820
rect 30760 38808 30788 38907
rect 30834 38904 30840 38956
rect 30892 38944 30898 38956
rect 31021 38947 31079 38953
rect 30892 38916 30937 38944
rect 30892 38904 30898 38916
rect 31021 38913 31033 38947
rect 31067 38944 31079 38947
rect 31294 38944 31300 38956
rect 31067 38916 31300 38944
rect 31067 38913 31079 38916
rect 31021 38907 31079 38913
rect 31294 38904 31300 38916
rect 31352 38944 31358 38956
rect 32766 38944 32772 38956
rect 31352 38916 32772 38944
rect 31352 38904 31358 38916
rect 32766 38904 32772 38916
rect 32824 38904 32830 38956
rect 33413 38947 33471 38953
rect 33413 38913 33425 38947
rect 33459 38913 33471 38947
rect 33413 38907 33471 38913
rect 33428 38876 33456 38907
rect 34422 38904 34428 38956
rect 34480 38953 34486 38956
rect 34480 38947 34529 38953
rect 34480 38913 34483 38947
rect 34517 38913 34529 38947
rect 34480 38907 34529 38913
rect 34606 38950 34664 38956
rect 34900 38953 34928 38984
rect 36170 38972 36176 38984
rect 36228 38972 36234 39024
rect 36385 39012 36413 39052
rect 36372 38984 36413 39012
rect 36485 39052 37657 39080
rect 36372 38956 36400 38984
rect 36485 38956 36513 39052
rect 37645 39049 37657 39052
rect 37691 39049 37703 39083
rect 46750 39080 46756 39092
rect 46711 39052 46756 39080
rect 37645 39043 37703 39049
rect 46750 39040 46756 39052
rect 46808 39040 46814 39092
rect 37458 39012 37464 39024
rect 37419 38984 37464 39012
rect 37458 38972 37464 38984
rect 37516 38972 37522 39024
rect 34606 38916 34618 38950
rect 34652 38916 34664 38950
rect 34606 38910 34664 38916
rect 34701 38947 34759 38953
rect 34701 38913 34713 38947
rect 34747 38913 34759 38947
rect 34701 38907 34759 38913
rect 34885 38947 34943 38953
rect 36265 38947 36323 38953
rect 34885 38913 34897 38947
rect 34931 38913 34943 38947
rect 34885 38907 34943 38913
rect 36260 38913 36277 38947
rect 36311 38913 36323 38947
rect 36260 38907 36323 38913
rect 36354 38950 36412 38956
rect 36354 38916 36366 38950
rect 36400 38916 36412 38950
rect 36354 38910 36412 38916
rect 36470 38950 36528 38956
rect 36470 38916 36482 38950
rect 36516 38916 36528 38950
rect 36630 38944 36636 38956
rect 36591 38916 36636 38944
rect 36470 38910 36528 38916
rect 34480 38904 34486 38907
rect 29328 38780 30788 38808
rect 31726 38848 33456 38876
rect 29328 38768 29334 38780
rect 31726 38740 31754 38848
rect 29196 38712 31754 38740
rect 33428 38740 33456 38848
rect 33781 38811 33839 38817
rect 33781 38777 33793 38811
rect 33827 38808 33839 38811
rect 34716 38808 34744 38907
rect 33827 38780 34744 38808
rect 36260 38808 36288 38907
rect 36630 38904 36636 38916
rect 36688 38904 36694 38956
rect 37274 38944 37280 38956
rect 37235 38916 37280 38944
rect 37274 38904 37280 38916
rect 37332 38904 37338 38956
rect 37366 38904 37372 38956
rect 37424 38944 37430 38956
rect 46661 38947 46719 38953
rect 46661 38944 46673 38947
rect 37424 38916 46673 38944
rect 37424 38904 37430 38916
rect 46661 38913 46673 38916
rect 46707 38913 46719 38947
rect 48130 38944 48136 38956
rect 48091 38916 48136 38944
rect 46661 38907 46719 38913
rect 48130 38904 48136 38916
rect 48188 38904 48194 38956
rect 45922 38876 45928 38888
rect 41386 38848 45928 38876
rect 41386 38808 41414 38848
rect 45922 38836 45928 38848
rect 45980 38836 45986 38888
rect 36260 38780 41414 38808
rect 33827 38777 33839 38780
rect 33781 38771 33839 38777
rect 34422 38740 34428 38752
rect 33428 38712 34428 38740
rect 24636 38700 24642 38712
rect 34422 38700 34428 38712
rect 34480 38700 34486 38752
rect 34514 38700 34520 38752
rect 34572 38740 34578 38752
rect 35710 38740 35716 38752
rect 34572 38712 35716 38740
rect 34572 38700 34578 38712
rect 35710 38700 35716 38712
rect 35768 38700 35774 38752
rect 35802 38700 35808 38752
rect 35860 38740 35866 38752
rect 37274 38740 37280 38752
rect 35860 38712 37280 38740
rect 35860 38700 35866 38712
rect 37274 38700 37280 38712
rect 37332 38700 37338 38752
rect 46750 38700 46756 38752
rect 46808 38740 46814 38752
rect 47949 38743 48007 38749
rect 47949 38740 47961 38743
rect 46808 38712 47961 38740
rect 46808 38700 46814 38712
rect 47949 38709 47961 38712
rect 47995 38709 48007 38743
rect 47949 38703 48007 38709
rect 1104 38650 48852 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 48852 38650
rect 1104 38576 48852 38598
rect 21729 38539 21787 38545
rect 21729 38505 21741 38539
rect 21775 38536 21787 38539
rect 22094 38536 22100 38548
rect 21775 38508 22100 38536
rect 21775 38505 21787 38508
rect 21729 38499 21787 38505
rect 22094 38496 22100 38508
rect 22152 38496 22158 38548
rect 22462 38496 22468 38548
rect 22520 38536 22526 38548
rect 24627 38539 24685 38545
rect 24627 38536 24639 38539
rect 22520 38508 24639 38536
rect 22520 38496 22526 38508
rect 24627 38505 24639 38508
rect 24673 38505 24685 38539
rect 25682 38536 25688 38548
rect 25643 38508 25688 38536
rect 24627 38499 24685 38505
rect 25682 38496 25688 38508
rect 25740 38496 25746 38548
rect 27798 38536 27804 38548
rect 26068 38508 27804 38536
rect 23014 38468 23020 38480
rect 22112 38440 23020 38468
rect 18598 38292 18604 38344
rect 18656 38332 18662 38344
rect 19245 38335 19303 38341
rect 19245 38332 19257 38335
rect 18656 38304 19257 38332
rect 18656 38292 18662 38304
rect 19245 38301 19257 38304
rect 19291 38332 19303 38335
rect 21818 38332 21824 38344
rect 19291 38304 21824 38332
rect 19291 38301 19303 38304
rect 19245 38295 19303 38301
rect 21818 38292 21824 38304
rect 21876 38292 21882 38344
rect 21910 38292 21916 38344
rect 21968 38332 21974 38344
rect 22112 38341 22140 38440
rect 23014 38428 23020 38440
rect 23072 38428 23078 38480
rect 23109 38471 23167 38477
rect 23109 38437 23121 38471
rect 23155 38468 23167 38471
rect 23934 38468 23940 38480
rect 23155 38440 23940 38468
rect 23155 38437 23167 38440
rect 23109 38431 23167 38437
rect 22005 38335 22063 38341
rect 22005 38332 22017 38335
rect 21968 38304 22017 38332
rect 21968 38292 21974 38304
rect 22005 38301 22017 38304
rect 22051 38301 22063 38335
rect 22005 38295 22063 38301
rect 22097 38335 22155 38341
rect 22097 38301 22109 38335
rect 22143 38301 22155 38335
rect 22097 38295 22155 38301
rect 22186 38292 22192 38344
rect 22244 38332 22250 38344
rect 22373 38335 22431 38341
rect 22244 38304 22289 38332
rect 22244 38292 22250 38304
rect 22373 38301 22385 38335
rect 22419 38332 22431 38335
rect 23124 38332 23152 38431
rect 23934 38428 23940 38440
rect 23992 38428 23998 38480
rect 25774 38428 25780 38480
rect 25832 38468 25838 38480
rect 26068 38468 26096 38508
rect 27798 38496 27804 38508
rect 27856 38536 27862 38548
rect 27856 38508 31754 38536
rect 27856 38496 27862 38508
rect 27154 38468 27160 38480
rect 25832 38440 26096 38468
rect 25832 38428 25838 38440
rect 23474 38360 23480 38412
rect 23532 38400 23538 38412
rect 23532 38372 26004 38400
rect 23532 38360 23538 38372
rect 22419 38304 23152 38332
rect 24397 38335 24455 38341
rect 22419 38301 22431 38304
rect 22373 38295 22431 38301
rect 24397 38301 24409 38335
rect 24443 38332 24455 38335
rect 24670 38332 24676 38344
rect 24443 38304 24676 38332
rect 24443 38301 24455 38304
rect 24397 38295 24455 38301
rect 24670 38292 24676 38304
rect 24728 38292 24734 38344
rect 25976 38341 26004 38372
rect 26068 38341 26096 38440
rect 26160 38440 27160 38468
rect 26160 38341 26188 38440
rect 27154 38428 27160 38440
rect 27212 38428 27218 38480
rect 29270 38400 29276 38412
rect 26252 38372 28672 38400
rect 25961 38335 26019 38341
rect 25961 38301 25973 38335
rect 26007 38301 26019 38335
rect 25961 38295 26019 38301
rect 26053 38335 26111 38341
rect 26053 38301 26065 38335
rect 26099 38301 26111 38335
rect 26053 38295 26111 38301
rect 26145 38335 26203 38341
rect 26145 38301 26157 38335
rect 26191 38301 26203 38335
rect 26145 38295 26203 38301
rect 18690 38224 18696 38276
rect 18748 38264 18754 38276
rect 19490 38267 19548 38273
rect 19490 38264 19502 38267
rect 18748 38236 19502 38264
rect 18748 38224 18754 38236
rect 19490 38233 19502 38236
rect 19536 38233 19548 38267
rect 19490 38227 19548 38233
rect 21358 38224 21364 38276
rect 21416 38264 21422 38276
rect 22925 38267 22983 38273
rect 22925 38264 22937 38267
rect 21416 38236 22937 38264
rect 21416 38224 21422 38236
rect 22925 38233 22937 38236
rect 22971 38233 22983 38267
rect 22925 38227 22983 38233
rect 23014 38224 23020 38276
rect 23072 38264 23078 38276
rect 23658 38264 23664 38276
rect 23072 38236 23664 38264
rect 23072 38224 23078 38236
rect 23658 38224 23664 38236
rect 23716 38224 23722 38276
rect 26252 38264 26280 38372
rect 28644 38341 28672 38372
rect 28736 38372 29276 38400
rect 28736 38341 28764 38372
rect 29270 38360 29276 38372
rect 29328 38360 29334 38412
rect 31726 38400 31754 38508
rect 31726 38372 32812 38400
rect 26329 38335 26387 38341
rect 26329 38301 26341 38335
rect 26375 38301 26387 38335
rect 26329 38295 26387 38301
rect 28629 38335 28687 38341
rect 28629 38301 28641 38335
rect 28675 38301 28687 38335
rect 28629 38295 28687 38301
rect 28721 38335 28779 38341
rect 28721 38301 28733 38335
rect 28767 38301 28779 38335
rect 28721 38295 28779 38301
rect 25976 38236 26280 38264
rect 19978 38156 19984 38208
rect 20036 38196 20042 38208
rect 20625 38199 20683 38205
rect 20625 38196 20637 38199
rect 20036 38168 20637 38196
rect 20036 38156 20042 38168
rect 20625 38165 20637 38168
rect 20671 38196 20683 38199
rect 25976 38196 26004 38236
rect 20671 38168 26004 38196
rect 20671 38165 20683 38168
rect 20625 38159 20683 38165
rect 26050 38156 26056 38208
rect 26108 38196 26114 38208
rect 26344 38196 26372 38295
rect 28810 38292 28816 38344
rect 28868 38332 28874 38344
rect 28868 38304 28913 38332
rect 28868 38292 28874 38304
rect 28994 38292 29000 38344
rect 29052 38332 29058 38344
rect 29549 38335 29607 38341
rect 29052 38304 29097 38332
rect 29052 38292 29058 38304
rect 29549 38301 29561 38335
rect 29595 38332 29607 38335
rect 30282 38332 30288 38344
rect 29595 38304 30288 38332
rect 29595 38301 29607 38304
rect 29549 38295 29607 38301
rect 30282 38292 30288 38304
rect 30340 38292 30346 38344
rect 32784 38341 32812 38372
rect 32677 38335 32735 38341
rect 32677 38301 32689 38335
rect 32723 38301 32735 38335
rect 32677 38295 32735 38301
rect 32769 38335 32827 38341
rect 32769 38301 32781 38335
rect 32815 38301 32827 38335
rect 32769 38295 32827 38301
rect 28353 38267 28411 38273
rect 28353 38233 28365 38267
rect 28399 38264 28411 38267
rect 29794 38267 29852 38273
rect 29794 38264 29806 38267
rect 28399 38236 29806 38264
rect 28399 38233 28411 38236
rect 28353 38227 28411 38233
rect 29794 38233 29806 38236
rect 29840 38233 29852 38267
rect 32692 38264 32720 38295
rect 32858 38292 32864 38344
rect 32916 38332 32922 38344
rect 33045 38335 33103 38341
rect 32916 38304 32961 38332
rect 32916 38292 32922 38304
rect 33045 38301 33057 38335
rect 33091 38332 33103 38335
rect 33134 38332 33140 38344
rect 33091 38304 33140 38332
rect 33091 38301 33103 38304
rect 33045 38295 33103 38301
rect 33134 38292 33140 38304
rect 33192 38332 33198 38344
rect 33870 38332 33876 38344
rect 33192 38304 33876 38332
rect 33192 38292 33198 38304
rect 33870 38292 33876 38304
rect 33928 38292 33934 38344
rect 35621 38335 35679 38341
rect 35621 38332 35633 38335
rect 35360 38304 35633 38332
rect 35360 38264 35388 38304
rect 35621 38301 35633 38304
rect 35667 38301 35679 38335
rect 35621 38295 35679 38301
rect 29794 38227 29852 38233
rect 29932 38236 32628 38264
rect 32692 38236 35388 38264
rect 35437 38267 35495 38273
rect 29932 38196 29960 38236
rect 26108 38168 29960 38196
rect 26108 38156 26114 38168
rect 30374 38156 30380 38208
rect 30432 38196 30438 38208
rect 30929 38199 30987 38205
rect 30929 38196 30941 38199
rect 30432 38168 30941 38196
rect 30432 38156 30438 38168
rect 30929 38165 30941 38168
rect 30975 38165 30987 38199
rect 30929 38159 30987 38165
rect 32401 38199 32459 38205
rect 32401 38165 32413 38199
rect 32447 38196 32459 38199
rect 32490 38196 32496 38208
rect 32447 38168 32496 38196
rect 32447 38165 32459 38168
rect 32401 38159 32459 38165
rect 32490 38156 32496 38168
rect 32548 38156 32554 38208
rect 32600 38196 32628 38236
rect 35437 38233 35449 38267
rect 35483 38233 35495 38267
rect 35636 38264 35664 38295
rect 35894 38292 35900 38344
rect 35952 38332 35958 38344
rect 36265 38335 36323 38341
rect 36265 38332 36277 38335
rect 35952 38304 36277 38332
rect 35952 38292 35958 38304
rect 36265 38301 36277 38304
rect 36311 38301 36323 38335
rect 47854 38332 47860 38344
rect 47815 38304 47860 38332
rect 36265 38295 36323 38301
rect 47854 38292 47860 38304
rect 47912 38292 47918 38344
rect 35636 38236 35940 38264
rect 35437 38227 35495 38233
rect 33134 38196 33140 38208
rect 32600 38168 33140 38196
rect 33134 38156 33140 38168
rect 33192 38156 33198 38208
rect 34514 38156 34520 38208
rect 34572 38196 34578 38208
rect 35452 38196 35480 38227
rect 35618 38196 35624 38208
rect 34572 38168 35624 38196
rect 34572 38156 34578 38168
rect 35618 38156 35624 38168
rect 35676 38156 35682 38208
rect 35802 38196 35808 38208
rect 35763 38168 35808 38196
rect 35802 38156 35808 38168
rect 35860 38156 35866 38208
rect 35912 38196 35940 38236
rect 36078 38224 36084 38276
rect 36136 38264 36142 38276
rect 36510 38267 36568 38273
rect 36510 38264 36522 38267
rect 36136 38236 36522 38264
rect 36136 38224 36142 38236
rect 36510 38233 36522 38236
rect 36556 38233 36568 38267
rect 36510 38227 36568 38233
rect 37645 38199 37703 38205
rect 37645 38196 37657 38199
rect 35912 38168 37657 38196
rect 37645 38165 37657 38168
rect 37691 38165 37703 38199
rect 37645 38159 37703 38165
rect 47118 38156 47124 38208
rect 47176 38196 47182 38208
rect 48041 38199 48099 38205
rect 48041 38196 48053 38199
rect 47176 38168 48053 38196
rect 47176 38156 47182 38168
rect 48041 38165 48053 38168
rect 48087 38165 48099 38199
rect 48041 38159 48099 38165
rect 1104 38106 48852 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 48852 38106
rect 1104 38032 48852 38054
rect 18601 37995 18659 38001
rect 18601 37961 18613 37995
rect 18647 37992 18659 37995
rect 18690 37992 18696 38004
rect 18647 37964 18696 37992
rect 18647 37961 18659 37964
rect 18601 37955 18659 37961
rect 18690 37952 18696 37964
rect 18748 37952 18754 38004
rect 22002 37992 22008 38004
rect 21963 37964 22008 37992
rect 22002 37952 22008 37964
rect 22060 37952 22066 38004
rect 25685 37995 25743 38001
rect 25685 37961 25697 37995
rect 25731 37992 25743 37995
rect 25774 37992 25780 38004
rect 25731 37964 25780 37992
rect 25731 37961 25743 37964
rect 25685 37955 25743 37961
rect 25774 37952 25780 37964
rect 25832 37952 25838 38004
rect 27430 37952 27436 38004
rect 27488 37992 27494 38004
rect 27525 37995 27583 38001
rect 27525 37992 27537 37995
rect 27488 37964 27537 37992
rect 27488 37952 27494 37964
rect 27525 37961 27537 37964
rect 27571 37961 27583 37995
rect 27525 37955 27583 37961
rect 28810 37952 28816 38004
rect 28868 37992 28874 38004
rect 29181 37995 29239 38001
rect 29181 37992 29193 37995
rect 28868 37964 29193 37992
rect 28868 37952 28874 37964
rect 29181 37961 29193 37964
rect 29227 37961 29239 37995
rect 36078 37992 36084 38004
rect 36039 37964 36084 37992
rect 29181 37955 29239 37961
rect 36078 37952 36084 37964
rect 36136 37952 36142 38004
rect 36372 37964 41414 37992
rect 19794 37924 19800 37936
rect 19260 37896 19800 37924
rect 1854 37856 1860 37868
rect 1815 37828 1860 37856
rect 1854 37816 1860 37828
rect 1912 37816 1918 37868
rect 18874 37856 18880 37868
rect 18835 37828 18880 37856
rect 18874 37816 18880 37828
rect 18932 37816 18938 37868
rect 19260 37865 19288 37896
rect 19794 37884 19800 37896
rect 19852 37884 19858 37936
rect 19889 37927 19947 37933
rect 19889 37893 19901 37927
rect 19935 37924 19947 37927
rect 19978 37924 19984 37936
rect 19935 37896 19984 37924
rect 19935 37893 19947 37896
rect 19889 37887 19947 37893
rect 19978 37884 19984 37896
rect 20036 37884 20042 37936
rect 23201 37927 23259 37933
rect 23201 37893 23213 37927
rect 23247 37924 23259 37927
rect 24578 37924 24584 37936
rect 23247 37896 24584 37924
rect 23247 37893 23259 37896
rect 23201 37887 23259 37893
rect 24578 37884 24584 37896
rect 24636 37884 24642 37936
rect 24670 37884 24676 37936
rect 24728 37924 24734 37936
rect 26234 37924 26240 37936
rect 24728 37896 26240 37924
rect 24728 37884 24734 37896
rect 26234 37884 26240 37896
rect 26292 37884 26298 37936
rect 29086 37924 29092 37936
rect 28828 37896 29092 37924
rect 18969 37859 19027 37865
rect 18969 37825 18981 37859
rect 19015 37825 19027 37859
rect 18969 37819 19027 37825
rect 19061 37859 19119 37865
rect 19061 37825 19073 37859
rect 19107 37825 19119 37859
rect 19061 37819 19119 37825
rect 19245 37859 19303 37865
rect 19245 37825 19257 37859
rect 19291 37825 19303 37859
rect 19245 37819 19303 37825
rect 19705 37859 19763 37865
rect 19705 37825 19717 37859
rect 19751 37856 19763 37859
rect 20346 37856 20352 37868
rect 19751 37828 20352 37856
rect 19751 37825 19763 37828
rect 19705 37819 19763 37825
rect 2041 37723 2099 37729
rect 2041 37689 2053 37723
rect 2087 37720 2099 37723
rect 2590 37720 2596 37732
rect 2087 37692 2596 37720
rect 2087 37689 2099 37692
rect 2041 37683 2099 37689
rect 2590 37680 2596 37692
rect 2648 37680 2654 37732
rect 18984 37720 19012 37819
rect 19076 37788 19104 37819
rect 20346 37816 20352 37828
rect 20404 37856 20410 37868
rect 20530 37856 20536 37868
rect 20404 37828 20536 37856
rect 20404 37816 20410 37828
rect 20530 37816 20536 37828
rect 20588 37816 20594 37868
rect 20625 37859 20683 37865
rect 20625 37825 20637 37859
rect 20671 37856 20683 37859
rect 21358 37856 21364 37868
rect 20671 37828 21364 37856
rect 20671 37825 20683 37828
rect 20625 37819 20683 37825
rect 21358 37816 21364 37828
rect 21416 37856 21422 37868
rect 21821 37859 21879 37865
rect 21821 37856 21833 37859
rect 21416 37828 21833 37856
rect 21416 37816 21422 37828
rect 21821 37825 21833 37828
rect 21867 37825 21879 37859
rect 21821 37819 21879 37825
rect 23017 37859 23075 37865
rect 23017 37825 23029 37859
rect 23063 37856 23075 37859
rect 23661 37859 23719 37865
rect 23661 37856 23673 37859
rect 23063 37828 23673 37856
rect 23063 37825 23075 37828
rect 23017 37819 23075 37825
rect 23661 37825 23673 37828
rect 23707 37856 23719 37859
rect 24688 37856 24716 37884
rect 23707 37828 24716 37856
rect 25593 37859 25651 37865
rect 23707 37825 23719 37828
rect 23661 37819 23719 37825
rect 25593 37825 25605 37859
rect 25639 37856 25651 37859
rect 26418 37856 26424 37868
rect 25639 37828 26424 37856
rect 25639 37825 25651 37828
rect 25593 37819 25651 37825
rect 26418 37816 26424 37828
rect 26476 37856 26482 37868
rect 27338 37856 27344 37868
rect 26476 37828 27344 37856
rect 26476 37816 26482 37828
rect 27338 37816 27344 37828
rect 27396 37816 27402 37868
rect 27433 37859 27491 37865
rect 27433 37825 27445 37859
rect 27479 37856 27491 37859
rect 28074 37856 28080 37868
rect 27479 37828 28080 37856
rect 27479 37825 27491 37828
rect 27433 37819 27491 37825
rect 28074 37816 28080 37828
rect 28132 37816 28138 37868
rect 28828 37865 28856 37896
rect 29086 37884 29092 37896
rect 29144 37884 29150 37936
rect 28813 37859 28871 37865
rect 28813 37825 28825 37859
rect 28859 37825 28871 37859
rect 28813 37819 28871 37825
rect 28997 37859 29055 37865
rect 28997 37825 29009 37859
rect 29043 37856 29055 37859
rect 29730 37856 29736 37868
rect 29043 37828 29736 37856
rect 29043 37825 29055 37828
rect 28997 37819 29055 37825
rect 29730 37816 29736 37828
rect 29788 37816 29794 37868
rect 30282 37816 30288 37868
rect 30340 37856 30346 37868
rect 31754 37856 31760 37868
rect 30340 37828 31760 37856
rect 30340 37816 30346 37828
rect 31754 37816 31760 37828
rect 31812 37856 31818 37868
rect 32401 37859 32459 37865
rect 32401 37856 32413 37859
rect 31812 37828 32413 37856
rect 31812 37816 31818 37828
rect 32401 37825 32413 37828
rect 32447 37825 32459 37859
rect 32401 37819 32459 37825
rect 32490 37816 32496 37868
rect 32548 37856 32554 37868
rect 36372 37865 36400 37964
rect 32657 37859 32715 37865
rect 32657 37856 32669 37859
rect 32548 37828 32669 37856
rect 32548 37816 32554 37828
rect 32657 37825 32669 37828
rect 32703 37825 32715 37859
rect 32657 37819 32715 37825
rect 36337 37859 36400 37865
rect 36337 37825 36349 37859
rect 36383 37828 36400 37859
rect 36462 37859 36520 37865
rect 36383 37825 36395 37828
rect 36337 37819 36395 37825
rect 36462 37825 36474 37859
rect 36508 37825 36520 37859
rect 36462 37819 36520 37825
rect 36562 37859 36620 37865
rect 36562 37825 36574 37859
rect 36608 37856 36620 37859
rect 36608 37828 36676 37856
rect 36608 37825 36620 37828
rect 36562 37819 36620 37825
rect 20073 37791 20131 37797
rect 20073 37788 20085 37791
rect 19076 37760 20085 37788
rect 20073 37757 20085 37760
rect 20119 37757 20131 37791
rect 23934 37788 23940 37800
rect 23895 37760 23940 37788
rect 20073 37751 20131 37757
rect 23934 37748 23940 37760
rect 23992 37748 23998 37800
rect 27522 37748 27528 37800
rect 27580 37788 27586 37800
rect 27709 37791 27767 37797
rect 27709 37788 27721 37791
rect 27580 37760 27721 37788
rect 27580 37748 27586 37760
rect 27709 37757 27721 37760
rect 27755 37788 27767 37791
rect 29822 37788 29828 37800
rect 27755 37760 29828 37788
rect 27755 37757 27767 37760
rect 27709 37751 27767 37757
rect 29822 37748 29828 37760
rect 29880 37748 29886 37800
rect 36170 37748 36176 37800
rect 36228 37788 36234 37800
rect 36464 37788 36492 37819
rect 36228 37760 36492 37788
rect 36228 37748 36234 37760
rect 19610 37720 19616 37732
rect 18984 37692 19616 37720
rect 19610 37680 19616 37692
rect 19668 37720 19674 37732
rect 20530 37720 20536 37732
rect 19668 37692 20536 37720
rect 19668 37680 19674 37692
rect 20530 37680 20536 37692
rect 20588 37680 20594 37732
rect 35802 37680 35808 37732
rect 35860 37720 35866 37732
rect 36648 37720 36676 37828
rect 36722 37816 36728 37868
rect 36780 37856 36786 37868
rect 41386 37856 41414 37964
rect 46750 37856 46756 37868
rect 36780 37828 36825 37856
rect 41386 37828 46756 37856
rect 36780 37816 36786 37828
rect 46750 37816 46756 37828
rect 46808 37816 46814 37868
rect 35860 37692 36676 37720
rect 35860 37680 35866 37692
rect 20809 37655 20867 37661
rect 20809 37621 20821 37655
rect 20855 37652 20867 37655
rect 21174 37652 21180 37664
rect 20855 37624 21180 37652
rect 20855 37621 20867 37624
rect 20809 37615 20867 37621
rect 21174 37612 21180 37624
rect 21232 37612 21238 37664
rect 26326 37612 26332 37664
rect 26384 37652 26390 37664
rect 27065 37655 27123 37661
rect 27065 37652 27077 37655
rect 26384 37624 27077 37652
rect 26384 37612 26390 37624
rect 27065 37621 27077 37624
rect 27111 37621 27123 37655
rect 27065 37615 27123 37621
rect 32674 37612 32680 37664
rect 32732 37652 32738 37664
rect 33781 37655 33839 37661
rect 33781 37652 33793 37655
rect 32732 37624 33793 37652
rect 32732 37612 32738 37624
rect 33781 37621 33793 37624
rect 33827 37621 33839 37655
rect 33781 37615 33839 37621
rect 1104 37562 48852 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 48852 37562
rect 1104 37488 48852 37510
rect 21910 37448 21916 37460
rect 12406 37420 21916 37448
rect 2041 37315 2099 37321
rect 2041 37281 2053 37315
rect 2087 37312 2099 37315
rect 12406 37312 12434 37420
rect 21910 37408 21916 37420
rect 21968 37408 21974 37460
rect 28994 37408 29000 37460
rect 29052 37448 29058 37460
rect 31294 37448 31300 37460
rect 29052 37420 31300 37448
rect 29052 37408 29058 37420
rect 31294 37408 31300 37420
rect 31352 37408 31358 37460
rect 32217 37451 32275 37457
rect 32217 37417 32229 37451
rect 32263 37448 32275 37451
rect 32858 37448 32864 37460
rect 32263 37420 32864 37448
rect 32263 37417 32275 37420
rect 32217 37411 32275 37417
rect 32858 37408 32864 37420
rect 32916 37408 32922 37460
rect 19610 37340 19616 37392
rect 19668 37340 19674 37392
rect 21542 37380 21548 37392
rect 21503 37352 21548 37380
rect 21542 37340 21548 37352
rect 21600 37340 21606 37392
rect 28813 37383 28871 37389
rect 28813 37349 28825 37383
rect 28859 37380 28871 37383
rect 29270 37380 29276 37392
rect 28859 37352 29276 37380
rect 28859 37349 28871 37352
rect 28813 37343 28871 37349
rect 29270 37340 29276 37352
rect 29328 37340 29334 37392
rect 29748 37352 31524 37380
rect 2087 37284 12434 37312
rect 2087 37281 2099 37284
rect 2041 37275 2099 37281
rect 19426 37204 19432 37256
rect 19484 37244 19490 37256
rect 19628 37253 19656 37340
rect 29086 37272 29092 37324
rect 29144 37312 29150 37324
rect 29748 37312 29776 37352
rect 29144 37284 29776 37312
rect 29144 37272 29150 37284
rect 29822 37272 29828 37324
rect 29880 37312 29886 37324
rect 30929 37315 30987 37321
rect 30929 37312 30941 37315
rect 29880 37284 30941 37312
rect 29880 37272 29886 37284
rect 30929 37281 30941 37284
rect 30975 37281 30987 37315
rect 30929 37275 30987 37281
rect 19521 37247 19579 37253
rect 19521 37244 19533 37247
rect 19484 37216 19533 37244
rect 19484 37204 19490 37216
rect 19521 37213 19533 37216
rect 19567 37213 19579 37247
rect 19521 37207 19579 37213
rect 19610 37247 19668 37253
rect 19610 37213 19622 37247
rect 19656 37213 19668 37247
rect 19610 37207 19668 37213
rect 19705 37247 19763 37253
rect 19705 37213 19717 37247
rect 19751 37213 19763 37247
rect 19705 37207 19763 37213
rect 1854 37176 1860 37188
rect 1815 37148 1860 37176
rect 1854 37136 1860 37148
rect 1912 37136 1918 37188
rect 19242 37108 19248 37120
rect 19203 37080 19248 37108
rect 19242 37068 19248 37080
rect 19300 37068 19306 37120
rect 19720 37108 19748 37207
rect 19794 37204 19800 37256
rect 19852 37244 19858 37256
rect 19889 37247 19947 37253
rect 19889 37244 19901 37247
rect 19852 37216 19901 37244
rect 19852 37204 19858 37216
rect 19889 37213 19901 37216
rect 19935 37244 19947 37247
rect 20717 37247 20775 37253
rect 19935 37216 20668 37244
rect 19935 37213 19947 37216
rect 19889 37207 19947 37213
rect 19978 37136 19984 37188
rect 20036 37176 20042 37188
rect 20533 37179 20591 37185
rect 20533 37176 20545 37179
rect 20036 37148 20545 37176
rect 20036 37136 20042 37148
rect 20533 37145 20545 37148
rect 20579 37145 20591 37179
rect 20640 37176 20668 37216
rect 20717 37213 20729 37247
rect 20763 37244 20775 37247
rect 21818 37244 21824 37256
rect 20763 37216 21824 37244
rect 20763 37213 20775 37216
rect 20717 37207 20775 37213
rect 21818 37204 21824 37216
rect 21876 37204 21882 37256
rect 23934 37244 23940 37256
rect 22664 37216 23940 37244
rect 22664 37188 22692 37216
rect 23934 37204 23940 37216
rect 23992 37244 23998 37256
rect 24397 37247 24455 37253
rect 24397 37244 24409 37247
rect 23992 37216 24409 37244
rect 23992 37204 23998 37216
rect 24397 37213 24409 37216
rect 24443 37213 24455 37247
rect 24397 37207 24455 37213
rect 24762 37204 24768 37256
rect 24820 37244 24826 37256
rect 26694 37244 26700 37256
rect 24820 37216 26700 37244
rect 24820 37204 24826 37216
rect 26694 37204 26700 37216
rect 26752 37204 26758 37256
rect 27338 37204 27344 37256
rect 27396 37244 27402 37256
rect 28629 37247 28687 37253
rect 28629 37244 28641 37247
rect 27396 37216 28641 37244
rect 27396 37204 27402 37216
rect 28629 37213 28641 37216
rect 28675 37213 28687 37247
rect 28629 37207 28687 37213
rect 29549 37247 29607 37253
rect 29549 37213 29561 37247
rect 29595 37244 29607 37247
rect 31496 37244 31524 37352
rect 32398 37340 32404 37392
rect 32456 37380 32462 37392
rect 36170 37380 36176 37392
rect 32456 37352 36176 37380
rect 32456 37340 32462 37352
rect 36170 37340 36176 37352
rect 36228 37340 36234 37392
rect 33318 37272 33324 37324
rect 33376 37312 33382 37324
rect 33376 37284 33548 37312
rect 33376 37272 33382 37284
rect 32398 37244 32404 37256
rect 29595 37216 30420 37244
rect 31496 37216 32404 37244
rect 29595 37213 29607 37216
rect 29549 37207 29607 37213
rect 21358 37176 21364 37188
rect 20640 37148 20944 37176
rect 21319 37148 21364 37176
rect 20533 37139 20591 37145
rect 20806 37108 20812 37120
rect 19720 37080 20812 37108
rect 20806 37068 20812 37080
rect 20864 37068 20870 37120
rect 20916 37108 20944 37148
rect 21358 37136 21364 37148
rect 21416 37136 21422 37188
rect 22646 37176 22652 37188
rect 22607 37148 22652 37176
rect 22646 37136 22652 37148
rect 22704 37136 22710 37188
rect 22833 37179 22891 37185
rect 22833 37145 22845 37179
rect 22879 37176 22891 37179
rect 23290 37176 23296 37188
rect 22879 37148 23296 37176
rect 22879 37145 22891 37148
rect 22833 37139 22891 37145
rect 23290 37136 23296 37148
rect 23348 37136 23354 37188
rect 24578 37176 24584 37188
rect 24539 37148 24584 37176
rect 24578 37136 24584 37148
rect 24636 37136 24642 37188
rect 25774 37176 25780 37188
rect 24688 37148 25780 37176
rect 21542 37108 21548 37120
rect 20916 37080 21548 37108
rect 21542 37068 21548 37080
rect 21600 37068 21606 37120
rect 22922 37068 22928 37120
rect 22980 37108 22986 37120
rect 23017 37111 23075 37117
rect 23017 37108 23029 37111
rect 22980 37080 23029 37108
rect 22980 37068 22986 37080
rect 23017 37077 23029 37080
rect 23063 37077 23075 37111
rect 23017 37071 23075 37077
rect 24394 37068 24400 37120
rect 24452 37108 24458 37120
rect 24688 37108 24716 37148
rect 25774 37136 25780 37148
rect 25832 37136 25838 37188
rect 25869 37179 25927 37185
rect 25869 37145 25881 37179
rect 25915 37145 25927 37179
rect 26050 37176 26056 37188
rect 26011 37148 26056 37176
rect 25869 37139 25927 37145
rect 24452 37080 24716 37108
rect 24765 37111 24823 37117
rect 24452 37068 24458 37080
rect 24765 37077 24777 37111
rect 24811 37108 24823 37111
rect 24854 37108 24860 37120
rect 24811 37080 24860 37108
rect 24811 37077 24823 37080
rect 24765 37071 24823 37077
rect 24854 37068 24860 37080
rect 24912 37068 24918 37120
rect 25884 37108 25912 37139
rect 26050 37136 26056 37148
rect 26108 37136 26114 37188
rect 26326 37176 26332 37188
rect 26160 37148 26332 37176
rect 26160 37108 26188 37148
rect 26326 37136 26332 37148
rect 26384 37136 26390 37188
rect 26970 37185 26976 37188
rect 26964 37139 26976 37185
rect 27028 37176 27034 37188
rect 27028 37148 27064 37176
rect 26970 37136 26976 37139
rect 27028 37136 27034 37148
rect 27982 37136 27988 37188
rect 28040 37176 28046 37188
rect 28994 37176 29000 37188
rect 28040 37148 29000 37176
rect 28040 37136 28046 37148
rect 28994 37136 29000 37148
rect 29052 37136 29058 37188
rect 29730 37176 29736 37188
rect 29691 37148 29736 37176
rect 29730 37136 29736 37148
rect 29788 37136 29794 37188
rect 25884 37080 26188 37108
rect 26237 37111 26295 37117
rect 26237 37077 26249 37111
rect 26283 37108 26295 37111
rect 27430 37108 27436 37120
rect 26283 37080 27436 37108
rect 26283 37077 26295 37080
rect 26237 37071 26295 37077
rect 27430 37068 27436 37080
rect 27488 37068 27494 37120
rect 28074 37108 28080 37120
rect 27987 37080 28080 37108
rect 28074 37068 28080 37080
rect 28132 37108 28138 37120
rect 28534 37108 28540 37120
rect 28132 37080 28540 37108
rect 28132 37068 28138 37080
rect 28534 37068 28540 37080
rect 28592 37068 28598 37120
rect 29362 37068 29368 37120
rect 29420 37108 29426 37120
rect 30392 37117 30420 37216
rect 32398 37204 32404 37216
rect 32456 37204 32462 37256
rect 32674 37244 32680 37256
rect 32635 37216 32680 37244
rect 32674 37204 32680 37216
rect 32732 37204 32738 37256
rect 33520 37253 33548 37284
rect 33413 37247 33471 37253
rect 33413 37213 33425 37247
rect 33459 37213 33471 37247
rect 33413 37207 33471 37213
rect 33505 37247 33563 37253
rect 33505 37213 33517 37247
rect 33551 37213 33563 37247
rect 33505 37207 33563 37213
rect 30837 37179 30895 37185
rect 30837 37145 30849 37179
rect 30883 37176 30895 37179
rect 32692 37176 32720 37204
rect 33226 37176 33232 37188
rect 30883 37148 32720 37176
rect 32968 37148 33232 37176
rect 30883 37145 30895 37148
rect 30837 37139 30895 37145
rect 29917 37111 29975 37117
rect 29917 37108 29929 37111
rect 29420 37080 29929 37108
rect 29420 37068 29426 37080
rect 29917 37077 29929 37080
rect 29963 37077 29975 37111
rect 29917 37071 29975 37077
rect 30377 37111 30435 37117
rect 30377 37077 30389 37111
rect 30423 37077 30435 37111
rect 30742 37108 30748 37120
rect 30703 37080 30748 37108
rect 30377 37071 30435 37077
rect 30742 37068 30748 37080
rect 30800 37068 30806 37120
rect 32585 37111 32643 37117
rect 32585 37077 32597 37111
rect 32631 37108 32643 37111
rect 32968 37108 32996 37148
rect 33226 37136 33232 37148
rect 33284 37136 33290 37188
rect 33428 37176 33456 37207
rect 33594 37204 33600 37256
rect 33652 37244 33658 37256
rect 33781 37247 33839 37253
rect 33652 37216 33697 37244
rect 33652 37204 33658 37216
rect 33781 37213 33793 37247
rect 33827 37244 33839 37247
rect 33870 37244 33876 37256
rect 33827 37216 33876 37244
rect 33827 37213 33839 37216
rect 33781 37207 33839 37213
rect 33870 37204 33876 37216
rect 33928 37204 33934 37256
rect 36078 37244 36084 37256
rect 36039 37216 36084 37244
rect 36078 37204 36084 37216
rect 36136 37204 36142 37256
rect 36188 37253 36216 37340
rect 40678 37272 40684 37324
rect 40736 37312 40742 37324
rect 46842 37312 46848 37324
rect 40736 37284 46848 37312
rect 40736 37272 40742 37284
rect 46842 37272 46848 37284
rect 46900 37272 46906 37324
rect 36173 37247 36231 37253
rect 36449 37247 36507 37253
rect 36173 37213 36185 37247
rect 36219 37213 36231 37247
rect 36173 37207 36231 37213
rect 36265 37241 36323 37247
rect 36265 37207 36277 37241
rect 36311 37207 36323 37241
rect 36449 37213 36461 37247
rect 36495 37244 36507 37247
rect 36630 37244 36636 37256
rect 36495 37216 36636 37244
rect 36495 37213 36507 37216
rect 36449 37207 36507 37213
rect 36265 37201 36323 37207
rect 36630 37204 36636 37216
rect 36688 37204 36694 37256
rect 42794 37244 42800 37256
rect 41386 37216 42800 37244
rect 35526 37176 35532 37188
rect 33428 37148 35532 37176
rect 35526 37136 35532 37148
rect 35584 37136 35590 37188
rect 33134 37108 33140 37120
rect 32631 37080 32996 37108
rect 33095 37080 33140 37108
rect 32631 37077 32643 37080
rect 32585 37071 32643 37077
rect 33134 37068 33140 37080
rect 33192 37068 33198 37120
rect 35710 37068 35716 37120
rect 35768 37108 35774 37120
rect 35805 37111 35863 37117
rect 35805 37108 35817 37111
rect 35768 37080 35817 37108
rect 35768 37068 35774 37080
rect 35805 37077 35817 37080
rect 35851 37077 35863 37111
rect 35805 37071 35863 37077
rect 35986 37068 35992 37120
rect 36044 37108 36050 37120
rect 36280 37108 36308 37201
rect 36354 37136 36360 37188
rect 36412 37176 36418 37188
rect 41386 37176 41414 37216
rect 42794 37204 42800 37216
rect 42852 37204 42858 37256
rect 36412 37148 41414 37176
rect 36412 37136 36418 37148
rect 36044 37080 36308 37108
rect 36044 37068 36050 37080
rect 1104 37018 48852 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 48852 37018
rect 1104 36944 48852 36966
rect 17402 36864 17408 36916
rect 17460 36904 17466 36916
rect 24394 36904 24400 36916
rect 17460 36876 24400 36904
rect 17460 36864 17466 36876
rect 24394 36864 24400 36876
rect 24452 36864 24458 36916
rect 24578 36864 24584 36916
rect 24636 36904 24642 36916
rect 25225 36907 25283 36913
rect 25225 36904 25237 36907
rect 24636 36876 25237 36904
rect 24636 36864 24642 36876
rect 25225 36873 25237 36876
rect 25271 36873 25283 36907
rect 25225 36867 25283 36873
rect 18868 36839 18926 36845
rect 18868 36805 18880 36839
rect 18914 36836 18926 36839
rect 19242 36836 19248 36848
rect 18914 36808 19248 36836
rect 18914 36805 18926 36808
rect 18868 36799 18926 36805
rect 19242 36796 19248 36808
rect 19300 36796 19306 36848
rect 20346 36796 20352 36848
rect 20404 36836 20410 36848
rect 20441 36839 20499 36845
rect 20441 36836 20453 36839
rect 20404 36808 20453 36836
rect 20404 36796 20410 36808
rect 20441 36805 20453 36808
rect 20487 36836 20499 36839
rect 22646 36836 22652 36848
rect 20487 36808 22652 36836
rect 20487 36805 20499 36808
rect 20441 36799 20499 36805
rect 22646 36796 22652 36808
rect 22704 36796 22710 36848
rect 23934 36836 23940 36848
rect 23847 36808 23940 36836
rect 18598 36768 18604 36780
rect 18559 36740 18604 36768
rect 18598 36728 18604 36740
rect 18656 36728 18662 36780
rect 20625 36771 20683 36777
rect 20625 36737 20637 36771
rect 20671 36768 20683 36771
rect 22180 36771 22238 36777
rect 20671 36740 20944 36768
rect 20671 36737 20683 36740
rect 20625 36731 20683 36737
rect 20806 36700 20812 36712
rect 20767 36672 20812 36700
rect 20806 36660 20812 36672
rect 20864 36660 20870 36712
rect 19981 36635 20039 36641
rect 19981 36601 19993 36635
rect 20027 36632 20039 36635
rect 20916 36632 20944 36740
rect 22180 36737 22192 36771
rect 22226 36768 22238 36771
rect 22462 36768 22468 36780
rect 22226 36740 22468 36768
rect 22226 36737 22238 36740
rect 22180 36731 22238 36737
rect 22462 36728 22468 36740
rect 22520 36728 22526 36780
rect 23860 36777 23888 36808
rect 23934 36796 23940 36808
rect 23992 36836 23998 36848
rect 24762 36836 24768 36848
rect 23992 36808 24768 36836
rect 23992 36796 23998 36808
rect 24762 36796 24768 36808
rect 24820 36796 24826 36848
rect 23845 36771 23903 36777
rect 23845 36737 23857 36771
rect 23891 36737 23903 36771
rect 23845 36731 23903 36737
rect 24112 36771 24170 36777
rect 24112 36737 24124 36771
rect 24158 36768 24170 36771
rect 24394 36768 24400 36780
rect 24158 36740 24400 36768
rect 24158 36737 24170 36740
rect 24112 36731 24170 36737
rect 24394 36728 24400 36740
rect 24452 36728 24458 36780
rect 25240 36768 25268 36867
rect 26694 36864 26700 36916
rect 26752 36904 26758 36916
rect 28261 36907 28319 36913
rect 28261 36904 28273 36907
rect 26752 36876 28273 36904
rect 26752 36864 26758 36876
rect 28261 36873 28273 36876
rect 28307 36873 28319 36907
rect 28261 36867 28319 36873
rect 28905 36907 28963 36913
rect 28905 36873 28917 36907
rect 28951 36904 28963 36907
rect 32861 36907 32919 36913
rect 28951 36876 30144 36904
rect 28951 36873 28963 36876
rect 28905 36867 28963 36873
rect 26970 36836 26976 36848
rect 26931 36808 26976 36836
rect 26970 36796 26976 36808
rect 27028 36796 27034 36848
rect 27062 36796 27068 36848
rect 27120 36836 27126 36848
rect 27982 36836 27988 36848
rect 27120 36808 27988 36836
rect 27120 36796 27126 36808
rect 27249 36771 27307 36777
rect 27249 36768 27261 36771
rect 25240 36740 27261 36768
rect 27249 36737 27261 36740
rect 27295 36737 27307 36771
rect 27249 36731 27307 36737
rect 27341 36771 27399 36777
rect 27341 36737 27353 36771
rect 27387 36737 27399 36771
rect 27341 36731 27399 36737
rect 21818 36660 21824 36712
rect 21876 36700 21882 36712
rect 21913 36703 21971 36709
rect 21913 36700 21925 36703
rect 21876 36672 21925 36700
rect 21876 36660 21882 36672
rect 21913 36669 21925 36672
rect 21959 36669 21971 36703
rect 21913 36663 21971 36669
rect 26878 36660 26884 36712
rect 26936 36700 26942 36712
rect 27356 36700 27384 36731
rect 27430 36728 27436 36780
rect 27488 36768 27494 36780
rect 27632 36777 27660 36808
rect 27982 36796 27988 36808
rect 28040 36796 28046 36848
rect 28166 36836 28172 36848
rect 28127 36808 28172 36836
rect 28166 36796 28172 36808
rect 28224 36796 28230 36848
rect 28276 36836 28304 36867
rect 30116 36836 30144 36876
rect 32861 36873 32873 36907
rect 32907 36904 32919 36907
rect 33594 36904 33600 36916
rect 32907 36876 33600 36904
rect 32907 36873 32919 36876
rect 32861 36867 32919 36873
rect 33594 36864 33600 36876
rect 33652 36864 33658 36916
rect 35986 36904 35992 36916
rect 35947 36876 35992 36904
rect 35986 36864 35992 36876
rect 36044 36864 36050 36916
rect 30254 36839 30312 36845
rect 30254 36836 30266 36839
rect 28276 36808 30052 36836
rect 30116 36808 30266 36836
rect 27617 36771 27675 36777
rect 27488 36740 27533 36768
rect 27488 36728 27494 36740
rect 27617 36737 27629 36771
rect 27663 36737 27675 36771
rect 27617 36731 27675 36737
rect 28810 36728 28816 36780
rect 28868 36768 28874 36780
rect 29181 36771 29239 36777
rect 29181 36768 29193 36771
rect 28868 36740 29193 36768
rect 28868 36728 28874 36740
rect 29181 36737 29193 36740
rect 29227 36737 29239 36771
rect 29181 36731 29239 36737
rect 29273 36771 29331 36777
rect 29273 36737 29285 36771
rect 29319 36737 29331 36771
rect 29273 36731 29331 36737
rect 29288 36700 29316 36731
rect 29362 36728 29368 36780
rect 29420 36777 29426 36780
rect 29420 36768 29428 36777
rect 29420 36740 29465 36768
rect 29420 36731 29428 36740
rect 29420 36728 29426 36731
rect 29546 36728 29552 36780
rect 29604 36768 29610 36780
rect 30024 36777 30052 36808
rect 30254 36805 30266 36808
rect 30300 36805 30312 36839
rect 30254 36799 30312 36805
rect 33134 36796 33140 36848
rect 33192 36836 33198 36848
rect 34026 36839 34084 36845
rect 34026 36836 34038 36839
rect 33192 36808 34038 36836
rect 33192 36796 33198 36808
rect 34026 36805 34038 36808
rect 34072 36805 34084 36839
rect 34026 36799 34084 36805
rect 35526 36796 35532 36848
rect 35584 36836 35590 36848
rect 35805 36839 35863 36845
rect 35805 36836 35817 36839
rect 35584 36808 35817 36836
rect 35584 36796 35590 36808
rect 35805 36805 35817 36808
rect 35851 36836 35863 36839
rect 36998 36836 37004 36848
rect 35851 36808 37004 36836
rect 35851 36805 35863 36808
rect 35805 36799 35863 36805
rect 36998 36796 37004 36808
rect 37056 36796 37062 36848
rect 30009 36771 30067 36777
rect 29604 36740 29649 36768
rect 29604 36728 29610 36740
rect 30009 36737 30021 36771
rect 30055 36737 30067 36771
rect 30009 36731 30067 36737
rect 30098 36728 30104 36780
rect 30156 36768 30162 36780
rect 31386 36768 31392 36780
rect 30156 36740 31392 36768
rect 30156 36728 30162 36740
rect 31386 36728 31392 36740
rect 31444 36728 31450 36780
rect 31938 36728 31944 36780
rect 31996 36768 32002 36780
rect 32217 36771 32275 36777
rect 32217 36768 32229 36771
rect 31996 36740 32229 36768
rect 31996 36728 32002 36740
rect 32217 36737 32229 36740
rect 32263 36768 32275 36771
rect 32306 36768 32312 36780
rect 32263 36740 32312 36768
rect 32263 36737 32275 36740
rect 32217 36731 32275 36737
rect 32306 36728 32312 36740
rect 32364 36728 32370 36780
rect 32398 36728 32404 36780
rect 32456 36768 32462 36780
rect 33045 36771 33103 36777
rect 33045 36768 33057 36771
rect 32456 36740 33057 36768
rect 32456 36728 32462 36740
rect 33045 36737 33057 36740
rect 33091 36737 33103 36771
rect 33226 36768 33232 36780
rect 33187 36740 33232 36768
rect 33045 36731 33103 36737
rect 33226 36728 33232 36740
rect 33284 36728 33290 36780
rect 33318 36728 33324 36780
rect 33376 36768 33382 36780
rect 35618 36768 35624 36780
rect 33376 36740 33421 36768
rect 35579 36740 35624 36768
rect 33376 36728 33382 36740
rect 35618 36728 35624 36740
rect 35676 36728 35682 36780
rect 30116 36700 30144 36728
rect 26936 36672 30144 36700
rect 26936 36660 26942 36672
rect 31754 36660 31760 36712
rect 31812 36700 31818 36712
rect 33781 36703 33839 36709
rect 33781 36700 33793 36703
rect 31812 36672 33793 36700
rect 31812 36660 31818 36672
rect 33781 36669 33793 36672
rect 33827 36669 33839 36703
rect 33781 36663 33839 36669
rect 20027 36604 20944 36632
rect 20027 36601 20039 36604
rect 19981 36595 20039 36601
rect 20916 36564 20944 36604
rect 32401 36635 32459 36641
rect 32401 36601 32413 36635
rect 32447 36632 32459 36635
rect 33226 36632 33232 36644
rect 32447 36604 33232 36632
rect 32447 36601 32459 36604
rect 32401 36595 32459 36601
rect 33226 36592 33232 36604
rect 33284 36592 33290 36644
rect 23198 36564 23204 36576
rect 20916 36536 23204 36564
rect 23198 36524 23204 36536
rect 23256 36524 23262 36576
rect 23290 36524 23296 36576
rect 23348 36564 23354 36576
rect 28810 36564 28816 36576
rect 23348 36536 28816 36564
rect 23348 36524 23354 36536
rect 28810 36524 28816 36536
rect 28868 36524 28874 36576
rect 30742 36524 30748 36576
rect 30800 36564 30806 36576
rect 31389 36567 31447 36573
rect 31389 36564 31401 36567
rect 30800 36536 31401 36564
rect 30800 36524 30806 36536
rect 31389 36533 31401 36536
rect 31435 36533 31447 36567
rect 31389 36527 31447 36533
rect 33318 36524 33324 36576
rect 33376 36564 33382 36576
rect 35161 36567 35219 36573
rect 35161 36564 35173 36567
rect 33376 36536 35173 36564
rect 33376 36524 33382 36536
rect 35161 36533 35173 36536
rect 35207 36533 35219 36567
rect 35161 36527 35219 36533
rect 46290 36524 46296 36576
rect 46348 36564 46354 36576
rect 47765 36567 47823 36573
rect 47765 36564 47777 36567
rect 46348 36536 47777 36564
rect 46348 36524 46354 36536
rect 47765 36533 47777 36536
rect 47811 36533 47823 36567
rect 47765 36527 47823 36533
rect 1104 36474 48852 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 48852 36474
rect 1104 36400 48852 36422
rect 20530 36320 20536 36372
rect 20588 36360 20594 36372
rect 21085 36363 21143 36369
rect 21085 36360 21097 36363
rect 20588 36332 21097 36360
rect 20588 36320 20594 36332
rect 21085 36329 21097 36332
rect 21131 36360 21143 36363
rect 22462 36360 22468 36372
rect 21131 36332 22324 36360
rect 22423 36332 22468 36360
rect 21131 36329 21143 36332
rect 21085 36323 21143 36329
rect 21542 36252 21548 36304
rect 21600 36292 21606 36304
rect 22296 36292 22324 36332
rect 22462 36320 22468 36332
rect 22520 36320 22526 36372
rect 22738 36320 22744 36372
rect 22796 36360 22802 36372
rect 23290 36360 23296 36372
rect 22796 36332 23296 36360
rect 22796 36320 22802 36332
rect 23290 36320 23296 36332
rect 23348 36320 23354 36372
rect 24394 36360 24400 36372
rect 24355 36332 24400 36360
rect 24394 36320 24400 36332
rect 24452 36320 24458 36372
rect 26050 36320 26056 36372
rect 26108 36360 26114 36372
rect 28074 36360 28080 36372
rect 26108 36332 28080 36360
rect 26108 36320 26114 36332
rect 28074 36320 28080 36332
rect 28132 36320 28138 36372
rect 28166 36320 28172 36372
rect 28224 36360 28230 36372
rect 30837 36363 30895 36369
rect 30837 36360 30849 36363
rect 28224 36332 30849 36360
rect 28224 36320 28230 36332
rect 30837 36329 30849 36332
rect 30883 36329 30895 36363
rect 30837 36323 30895 36329
rect 23014 36292 23020 36304
rect 21600 36264 22094 36292
rect 22296 36264 23020 36292
rect 21600 36252 21606 36264
rect 20438 36224 20444 36236
rect 19536 36196 20444 36224
rect 2038 36116 2044 36168
rect 2096 36156 2102 36168
rect 2225 36159 2283 36165
rect 2225 36156 2237 36159
rect 2096 36128 2237 36156
rect 2096 36116 2102 36128
rect 2225 36125 2237 36128
rect 2271 36125 2283 36159
rect 2225 36119 2283 36125
rect 2869 36159 2927 36165
rect 2869 36125 2881 36159
rect 2915 36156 2927 36159
rect 16666 36156 16672 36168
rect 2915 36128 16672 36156
rect 2915 36125 2927 36128
rect 2869 36119 2927 36125
rect 16666 36116 16672 36128
rect 16724 36116 16730 36168
rect 19536 36165 19564 36196
rect 20438 36184 20444 36196
rect 20496 36184 20502 36236
rect 21560 36224 21588 36252
rect 20548 36196 21588 36224
rect 22066 36224 22094 36264
rect 23014 36252 23020 36264
rect 23072 36252 23078 36304
rect 23198 36252 23204 36304
rect 23256 36292 23262 36304
rect 28353 36295 28411 36301
rect 28353 36292 28365 36295
rect 23256 36264 25176 36292
rect 23256 36252 23262 36264
rect 22066 36196 25084 36224
rect 19521 36159 19579 36165
rect 19521 36125 19533 36159
rect 19567 36125 19579 36159
rect 19521 36119 19579 36125
rect 19613 36159 19671 36165
rect 19613 36125 19625 36159
rect 19659 36125 19671 36159
rect 19613 36119 19671 36125
rect 19705 36159 19763 36165
rect 19705 36125 19717 36159
rect 19751 36125 19763 36159
rect 19705 36119 19763 36125
rect 19889 36159 19947 36165
rect 19889 36125 19901 36159
rect 19935 36156 19947 36159
rect 20548 36156 20576 36196
rect 19935 36128 20576 36156
rect 20901 36159 20959 36165
rect 19935 36125 19947 36128
rect 19889 36119 19947 36125
rect 20901 36125 20913 36159
rect 20947 36156 20959 36159
rect 22738 36156 22744 36168
rect 20947 36128 21680 36156
rect 22699 36128 22744 36156
rect 20947 36125 20959 36128
rect 20901 36119 20959 36125
rect 19150 36048 19156 36100
rect 19208 36088 19214 36100
rect 19628 36088 19656 36119
rect 19208 36060 19656 36088
rect 19720 36088 19748 36119
rect 21652 36100 21680 36128
rect 22738 36116 22744 36128
rect 22796 36116 22802 36168
rect 22833 36159 22891 36165
rect 22833 36125 22845 36159
rect 22879 36125 22891 36159
rect 22833 36119 22891 36125
rect 20806 36088 20812 36100
rect 19720 36060 20812 36088
rect 19208 36048 19214 36060
rect 2958 36020 2964 36032
rect 2919 35992 2964 36020
rect 2958 35980 2964 35992
rect 3016 35980 3022 36032
rect 19242 36020 19248 36032
rect 19203 35992 19248 36020
rect 19242 35980 19248 35992
rect 19300 35980 19306 36032
rect 19628 36020 19656 36060
rect 20806 36048 20812 36060
rect 20864 36048 20870 36100
rect 21634 36048 21640 36100
rect 21692 36088 21698 36100
rect 21729 36091 21787 36097
rect 21729 36088 21741 36091
rect 21692 36060 21741 36088
rect 21692 36048 21698 36060
rect 21729 36057 21741 36060
rect 21775 36057 21787 36091
rect 21729 36051 21787 36057
rect 21821 36023 21879 36029
rect 21821 36020 21833 36023
rect 19628 35992 21833 36020
rect 21821 35989 21833 35992
rect 21867 36020 21879 36023
rect 21910 36020 21916 36032
rect 21867 35992 21916 36020
rect 21867 35989 21879 35992
rect 21821 35983 21879 35989
rect 21910 35980 21916 35992
rect 21968 36020 21974 36032
rect 22848 36020 22876 36119
rect 22922 36116 22928 36168
rect 22980 36156 22986 36168
rect 23124 36165 23152 36196
rect 23109 36159 23167 36165
rect 22980 36128 23025 36156
rect 22980 36116 22986 36128
rect 23109 36125 23121 36159
rect 23155 36125 23167 36159
rect 24670 36156 24676 36168
rect 24631 36128 24676 36156
rect 23109 36119 23167 36125
rect 24670 36116 24676 36128
rect 24728 36116 24734 36168
rect 24765 36159 24823 36165
rect 24765 36125 24777 36159
rect 24811 36125 24823 36159
rect 24765 36119 24823 36125
rect 23014 36048 23020 36100
rect 23072 36088 23078 36100
rect 24780 36088 24808 36119
rect 24854 36116 24860 36168
rect 24912 36156 24918 36168
rect 25056 36165 25084 36196
rect 25041 36159 25099 36165
rect 24912 36128 24957 36156
rect 24912 36116 24918 36128
rect 25041 36125 25053 36159
rect 25087 36125 25099 36159
rect 25148 36156 25176 36264
rect 26160 36264 28365 36292
rect 26160 36165 26188 36264
rect 28353 36261 28365 36264
rect 28399 36261 28411 36295
rect 28353 36255 28411 36261
rect 29546 36252 29552 36304
rect 29604 36292 29610 36304
rect 29604 36264 30236 36292
rect 29604 36252 29610 36264
rect 27246 36224 27252 36236
rect 27207 36196 27252 36224
rect 27246 36184 27252 36196
rect 27304 36184 27310 36236
rect 27433 36227 27491 36233
rect 27433 36193 27445 36227
rect 27479 36224 27491 36227
rect 27522 36224 27528 36236
rect 27479 36196 27528 36224
rect 27479 36193 27491 36196
rect 27433 36187 27491 36193
rect 27522 36184 27528 36196
rect 27580 36184 27586 36236
rect 27982 36184 27988 36236
rect 28040 36224 28046 36236
rect 28040 36196 28948 36224
rect 28040 36184 28046 36196
rect 25961 36159 26019 36165
rect 25961 36156 25973 36159
rect 25148 36128 25973 36156
rect 25041 36119 25099 36125
rect 25961 36125 25973 36128
rect 26007 36125 26019 36159
rect 25961 36119 26019 36125
rect 26053 36159 26111 36165
rect 26053 36125 26065 36159
rect 26099 36125 26111 36159
rect 26053 36119 26111 36125
rect 26145 36159 26203 36165
rect 26145 36125 26157 36159
rect 26191 36125 26203 36159
rect 26145 36119 26203 36125
rect 26329 36159 26387 36165
rect 26329 36125 26341 36159
rect 26375 36156 26387 36159
rect 27062 36156 27068 36168
rect 26375 36128 27068 36156
rect 26375 36125 26387 36128
rect 26329 36119 26387 36125
rect 24946 36088 24952 36100
rect 23072 36060 24952 36088
rect 23072 36048 23078 36060
rect 24946 36048 24952 36060
rect 25004 36048 25010 36100
rect 26068 36088 26096 36119
rect 27062 36116 27068 36128
rect 27120 36116 27126 36168
rect 27157 36159 27215 36165
rect 27157 36125 27169 36159
rect 27203 36156 27215 36159
rect 28350 36156 28356 36168
rect 27203 36128 28356 36156
rect 27203 36125 27215 36128
rect 27157 36119 27215 36125
rect 28350 36116 28356 36128
rect 28408 36116 28414 36168
rect 28920 36156 28948 36196
rect 29805 36159 29863 36165
rect 28920 36153 29776 36156
rect 29805 36153 29817 36159
rect 28920 36128 29817 36153
rect 29748 36125 29817 36128
rect 29851 36125 29863 36159
rect 29805 36119 29863 36125
rect 29914 36153 29972 36159
rect 29914 36119 29926 36153
rect 29960 36150 29972 36153
rect 29960 36119 29973 36150
rect 29914 36113 29973 36119
rect 30006 36116 30012 36168
rect 30064 36165 30070 36168
rect 30208 36165 30236 36264
rect 30064 36156 30072 36165
rect 30193 36159 30251 36165
rect 30064 36128 30109 36156
rect 30064 36119 30072 36128
rect 30193 36125 30205 36159
rect 30239 36156 30251 36159
rect 30558 36156 30564 36168
rect 30239 36128 30564 36156
rect 30239 36125 30251 36128
rect 30193 36119 30251 36125
rect 30064 36116 30070 36119
rect 30558 36116 30564 36128
rect 30616 36116 30622 36168
rect 30852 36156 30880 36323
rect 33226 36320 33232 36372
rect 33284 36360 33290 36372
rect 34698 36360 34704 36372
rect 33284 36332 34704 36360
rect 33284 36320 33290 36332
rect 34698 36320 34704 36332
rect 34756 36320 34762 36372
rect 35894 36360 35900 36372
rect 35636 36332 35900 36360
rect 31665 36295 31723 36301
rect 31665 36261 31677 36295
rect 31711 36292 31723 36295
rect 31754 36292 31760 36304
rect 31711 36264 31760 36292
rect 31711 36261 31723 36264
rect 31665 36255 31723 36261
rect 31754 36252 31760 36264
rect 31812 36252 31818 36304
rect 35636 36233 35664 36332
rect 35894 36320 35900 36332
rect 35952 36320 35958 36372
rect 36998 36360 37004 36372
rect 36959 36332 37004 36360
rect 36998 36320 37004 36332
rect 37056 36320 37062 36372
rect 35621 36227 35679 36233
rect 35621 36193 35633 36227
rect 35667 36193 35679 36227
rect 46290 36224 46296 36236
rect 46251 36196 46296 36224
rect 35621 36187 35679 36193
rect 46290 36184 46296 36196
rect 46348 36184 46354 36236
rect 48130 36224 48136 36236
rect 48091 36196 48136 36224
rect 48130 36184 48136 36196
rect 48188 36184 48194 36236
rect 31481 36159 31539 36165
rect 31481 36156 31493 36159
rect 30852 36128 31493 36156
rect 31481 36125 31493 36128
rect 31527 36125 31539 36159
rect 31481 36119 31539 36125
rect 35710 36116 35716 36168
rect 35768 36156 35774 36168
rect 35877 36159 35935 36165
rect 35877 36156 35889 36159
rect 35768 36128 35889 36156
rect 35768 36116 35774 36128
rect 35877 36125 35889 36128
rect 35923 36125 35935 36159
rect 35877 36119 35935 36125
rect 26234 36088 26240 36100
rect 26068 36060 26240 36088
rect 26234 36048 26240 36060
rect 26292 36048 26298 36100
rect 27985 36091 28043 36097
rect 27985 36088 27997 36091
rect 26804 36060 27997 36088
rect 21968 35992 22876 36020
rect 25685 36023 25743 36029
rect 21968 35980 21974 35992
rect 25685 35989 25697 36023
rect 25731 36020 25743 36023
rect 26602 36020 26608 36032
rect 25731 35992 26608 36020
rect 25731 35989 25743 35992
rect 25685 35983 25743 35989
rect 26602 35980 26608 35992
rect 26660 35980 26666 36032
rect 26804 36029 26832 36060
rect 27985 36057 27997 36060
rect 28031 36057 28043 36091
rect 28166 36088 28172 36100
rect 28127 36060 28172 36088
rect 27985 36051 28043 36057
rect 28166 36048 28172 36060
rect 28224 36048 28230 36100
rect 29945 36088 29973 36113
rect 30098 36088 30104 36100
rect 29945 36060 30104 36088
rect 30098 36048 30104 36060
rect 30156 36048 30162 36100
rect 30742 36088 30748 36100
rect 30703 36060 30748 36088
rect 30742 36048 30748 36060
rect 30800 36048 30806 36100
rect 46477 36091 46535 36097
rect 46477 36057 46489 36091
rect 46523 36088 46535 36091
rect 47670 36088 47676 36100
rect 46523 36060 47676 36088
rect 46523 36057 46535 36060
rect 46477 36051 46535 36057
rect 47670 36048 47676 36060
rect 47728 36048 47734 36100
rect 26789 36023 26847 36029
rect 26789 35989 26801 36023
rect 26835 35989 26847 36023
rect 26789 35983 26847 35989
rect 29549 36023 29607 36029
rect 29549 35989 29561 36023
rect 29595 36020 29607 36023
rect 29822 36020 29828 36032
rect 29595 35992 29828 36020
rect 29595 35989 29607 35992
rect 29549 35983 29607 35989
rect 29822 35980 29828 35992
rect 29880 35980 29886 36032
rect 30190 35980 30196 36032
rect 30248 36020 30254 36032
rect 33318 36020 33324 36032
rect 30248 35992 33324 36020
rect 30248 35980 30254 35992
rect 33318 35980 33324 35992
rect 33376 35980 33382 36032
rect 1104 35930 48852 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 48852 35930
rect 1104 35856 48852 35878
rect 19981 35819 20039 35825
rect 19981 35785 19993 35819
rect 20027 35785 20039 35819
rect 20806 35816 20812 35828
rect 20767 35788 20812 35816
rect 19981 35779 20039 35785
rect 2225 35751 2283 35757
rect 2225 35717 2237 35751
rect 2271 35748 2283 35751
rect 2958 35748 2964 35760
rect 2271 35720 2964 35748
rect 2271 35717 2283 35720
rect 2225 35711 2283 35717
rect 2958 35708 2964 35720
rect 3016 35708 3022 35760
rect 18868 35751 18926 35757
rect 18868 35717 18880 35751
rect 18914 35748 18926 35751
rect 19242 35748 19248 35760
rect 18914 35720 19248 35748
rect 18914 35717 18926 35720
rect 18868 35711 18926 35717
rect 19242 35708 19248 35720
rect 19300 35708 19306 35760
rect 19996 35748 20024 35779
rect 20806 35776 20812 35788
rect 20864 35776 20870 35828
rect 27982 35816 27988 35828
rect 22066 35788 27988 35816
rect 20625 35751 20683 35757
rect 20625 35748 20637 35751
rect 19996 35720 20637 35748
rect 20625 35717 20637 35720
rect 20671 35748 20683 35751
rect 22066 35748 22094 35788
rect 27982 35776 27988 35788
rect 28040 35776 28046 35828
rect 28350 35816 28356 35828
rect 28311 35788 28356 35816
rect 28350 35776 28356 35788
rect 28408 35776 28414 35828
rect 29825 35819 29883 35825
rect 29825 35816 29837 35819
rect 29012 35788 29837 35816
rect 20671 35720 22094 35748
rect 24673 35751 24731 35757
rect 20671 35717 20683 35720
rect 20625 35711 20683 35717
rect 24673 35717 24685 35751
rect 24719 35748 24731 35751
rect 26237 35751 26295 35757
rect 26237 35748 26249 35751
rect 24719 35720 26249 35748
rect 24719 35717 24731 35720
rect 24673 35711 24731 35717
rect 26237 35717 26249 35720
rect 26283 35748 26295 35751
rect 26418 35748 26424 35760
rect 26283 35720 26424 35748
rect 26283 35717 26295 35720
rect 26237 35711 26295 35717
rect 26418 35708 26424 35720
rect 26476 35708 26482 35760
rect 26602 35708 26608 35760
rect 26660 35748 26666 35760
rect 29012 35757 29040 35788
rect 29825 35785 29837 35788
rect 29871 35785 29883 35819
rect 29825 35779 29883 35785
rect 29914 35776 29920 35828
rect 29972 35816 29978 35828
rect 30193 35819 30251 35825
rect 30193 35816 30205 35819
rect 29972 35788 30205 35816
rect 29972 35776 29978 35788
rect 30193 35785 30205 35788
rect 30239 35785 30251 35819
rect 30193 35779 30251 35785
rect 27218 35751 27276 35757
rect 27218 35748 27230 35751
rect 26660 35720 27230 35748
rect 26660 35708 26666 35720
rect 27218 35717 27230 35720
rect 27264 35717 27276 35751
rect 27218 35711 27276 35717
rect 28997 35751 29055 35757
rect 28997 35717 29009 35751
rect 29043 35717 29055 35751
rect 28997 35711 29055 35717
rect 29365 35751 29423 35757
rect 29365 35717 29377 35751
rect 29411 35748 29423 35751
rect 30098 35748 30104 35760
rect 29411 35720 30104 35748
rect 29411 35717 29423 35720
rect 29365 35711 29423 35717
rect 30098 35708 30104 35720
rect 30156 35708 30162 35760
rect 31113 35751 31171 35757
rect 31113 35748 31125 35751
rect 30484 35720 31125 35748
rect 2038 35680 2044 35692
rect 1999 35652 2044 35680
rect 2038 35640 2044 35652
rect 2096 35640 2102 35692
rect 11698 35640 11704 35692
rect 11756 35680 11762 35692
rect 19426 35680 19432 35692
rect 11756 35652 19432 35680
rect 11756 35640 11762 35652
rect 19426 35640 19432 35652
rect 19484 35640 19490 35692
rect 20438 35680 20444 35692
rect 20399 35652 20444 35680
rect 20438 35640 20444 35652
rect 20496 35640 20502 35692
rect 21450 35640 21456 35692
rect 21508 35680 21514 35692
rect 21821 35683 21879 35689
rect 21821 35680 21833 35683
rect 21508 35652 21833 35680
rect 21508 35640 21514 35652
rect 21821 35649 21833 35652
rect 21867 35680 21879 35683
rect 22557 35683 22615 35689
rect 22557 35680 22569 35683
rect 21867 35652 22569 35680
rect 21867 35649 21879 35652
rect 21821 35643 21879 35649
rect 22557 35649 22569 35652
rect 22603 35680 22615 35683
rect 24489 35683 24547 35689
rect 24489 35680 24501 35683
rect 22603 35652 24501 35680
rect 22603 35649 22615 35652
rect 22557 35643 22615 35649
rect 24489 35649 24501 35652
rect 24535 35649 24547 35683
rect 24489 35643 24547 35649
rect 26694 35640 26700 35692
rect 26752 35680 26758 35692
rect 26973 35683 27031 35689
rect 26973 35680 26985 35683
rect 26752 35652 26985 35680
rect 26752 35640 26758 35652
rect 26973 35649 26985 35652
rect 27019 35649 27031 35683
rect 26973 35643 27031 35649
rect 29181 35683 29239 35689
rect 29181 35649 29193 35683
rect 29227 35680 29239 35683
rect 29730 35680 29736 35692
rect 29227 35652 29736 35680
rect 29227 35649 29239 35652
rect 29181 35643 29239 35649
rect 2774 35612 2780 35624
rect 2735 35584 2780 35612
rect 2774 35572 2780 35584
rect 2832 35572 2838 35624
rect 18598 35612 18604 35624
rect 18559 35584 18604 35612
rect 18598 35572 18604 35584
rect 18656 35572 18662 35624
rect 26234 35572 26240 35624
rect 26292 35612 26298 35624
rect 26421 35615 26479 35621
rect 26421 35612 26433 35615
rect 26292 35584 26433 35612
rect 26292 35572 26298 35584
rect 26421 35581 26433 35584
rect 26467 35612 26479 35615
rect 26878 35612 26884 35624
rect 26467 35584 26884 35612
rect 26467 35581 26479 35584
rect 26421 35575 26479 35581
rect 26878 35572 26884 35584
rect 26936 35572 26942 35624
rect 28166 35572 28172 35624
rect 28224 35612 28230 35624
rect 29196 35612 29224 35643
rect 29730 35640 29736 35652
rect 29788 35640 29794 35692
rect 30484 35680 30512 35720
rect 31113 35717 31125 35720
rect 31159 35717 31171 35751
rect 31294 35748 31300 35760
rect 31255 35720 31300 35748
rect 31113 35711 31171 35717
rect 31294 35708 31300 35720
rect 31352 35708 31358 35760
rect 31386 35708 31392 35760
rect 31444 35748 31450 35760
rect 31444 35720 32536 35748
rect 31444 35708 31450 35720
rect 30024 35652 30512 35680
rect 28224 35584 29224 35612
rect 28224 35572 28230 35584
rect 22741 35547 22799 35553
rect 22741 35513 22753 35547
rect 22787 35544 22799 35547
rect 22830 35544 22836 35556
rect 22787 35516 22836 35544
rect 22787 35513 22799 35516
rect 22741 35507 22799 35513
rect 22830 35504 22836 35516
rect 22888 35504 22894 35556
rect 28902 35504 28908 35556
rect 28960 35544 28966 35556
rect 30024 35544 30052 35652
rect 31478 35640 31484 35692
rect 31536 35680 31542 35692
rect 32508 35689 32536 35720
rect 32355 35683 32413 35689
rect 32355 35680 32367 35683
rect 31536 35652 32367 35680
rect 31536 35640 31542 35652
rect 32355 35649 32367 35652
rect 32401 35649 32413 35683
rect 32355 35643 32413 35649
rect 32493 35683 32551 35689
rect 32493 35649 32505 35683
rect 32539 35649 32551 35683
rect 32606 35683 32664 35689
rect 32606 35680 32618 35683
rect 32493 35643 32551 35649
rect 32600 35649 32618 35680
rect 32652 35649 32664 35683
rect 32600 35643 32664 35649
rect 32769 35683 32827 35689
rect 32769 35649 32781 35683
rect 32815 35649 32827 35683
rect 47854 35680 47860 35692
rect 47815 35652 47860 35680
rect 32769 35643 32827 35649
rect 30190 35572 30196 35624
rect 30248 35612 30254 35624
rect 30285 35615 30343 35621
rect 30285 35612 30297 35615
rect 30248 35584 30297 35612
rect 30248 35572 30254 35584
rect 30285 35581 30297 35584
rect 30331 35581 30343 35615
rect 30466 35612 30472 35624
rect 30427 35584 30472 35612
rect 30285 35575 30343 35581
rect 30466 35572 30472 35584
rect 30524 35572 30530 35624
rect 32030 35572 32036 35624
rect 32088 35612 32094 35624
rect 32600 35612 32628 35643
rect 32088 35584 32628 35612
rect 32088 35572 32094 35584
rect 28960 35516 30052 35544
rect 28960 35504 28966 35516
rect 30558 35504 30564 35556
rect 30616 35544 30622 35556
rect 32582 35544 32588 35556
rect 30616 35516 32588 35544
rect 30616 35504 30622 35516
rect 32582 35504 32588 35516
rect 32640 35544 32646 35556
rect 32784 35544 32812 35643
rect 47854 35640 47860 35652
rect 47912 35640 47918 35692
rect 32640 35516 32812 35544
rect 32640 35504 32646 35516
rect 1578 35436 1584 35488
rect 1636 35476 1642 35488
rect 2590 35476 2596 35488
rect 1636 35448 2596 35476
rect 1636 35436 1642 35448
rect 2590 35436 2596 35448
rect 2648 35436 2654 35488
rect 15838 35436 15844 35488
rect 15896 35476 15902 35488
rect 20806 35476 20812 35488
rect 15896 35448 20812 35476
rect 15896 35436 15902 35448
rect 20806 35436 20812 35448
rect 20864 35436 20870 35488
rect 21542 35436 21548 35488
rect 21600 35476 21606 35488
rect 22002 35476 22008 35488
rect 21600 35448 22008 35476
rect 21600 35436 21606 35448
rect 22002 35436 22008 35448
rect 22060 35436 22066 35488
rect 32122 35476 32128 35488
rect 32083 35448 32128 35476
rect 32122 35436 32128 35448
rect 32180 35436 32186 35488
rect 46290 35436 46296 35488
rect 46348 35476 46354 35488
rect 46385 35479 46443 35485
rect 46385 35476 46397 35479
rect 46348 35448 46397 35476
rect 46348 35436 46354 35448
rect 46385 35445 46397 35448
rect 46431 35445 46443 35479
rect 47026 35476 47032 35488
rect 46987 35448 47032 35476
rect 46385 35439 46443 35445
rect 47026 35436 47032 35448
rect 47084 35436 47090 35488
rect 48038 35476 48044 35488
rect 47999 35448 48044 35476
rect 48038 35436 48044 35448
rect 48096 35436 48102 35488
rect 1104 35386 48852 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 48852 35386
rect 1104 35312 48852 35334
rect 17770 35232 17776 35284
rect 17828 35272 17834 35284
rect 17828 35244 20760 35272
rect 17828 35232 17834 35244
rect 5350 35164 5356 35216
rect 5408 35204 5414 35216
rect 15838 35204 15844 35216
rect 5408 35176 15844 35204
rect 5408 35164 5414 35176
rect 15838 35164 15844 35176
rect 15896 35164 15902 35216
rect 1673 35139 1731 35145
rect 1673 35105 1685 35139
rect 1719 35136 1731 35139
rect 11698 35136 11704 35148
rect 1719 35108 11704 35136
rect 1719 35105 1731 35108
rect 1673 35099 1731 35105
rect 11698 35096 11704 35108
rect 11756 35096 11762 35148
rect 20732 35136 20760 35244
rect 20806 35232 20812 35284
rect 20864 35272 20870 35284
rect 20864 35244 22094 35272
rect 20864 35232 20870 35244
rect 22066 35204 22094 35244
rect 27522 35232 27528 35284
rect 27580 35272 27586 35284
rect 28445 35275 28503 35281
rect 28445 35272 28457 35275
rect 27580 35244 28457 35272
rect 27580 35232 27586 35244
rect 28445 35241 28457 35244
rect 28491 35241 28503 35275
rect 31941 35275 31999 35281
rect 28445 35235 28503 35241
rect 29564 35244 31708 35272
rect 29362 35204 29368 35216
rect 22066 35176 29368 35204
rect 29362 35164 29368 35176
rect 29420 35164 29426 35216
rect 21450 35136 21456 35148
rect 20732 35108 21456 35136
rect 21450 35096 21456 35108
rect 21508 35096 21514 35148
rect 26881 35139 26939 35145
rect 26881 35105 26893 35139
rect 26927 35136 26939 35139
rect 28166 35136 28172 35148
rect 26927 35108 28172 35136
rect 26927 35105 26939 35108
rect 26881 35099 26939 35105
rect 28166 35096 28172 35108
rect 28224 35096 28230 35148
rect 1394 35068 1400 35080
rect 1355 35040 1400 35068
rect 1394 35028 1400 35040
rect 1452 35028 1458 35080
rect 15194 35028 15200 35080
rect 15252 35068 15258 35080
rect 17957 35071 18015 35077
rect 17957 35068 17969 35071
rect 15252 35040 17969 35068
rect 15252 35028 15258 35040
rect 17957 35037 17969 35040
rect 18003 35068 18015 35071
rect 18598 35068 18604 35080
rect 18003 35040 18604 35068
rect 18003 35037 18015 35040
rect 17957 35031 18015 35037
rect 18598 35028 18604 35040
rect 18656 35068 18662 35080
rect 19150 35068 19156 35080
rect 18656 35040 19156 35068
rect 18656 35028 18662 35040
rect 19150 35028 19156 35040
rect 19208 35068 19214 35080
rect 19245 35071 19303 35077
rect 19245 35068 19257 35071
rect 19208 35040 19257 35068
rect 19208 35028 19214 35040
rect 19245 35037 19257 35040
rect 19291 35037 19303 35071
rect 19978 35068 19984 35080
rect 19245 35031 19303 35037
rect 19444 35040 19984 35068
rect 17773 35003 17831 35009
rect 17773 34969 17785 35003
rect 17819 35000 17831 35003
rect 19444 35000 19472 35040
rect 19978 35028 19984 35040
rect 20036 35028 20042 35080
rect 21634 35028 21640 35080
rect 21692 35068 21698 35080
rect 21729 35071 21787 35077
rect 21729 35068 21741 35071
rect 21692 35040 21741 35068
rect 21692 35028 21698 35040
rect 21729 35037 21741 35040
rect 21775 35068 21787 35071
rect 22554 35068 22560 35080
rect 21775 35040 22560 35068
rect 21775 35037 21787 35040
rect 21729 35031 21787 35037
rect 22554 35028 22560 35040
rect 22612 35028 22618 35080
rect 23474 35068 23480 35080
rect 23435 35040 23480 35068
rect 23474 35028 23480 35040
rect 23532 35068 23538 35080
rect 23842 35068 23848 35080
rect 23532 35040 23848 35068
rect 23532 35028 23538 35040
rect 23842 35028 23848 35040
rect 23900 35028 23906 35080
rect 26234 35068 26240 35080
rect 24872 35040 26240 35068
rect 17819 34972 19472 35000
rect 19512 35003 19570 35009
rect 17819 34969 17831 34972
rect 17773 34963 17831 34969
rect 19512 34969 19524 35003
rect 19558 34969 19570 35003
rect 19512 34963 19570 34969
rect 18690 34892 18696 34944
rect 18748 34932 18754 34944
rect 19536 34932 19564 34963
rect 22646 34960 22652 35012
rect 22704 35000 22710 35012
rect 24872 35009 24900 35040
rect 26234 35028 26240 35040
rect 26292 35068 26298 35080
rect 29564 35077 29592 35244
rect 31680 35136 31708 35244
rect 31941 35241 31953 35275
rect 31987 35272 31999 35275
rect 32030 35272 32036 35284
rect 31987 35244 32036 35272
rect 31987 35241 31999 35244
rect 31941 35235 31999 35241
rect 32030 35232 32036 35244
rect 32088 35232 32094 35284
rect 31754 35136 31760 35148
rect 31680 35108 31760 35136
rect 31754 35096 31760 35108
rect 31812 35136 31818 35148
rect 32401 35139 32459 35145
rect 32401 35136 32413 35139
rect 31812 35108 32413 35136
rect 31812 35096 31818 35108
rect 32401 35105 32413 35108
rect 32447 35105 32459 35139
rect 46290 35136 46296 35148
rect 46251 35108 46296 35136
rect 32401 35099 32459 35105
rect 46290 35096 46296 35108
rect 46348 35096 46354 35148
rect 48130 35136 48136 35148
rect 48091 35108 48136 35136
rect 48130 35096 48136 35108
rect 48188 35096 48194 35148
rect 26605 35071 26663 35077
rect 26605 35068 26617 35071
rect 26292 35040 26617 35068
rect 26292 35028 26298 35040
rect 26605 35037 26617 35040
rect 26651 35037 26663 35071
rect 26605 35031 26663 35037
rect 28261 35071 28319 35077
rect 28261 35037 28273 35071
rect 28307 35037 28319 35071
rect 28261 35031 28319 35037
rect 29549 35071 29607 35077
rect 29549 35037 29561 35071
rect 29595 35037 29607 35071
rect 29549 35031 29607 35037
rect 23293 35003 23351 35009
rect 23293 35000 23305 35003
rect 22704 34972 23305 35000
rect 22704 34960 22710 34972
rect 23293 34969 23305 34972
rect 23339 35000 23351 35003
rect 24857 35003 24915 35009
rect 24857 35000 24869 35003
rect 23339 34972 24869 35000
rect 23339 34969 23351 34972
rect 23293 34963 23351 34969
rect 24857 34969 24869 34972
rect 24903 34969 24915 35003
rect 24857 34963 24915 34969
rect 25041 35003 25099 35009
rect 25041 34969 25053 35003
rect 25087 35000 25099 35003
rect 26326 35000 26332 35012
rect 25087 34972 26332 35000
rect 25087 34969 25099 34972
rect 25041 34963 25099 34969
rect 26326 34960 26332 34972
rect 26384 35000 26390 35012
rect 26970 35000 26976 35012
rect 26384 34972 26976 35000
rect 26384 34960 26390 34972
rect 26970 34960 26976 34972
rect 27028 34960 27034 35012
rect 28276 35000 28304 35031
rect 32122 35028 32128 35080
rect 32180 35068 32186 35080
rect 32657 35071 32715 35077
rect 32657 35068 32669 35071
rect 32180 35040 32669 35068
rect 32180 35028 32186 35040
rect 32657 35037 32669 35040
rect 32703 35037 32715 35071
rect 32657 35031 32715 35037
rect 45554 35028 45560 35080
rect 45612 35068 45618 35080
rect 45649 35071 45707 35077
rect 45649 35068 45661 35071
rect 45612 35040 45661 35068
rect 45612 35028 45618 35040
rect 45649 35037 45661 35040
rect 45695 35037 45707 35071
rect 45649 35031 45707 35037
rect 28718 35000 28724 35012
rect 28276 34972 28724 35000
rect 28718 34960 28724 34972
rect 28776 35000 28782 35012
rect 29638 35000 29644 35012
rect 28776 34972 29644 35000
rect 28776 34960 28782 34972
rect 29638 34960 29644 34972
rect 29696 34960 29702 35012
rect 29822 35009 29828 35012
rect 29816 35000 29828 35009
rect 29783 34972 29828 35000
rect 29816 34963 29828 34972
rect 29822 34960 29828 34963
rect 29880 34960 29886 35012
rect 31570 35000 31576 35012
rect 31531 34972 31576 35000
rect 31570 34960 31576 34972
rect 31628 34960 31634 35012
rect 31757 35003 31815 35009
rect 31757 34969 31769 35003
rect 31803 35000 31815 35003
rect 32030 35000 32036 35012
rect 31803 34972 32036 35000
rect 31803 34969 31815 34972
rect 31757 34963 31815 34969
rect 32030 34960 32036 34972
rect 32088 34960 32094 35012
rect 45741 35003 45799 35009
rect 45741 34969 45753 35003
rect 45787 35000 45799 35003
rect 46477 35003 46535 35009
rect 46477 35000 46489 35003
rect 45787 34972 46489 35000
rect 45787 34969 45799 34972
rect 45741 34963 45799 34969
rect 46477 34969 46489 34972
rect 46523 34969 46535 35003
rect 46477 34963 46535 34969
rect 20622 34932 20628 34944
rect 18748 34904 19564 34932
rect 20535 34904 20628 34932
rect 18748 34892 18754 34904
rect 20622 34892 20628 34904
rect 20680 34932 20686 34944
rect 23198 34932 23204 34944
rect 20680 34904 23204 34932
rect 20680 34892 20686 34904
rect 23198 34892 23204 34904
rect 23256 34892 23262 34944
rect 29546 34892 29552 34944
rect 29604 34932 29610 34944
rect 29914 34932 29920 34944
rect 29604 34904 29920 34932
rect 29604 34892 29610 34904
rect 29914 34892 29920 34904
rect 29972 34932 29978 34944
rect 30929 34935 30987 34941
rect 30929 34932 30941 34935
rect 29972 34904 30941 34932
rect 29972 34892 29978 34904
rect 30929 34901 30941 34904
rect 30975 34901 30987 34935
rect 30929 34895 30987 34901
rect 33226 34892 33232 34944
rect 33284 34932 33290 34944
rect 33781 34935 33839 34941
rect 33781 34932 33793 34935
rect 33284 34904 33793 34932
rect 33284 34892 33290 34904
rect 33781 34901 33793 34904
rect 33827 34901 33839 34935
rect 33781 34895 33839 34901
rect 1104 34842 48852 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 48852 34842
rect 1104 34768 48852 34790
rect 12986 34688 12992 34740
rect 13044 34728 13050 34740
rect 18690 34728 18696 34740
rect 13044 34700 17908 34728
rect 18651 34700 18696 34728
rect 13044 34688 13050 34700
rect 15838 34660 15844 34672
rect 15799 34632 15844 34660
rect 15838 34620 15844 34632
rect 15896 34620 15902 34672
rect 2038 34592 2044 34604
rect 1951 34564 2044 34592
rect 2038 34552 2044 34564
rect 2096 34592 2102 34604
rect 3050 34592 3056 34604
rect 2096 34564 3056 34592
rect 2096 34552 2102 34564
rect 3050 34552 3056 34564
rect 3108 34552 3114 34604
rect 14185 34595 14243 34601
rect 14185 34561 14197 34595
rect 14231 34592 14243 34595
rect 15194 34592 15200 34604
rect 14231 34564 15200 34592
rect 14231 34561 14243 34564
rect 14185 34555 14243 34561
rect 15194 34552 15200 34564
rect 15252 34552 15258 34604
rect 16945 34595 17003 34601
rect 16945 34561 16957 34595
rect 16991 34592 17003 34595
rect 17589 34595 17647 34601
rect 17589 34592 17601 34595
rect 16991 34564 17601 34592
rect 16991 34561 17003 34564
rect 16945 34555 17003 34561
rect 17589 34561 17601 34564
rect 17635 34592 17647 34595
rect 17678 34592 17684 34604
rect 17635 34564 17684 34592
rect 17635 34561 17647 34564
rect 17589 34555 17647 34561
rect 17678 34552 17684 34564
rect 17736 34552 17742 34604
rect 17773 34595 17831 34601
rect 17773 34561 17785 34595
rect 17819 34561 17831 34595
rect 17880 34592 17908 34700
rect 18690 34688 18696 34700
rect 18748 34688 18754 34740
rect 19058 34688 19064 34740
rect 19116 34728 19122 34740
rect 22278 34728 22284 34740
rect 19116 34700 22284 34728
rect 19116 34688 19122 34700
rect 19242 34660 19248 34672
rect 19076 34632 19248 34660
rect 19076 34601 19104 34632
rect 19242 34620 19248 34632
rect 19300 34620 19306 34672
rect 19352 34601 19380 34700
rect 22278 34688 22284 34700
rect 22336 34688 22342 34740
rect 23198 34688 23204 34740
rect 23256 34728 23262 34740
rect 31478 34728 31484 34740
rect 23256 34700 31484 34728
rect 23256 34688 23262 34700
rect 31478 34688 31484 34700
rect 31536 34688 31542 34740
rect 31570 34688 31576 34740
rect 31628 34728 31634 34740
rect 32769 34731 32827 34737
rect 32769 34728 32781 34731
rect 31628 34700 32781 34728
rect 31628 34688 31634 34700
rect 32769 34697 32781 34700
rect 32815 34697 32827 34731
rect 47670 34728 47676 34740
rect 47631 34700 47676 34728
rect 32769 34691 32827 34697
rect 47670 34688 47676 34700
rect 47728 34688 47734 34740
rect 19981 34663 20039 34669
rect 19981 34629 19993 34663
rect 20027 34660 20039 34663
rect 20622 34660 20628 34672
rect 20027 34632 20628 34660
rect 20027 34629 20039 34632
rect 19981 34623 20039 34629
rect 20622 34620 20628 34632
rect 20680 34620 20686 34672
rect 21085 34663 21143 34669
rect 21085 34629 21097 34663
rect 21131 34660 21143 34663
rect 26421 34663 26479 34669
rect 21131 34632 23244 34660
rect 21131 34629 21143 34632
rect 21085 34623 21143 34629
rect 18969 34595 19027 34601
rect 18969 34592 18981 34595
rect 17880 34564 18981 34592
rect 17773 34555 17831 34561
rect 18969 34561 18981 34564
rect 19015 34561 19027 34595
rect 18969 34555 19027 34561
rect 19061 34595 19119 34601
rect 19061 34561 19073 34595
rect 19107 34561 19119 34595
rect 19061 34555 19119 34561
rect 19153 34595 19211 34601
rect 19153 34561 19165 34595
rect 19199 34561 19211 34595
rect 19153 34555 19211 34561
rect 19337 34595 19395 34601
rect 19337 34561 19349 34595
rect 19383 34561 19395 34595
rect 19337 34555 19395 34561
rect 1762 34484 1768 34536
rect 1820 34524 1826 34536
rect 2685 34527 2743 34533
rect 2685 34524 2697 34527
rect 1820 34496 2697 34524
rect 1820 34484 1826 34496
rect 2685 34493 2697 34496
rect 2731 34493 2743 34527
rect 14458 34524 14464 34536
rect 14419 34496 14464 34524
rect 2685 34487 2743 34493
rect 14458 34484 14464 34496
rect 14516 34484 14522 34536
rect 16574 34484 16580 34536
rect 16632 34524 16638 34536
rect 16761 34527 16819 34533
rect 16761 34524 16773 34527
rect 16632 34496 16773 34524
rect 16632 34484 16638 34496
rect 16761 34493 16773 34496
rect 16807 34524 16819 34527
rect 17788 34524 17816 34555
rect 16807 34496 17816 34524
rect 19168 34524 19196 34555
rect 19426 34552 19432 34604
rect 19484 34592 19490 34604
rect 19797 34595 19855 34601
rect 19797 34592 19809 34595
rect 19484 34564 19809 34592
rect 19484 34552 19490 34564
rect 19797 34561 19809 34564
rect 19843 34592 19855 34595
rect 20438 34592 20444 34604
rect 19843 34564 20444 34592
rect 19843 34561 19855 34564
rect 19797 34555 19855 34561
rect 20438 34552 20444 34564
rect 20496 34592 20502 34604
rect 22094 34601 22100 34604
rect 20901 34595 20959 34601
rect 20901 34592 20913 34595
rect 20496 34564 20913 34592
rect 20496 34552 20502 34564
rect 20901 34561 20913 34564
rect 20947 34561 20959 34595
rect 20901 34555 20959 34561
rect 22088 34555 22100 34601
rect 22152 34592 22158 34604
rect 22152 34564 22188 34592
rect 20165 34527 20223 34533
rect 20165 34524 20177 34527
rect 19168 34496 20177 34524
rect 16807 34493 16819 34496
rect 16761 34487 16819 34493
rect 20165 34493 20177 34496
rect 20211 34493 20223 34527
rect 20165 34487 20223 34493
rect 17681 34459 17739 34465
rect 17681 34425 17693 34459
rect 17727 34456 17739 34459
rect 17770 34456 17776 34468
rect 17727 34428 17776 34456
rect 17727 34425 17739 34428
rect 17681 34419 17739 34425
rect 17770 34416 17776 34428
rect 17828 34416 17834 34468
rect 20916 34456 20944 34555
rect 22094 34552 22100 34555
rect 22152 34552 22158 34564
rect 21818 34524 21824 34536
rect 21779 34496 21824 34524
rect 21818 34484 21824 34496
rect 21876 34484 21882 34536
rect 23216 34524 23244 34632
rect 24044 34632 26372 34660
rect 23934 34592 23940 34604
rect 23895 34564 23940 34592
rect 23934 34552 23940 34564
rect 23992 34552 23998 34604
rect 24044 34524 24072 34632
rect 24210 34601 24216 34604
rect 24204 34555 24216 34601
rect 24268 34592 24274 34604
rect 26234 34592 26240 34604
rect 24268 34564 24304 34592
rect 26195 34564 26240 34592
rect 24210 34552 24216 34555
rect 24268 34552 24274 34564
rect 26234 34552 26240 34564
rect 26292 34552 26298 34604
rect 26344 34592 26372 34632
rect 26421 34629 26433 34663
rect 26467 34660 26479 34663
rect 26510 34660 26516 34672
rect 26467 34632 26516 34660
rect 26467 34629 26479 34632
rect 26421 34623 26479 34629
rect 26510 34620 26516 34632
rect 26568 34620 26574 34672
rect 28721 34663 28779 34669
rect 26620 34632 28672 34660
rect 26620 34592 26648 34632
rect 28534 34592 28540 34604
rect 26344 34564 26648 34592
rect 28495 34564 28540 34592
rect 28534 34552 28540 34564
rect 28592 34552 28598 34604
rect 28644 34592 28672 34632
rect 28721 34629 28733 34663
rect 28767 34660 28779 34663
rect 30742 34660 30748 34672
rect 28767 34632 30748 34660
rect 28767 34629 28779 34632
rect 28721 34623 28779 34629
rect 30742 34620 30748 34632
rect 30800 34620 30806 34672
rect 33137 34663 33195 34669
rect 33137 34629 33149 34663
rect 33183 34660 33195 34663
rect 33226 34660 33232 34672
rect 33183 34632 33232 34660
rect 33183 34629 33195 34632
rect 33137 34623 33195 34629
rect 33226 34620 33232 34632
rect 33284 34620 33290 34672
rect 39850 34620 39856 34672
rect 39908 34660 39914 34672
rect 39908 34632 46612 34660
rect 39908 34620 39914 34632
rect 46584 34604 46612 34632
rect 28644 34564 29592 34592
rect 23216 34496 24072 34524
rect 26252 34524 26280 34552
rect 26973 34527 27031 34533
rect 26973 34524 26985 34527
rect 26252 34496 26985 34524
rect 23216 34465 23244 34496
rect 26973 34493 26985 34496
rect 27019 34493 27031 34527
rect 26973 34487 27031 34493
rect 27249 34527 27307 34533
rect 27249 34493 27261 34527
rect 27295 34524 27307 34527
rect 28166 34524 28172 34536
rect 27295 34496 28172 34524
rect 27295 34493 27307 34496
rect 27249 34487 27307 34493
rect 28166 34484 28172 34496
rect 28224 34484 28230 34536
rect 28902 34484 28908 34536
rect 28960 34524 28966 34536
rect 29181 34527 29239 34533
rect 29181 34524 29193 34527
rect 28960 34496 29193 34524
rect 28960 34484 28966 34496
rect 29181 34493 29193 34496
rect 29227 34493 29239 34527
rect 29181 34487 29239 34493
rect 29457 34527 29515 34533
rect 29457 34493 29469 34527
rect 29503 34493 29515 34527
rect 29564 34524 29592 34564
rect 29638 34552 29644 34604
rect 29696 34592 29702 34604
rect 30561 34595 30619 34601
rect 30561 34592 30573 34595
rect 29696 34564 30573 34592
rect 29696 34552 29702 34564
rect 30561 34561 30573 34564
rect 30607 34561 30619 34595
rect 46106 34592 46112 34604
rect 46067 34564 46112 34592
rect 30561 34555 30619 34561
rect 46106 34552 46112 34564
rect 46164 34552 46170 34604
rect 46566 34552 46572 34604
rect 46624 34592 46630 34604
rect 46753 34595 46811 34601
rect 46753 34592 46765 34595
rect 46624 34564 46765 34592
rect 46624 34552 46630 34564
rect 46753 34561 46765 34564
rect 46799 34561 46811 34595
rect 47578 34592 47584 34604
rect 47539 34564 47584 34592
rect 46753 34555 46811 34561
rect 47578 34552 47584 34564
rect 47636 34552 47642 34604
rect 32214 34524 32220 34536
rect 29564 34496 32220 34524
rect 29457 34487 29515 34493
rect 23201 34459 23259 34465
rect 20916 34428 21404 34456
rect 1394 34348 1400 34400
rect 1452 34388 1458 34400
rect 1581 34391 1639 34397
rect 1581 34388 1593 34391
rect 1452 34360 1593 34388
rect 1452 34348 1458 34360
rect 1581 34357 1593 34360
rect 1627 34357 1639 34391
rect 2130 34388 2136 34400
rect 2091 34360 2136 34388
rect 1581 34351 1639 34357
rect 2130 34348 2136 34360
rect 2188 34348 2194 34400
rect 17129 34391 17187 34397
rect 17129 34357 17141 34391
rect 17175 34388 17187 34391
rect 17494 34388 17500 34400
rect 17175 34360 17500 34388
rect 17175 34357 17187 34360
rect 17129 34351 17187 34357
rect 17494 34348 17500 34360
rect 17552 34348 17558 34400
rect 21266 34388 21272 34400
rect 21227 34360 21272 34388
rect 21266 34348 21272 34360
rect 21324 34348 21330 34400
rect 21376 34388 21404 34428
rect 23201 34425 23213 34459
rect 23247 34425 23259 34459
rect 29472 34456 29500 34487
rect 32214 34484 32220 34496
rect 32272 34484 32278 34536
rect 33229 34527 33287 34533
rect 33229 34493 33241 34527
rect 33275 34524 33287 34527
rect 33318 34524 33324 34536
rect 33275 34496 33324 34524
rect 33275 34493 33287 34496
rect 33229 34487 33287 34493
rect 33318 34484 33324 34496
rect 33376 34484 33382 34536
rect 33413 34527 33471 34533
rect 33413 34493 33425 34527
rect 33459 34524 33471 34527
rect 33502 34524 33508 34536
rect 33459 34496 33508 34524
rect 33459 34493 33471 34496
rect 33413 34487 33471 34493
rect 33502 34484 33508 34496
rect 33560 34484 33566 34536
rect 46842 34524 46848 34536
rect 46803 34496 46848 34524
rect 46842 34484 46848 34496
rect 46900 34484 46906 34536
rect 47670 34484 47676 34536
rect 47728 34524 47734 34536
rect 48038 34524 48044 34536
rect 47728 34496 48044 34524
rect 47728 34484 47734 34496
rect 48038 34484 48044 34496
rect 48096 34484 48102 34536
rect 30558 34456 30564 34468
rect 29472 34428 30564 34456
rect 23201 34419 23259 34425
rect 30558 34416 30564 34428
rect 30616 34416 30622 34468
rect 23106 34388 23112 34400
rect 21376 34360 23112 34388
rect 23106 34348 23112 34360
rect 23164 34348 23170 34400
rect 25317 34391 25375 34397
rect 25317 34357 25329 34391
rect 25363 34388 25375 34391
rect 25682 34388 25688 34400
rect 25363 34360 25688 34388
rect 25363 34357 25375 34360
rect 25317 34351 25375 34357
rect 25682 34348 25688 34360
rect 25740 34348 25746 34400
rect 30466 34348 30472 34400
rect 30524 34388 30530 34400
rect 30653 34391 30711 34397
rect 30653 34388 30665 34391
rect 30524 34360 30665 34388
rect 30524 34348 30530 34360
rect 30653 34357 30665 34360
rect 30699 34357 30711 34391
rect 30653 34351 30711 34357
rect 46201 34391 46259 34397
rect 46201 34357 46213 34391
rect 46247 34388 46259 34391
rect 46474 34388 46480 34400
rect 46247 34360 46480 34388
rect 46247 34357 46259 34360
rect 46201 34351 46259 34357
rect 46474 34348 46480 34360
rect 46532 34348 46538 34400
rect 1104 34298 48852 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 48852 34298
rect 1104 34224 48852 34246
rect 17678 34184 17684 34196
rect 12406 34156 16528 34184
rect 17639 34156 17684 34184
rect 1394 34048 1400 34060
rect 1355 34020 1400 34048
rect 1394 34008 1400 34020
rect 1452 34008 1458 34060
rect 1581 34051 1639 34057
rect 1581 34017 1593 34051
rect 1627 34048 1639 34051
rect 2130 34048 2136 34060
rect 1627 34020 2136 34048
rect 1627 34017 1639 34020
rect 1581 34011 1639 34017
rect 2130 34008 2136 34020
rect 2188 34008 2194 34060
rect 2774 34048 2780 34060
rect 2735 34020 2780 34048
rect 2774 34008 2780 34020
rect 2832 34008 2838 34060
rect 11701 34051 11759 34057
rect 11701 34017 11713 34051
rect 11747 34048 11759 34051
rect 12406 34048 12434 34156
rect 16500 34116 16528 34156
rect 17678 34144 17684 34156
rect 17736 34144 17742 34196
rect 21453 34187 21511 34193
rect 21453 34153 21465 34187
rect 21499 34184 21511 34187
rect 22094 34184 22100 34196
rect 21499 34156 22100 34184
rect 21499 34153 21511 34156
rect 21453 34147 21511 34153
rect 22094 34144 22100 34156
rect 22152 34144 22158 34196
rect 22186 34144 22192 34196
rect 22244 34184 22250 34196
rect 22741 34187 22799 34193
rect 22741 34184 22753 34187
rect 22244 34156 22753 34184
rect 22244 34144 22250 34156
rect 22741 34153 22753 34156
rect 22787 34184 22799 34187
rect 23014 34184 23020 34196
rect 22787 34156 23020 34184
rect 22787 34153 22799 34156
rect 22741 34147 22799 34153
rect 23014 34144 23020 34156
rect 23072 34144 23078 34196
rect 24210 34144 24216 34196
rect 24268 34184 24274 34196
rect 24397 34187 24455 34193
rect 24397 34184 24409 34187
rect 24268 34156 24409 34184
rect 24268 34144 24274 34156
rect 24397 34153 24409 34156
rect 24443 34153 24455 34187
rect 24397 34147 24455 34153
rect 30466 34144 30472 34196
rect 30524 34184 30530 34196
rect 30524 34156 32720 34184
rect 30524 34144 30530 34156
rect 18138 34116 18144 34128
rect 16500 34088 18144 34116
rect 18138 34076 18144 34088
rect 18196 34076 18202 34128
rect 19978 34116 19984 34128
rect 19939 34088 19984 34116
rect 19978 34076 19984 34088
rect 20036 34076 20042 34128
rect 21910 34076 21916 34128
rect 21968 34116 21974 34128
rect 21968 34088 23796 34116
rect 21968 34076 21974 34088
rect 11747 34020 12434 34048
rect 13081 34051 13139 34057
rect 11747 34017 11759 34020
rect 11701 34011 11759 34017
rect 13081 34017 13093 34051
rect 13127 34017 13139 34051
rect 13081 34011 13139 34017
rect 11882 33912 11888 33924
rect 11843 33884 11888 33912
rect 11882 33872 11888 33884
rect 11940 33872 11946 33924
rect 9858 33804 9864 33856
rect 9916 33844 9922 33856
rect 13096 33844 13124 34011
rect 15194 34008 15200 34060
rect 15252 34048 15258 34060
rect 15565 34051 15623 34057
rect 15565 34048 15577 34051
rect 15252 34020 15577 34048
rect 15252 34008 15258 34020
rect 15565 34017 15577 34020
rect 15611 34017 15623 34051
rect 15565 34011 15623 34017
rect 21266 34008 21272 34060
rect 21324 34048 21330 34060
rect 21324 34020 21956 34048
rect 21324 34008 21330 34020
rect 17405 33983 17463 33989
rect 17405 33980 17417 33983
rect 16960 33952 17417 33980
rect 15832 33915 15890 33921
rect 15832 33881 15844 33915
rect 15878 33912 15890 33915
rect 16666 33912 16672 33924
rect 15878 33884 16672 33912
rect 15878 33881 15890 33884
rect 15832 33875 15890 33881
rect 16666 33872 16672 33884
rect 16724 33872 16730 33924
rect 9916 33816 13124 33844
rect 9916 33804 9922 33816
rect 16574 33804 16580 33856
rect 16632 33844 16638 33856
rect 16960 33853 16988 33952
rect 17405 33949 17417 33952
rect 17451 33949 17463 33983
rect 17405 33943 17463 33949
rect 18601 33983 18659 33989
rect 18601 33949 18613 33983
rect 18647 33980 18659 33983
rect 21726 33980 21732 33992
rect 18647 33952 21588 33980
rect 21687 33952 21732 33980
rect 18647 33949 18659 33952
rect 18601 33943 18659 33949
rect 17494 33872 17500 33924
rect 17552 33912 17558 33924
rect 18417 33915 18475 33921
rect 18417 33912 18429 33915
rect 17552 33884 18429 33912
rect 17552 33872 17558 33884
rect 18417 33881 18429 33884
rect 18463 33881 18475 33915
rect 18417 33875 18475 33881
rect 19797 33915 19855 33921
rect 19797 33881 19809 33915
rect 19843 33912 19855 33915
rect 20898 33912 20904 33924
rect 19843 33884 20904 33912
rect 19843 33881 19855 33884
rect 19797 33875 19855 33881
rect 20898 33872 20904 33884
rect 20956 33872 20962 33924
rect 16945 33847 17003 33853
rect 16945 33844 16957 33847
rect 16632 33816 16957 33844
rect 16632 33804 16638 33816
rect 16945 33813 16957 33816
rect 16991 33813 17003 33847
rect 17862 33844 17868 33856
rect 17823 33816 17868 33844
rect 16945 33807 17003 33813
rect 17862 33804 17868 33816
rect 17920 33804 17926 33856
rect 21560 33844 21588 33952
rect 21726 33940 21732 33952
rect 21784 33940 21790 33992
rect 21928 33989 21956 34020
rect 21821 33983 21879 33989
rect 21821 33949 21833 33983
rect 21867 33949 21879 33983
rect 21821 33943 21879 33949
rect 21913 33983 21971 33989
rect 21913 33949 21925 33983
rect 21959 33949 21971 33983
rect 21913 33943 21971 33949
rect 21836 33912 21864 33943
rect 22020 33912 22048 34088
rect 22278 34048 22284 34060
rect 22112 34020 22284 34048
rect 22112 33989 22140 34020
rect 22278 34008 22284 34020
rect 22336 34008 22342 34060
rect 22097 33983 22155 33989
rect 22097 33949 22109 33983
rect 22143 33949 22155 33983
rect 22554 33980 22560 33992
rect 22515 33952 22560 33980
rect 22097 33943 22155 33949
rect 22554 33940 22560 33952
rect 22612 33940 22618 33992
rect 23106 33940 23112 33992
rect 23164 33980 23170 33992
rect 23477 33983 23535 33989
rect 23477 33980 23489 33983
rect 23164 33952 23489 33980
rect 23164 33940 23170 33952
rect 23477 33949 23489 33952
rect 23523 33949 23535 33983
rect 23477 33943 23535 33949
rect 21836 33884 22048 33912
rect 23661 33915 23719 33921
rect 23661 33881 23673 33915
rect 23707 33881 23719 33915
rect 23768 33912 23796 34088
rect 24762 34076 24768 34128
rect 24820 34116 24826 34128
rect 24820 34088 25176 34116
rect 24820 34076 24826 34088
rect 23845 34051 23903 34057
rect 23845 34017 23857 34051
rect 23891 34048 23903 34051
rect 23891 34020 24900 34048
rect 23891 34017 23903 34020
rect 23845 34011 23903 34017
rect 23934 33940 23940 33992
rect 23992 33980 23998 33992
rect 24872 33989 24900 34020
rect 24673 33983 24731 33989
rect 24673 33980 24685 33983
rect 23992 33952 24685 33980
rect 23992 33940 23998 33952
rect 24673 33949 24685 33952
rect 24719 33949 24731 33983
rect 24673 33943 24731 33949
rect 24765 33983 24823 33989
rect 24765 33949 24777 33983
rect 24811 33949 24823 33983
rect 24765 33943 24823 33949
rect 24857 33983 24915 33989
rect 24857 33949 24869 33983
rect 24903 33949 24915 33983
rect 25038 33980 25044 33992
rect 24999 33952 25044 33980
rect 24857 33943 24915 33949
rect 24780 33912 24808 33943
rect 25038 33940 25044 33952
rect 25096 33940 25102 33992
rect 25148 33980 25176 34088
rect 25682 34076 25688 34128
rect 25740 34116 25746 34128
rect 25740 34088 31432 34116
rect 25740 34076 25746 34088
rect 26878 34008 26884 34060
rect 26936 34048 26942 34060
rect 28353 34051 28411 34057
rect 28353 34048 28365 34051
rect 26936 34020 27289 34048
rect 26936 34008 26942 34020
rect 27261 33989 27289 34020
rect 27356 34020 28365 34048
rect 27356 33989 27384 34020
rect 28353 34017 28365 34020
rect 28399 34017 28411 34051
rect 28353 34011 28411 34017
rect 27157 33983 27215 33989
rect 27157 33980 27169 33983
rect 25148 33952 27169 33980
rect 27157 33949 27169 33952
rect 27203 33949 27215 33983
rect 27157 33943 27215 33949
rect 27246 33983 27304 33989
rect 27246 33949 27258 33983
rect 27292 33949 27304 33983
rect 27246 33943 27304 33949
rect 27341 33983 27399 33989
rect 27341 33949 27353 33983
rect 27387 33949 27399 33983
rect 27341 33943 27399 33949
rect 27525 33983 27583 33989
rect 27525 33949 27537 33983
rect 27571 33980 27583 33983
rect 27706 33980 27712 33992
rect 27571 33952 27712 33980
rect 27571 33949 27583 33952
rect 27525 33943 27583 33949
rect 27706 33940 27712 33952
rect 27764 33940 27770 33992
rect 28166 33980 28172 33992
rect 28079 33952 28172 33980
rect 28166 33940 28172 33952
rect 28224 33980 28230 33992
rect 31404 33989 31432 34088
rect 31478 34076 31484 34128
rect 31536 34076 31542 34128
rect 32692 34116 32720 34156
rect 47026 34116 47032 34128
rect 32692 34088 32812 34116
rect 31496 33989 31524 34076
rect 31662 34008 31668 34060
rect 31720 34048 31726 34060
rect 32784 34057 32812 34088
rect 46308 34088 47032 34116
rect 32677 34051 32735 34057
rect 32677 34048 32689 34051
rect 31720 34020 32689 34048
rect 31720 34008 31726 34020
rect 32677 34017 32689 34020
rect 32723 34017 32735 34051
rect 32677 34011 32735 34017
rect 32769 34051 32827 34057
rect 32769 34017 32781 34051
rect 32815 34048 32827 34051
rect 33502 34048 33508 34060
rect 32815 34020 33508 34048
rect 32815 34017 32827 34020
rect 32769 34011 32827 34017
rect 33502 34008 33508 34020
rect 33560 34048 33566 34060
rect 46308 34057 46336 34088
rect 47026 34076 47032 34088
rect 47084 34076 47090 34128
rect 33965 34051 34023 34057
rect 33965 34048 33977 34051
rect 33560 34020 33977 34048
rect 33560 34008 33566 34020
rect 33965 34017 33977 34020
rect 34011 34017 34023 34051
rect 33965 34011 34023 34017
rect 46293 34051 46351 34057
rect 46293 34017 46305 34051
rect 46339 34017 46351 34051
rect 46474 34048 46480 34060
rect 46435 34020 46480 34048
rect 46293 34011 46351 34017
rect 46474 34008 46480 34020
rect 46532 34008 46538 34060
rect 48130 34048 48136 34060
rect 48091 34020 48136 34048
rect 48130 34008 48136 34020
rect 48188 34008 48194 34060
rect 31389 33983 31447 33989
rect 28224 33952 29868 33980
rect 28224 33940 28230 33952
rect 23768 33884 24808 33912
rect 23661 33875 23719 33881
rect 22646 33844 22652 33856
rect 21560 33816 22652 33844
rect 22646 33804 22652 33816
rect 22704 33804 22710 33856
rect 23676 33844 23704 33875
rect 27430 33872 27436 33924
rect 27488 33912 27494 33924
rect 27985 33915 28043 33921
rect 27985 33912 27997 33915
rect 27488 33884 27997 33912
rect 27488 33872 27494 33884
rect 27985 33881 27997 33884
rect 28031 33881 28043 33915
rect 29638 33912 29644 33924
rect 29599 33884 29644 33912
rect 27985 33875 28043 33881
rect 29638 33872 29644 33884
rect 29696 33872 29702 33924
rect 29840 33921 29868 33952
rect 31389 33949 31401 33983
rect 31435 33949 31447 33983
rect 31389 33943 31447 33949
rect 31481 33983 31539 33989
rect 31481 33949 31493 33983
rect 31527 33949 31539 33983
rect 31481 33943 31539 33949
rect 31570 33940 31576 33992
rect 31628 33980 31634 33992
rect 31757 33983 31815 33989
rect 31628 33952 31673 33980
rect 31628 33940 31634 33952
rect 31757 33949 31769 33983
rect 31803 33980 31815 33983
rect 32490 33980 32496 33992
rect 31803 33952 32496 33980
rect 31803 33949 31815 33952
rect 31757 33943 31815 33949
rect 32490 33940 32496 33952
rect 32548 33940 32554 33992
rect 32585 33983 32643 33989
rect 32585 33949 32597 33983
rect 32631 33980 32643 33983
rect 34422 33980 34428 33992
rect 32631 33952 34428 33980
rect 32631 33949 32643 33952
rect 32585 33943 32643 33949
rect 34422 33940 34428 33952
rect 34480 33940 34486 33992
rect 29825 33915 29883 33921
rect 29825 33881 29837 33915
rect 29871 33912 29883 33915
rect 31113 33915 31171 33921
rect 29871 33884 30144 33912
rect 29871 33881 29883 33884
rect 29825 33875 29883 33881
rect 25682 33844 25688 33856
rect 23676 33816 25688 33844
rect 25682 33804 25688 33816
rect 25740 33804 25746 33856
rect 26881 33847 26939 33853
rect 26881 33813 26893 33847
rect 26927 33844 26939 33847
rect 27154 33844 27160 33856
rect 26927 33816 27160 33844
rect 26927 33813 26939 33816
rect 26881 33807 26939 33813
rect 27154 33804 27160 33816
rect 27212 33804 27218 33856
rect 29914 33804 29920 33856
rect 29972 33844 29978 33856
rect 30009 33847 30067 33853
rect 30009 33844 30021 33847
rect 29972 33816 30021 33844
rect 29972 33804 29978 33816
rect 30009 33813 30021 33816
rect 30055 33813 30067 33847
rect 30116 33844 30144 33884
rect 31113 33881 31125 33915
rect 31159 33912 31171 33915
rect 33318 33912 33324 33924
rect 31159 33884 33324 33912
rect 31159 33881 31171 33884
rect 31113 33875 31171 33881
rect 33318 33872 33324 33884
rect 33376 33872 33382 33924
rect 33870 33912 33876 33924
rect 33831 33884 33876 33912
rect 33870 33872 33876 33884
rect 33928 33872 33934 33924
rect 32030 33844 32036 33856
rect 30116 33816 32036 33844
rect 30009 33807 30067 33813
rect 32030 33804 32036 33816
rect 32088 33804 32094 33856
rect 32122 33804 32128 33856
rect 32180 33844 32186 33856
rect 32217 33847 32275 33853
rect 32217 33844 32229 33847
rect 32180 33816 32229 33844
rect 32180 33804 32186 33816
rect 32217 33813 32229 33816
rect 32263 33813 32275 33847
rect 32217 33807 32275 33813
rect 33134 33804 33140 33856
rect 33192 33844 33198 33856
rect 33413 33847 33471 33853
rect 33413 33844 33425 33847
rect 33192 33816 33425 33844
rect 33192 33804 33198 33816
rect 33413 33813 33425 33816
rect 33459 33813 33471 33847
rect 33778 33844 33784 33856
rect 33739 33816 33784 33844
rect 33413 33807 33471 33813
rect 33778 33804 33784 33816
rect 33836 33804 33842 33856
rect 1104 33754 48852 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 48852 33754
rect 1104 33680 48852 33702
rect 11882 33640 11888 33652
rect 11843 33612 11888 33640
rect 11882 33600 11888 33612
rect 11940 33600 11946 33652
rect 14458 33600 14464 33652
rect 14516 33640 14522 33652
rect 14737 33643 14795 33649
rect 14737 33640 14749 33643
rect 14516 33612 14749 33640
rect 14516 33600 14522 33612
rect 14737 33609 14749 33612
rect 14783 33609 14795 33643
rect 14737 33603 14795 33609
rect 15289 33643 15347 33649
rect 15289 33609 15301 33643
rect 15335 33609 15347 33643
rect 15289 33603 15347 33609
rect 15473 33643 15531 33649
rect 15473 33609 15485 33643
rect 15519 33640 15531 33643
rect 16758 33640 16764 33652
rect 15519 33612 16764 33640
rect 15519 33609 15531 33612
rect 15473 33603 15531 33609
rect 15304 33572 15332 33603
rect 16758 33600 16764 33612
rect 16816 33600 16822 33652
rect 23106 33600 23112 33652
rect 23164 33640 23170 33652
rect 27430 33640 27436 33652
rect 23164 33612 24072 33640
rect 27391 33612 27436 33640
rect 23164 33600 23170 33612
rect 14660 33544 15332 33572
rect 1762 33504 1768 33516
rect 1723 33476 1768 33504
rect 1762 33464 1768 33476
rect 1820 33464 1826 33516
rect 11698 33464 11704 33516
rect 11756 33504 11762 33516
rect 14660 33513 14688 33544
rect 16022 33532 16028 33584
rect 16080 33572 16086 33584
rect 16853 33575 16911 33581
rect 16853 33572 16865 33575
rect 16080 33544 16865 33572
rect 16080 33532 16086 33544
rect 16853 33541 16865 33544
rect 16899 33541 16911 33575
rect 16853 33535 16911 33541
rect 22278 33532 22284 33584
rect 22336 33572 22342 33584
rect 24044 33581 24072 33612
rect 27430 33600 27436 33612
rect 27488 33600 27494 33652
rect 27893 33643 27951 33649
rect 27893 33609 27905 33643
rect 27939 33640 27951 33643
rect 28350 33640 28356 33652
rect 27939 33612 28356 33640
rect 27939 33609 27951 33612
rect 27893 33603 27951 33609
rect 28350 33600 28356 33612
rect 28408 33600 28414 33652
rect 29638 33600 29644 33652
rect 29696 33640 29702 33652
rect 29917 33643 29975 33649
rect 29917 33640 29929 33643
rect 29696 33612 29929 33640
rect 29696 33600 29702 33612
rect 29917 33609 29929 33612
rect 29963 33609 29975 33643
rect 30374 33640 30380 33652
rect 30335 33612 30380 33640
rect 29917 33603 29975 33609
rect 30374 33600 30380 33612
rect 30432 33600 30438 33652
rect 31570 33600 31576 33652
rect 31628 33640 31634 33652
rect 32493 33643 32551 33649
rect 32493 33640 32505 33643
rect 31628 33612 32505 33640
rect 31628 33600 31634 33612
rect 32493 33609 32505 33612
rect 32539 33609 32551 33643
rect 32493 33603 32551 33609
rect 33778 33600 33784 33652
rect 33836 33640 33842 33652
rect 36265 33643 36323 33649
rect 36265 33640 36277 33643
rect 33836 33612 36277 33640
rect 33836 33600 33842 33612
rect 36265 33609 36277 33612
rect 36311 33609 36323 33643
rect 36265 33603 36323 33609
rect 23293 33575 23351 33581
rect 23293 33572 23305 33575
rect 22336 33544 23305 33572
rect 22336 33532 22342 33544
rect 23293 33541 23305 33544
rect 23339 33541 23351 33575
rect 23293 33535 23351 33541
rect 24029 33575 24087 33581
rect 24029 33541 24041 33575
rect 24075 33541 24087 33575
rect 24486 33572 24492 33584
rect 24029 33535 24087 33541
rect 24136 33544 24492 33572
rect 11793 33507 11851 33513
rect 11793 33504 11805 33507
rect 11756 33476 11805 33504
rect 11756 33464 11762 33476
rect 11793 33473 11805 33476
rect 11839 33473 11851 33507
rect 11793 33467 11851 33473
rect 14645 33507 14703 33513
rect 14645 33473 14657 33507
rect 14691 33473 14703 33507
rect 14645 33467 14703 33473
rect 14829 33507 14887 33513
rect 14829 33473 14841 33507
rect 14875 33473 14887 33507
rect 14829 33467 14887 33473
rect 15470 33507 15528 33513
rect 15470 33473 15482 33507
rect 15516 33504 15528 33507
rect 15746 33504 15752 33516
rect 15516 33476 15752 33504
rect 15516 33473 15528 33476
rect 15470 33467 15528 33473
rect 1946 33436 1952 33448
rect 1907 33408 1952 33436
rect 1946 33396 1952 33408
rect 2004 33396 2010 33448
rect 2774 33436 2780 33448
rect 2735 33408 2780 33436
rect 2774 33396 2780 33408
rect 2832 33396 2838 33448
rect 14844 33368 14872 33467
rect 15746 33464 15752 33476
rect 15804 33464 15810 33516
rect 15841 33507 15899 33513
rect 15841 33473 15853 33507
rect 15887 33504 15899 33507
rect 16574 33504 16580 33516
rect 15887 33476 16580 33504
rect 15887 33473 15899 33476
rect 15841 33467 15899 33473
rect 16574 33464 16580 33476
rect 16632 33464 16638 33516
rect 16669 33507 16727 33513
rect 16669 33473 16681 33507
rect 16715 33473 16727 33507
rect 16669 33467 16727 33473
rect 16945 33507 17003 33513
rect 16945 33473 16957 33507
rect 16991 33504 17003 33507
rect 17862 33504 17868 33516
rect 16991 33476 17868 33504
rect 16991 33473 17003 33476
rect 16945 33467 17003 33473
rect 15930 33436 15936 33448
rect 15891 33408 15936 33436
rect 15930 33396 15936 33408
rect 15988 33396 15994 33448
rect 16684 33436 16712 33467
rect 17862 33464 17868 33476
rect 17920 33464 17926 33516
rect 19337 33507 19395 33513
rect 19337 33473 19349 33507
rect 19383 33504 19395 33507
rect 19426 33504 19432 33516
rect 19383 33476 19432 33504
rect 19383 33473 19395 33476
rect 19337 33467 19395 33473
rect 19426 33464 19432 33476
rect 19484 33464 19490 33516
rect 23106 33464 23112 33516
rect 23164 33504 23170 33516
rect 23308 33504 23336 33535
rect 24136 33504 24164 33544
rect 24486 33532 24492 33544
rect 24544 33572 24550 33584
rect 25038 33572 25044 33584
rect 24544 33544 25044 33572
rect 24544 33532 24550 33544
rect 25038 33532 25044 33544
rect 25096 33532 25102 33584
rect 26237 33575 26295 33581
rect 26237 33541 26249 33575
rect 26283 33572 26295 33575
rect 26418 33572 26424 33584
rect 26283 33544 26424 33572
rect 26283 33541 26295 33544
rect 26237 33535 26295 33541
rect 26418 33532 26424 33544
rect 26476 33532 26482 33584
rect 27706 33532 27712 33584
rect 27764 33572 27770 33584
rect 28905 33575 28963 33581
rect 28905 33572 28917 33575
rect 27764 33544 28917 33572
rect 27764 33532 27770 33544
rect 28905 33541 28917 33544
rect 28951 33541 28963 33575
rect 32122 33572 32128 33584
rect 32083 33544 32128 33572
rect 28905 33535 28963 33541
rect 32122 33532 32128 33544
rect 32180 33532 32186 33584
rect 33060 33544 34928 33572
rect 33060 33516 33088 33544
rect 23164 33476 23244 33504
rect 23308 33476 24164 33504
rect 24213 33507 24271 33513
rect 23164 33464 23170 33476
rect 17494 33436 17500 33448
rect 16040 33408 16712 33436
rect 17455 33408 17500 33436
rect 15286 33368 15292 33380
rect 14844 33340 15292 33368
rect 15286 33328 15292 33340
rect 15344 33368 15350 33380
rect 16040 33368 16068 33408
rect 17494 33396 17500 33408
rect 17552 33396 17558 33448
rect 17773 33439 17831 33445
rect 17773 33405 17785 33439
rect 17819 33436 17831 33439
rect 18046 33436 18052 33448
rect 17819 33408 18052 33436
rect 17819 33405 17831 33408
rect 17773 33399 17831 33405
rect 18046 33396 18052 33408
rect 18104 33436 18110 33448
rect 19061 33439 19119 33445
rect 19061 33436 19073 33439
rect 18104 33408 19073 33436
rect 18104 33396 18110 33408
rect 19061 33405 19073 33408
rect 19107 33405 19119 33439
rect 23216 33436 23244 33476
rect 24213 33473 24225 33507
rect 24259 33504 24271 33507
rect 25774 33504 25780 33516
rect 24259 33476 25780 33504
rect 24259 33473 24271 33476
rect 24213 33467 24271 33473
rect 25774 33464 25780 33476
rect 25832 33464 25838 33516
rect 27801 33507 27859 33513
rect 27801 33473 27813 33507
rect 27847 33504 27859 33507
rect 27982 33504 27988 33516
rect 27847 33476 27988 33504
rect 27847 33473 27859 33476
rect 27801 33467 27859 33473
rect 27982 33464 27988 33476
rect 28040 33464 28046 33516
rect 28166 33464 28172 33516
rect 28224 33504 28230 33516
rect 28721 33507 28779 33513
rect 28721 33504 28733 33507
rect 28224 33476 28733 33504
rect 28224 33464 28230 33476
rect 28721 33473 28733 33476
rect 28767 33504 28779 33507
rect 28810 33504 28816 33516
rect 28767 33476 28816 33504
rect 28767 33473 28779 33476
rect 28721 33467 28779 33473
rect 28810 33464 28816 33476
rect 28868 33464 28874 33516
rect 30285 33507 30343 33513
rect 30285 33473 30297 33507
rect 30331 33504 30343 33507
rect 31386 33504 31392 33516
rect 30331 33476 31392 33504
rect 30331 33473 30343 33476
rect 30285 33467 30343 33473
rect 31386 33464 31392 33476
rect 31444 33464 31450 33516
rect 32030 33464 32036 33516
rect 32088 33504 32094 33516
rect 32309 33507 32367 33513
rect 32309 33504 32321 33507
rect 32088 33476 32321 33504
rect 32088 33464 32094 33476
rect 32309 33473 32321 33476
rect 32355 33504 32367 33507
rect 32490 33504 32496 33516
rect 32355 33476 32496 33504
rect 32355 33473 32367 33476
rect 32309 33467 32367 33473
rect 32490 33464 32496 33476
rect 32548 33464 32554 33516
rect 33042 33504 33048 33516
rect 32955 33476 33048 33504
rect 33042 33464 33048 33476
rect 33100 33464 33106 33516
rect 33318 33513 33324 33516
rect 33312 33467 33324 33513
rect 33376 33504 33382 33516
rect 34900 33513 34928 33544
rect 34885 33507 34943 33513
rect 33376 33476 33412 33504
rect 33318 33464 33324 33467
rect 33376 33464 33382 33476
rect 34885 33473 34897 33507
rect 34931 33473 34943 33507
rect 35141 33507 35199 33513
rect 35141 33504 35153 33507
rect 34885 33467 34943 33473
rect 34992 33476 35153 33504
rect 23382 33436 23388 33448
rect 23216 33408 23388 33436
rect 19061 33399 19119 33405
rect 23382 33396 23388 33408
rect 23440 33396 23446 33448
rect 28074 33436 28080 33448
rect 28035 33408 28080 33436
rect 28074 33396 28080 33408
rect 28132 33396 28138 33448
rect 30466 33436 30472 33448
rect 30427 33408 30472 33436
rect 30466 33396 30472 33408
rect 30524 33396 30530 33448
rect 34238 33396 34244 33448
rect 34296 33436 34302 33448
rect 34992 33436 35020 33476
rect 35141 33473 35153 33476
rect 35187 33473 35199 33507
rect 46477 33507 46535 33513
rect 46477 33504 46489 33507
rect 35141 33467 35199 33473
rect 45526 33476 46489 33504
rect 34296 33408 35020 33436
rect 34296 33396 34302 33408
rect 42794 33396 42800 33448
rect 42852 33436 42858 33448
rect 45526 33436 45554 33476
rect 46477 33473 46489 33476
rect 46523 33473 46535 33507
rect 46477 33467 46535 33473
rect 46198 33436 46204 33448
rect 42852 33408 45554 33436
rect 46159 33408 46204 33436
rect 42852 33396 42858 33408
rect 46198 33396 46204 33408
rect 46256 33396 46262 33448
rect 16666 33368 16672 33380
rect 15344 33340 16068 33368
rect 16627 33340 16672 33368
rect 15344 33328 15350 33340
rect 16666 33328 16672 33340
rect 16724 33328 16730 33380
rect 26421 33371 26479 33377
rect 26421 33337 26433 33371
rect 26467 33368 26479 33371
rect 26878 33368 26884 33380
rect 26467 33340 26884 33368
rect 26467 33337 26479 33340
rect 26421 33331 26479 33337
rect 26878 33328 26884 33340
rect 26936 33328 26942 33380
rect 34422 33368 34428 33380
rect 34383 33340 34428 33368
rect 34422 33328 34428 33340
rect 34480 33328 34486 33380
rect 2590 33260 2596 33312
rect 2648 33300 2654 33312
rect 2774 33300 2780 33312
rect 2648 33272 2780 33300
rect 2648 33260 2654 33272
rect 2774 33260 2780 33272
rect 2832 33260 2838 33312
rect 11698 33260 11704 33312
rect 11756 33300 11762 33312
rect 20530 33300 20536 33312
rect 11756 33272 20536 33300
rect 11756 33260 11762 33272
rect 20530 33260 20536 33272
rect 20588 33260 20594 33312
rect 24302 33260 24308 33312
rect 24360 33300 24366 33312
rect 24397 33303 24455 33309
rect 24397 33300 24409 33303
rect 24360 33272 24409 33300
rect 24360 33260 24366 33272
rect 24397 33269 24409 33272
rect 24443 33269 24455 33303
rect 47762 33300 47768 33312
rect 47723 33272 47768 33300
rect 24397 33263 24455 33269
rect 47762 33260 47768 33272
rect 47820 33260 47826 33312
rect 1104 33210 48852 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 48852 33210
rect 1104 33136 48852 33158
rect 1946 33056 1952 33108
rect 2004 33096 2010 33108
rect 2225 33099 2283 33105
rect 2225 33096 2237 33099
rect 2004 33068 2237 33096
rect 2004 33056 2010 33068
rect 2225 33065 2237 33068
rect 2271 33065 2283 33099
rect 2225 33059 2283 33065
rect 2590 33056 2596 33108
rect 2648 33096 2654 33108
rect 23750 33096 23756 33108
rect 2648 33068 22094 33096
rect 23663 33068 23756 33096
rect 2648 33056 2654 33068
rect 15933 33031 15991 33037
rect 15933 32997 15945 33031
rect 15979 33028 15991 33031
rect 16022 33028 16028 33040
rect 15979 33000 16028 33028
rect 15979 32997 15991 33000
rect 15933 32991 15991 32997
rect 16022 32988 16028 33000
rect 16080 32988 16086 33040
rect 18049 33031 18107 33037
rect 18049 32997 18061 33031
rect 18095 33028 18107 33031
rect 22066 33028 22094 33068
rect 23750 33056 23756 33068
rect 23808 33096 23814 33108
rect 28534 33096 28540 33108
rect 23808 33068 28540 33096
rect 23808 33056 23814 33068
rect 28534 33056 28540 33068
rect 28592 33056 28598 33108
rect 30374 33096 30380 33108
rect 28644 33068 30380 33096
rect 24118 33028 24124 33040
rect 18095 33000 19196 33028
rect 22066 33000 24124 33028
rect 18095 32997 18107 33000
rect 18049 32991 18107 32997
rect 9030 32960 9036 32972
rect 2148 32932 9036 32960
rect 2148 32901 2176 32932
rect 9030 32920 9036 32932
rect 9088 32920 9094 32972
rect 2133 32895 2191 32901
rect 2133 32861 2145 32895
rect 2179 32861 2191 32895
rect 2133 32855 2191 32861
rect 2961 32895 3019 32901
rect 2961 32861 2973 32895
rect 3007 32861 3019 32895
rect 2961 32855 3019 32861
rect 15749 32895 15807 32901
rect 15749 32861 15761 32895
rect 15795 32892 15807 32895
rect 15930 32892 15936 32904
rect 15795 32864 15936 32892
rect 15795 32861 15807 32864
rect 15749 32855 15807 32861
rect 2038 32784 2044 32836
rect 2096 32824 2102 32836
rect 2976 32824 3004 32855
rect 15930 32852 15936 32864
rect 15988 32852 15994 32904
rect 18322 32892 18328 32904
rect 18283 32864 18328 32892
rect 18322 32852 18328 32864
rect 18380 32852 18386 32904
rect 18414 32889 18472 32895
rect 18414 32855 18426 32889
rect 18460 32855 18472 32889
rect 18414 32849 18472 32855
rect 18506 32852 18512 32904
rect 18564 32901 18570 32904
rect 18564 32892 18572 32901
rect 18693 32895 18751 32901
rect 18564 32864 18609 32892
rect 18564 32855 18572 32864
rect 18693 32861 18705 32895
rect 18739 32892 18751 32895
rect 19058 32892 19064 32904
rect 18739 32864 19064 32892
rect 18739 32861 18751 32864
rect 18693 32855 18751 32861
rect 18564 32852 18570 32855
rect 19058 32852 19064 32864
rect 19116 32852 19122 32904
rect 2096 32796 3004 32824
rect 2096 32784 2102 32796
rect 18429 32756 18457 32849
rect 19168 32824 19196 33000
rect 24118 32988 24124 33000
rect 24176 32988 24182 33040
rect 19242 32920 19248 32972
rect 19300 32960 19306 32972
rect 19300 32932 19345 32960
rect 19300 32920 19306 32932
rect 24397 32895 24455 32901
rect 24397 32861 24409 32895
rect 24443 32892 24455 32895
rect 27062 32892 27068 32904
rect 24443 32864 27068 32892
rect 24443 32861 24455 32864
rect 24397 32855 24455 32861
rect 27062 32852 27068 32864
rect 27120 32852 27126 32904
rect 27154 32852 27160 32904
rect 27212 32892 27218 32904
rect 27321 32895 27379 32901
rect 27321 32892 27333 32895
rect 27212 32864 27333 32892
rect 27212 32852 27218 32864
rect 27321 32861 27333 32864
rect 27367 32861 27379 32895
rect 27321 32855 27379 32861
rect 27614 32852 27620 32904
rect 27672 32892 27678 32904
rect 28644 32892 28672 33068
rect 30374 33056 30380 33068
rect 30432 33056 30438 33108
rect 31386 33096 31392 33108
rect 31347 33068 31392 33096
rect 31386 33056 31392 33068
rect 31444 33056 31450 33108
rect 31941 33099 31999 33105
rect 31941 33065 31953 33099
rect 31987 33096 31999 33099
rect 34238 33096 34244 33108
rect 31987 33068 34244 33096
rect 31987 33065 31999 33068
rect 31941 33059 31999 33065
rect 34238 33056 34244 33068
rect 34296 33056 34302 33108
rect 31478 32920 31484 32972
rect 31536 32960 31542 32972
rect 33413 32963 33471 32969
rect 33413 32960 33425 32963
rect 31536 32932 32352 32960
rect 31536 32920 31542 32932
rect 27672 32864 28672 32892
rect 30009 32895 30067 32901
rect 27672 32852 27678 32864
rect 30009 32861 30021 32895
rect 30055 32892 30067 32895
rect 31754 32892 31760 32904
rect 30055 32864 31760 32892
rect 30055 32861 30067 32864
rect 30009 32855 30067 32861
rect 31754 32852 31760 32864
rect 31812 32852 31818 32904
rect 32214 32892 32220 32904
rect 32175 32864 32220 32892
rect 32214 32852 32220 32864
rect 32272 32852 32278 32904
rect 32324 32901 32352 32932
rect 32416 32932 33425 32960
rect 32416 32901 32444 32932
rect 33413 32929 33425 32932
rect 33459 32929 33471 32963
rect 33413 32923 33471 32929
rect 46293 32963 46351 32969
rect 46293 32929 46305 32963
rect 46339 32960 46351 32963
rect 47762 32960 47768 32972
rect 46339 32932 47768 32960
rect 46339 32929 46351 32932
rect 46293 32923 46351 32929
rect 47762 32920 47768 32932
rect 47820 32920 47826 32972
rect 48038 32960 48044 32972
rect 47999 32932 48044 32960
rect 48038 32920 48044 32932
rect 48096 32920 48102 32972
rect 32309 32895 32367 32901
rect 32309 32861 32321 32895
rect 32355 32861 32367 32895
rect 32309 32855 32367 32861
rect 32401 32895 32459 32901
rect 32401 32861 32413 32895
rect 32447 32861 32459 32895
rect 32582 32892 32588 32904
rect 32543 32864 32588 32892
rect 32401 32855 32459 32861
rect 32582 32852 32588 32864
rect 32640 32852 32646 32904
rect 33045 32895 33103 32901
rect 33045 32861 33057 32895
rect 33091 32892 33103 32895
rect 33134 32892 33140 32904
rect 33091 32864 33140 32892
rect 33091 32861 33103 32864
rect 33045 32855 33103 32861
rect 33134 32852 33140 32864
rect 33192 32852 33198 32904
rect 19490 32827 19548 32833
rect 19490 32824 19502 32827
rect 19168 32796 19502 32824
rect 19490 32793 19502 32796
rect 19536 32793 19548 32827
rect 19490 32787 19548 32793
rect 23382 32784 23388 32836
rect 23440 32824 23446 32836
rect 23661 32827 23719 32833
rect 23661 32824 23673 32827
rect 23440 32796 23673 32824
rect 23440 32784 23446 32796
rect 23661 32793 23673 32796
rect 23707 32793 23719 32827
rect 23661 32787 23719 32793
rect 23842 32784 23848 32836
rect 23900 32824 23906 32836
rect 24642 32827 24700 32833
rect 24642 32824 24654 32827
rect 23900 32796 24654 32824
rect 23900 32784 23906 32796
rect 24642 32793 24654 32796
rect 24688 32793 24700 32827
rect 24642 32787 24700 32793
rect 29362 32784 29368 32836
rect 29420 32824 29426 32836
rect 30254 32827 30312 32833
rect 30254 32824 30266 32827
rect 29420 32796 30266 32824
rect 29420 32784 29426 32796
rect 30254 32793 30266 32796
rect 30300 32793 30312 32827
rect 30254 32787 30312 32793
rect 32490 32784 32496 32836
rect 32548 32824 32554 32836
rect 33229 32827 33287 32833
rect 33229 32824 33241 32827
rect 32548 32796 33241 32824
rect 32548 32784 32554 32796
rect 33229 32793 33241 32796
rect 33275 32793 33287 32827
rect 33229 32787 33287 32793
rect 46477 32827 46535 32833
rect 46477 32793 46489 32827
rect 46523 32824 46535 32827
rect 46842 32824 46848 32836
rect 46523 32796 46848 32824
rect 46523 32793 46535 32796
rect 46477 32787 46535 32793
rect 46842 32784 46848 32796
rect 46900 32784 46906 32836
rect 19150 32756 19156 32768
rect 18429 32728 19156 32756
rect 19150 32716 19156 32728
rect 19208 32716 19214 32768
rect 20622 32756 20628 32768
rect 20535 32728 20628 32756
rect 20622 32716 20628 32728
rect 20680 32756 20686 32768
rect 24762 32756 24768 32768
rect 20680 32728 24768 32756
rect 20680 32716 20686 32728
rect 24762 32716 24768 32728
rect 24820 32716 24826 32768
rect 25774 32756 25780 32768
rect 25735 32728 25780 32756
rect 25774 32716 25780 32728
rect 25832 32716 25838 32768
rect 27982 32716 27988 32768
rect 28040 32756 28046 32768
rect 28445 32759 28503 32765
rect 28445 32756 28457 32759
rect 28040 32728 28457 32756
rect 28040 32716 28046 32728
rect 28445 32725 28457 32728
rect 28491 32756 28503 32759
rect 28810 32756 28816 32768
rect 28491 32728 28816 32756
rect 28491 32725 28503 32728
rect 28445 32719 28503 32725
rect 28810 32716 28816 32728
rect 28868 32716 28874 32768
rect 1104 32666 48852 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 48852 32666
rect 1104 32592 48852 32614
rect 15657 32555 15715 32561
rect 6886 32524 15608 32552
rect 2682 32444 2688 32496
rect 2740 32484 2746 32496
rect 6886 32484 6914 32524
rect 15194 32484 15200 32496
rect 2740 32456 6914 32484
rect 13372 32456 15200 32484
rect 2740 32444 2746 32456
rect 2038 32416 2044 32428
rect 1999 32388 2044 32416
rect 2038 32376 2044 32388
rect 2096 32376 2102 32428
rect 13372 32425 13400 32456
rect 15194 32444 15200 32456
rect 15252 32444 15258 32496
rect 15580 32484 15608 32524
rect 15657 32521 15669 32555
rect 15703 32552 15715 32555
rect 15930 32552 15936 32564
rect 15703 32524 15936 32552
rect 15703 32521 15715 32524
rect 15657 32515 15715 32521
rect 15930 32512 15936 32524
rect 15988 32512 15994 32564
rect 16758 32552 16764 32564
rect 16719 32524 16764 32552
rect 16758 32512 16764 32524
rect 16816 32512 16822 32564
rect 18506 32512 18512 32564
rect 18564 32552 18570 32564
rect 20257 32555 20315 32561
rect 20257 32552 20269 32555
rect 18564 32524 20269 32552
rect 18564 32512 18570 32524
rect 20257 32521 20269 32524
rect 20303 32521 20315 32555
rect 22646 32552 22652 32564
rect 20257 32515 20315 32521
rect 21652 32524 22652 32552
rect 20073 32487 20131 32493
rect 15580 32456 17954 32484
rect 13357 32419 13415 32425
rect 13357 32385 13369 32419
rect 13403 32385 13415 32419
rect 13357 32379 13415 32385
rect 13624 32419 13682 32425
rect 13624 32385 13636 32419
rect 13670 32416 13682 32419
rect 14090 32416 14096 32428
rect 13670 32388 14096 32416
rect 13670 32385 13682 32388
rect 13624 32379 13682 32385
rect 14090 32376 14096 32388
rect 14148 32376 14154 32428
rect 15378 32416 15384 32428
rect 15339 32388 15384 32416
rect 15378 32376 15384 32388
rect 15436 32376 15442 32428
rect 16669 32419 16727 32425
rect 16669 32385 16681 32419
rect 16715 32385 16727 32419
rect 16850 32416 16856 32428
rect 16811 32388 16856 32416
rect 16669 32379 16727 32385
rect 2225 32351 2283 32357
rect 2225 32317 2237 32351
rect 2271 32348 2283 32351
rect 2958 32348 2964 32360
rect 2271 32320 2964 32348
rect 2271 32317 2283 32320
rect 2225 32311 2283 32317
rect 2958 32308 2964 32320
rect 3016 32308 3022 32360
rect 3050 32308 3056 32360
rect 3108 32348 3114 32360
rect 3108 32320 3153 32348
rect 3108 32308 3114 32320
rect 15562 32308 15568 32360
rect 15620 32348 15626 32360
rect 15657 32351 15715 32357
rect 15657 32348 15669 32351
rect 15620 32320 15669 32348
rect 15620 32308 15626 32320
rect 15657 32317 15669 32320
rect 15703 32317 15715 32351
rect 16684 32348 16712 32379
rect 16850 32376 16856 32388
rect 16908 32376 16914 32428
rect 17926 32416 17954 32456
rect 19168 32456 19748 32484
rect 19168 32428 19196 32456
rect 19015 32419 19073 32425
rect 19015 32416 19027 32419
rect 17926 32388 19027 32416
rect 19015 32385 19027 32388
rect 19061 32385 19073 32419
rect 19150 32416 19156 32428
rect 19111 32388 19156 32416
rect 19015 32379 19073 32385
rect 19150 32376 19156 32388
rect 19208 32376 19214 32428
rect 19245 32419 19303 32425
rect 19245 32385 19257 32419
rect 19291 32385 19303 32419
rect 19426 32416 19432 32428
rect 19387 32388 19432 32416
rect 19245 32379 19303 32385
rect 18046 32348 18052 32360
rect 16684 32320 18052 32348
rect 15657 32311 15715 32317
rect 18046 32308 18052 32320
rect 18104 32308 18110 32360
rect 18690 32308 18696 32360
rect 18748 32348 18754 32360
rect 19260 32348 19288 32379
rect 19426 32376 19432 32388
rect 19484 32376 19490 32428
rect 18748 32320 19288 32348
rect 19720 32348 19748 32456
rect 20073 32453 20085 32487
rect 20119 32484 20131 32487
rect 20622 32484 20628 32496
rect 20119 32456 20628 32484
rect 20119 32453 20131 32456
rect 20073 32447 20131 32453
rect 20622 32444 20628 32456
rect 20680 32444 20686 32496
rect 20809 32487 20867 32493
rect 20809 32453 20821 32487
rect 20855 32484 20867 32487
rect 21542 32484 21548 32496
rect 20855 32456 21548 32484
rect 20855 32453 20867 32456
rect 20809 32447 20867 32453
rect 21542 32444 21548 32456
rect 21600 32444 21606 32496
rect 19886 32416 19892 32428
rect 19847 32388 19892 32416
rect 19886 32376 19892 32388
rect 19944 32416 19950 32428
rect 21652 32416 21680 32524
rect 22646 32512 22652 32524
rect 22704 32552 22710 32564
rect 23014 32552 23020 32564
rect 22704 32524 23020 32552
rect 22704 32512 22710 32524
rect 23014 32512 23020 32524
rect 23072 32512 23078 32564
rect 23842 32552 23848 32564
rect 23803 32524 23848 32552
rect 23842 32512 23848 32524
rect 23900 32512 23906 32564
rect 24118 32512 24124 32564
rect 24176 32552 24182 32564
rect 27614 32552 27620 32564
rect 24176 32524 27620 32552
rect 24176 32512 24182 32524
rect 27614 32512 27620 32524
rect 27672 32512 27678 32564
rect 28074 32512 28080 32564
rect 28132 32552 28138 32564
rect 28534 32552 28540 32564
rect 28132 32524 28540 32552
rect 28132 32512 28138 32524
rect 28534 32512 28540 32524
rect 28592 32552 28598 32564
rect 28813 32555 28871 32561
rect 28813 32552 28825 32555
rect 28592 32524 28825 32552
rect 28592 32512 28598 32524
rect 28813 32521 28825 32524
rect 28859 32521 28871 32555
rect 29362 32552 29368 32564
rect 29323 32524 29368 32552
rect 28813 32515 28871 32521
rect 29362 32512 29368 32524
rect 29420 32512 29426 32564
rect 29730 32512 29736 32564
rect 29788 32512 29794 32564
rect 29914 32512 29920 32564
rect 29972 32512 29978 32564
rect 21726 32444 21732 32496
rect 21784 32484 21790 32496
rect 23750 32484 23756 32496
rect 21784 32456 23756 32484
rect 21784 32444 21790 32456
rect 23750 32444 23756 32456
rect 23808 32444 23814 32496
rect 23952 32456 24237 32484
rect 19944 32388 21680 32416
rect 19944 32376 19950 32388
rect 21910 32376 21916 32428
rect 21968 32416 21974 32428
rect 22281 32419 22339 32425
rect 22281 32416 22293 32419
rect 21968 32388 22293 32416
rect 21968 32376 21974 32388
rect 22281 32385 22293 32388
rect 22327 32416 22339 32419
rect 22554 32416 22560 32428
rect 22327 32388 22560 32416
rect 22327 32385 22339 32388
rect 22281 32379 22339 32385
rect 22554 32376 22560 32388
rect 22612 32376 22618 32428
rect 23014 32416 23020 32428
rect 22975 32388 23020 32416
rect 23014 32376 23020 32388
rect 23072 32376 23078 32428
rect 23198 32416 23204 32428
rect 23159 32388 23204 32416
rect 23198 32376 23204 32388
rect 23256 32376 23262 32428
rect 22462 32348 22468 32360
rect 19720 32320 22468 32348
rect 18748 32308 18754 32320
rect 22462 32308 22468 32320
rect 22520 32348 22526 32360
rect 22830 32348 22836 32360
rect 22520 32320 22836 32348
rect 22520 32308 22526 32320
rect 22830 32308 22836 32320
rect 22888 32348 22894 32360
rect 23952 32348 23980 32456
rect 24209 32428 24237 32456
rect 25774 32444 25780 32496
rect 25832 32484 25838 32496
rect 25832 32456 28948 32484
rect 25832 32444 25838 32456
rect 24101 32419 24159 32425
rect 24101 32385 24113 32419
rect 24147 32385 24159 32419
rect 24101 32379 24159 32385
rect 24194 32422 24252 32428
rect 24194 32388 24206 32422
rect 24240 32388 24252 32422
rect 24194 32382 24252 32388
rect 22888 32320 23980 32348
rect 22888 32308 22894 32320
rect 22370 32280 22376 32292
rect 14292 32252 22376 32280
rect 12158 32172 12164 32224
rect 12216 32212 12222 32224
rect 14292 32212 14320 32252
rect 22370 32240 22376 32252
rect 22428 32240 22434 32292
rect 24116 32280 24144 32379
rect 24302 32376 24308 32428
rect 24360 32416 24366 32428
rect 24360 32388 24405 32416
rect 24360 32376 24366 32388
rect 24486 32376 24492 32428
rect 24544 32416 24550 32428
rect 26237 32419 26295 32425
rect 24544 32388 24589 32416
rect 24544 32376 24550 32388
rect 26237 32385 26249 32419
rect 26283 32416 26295 32419
rect 26418 32416 26424 32428
rect 26283 32388 26424 32416
rect 26283 32385 26295 32388
rect 26237 32379 26295 32385
rect 26418 32376 26424 32388
rect 26476 32376 26482 32428
rect 27338 32416 27344 32428
rect 27299 32388 27344 32416
rect 27338 32376 27344 32388
rect 27396 32376 27402 32428
rect 27430 32419 27488 32425
rect 27430 32385 27442 32419
rect 27476 32385 27488 32419
rect 27430 32379 27488 32385
rect 27546 32419 27604 32425
rect 27546 32385 27558 32419
rect 27592 32416 27604 32419
rect 27706 32416 27712 32428
rect 27592 32385 27614 32416
rect 27667 32388 27712 32416
rect 27546 32379 27614 32385
rect 26878 32308 26884 32360
rect 26936 32348 26942 32360
rect 27445 32348 27473 32379
rect 26936 32320 27473 32348
rect 27586 32348 27614 32379
rect 27706 32376 27712 32388
rect 27764 32416 27770 32428
rect 27764 32388 28672 32416
rect 27764 32376 27770 32388
rect 28350 32348 28356 32360
rect 27586 32320 28356 32348
rect 26936 32308 26942 32320
rect 28350 32308 28356 32320
rect 28408 32308 28414 32360
rect 28644 32348 28672 32388
rect 28718 32376 28724 32428
rect 28776 32416 28782 32428
rect 28920 32416 28948 32456
rect 29748 32431 29776 32512
rect 29746 32425 29804 32431
rect 29595 32419 29653 32425
rect 29595 32416 29607 32419
rect 28776 32388 28821 32416
rect 28920 32388 29607 32416
rect 28776 32376 28782 32388
rect 29595 32385 29607 32388
rect 29641 32385 29653 32419
rect 29746 32391 29758 32425
rect 29792 32391 29804 32425
rect 29746 32385 29804 32391
rect 29846 32422 29904 32428
rect 29846 32388 29858 32422
rect 29892 32419 29904 32422
rect 29932 32419 29960 32512
rect 30561 32487 30619 32493
rect 30561 32453 30573 32487
rect 30607 32484 30619 32487
rect 30742 32484 30748 32496
rect 30607 32456 30748 32484
rect 30607 32453 30619 32456
rect 30561 32447 30619 32453
rect 30742 32444 30748 32456
rect 30800 32444 30806 32496
rect 29892 32391 29960 32419
rect 30009 32419 30067 32425
rect 29892 32388 29904 32391
rect 29595 32379 29653 32385
rect 29846 32382 29904 32388
rect 30009 32385 30021 32419
rect 30055 32385 30067 32419
rect 47670 32416 47676 32428
rect 47631 32388 47676 32416
rect 30009 32379 30067 32385
rect 30024 32348 30052 32379
rect 47670 32376 47676 32388
rect 47728 32376 47734 32428
rect 30190 32348 30196 32360
rect 28644 32320 30196 32348
rect 30190 32308 30196 32320
rect 30248 32308 30254 32360
rect 47486 32308 47492 32360
rect 47544 32348 47550 32360
rect 47857 32351 47915 32357
rect 47857 32348 47869 32351
rect 47544 32320 47869 32348
rect 47544 32308 47550 32320
rect 47857 32317 47869 32320
rect 47903 32317 47915 32351
rect 47857 32311 47915 32317
rect 24302 32280 24308 32292
rect 24116 32252 24308 32280
rect 24302 32240 24308 32252
rect 24360 32240 24366 32292
rect 25774 32240 25780 32292
rect 25832 32280 25838 32292
rect 39206 32280 39212 32292
rect 25832 32252 39212 32280
rect 25832 32240 25838 32252
rect 39206 32240 39212 32252
rect 39264 32240 39270 32292
rect 12216 32184 14320 32212
rect 14737 32215 14795 32221
rect 12216 32172 12222 32184
rect 14737 32181 14749 32215
rect 14783 32212 14795 32215
rect 15194 32212 15200 32224
rect 14783 32184 15200 32212
rect 14783 32181 14795 32184
rect 14737 32175 14795 32181
rect 15194 32172 15200 32184
rect 15252 32212 15258 32224
rect 15470 32212 15476 32224
rect 15252 32184 15476 32212
rect 15252 32172 15258 32184
rect 15470 32172 15476 32184
rect 15528 32172 15534 32224
rect 18782 32212 18788 32224
rect 18743 32184 18788 32212
rect 18782 32172 18788 32184
rect 18840 32172 18846 32224
rect 18874 32172 18880 32224
rect 18932 32212 18938 32224
rect 19886 32212 19892 32224
rect 18932 32184 19892 32212
rect 18932 32172 18938 32184
rect 19886 32172 19892 32184
rect 19944 32172 19950 32224
rect 20898 32212 20904 32224
rect 20859 32184 20904 32212
rect 20898 32172 20904 32184
rect 20956 32172 20962 32224
rect 23385 32215 23443 32221
rect 23385 32181 23397 32215
rect 23431 32212 23443 32215
rect 23750 32212 23756 32224
rect 23431 32184 23756 32212
rect 23431 32181 23443 32184
rect 23385 32175 23443 32181
rect 23750 32172 23756 32184
rect 23808 32172 23814 32224
rect 26142 32172 26148 32224
rect 26200 32212 26206 32224
rect 26329 32215 26387 32221
rect 26329 32212 26341 32215
rect 26200 32184 26341 32212
rect 26200 32172 26206 32184
rect 26329 32181 26341 32184
rect 26375 32212 26387 32215
rect 26878 32212 26884 32224
rect 26375 32184 26884 32212
rect 26375 32181 26387 32184
rect 26329 32175 26387 32181
rect 26878 32172 26884 32184
rect 26936 32172 26942 32224
rect 27065 32215 27123 32221
rect 27065 32181 27077 32215
rect 27111 32212 27123 32215
rect 27614 32212 27620 32224
rect 27111 32184 27620 32212
rect 27111 32181 27123 32184
rect 27065 32175 27123 32181
rect 27614 32172 27620 32184
rect 27672 32172 27678 32224
rect 28166 32172 28172 32224
rect 28224 32212 28230 32224
rect 28718 32212 28724 32224
rect 28224 32184 28724 32212
rect 28224 32172 28230 32184
rect 28718 32172 28724 32184
rect 28776 32172 28782 32224
rect 29454 32172 29460 32224
rect 29512 32212 29518 32224
rect 30282 32212 30288 32224
rect 29512 32184 30288 32212
rect 29512 32172 29518 32184
rect 30282 32172 30288 32184
rect 30340 32212 30346 32224
rect 30653 32215 30711 32221
rect 30653 32212 30665 32215
rect 30340 32184 30665 32212
rect 30340 32172 30346 32184
rect 30653 32181 30665 32184
rect 30699 32181 30711 32215
rect 30653 32175 30711 32181
rect 31754 32172 31760 32224
rect 31812 32212 31818 32224
rect 33042 32212 33048 32224
rect 31812 32184 33048 32212
rect 31812 32172 31818 32184
rect 33042 32172 33048 32184
rect 33100 32172 33106 32224
rect 1104 32122 48852 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 48852 32122
rect 1104 32048 48852 32070
rect 1581 32011 1639 32017
rect 1581 31977 1593 32011
rect 1627 32008 1639 32011
rect 2590 32008 2596 32020
rect 1627 31980 2596 32008
rect 1627 31977 1639 31980
rect 1581 31971 1639 31977
rect 2590 31968 2596 31980
rect 2648 31968 2654 32020
rect 2958 32008 2964 32020
rect 2919 31980 2964 32008
rect 2958 31968 2964 31980
rect 3016 31968 3022 32020
rect 14090 32008 14096 32020
rect 14051 31980 14096 32008
rect 14090 31968 14096 31980
rect 14148 31968 14154 32020
rect 17402 32008 17408 32020
rect 17363 31980 17408 32008
rect 17402 31968 17408 31980
rect 17460 31968 17466 32020
rect 18690 32008 18696 32020
rect 18651 31980 18696 32008
rect 18690 31968 18696 31980
rect 18748 31968 18754 32020
rect 20625 32011 20683 32017
rect 20625 32008 20637 32011
rect 19260 31980 20637 32008
rect 15286 31940 15292 31952
rect 14292 31912 15292 31940
rect 13170 31872 13176 31884
rect 12406 31844 13176 31872
rect 1394 31804 1400 31816
rect 1355 31776 1400 31804
rect 1394 31764 1400 31776
rect 1452 31764 1458 31816
rect 1946 31764 1952 31816
rect 2004 31804 2010 31816
rect 2317 31807 2375 31813
rect 2317 31804 2329 31807
rect 2004 31776 2329 31804
rect 2004 31764 2010 31776
rect 2317 31773 2329 31776
rect 2363 31773 2375 31807
rect 2317 31767 2375 31773
rect 2869 31807 2927 31813
rect 2869 31773 2881 31807
rect 2915 31804 2927 31807
rect 12158 31804 12164 31816
rect 2915 31776 12164 31804
rect 2915 31773 2927 31776
rect 2869 31767 2927 31773
rect 12158 31764 12164 31776
rect 12216 31764 12222 31816
rect 12250 31736 12256 31748
rect 12211 31708 12256 31736
rect 12250 31696 12256 31708
rect 12308 31696 12314 31748
rect 12406 31745 12434 31844
rect 13170 31832 13176 31844
rect 13228 31832 13234 31884
rect 14292 31813 14320 31912
rect 15286 31900 15292 31912
rect 15344 31900 15350 31952
rect 19260 31940 19288 31980
rect 20625 31977 20637 31980
rect 20671 31977 20683 32011
rect 20625 31971 20683 31977
rect 22097 32011 22155 32017
rect 22097 31977 22109 32011
rect 22143 32008 22155 32011
rect 23934 32008 23940 32020
rect 22143 31980 23940 32008
rect 22143 31977 22155 31980
rect 22097 31971 22155 31977
rect 18524 31912 19288 31940
rect 20640 31940 20668 31971
rect 23934 31968 23940 31980
rect 23992 31968 23998 32020
rect 25682 31968 25688 32020
rect 25740 32008 25746 32020
rect 25777 32011 25835 32017
rect 25777 32008 25789 32011
rect 25740 31980 25789 32008
rect 25740 31968 25746 31980
rect 25777 31977 25789 31980
rect 25823 32008 25835 32011
rect 29638 32008 29644 32020
rect 25823 31980 29644 32008
rect 25823 31977 25835 31980
rect 25777 31971 25835 31977
rect 29638 31968 29644 31980
rect 29696 31968 29702 32020
rect 22922 31940 22928 31952
rect 20640 31912 22928 31940
rect 15194 31872 15200 31884
rect 14476 31844 15200 31872
rect 14476 31813 14504 31844
rect 15194 31832 15200 31844
rect 15252 31832 15258 31884
rect 14277 31807 14335 31813
rect 14277 31773 14289 31807
rect 14323 31773 14335 31807
rect 14277 31767 14335 31773
rect 14461 31807 14519 31813
rect 14461 31773 14473 31807
rect 14507 31773 14519 31807
rect 14461 31767 14519 31773
rect 14550 31764 14556 31816
rect 14608 31804 14614 31816
rect 15381 31807 15439 31813
rect 15381 31804 15393 31807
rect 14608 31776 14653 31804
rect 14844 31776 15393 31804
rect 14608 31764 14614 31776
rect 12406 31739 12484 31745
rect 12406 31708 12438 31739
rect 12426 31705 12438 31708
rect 12472 31705 12484 31739
rect 14844 31736 14872 31776
rect 15381 31773 15393 31776
rect 15427 31804 15439 31807
rect 17126 31804 17132 31816
rect 15427 31776 17132 31804
rect 15427 31773 15439 31776
rect 15381 31767 15439 31773
rect 17126 31764 17132 31776
rect 17184 31764 17190 31816
rect 17221 31807 17279 31813
rect 17221 31773 17233 31807
rect 17267 31804 17279 31807
rect 18046 31804 18052 31816
rect 17267 31776 18052 31804
rect 17267 31773 17279 31776
rect 17221 31767 17279 31773
rect 18046 31764 18052 31776
rect 18104 31764 18110 31816
rect 18524 31813 18552 31912
rect 22922 31900 22928 31912
rect 22980 31900 22986 31952
rect 27617 31943 27675 31949
rect 23124 31912 24440 31940
rect 19242 31872 19248 31884
rect 19203 31844 19248 31872
rect 19242 31832 19248 31844
rect 19300 31832 19306 31884
rect 21818 31832 21824 31884
rect 21876 31872 21882 31884
rect 23124 31872 23152 31912
rect 24412 31881 24440 31912
rect 27617 31909 27629 31943
rect 27663 31909 27675 31943
rect 29546 31940 29552 31952
rect 27617 31903 27675 31909
rect 28092 31912 29552 31940
rect 21876 31844 23152 31872
rect 23201 31875 23259 31881
rect 21876 31832 21882 31844
rect 23201 31841 23213 31875
rect 23247 31872 23259 31875
rect 24397 31875 24455 31881
rect 23247 31844 23971 31872
rect 23247 31841 23259 31844
rect 23201 31835 23259 31841
rect 18509 31807 18567 31813
rect 18509 31773 18521 31807
rect 18555 31773 18567 31807
rect 18509 31767 18567 31773
rect 18782 31764 18788 31816
rect 18840 31804 18846 31816
rect 19501 31807 19559 31813
rect 19501 31804 19513 31807
rect 18840 31776 19513 31804
rect 18840 31764 18846 31776
rect 19501 31773 19513 31776
rect 19547 31773 19559 31807
rect 19501 31767 19559 31773
rect 21453 31807 21511 31813
rect 21453 31773 21465 31807
rect 21499 31804 21511 31807
rect 21910 31804 21916 31816
rect 21499 31776 21916 31804
rect 21499 31773 21511 31776
rect 21453 31767 21511 31773
rect 21910 31764 21916 31776
rect 21968 31764 21974 31816
rect 22353 31807 22411 31813
rect 22353 31804 22365 31807
rect 22296 31776 22365 31804
rect 12426 31699 12484 31705
rect 12544 31708 14872 31736
rect 15648 31739 15706 31745
rect 11514 31628 11520 31680
rect 11572 31668 11578 31680
rect 12544 31668 12572 31708
rect 15648 31705 15660 31739
rect 15694 31736 15706 31739
rect 15838 31736 15844 31748
rect 15694 31708 15844 31736
rect 15694 31705 15706 31708
rect 15648 31699 15706 31705
rect 15838 31696 15844 31708
rect 15896 31696 15902 31748
rect 18325 31739 18383 31745
rect 18325 31705 18337 31739
rect 18371 31736 18383 31739
rect 18874 31736 18880 31748
rect 18371 31708 18880 31736
rect 18371 31705 18383 31708
rect 18325 31699 18383 31705
rect 18874 31696 18880 31708
rect 18932 31696 18938 31748
rect 11572 31640 12572 31668
rect 11572 31628 11578 31640
rect 12618 31628 12624 31680
rect 12676 31668 12682 31680
rect 12676 31640 12721 31668
rect 12676 31628 12682 31640
rect 15562 31628 15568 31680
rect 15620 31668 15626 31680
rect 16761 31671 16819 31677
rect 16761 31668 16773 31671
rect 15620 31640 16773 31668
rect 15620 31628 15626 31640
rect 16761 31637 16773 31640
rect 16807 31637 16819 31671
rect 16761 31631 16819 31637
rect 19426 31628 19432 31680
rect 19484 31668 19490 31680
rect 21266 31668 21272 31680
rect 19484 31640 21272 31668
rect 19484 31628 19490 31640
rect 21266 31628 21272 31640
rect 21324 31628 21330 31680
rect 21450 31628 21456 31680
rect 21508 31668 21514 31680
rect 21545 31671 21603 31677
rect 21545 31668 21557 31671
rect 21508 31640 21557 31668
rect 21508 31628 21514 31640
rect 21545 31637 21557 31640
rect 21591 31637 21603 31671
rect 22296 31668 22324 31776
rect 22353 31773 22365 31776
rect 22399 31773 22411 31807
rect 22353 31767 22411 31773
rect 22446 31804 22504 31810
rect 22446 31770 22458 31804
rect 22492 31770 22504 31804
rect 22446 31764 22504 31770
rect 22461 31736 22489 31764
rect 22554 31758 22560 31810
rect 22612 31798 22618 31810
rect 22738 31804 22744 31816
rect 22612 31770 22657 31798
rect 22699 31776 22744 31804
rect 22612 31758 22618 31770
rect 22738 31764 22744 31776
rect 22796 31764 22802 31816
rect 23474 31804 23480 31816
rect 23435 31776 23480 31804
rect 23474 31764 23480 31776
rect 23532 31764 23538 31816
rect 23569 31807 23627 31813
rect 23569 31773 23581 31807
rect 23615 31773 23627 31807
rect 23569 31767 23627 31773
rect 23661 31807 23719 31813
rect 23661 31773 23673 31807
rect 23707 31801 23719 31807
rect 23750 31801 23756 31816
rect 23707 31773 23756 31801
rect 23661 31767 23719 31773
rect 22461 31708 22508 31736
rect 22480 31680 22508 31708
rect 22830 31696 22836 31748
rect 22888 31736 22894 31748
rect 23584 31736 23612 31767
rect 23750 31764 23756 31773
rect 23808 31764 23814 31816
rect 23845 31807 23903 31813
rect 23845 31773 23857 31807
rect 23891 31773 23903 31807
rect 23943 31804 23971 31844
rect 24397 31841 24409 31875
rect 24443 31841 24455 31875
rect 27632 31872 27660 31903
rect 28092 31881 28120 31912
rect 29546 31900 29552 31912
rect 29604 31900 29610 31952
rect 31021 31943 31079 31949
rect 31021 31940 31033 31943
rect 30024 31912 31033 31940
rect 24397 31835 24455 31841
rect 26804 31844 27660 31872
rect 28077 31875 28135 31881
rect 24653 31807 24711 31813
rect 24653 31804 24665 31807
rect 23943 31776 24665 31804
rect 23845 31767 23903 31773
rect 24653 31773 24665 31776
rect 24699 31773 24711 31807
rect 24653 31767 24711 31773
rect 23860 31736 23888 31767
rect 26804 31745 26832 31844
rect 28077 31841 28089 31875
rect 28123 31841 28135 31875
rect 28077 31835 28135 31841
rect 28261 31875 28319 31881
rect 28261 31841 28273 31875
rect 28307 31872 28319 31875
rect 28534 31872 28540 31884
rect 28307 31844 28540 31872
rect 28307 31841 28319 31844
rect 28261 31835 28319 31841
rect 28534 31832 28540 31844
rect 28592 31872 28598 31884
rect 28902 31872 28908 31884
rect 28592 31844 28908 31872
rect 28592 31832 28598 31844
rect 28902 31832 28908 31844
rect 28960 31832 28966 31884
rect 26878 31764 26884 31816
rect 26936 31804 26942 31816
rect 26936 31776 29592 31804
rect 26936 31764 26942 31776
rect 22888 31708 23612 31736
rect 23759 31708 23888 31736
rect 26789 31739 26847 31745
rect 22888 31696 22894 31708
rect 22370 31668 22376 31680
rect 22296 31640 22376 31668
rect 21545 31631 21603 31637
rect 22370 31628 22376 31640
rect 22428 31628 22434 31680
rect 22462 31628 22468 31680
rect 22520 31628 22526 31680
rect 22738 31628 22744 31680
rect 22796 31668 22802 31680
rect 23759 31668 23787 31708
rect 26789 31705 26801 31739
rect 26835 31705 26847 31739
rect 26789 31699 26847 31705
rect 26973 31739 27031 31745
rect 26973 31705 26985 31739
rect 27019 31736 27031 31739
rect 27522 31736 27528 31748
rect 27019 31708 27528 31736
rect 27019 31705 27031 31708
rect 26973 31699 27031 31705
rect 27522 31696 27528 31708
rect 27580 31736 27586 31748
rect 29362 31736 29368 31748
rect 27580 31708 29368 31736
rect 27580 31696 27586 31708
rect 29362 31696 29368 31708
rect 29420 31696 29426 31748
rect 29564 31736 29592 31776
rect 29638 31764 29644 31816
rect 29696 31804 29702 31816
rect 30024 31813 30052 31912
rect 31021 31909 31033 31912
rect 31067 31909 31079 31943
rect 31754 31940 31760 31952
rect 31715 31912 31760 31940
rect 31021 31903 31079 31909
rect 31754 31900 31760 31912
rect 31812 31900 31818 31952
rect 30282 31832 30288 31884
rect 30340 31872 30346 31884
rect 30340 31844 31616 31872
rect 30340 31832 30346 31844
rect 29779 31807 29837 31813
rect 29779 31804 29791 31807
rect 29696 31776 29791 31804
rect 29696 31764 29702 31776
rect 29779 31773 29791 31776
rect 29825 31773 29837 31807
rect 29779 31767 29837 31773
rect 29917 31807 29975 31813
rect 29917 31773 29929 31807
rect 29963 31773 29975 31807
rect 29917 31767 29975 31773
rect 30014 31807 30072 31813
rect 30014 31773 30026 31807
rect 30060 31773 30072 31807
rect 30190 31804 30196 31816
rect 30151 31776 30196 31804
rect 30014 31767 30072 31773
rect 29932 31736 29960 31767
rect 30190 31764 30196 31776
rect 30248 31764 30254 31816
rect 31588 31813 31616 31844
rect 45922 31832 45928 31884
rect 45980 31872 45986 31884
rect 47581 31875 47639 31881
rect 47581 31872 47593 31875
rect 45980 31844 47593 31872
rect 45980 31832 45986 31844
rect 47581 31841 47593 31844
rect 47627 31841 47639 31875
rect 47581 31835 47639 31841
rect 31573 31807 31631 31813
rect 31573 31773 31585 31807
rect 31619 31773 31631 31807
rect 31573 31767 31631 31773
rect 32490 31764 32496 31816
rect 32548 31801 32554 31816
rect 32585 31807 32643 31813
rect 32585 31801 32597 31807
rect 32548 31773 32597 31801
rect 32631 31773 32643 31807
rect 32677 31807 32735 31813
rect 32677 31804 32689 31807
rect 32548 31764 32554 31773
rect 32585 31767 32643 31773
rect 32673 31773 32689 31804
rect 32723 31773 32735 31807
rect 32673 31767 32735 31773
rect 29564 31708 29960 31736
rect 22796 31640 23787 31668
rect 22796 31628 22802 31640
rect 26234 31628 26240 31680
rect 26292 31668 26298 31680
rect 27157 31671 27215 31677
rect 27157 31668 27169 31671
rect 26292 31640 27169 31668
rect 26292 31628 26298 31640
rect 27157 31637 27169 31640
rect 27203 31637 27215 31671
rect 27157 31631 27215 31637
rect 27430 31628 27436 31680
rect 27488 31668 27494 31680
rect 27985 31671 28043 31677
rect 27985 31668 27997 31671
rect 27488 31640 27997 31668
rect 27488 31628 27494 31640
rect 27985 31637 27997 31640
rect 28031 31637 28043 31671
rect 27985 31631 28043 31637
rect 29549 31671 29607 31677
rect 29549 31637 29561 31671
rect 29595 31668 29607 31671
rect 29822 31668 29828 31680
rect 29595 31640 29828 31668
rect 29595 31637 29607 31640
rect 29549 31631 29607 31637
rect 29822 31628 29828 31640
rect 29880 31628 29886 31680
rect 29932 31668 29960 31708
rect 30374 31696 30380 31748
rect 30432 31736 30438 31748
rect 30653 31739 30711 31745
rect 30653 31736 30665 31739
rect 30432 31708 30665 31736
rect 30432 31696 30438 31708
rect 30653 31705 30665 31708
rect 30699 31705 30711 31739
rect 30653 31699 30711 31705
rect 30742 31696 30748 31748
rect 30800 31736 30806 31748
rect 30837 31739 30895 31745
rect 30837 31736 30849 31739
rect 30800 31708 30849 31736
rect 30800 31696 30806 31708
rect 30837 31705 30849 31708
rect 30883 31705 30895 31739
rect 32398 31736 32404 31748
rect 30837 31699 30895 31705
rect 32232 31708 32404 31736
rect 32232 31668 32260 31708
rect 32398 31696 32404 31708
rect 32456 31736 32462 31748
rect 32673 31736 32701 31767
rect 32766 31764 32772 31816
rect 32824 31804 32830 31816
rect 32953 31807 33011 31813
rect 32824 31776 32869 31804
rect 32824 31764 32830 31776
rect 32953 31773 32965 31807
rect 32999 31804 33011 31807
rect 33502 31804 33508 31816
rect 32999 31776 33508 31804
rect 32999 31773 33011 31776
rect 32953 31767 33011 31773
rect 33502 31764 33508 31776
rect 33560 31764 33566 31816
rect 47302 31804 47308 31816
rect 47263 31776 47308 31804
rect 47302 31764 47308 31776
rect 47360 31764 47366 31816
rect 32456 31708 32701 31736
rect 32456 31696 32462 31708
rect 29932 31640 32260 31668
rect 32309 31671 32367 31677
rect 32309 31637 32321 31671
rect 32355 31668 32367 31671
rect 33318 31668 33324 31680
rect 32355 31640 33324 31668
rect 32355 31637 32367 31640
rect 32309 31631 32367 31637
rect 33318 31628 33324 31640
rect 33376 31628 33382 31680
rect 1104 31578 48852 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 48852 31578
rect 1104 31504 48852 31526
rect 4798 31424 4804 31476
rect 4856 31464 4862 31476
rect 13170 31464 13176 31476
rect 4856 31436 12204 31464
rect 13131 31436 13176 31464
rect 4856 31424 4862 31436
rect 11514 31396 11520 31408
rect 9508 31368 11520 31396
rect 1946 31328 1952 31340
rect 1907 31300 1952 31328
rect 1946 31288 1952 31300
rect 2004 31288 2010 31340
rect 2133 31263 2191 31269
rect 2133 31229 2145 31263
rect 2179 31260 2191 31263
rect 2866 31260 2872 31272
rect 2179 31232 2872 31260
rect 2179 31229 2191 31232
rect 2133 31223 2191 31229
rect 2866 31220 2872 31232
rect 2924 31220 2930 31272
rect 3050 31260 3056 31272
rect 3011 31232 3056 31260
rect 3050 31220 3056 31232
rect 3108 31220 3114 31272
rect 8478 31220 8484 31272
rect 8536 31260 8542 31272
rect 9508 31269 9536 31368
rect 11514 31356 11520 31368
rect 11572 31396 11578 31408
rect 11572 31368 11836 31396
rect 11572 31356 11578 31368
rect 9760 31331 9818 31337
rect 9760 31297 9772 31331
rect 9806 31328 9818 31331
rect 10318 31328 10324 31340
rect 9806 31300 10324 31328
rect 9806 31297 9818 31300
rect 9760 31291 9818 31297
rect 10318 31288 10324 31300
rect 10376 31288 10382 31340
rect 11808 31337 11836 31368
rect 11793 31331 11851 31337
rect 11793 31297 11805 31331
rect 11839 31297 11851 31331
rect 11793 31291 11851 31297
rect 11882 31288 11888 31340
rect 11940 31328 11946 31340
rect 12049 31331 12107 31337
rect 12049 31328 12061 31331
rect 11940 31300 12061 31328
rect 11940 31288 11946 31300
rect 12049 31297 12061 31300
rect 12095 31297 12107 31331
rect 12176 31328 12204 31436
rect 13170 31424 13176 31436
rect 13228 31464 13234 31476
rect 14090 31464 14096 31476
rect 13228 31436 14096 31464
rect 13228 31424 13234 31436
rect 14090 31424 14096 31436
rect 14148 31424 14154 31476
rect 15378 31424 15384 31476
rect 15436 31464 15442 31476
rect 15930 31464 15936 31476
rect 15436 31436 15936 31464
rect 15436 31424 15442 31436
rect 15930 31424 15936 31436
rect 15988 31424 15994 31476
rect 16025 31467 16083 31473
rect 16025 31433 16037 31467
rect 16071 31464 16083 31467
rect 16850 31464 16856 31476
rect 16071 31436 16856 31464
rect 16071 31433 16083 31436
rect 16025 31427 16083 31433
rect 16850 31424 16856 31436
rect 16908 31464 16914 31476
rect 17037 31467 17095 31473
rect 17037 31464 17049 31467
rect 16908 31436 17049 31464
rect 16908 31424 16914 31436
rect 17037 31433 17049 31436
rect 17083 31433 17095 31467
rect 17037 31427 17095 31433
rect 18693 31467 18751 31473
rect 18693 31433 18705 31467
rect 18739 31464 18751 31467
rect 18874 31464 18880 31476
rect 18739 31436 18880 31464
rect 18739 31433 18751 31436
rect 18693 31427 18751 31433
rect 18874 31424 18880 31436
rect 18932 31424 18938 31476
rect 20625 31467 20683 31473
rect 20625 31433 20637 31467
rect 20671 31433 20683 31467
rect 20625 31427 20683 31433
rect 12250 31356 12256 31408
rect 12308 31396 12314 31408
rect 14366 31396 14372 31408
rect 12308 31368 14372 31396
rect 12308 31356 12314 31368
rect 14366 31356 14372 31368
rect 14424 31396 14430 31408
rect 14921 31399 14979 31405
rect 14921 31396 14933 31399
rect 14424 31368 14933 31396
rect 14424 31356 14430 31368
rect 14921 31365 14933 31368
rect 14967 31365 14979 31399
rect 14921 31359 14979 31365
rect 15286 31356 15292 31408
rect 15344 31396 15350 31408
rect 15841 31399 15899 31405
rect 15841 31396 15853 31399
rect 15344 31368 15853 31396
rect 15344 31356 15350 31368
rect 15841 31365 15853 31368
rect 15887 31396 15899 31399
rect 16206 31396 16212 31408
rect 15887 31368 16212 31396
rect 15887 31365 15899 31368
rect 15841 31359 15899 31365
rect 16206 31356 16212 31368
rect 16264 31356 16270 31408
rect 20640 31396 20668 31427
rect 21542 31424 21548 31476
rect 21600 31464 21606 31476
rect 23201 31467 23259 31473
rect 23201 31464 23213 31467
rect 21600 31436 23213 31464
rect 21600 31424 21606 31436
rect 23201 31433 23213 31436
rect 23247 31464 23259 31467
rect 23247 31436 26464 31464
rect 23247 31433 23259 31436
rect 23201 31427 23259 31433
rect 23934 31405 23940 31408
rect 23928 31396 23940 31405
rect 20640 31368 22120 31396
rect 23895 31368 23940 31396
rect 13354 31328 13360 31340
rect 12176 31300 13360 31328
rect 12049 31291 12107 31297
rect 13354 31288 13360 31300
rect 13412 31288 13418 31340
rect 15105 31331 15163 31337
rect 15105 31297 15117 31331
rect 15151 31328 15163 31331
rect 15562 31328 15568 31340
rect 15151 31300 15568 31328
rect 15151 31297 15163 31300
rect 15105 31291 15163 31297
rect 15562 31288 15568 31300
rect 15620 31328 15626 31340
rect 15746 31328 15752 31340
rect 15620 31300 15752 31328
rect 15620 31288 15626 31300
rect 15746 31288 15752 31300
rect 15804 31288 15810 31340
rect 16114 31288 16120 31340
rect 16172 31328 16178 31340
rect 16669 31331 16727 31337
rect 16172 31300 16217 31328
rect 16172 31288 16178 31300
rect 16669 31297 16681 31331
rect 16715 31297 16727 31331
rect 16669 31291 16727 31297
rect 9493 31263 9551 31269
rect 9493 31260 9505 31263
rect 8536 31232 9505 31260
rect 8536 31220 8542 31232
rect 9493 31229 9505 31232
rect 9539 31229 9551 31263
rect 15378 31260 15384 31272
rect 15339 31232 15384 31260
rect 9493 31223 9551 31229
rect 15378 31220 15384 31232
rect 15436 31220 15442 31272
rect 16684 31260 16712 31291
rect 18046 31288 18052 31340
rect 18104 31328 18110 31340
rect 18877 31331 18935 31337
rect 18877 31328 18889 31331
rect 18104 31300 18889 31328
rect 18104 31288 18110 31300
rect 18877 31297 18889 31300
rect 18923 31328 18935 31331
rect 19337 31331 19395 31337
rect 19337 31328 19349 31331
rect 18923 31300 19349 31328
rect 18923 31297 18935 31300
rect 18877 31291 18935 31297
rect 19337 31297 19349 31300
rect 19383 31297 19395 31331
rect 19337 31291 19395 31297
rect 20806 31288 20812 31340
rect 20864 31328 20870 31340
rect 20901 31331 20959 31337
rect 20901 31328 20913 31331
rect 20864 31300 20913 31328
rect 20864 31288 20870 31300
rect 20901 31297 20913 31300
rect 20947 31297 20959 31331
rect 20901 31291 20959 31297
rect 20993 31331 21051 31337
rect 20993 31297 21005 31331
rect 21039 31297 21051 31331
rect 20993 31291 21051 31297
rect 15672 31232 16712 31260
rect 16761 31263 16819 31269
rect 14550 31152 14556 31204
rect 14608 31192 14614 31204
rect 15672 31192 15700 31232
rect 16761 31229 16773 31263
rect 16807 31229 16819 31263
rect 16761 31223 16819 31229
rect 19613 31263 19671 31269
rect 19613 31229 19625 31263
rect 19659 31260 19671 31263
rect 20346 31260 20352 31272
rect 19659 31232 20352 31260
rect 19659 31229 19671 31232
rect 19613 31223 19671 31229
rect 15838 31192 15844 31204
rect 14608 31164 15700 31192
rect 15799 31164 15844 31192
rect 14608 31152 14614 31164
rect 15838 31152 15844 31164
rect 15896 31152 15902 31204
rect 15930 31152 15936 31204
rect 15988 31192 15994 31204
rect 16776 31192 16804 31223
rect 20346 31220 20352 31232
rect 20404 31220 20410 31272
rect 20070 31192 20076 31204
rect 15988 31164 20076 31192
rect 15988 31152 15994 31164
rect 20070 31152 20076 31164
rect 20128 31152 20134 31204
rect 21008 31192 21036 31291
rect 21082 31288 21088 31340
rect 21140 31328 21146 31340
rect 21266 31328 21272 31340
rect 21140 31300 21185 31328
rect 21227 31300 21272 31328
rect 21140 31288 21146 31300
rect 21266 31288 21272 31300
rect 21324 31288 21330 31340
rect 22092 31337 22120 31368
rect 23928 31359 23940 31368
rect 23934 31356 23940 31359
rect 23992 31356 23998 31408
rect 26436 31396 26464 31436
rect 28626 31424 28632 31476
rect 28684 31464 28690 31476
rect 28997 31467 29055 31473
rect 28997 31464 29009 31467
rect 28684 31436 29009 31464
rect 28684 31424 28690 31436
rect 28997 31433 29009 31436
rect 29043 31433 29055 31467
rect 28997 31427 29055 31433
rect 30285 31467 30343 31473
rect 30285 31433 30297 31467
rect 30331 31464 30343 31467
rect 30374 31464 30380 31476
rect 30331 31436 30380 31464
rect 30331 31433 30343 31436
rect 30285 31427 30343 31433
rect 30374 31424 30380 31436
rect 30432 31424 30438 31476
rect 30745 31467 30803 31473
rect 30745 31433 30757 31467
rect 30791 31464 30803 31467
rect 30834 31464 30840 31476
rect 30791 31436 30840 31464
rect 30791 31433 30803 31436
rect 30745 31427 30803 31433
rect 30834 31424 30840 31436
rect 30892 31424 30898 31476
rect 32585 31467 32643 31473
rect 32585 31433 32597 31467
rect 32631 31464 32643 31467
rect 32766 31464 32772 31476
rect 32631 31436 32772 31464
rect 32631 31433 32643 31436
rect 32585 31427 32643 31433
rect 32766 31424 32772 31436
rect 32824 31424 32830 31476
rect 32490 31396 32496 31408
rect 26436 31368 32496 31396
rect 32490 31356 32496 31368
rect 32548 31356 32554 31408
rect 33318 31405 33324 31408
rect 33312 31396 33324 31405
rect 33279 31368 33324 31396
rect 33312 31359 33324 31368
rect 33318 31356 33324 31359
rect 33376 31356 33382 31408
rect 22077 31331 22135 31337
rect 22077 31297 22089 31331
rect 22123 31297 22135 31331
rect 22077 31291 22135 31297
rect 22922 31288 22928 31340
rect 22980 31328 22986 31340
rect 26007 31331 26065 31337
rect 26007 31328 26019 31331
rect 22980 31300 26019 31328
rect 22980 31288 22986 31300
rect 26007 31297 26019 31300
rect 26053 31297 26065 31331
rect 26142 31328 26148 31340
rect 26103 31300 26148 31328
rect 26007 31291 26065 31297
rect 26142 31288 26148 31300
rect 26200 31288 26206 31340
rect 26234 31288 26240 31340
rect 26292 31328 26298 31340
rect 26421 31331 26479 31337
rect 26292 31300 26337 31328
rect 26292 31288 26298 31300
rect 26421 31297 26433 31331
rect 26467 31328 26479 31331
rect 27706 31328 27712 31340
rect 26467 31300 27712 31328
rect 26467 31297 26479 31300
rect 26421 31291 26479 31297
rect 27706 31288 27712 31300
rect 27764 31288 27770 31340
rect 28258 31288 28264 31340
rect 28316 31328 28322 31340
rect 28534 31328 28540 31340
rect 28316 31300 28540 31328
rect 28316 31288 28322 31300
rect 28534 31288 28540 31300
rect 28592 31288 28598 31340
rect 28718 31288 28724 31340
rect 28776 31328 28782 31340
rect 28905 31331 28963 31337
rect 28905 31328 28917 31331
rect 28776 31300 28917 31328
rect 28776 31288 28782 31300
rect 28905 31297 28917 31300
rect 28951 31297 28963 31331
rect 28905 31291 28963 31297
rect 30006 31288 30012 31340
rect 30064 31328 30070 31340
rect 30653 31331 30711 31337
rect 30653 31328 30665 31331
rect 30064 31300 30665 31328
rect 30064 31288 30070 31300
rect 30653 31297 30665 31300
rect 30699 31297 30711 31331
rect 30653 31291 30711 31297
rect 30742 31288 30748 31340
rect 30800 31328 30806 31340
rect 31938 31328 31944 31340
rect 30800 31300 31944 31328
rect 30800 31288 30806 31300
rect 31938 31288 31944 31300
rect 31996 31328 32002 31340
rect 32214 31328 32220 31340
rect 31996 31300 32076 31328
rect 32175 31300 32220 31328
rect 31996 31288 32002 31300
rect 21821 31263 21879 31269
rect 21821 31229 21833 31263
rect 21867 31229 21879 31263
rect 21821 31223 21879 31229
rect 23661 31263 23719 31269
rect 23661 31229 23673 31263
rect 23707 31229 23719 31263
rect 23661 31223 23719 31229
rect 21450 31192 21456 31204
rect 21008 31164 21456 31192
rect 21450 31152 21456 31164
rect 21508 31152 21514 31204
rect 21836 31136 21864 31223
rect 23676 31192 23704 31223
rect 26970 31220 26976 31272
rect 27028 31260 27034 31272
rect 27246 31260 27252 31272
rect 27028 31232 27252 31260
rect 27028 31220 27034 31232
rect 27246 31220 27252 31232
rect 27304 31220 27310 31272
rect 27522 31260 27528 31272
rect 27483 31232 27528 31260
rect 27522 31220 27528 31232
rect 27580 31220 27586 31272
rect 29089 31263 29147 31269
rect 29089 31229 29101 31263
rect 29135 31260 29147 31263
rect 30834 31260 30840 31272
rect 29135 31232 30840 31260
rect 29135 31229 29147 31232
rect 29089 31223 29147 31229
rect 25038 31192 25044 31204
rect 22848 31164 23704 31192
rect 24951 31164 25044 31192
rect 10134 31084 10140 31136
rect 10192 31124 10198 31136
rect 10873 31127 10931 31133
rect 10873 31124 10885 31127
rect 10192 31096 10885 31124
rect 10192 31084 10198 31096
rect 10873 31093 10885 31096
rect 10919 31093 10931 31127
rect 10873 31087 10931 31093
rect 15289 31127 15347 31133
rect 15289 31093 15301 31127
rect 15335 31124 15347 31127
rect 15470 31124 15476 31136
rect 15335 31096 15476 31124
rect 15335 31093 15347 31096
rect 15289 31087 15347 31093
rect 15470 31084 15476 31096
rect 15528 31124 15534 31136
rect 16669 31127 16727 31133
rect 16669 31124 16681 31127
rect 15528 31096 16681 31124
rect 15528 31084 15534 31096
rect 16669 31093 16681 31096
rect 16715 31093 16727 31127
rect 16669 31087 16727 31093
rect 18414 31084 18420 31136
rect 18472 31124 18478 31136
rect 20898 31124 20904 31136
rect 18472 31096 20904 31124
rect 18472 31084 18478 31096
rect 20898 31084 20904 31096
rect 20956 31084 20962 31136
rect 21818 31124 21824 31136
rect 21731 31096 21824 31124
rect 21818 31084 21824 31096
rect 21876 31124 21882 31136
rect 22848 31124 22876 31164
rect 25038 31152 25044 31164
rect 25096 31192 25102 31204
rect 27338 31192 27344 31204
rect 25096 31164 27344 31192
rect 25096 31152 25102 31164
rect 27338 31152 27344 31164
rect 27396 31152 27402 31204
rect 28902 31152 28908 31204
rect 28960 31192 28966 31204
rect 29104 31192 29132 31223
rect 30834 31220 30840 31232
rect 30892 31220 30898 31272
rect 32048 31260 32076 31300
rect 32214 31288 32220 31300
rect 32272 31288 32278 31340
rect 32401 31331 32459 31337
rect 32401 31297 32413 31331
rect 32447 31297 32459 31331
rect 33042 31328 33048 31340
rect 33003 31300 33048 31328
rect 32401 31291 32459 31297
rect 32416 31260 32444 31291
rect 33042 31288 33048 31300
rect 33100 31288 33106 31340
rect 32048 31232 32444 31260
rect 28960 31164 29132 31192
rect 28960 31152 28966 31164
rect 25774 31124 25780 31136
rect 21876 31096 22876 31124
rect 25735 31096 25780 31124
rect 21876 31084 21882 31096
rect 25774 31084 25780 31096
rect 25832 31084 25838 31136
rect 28166 31084 28172 31136
rect 28224 31124 28230 31136
rect 28537 31127 28595 31133
rect 28537 31124 28549 31127
rect 28224 31096 28549 31124
rect 28224 31084 28230 31096
rect 28537 31093 28549 31096
rect 28583 31093 28595 31127
rect 28537 31087 28595 31093
rect 33410 31084 33416 31136
rect 33468 31124 33474 31136
rect 34425 31127 34483 31133
rect 34425 31124 34437 31127
rect 33468 31096 34437 31124
rect 33468 31084 33474 31096
rect 34425 31093 34437 31096
rect 34471 31093 34483 31127
rect 34425 31087 34483 31093
rect 1104 31034 48852 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 48852 31034
rect 1104 30960 48852 30982
rect 2866 30920 2872 30932
rect 2827 30892 2872 30920
rect 2866 30880 2872 30892
rect 2924 30880 2930 30932
rect 10318 30880 10324 30932
rect 10376 30920 10382 30932
rect 10413 30923 10471 30929
rect 10413 30920 10425 30923
rect 10376 30892 10425 30920
rect 10376 30880 10382 30892
rect 10413 30889 10425 30892
rect 10459 30889 10471 30923
rect 10413 30883 10471 30889
rect 11793 30923 11851 30929
rect 11793 30889 11805 30923
rect 11839 30920 11851 30923
rect 11882 30920 11888 30932
rect 11839 30892 11888 30920
rect 11839 30889 11851 30892
rect 11793 30883 11851 30889
rect 11882 30880 11888 30892
rect 11940 30880 11946 30932
rect 16114 30880 16120 30932
rect 16172 30920 16178 30932
rect 16393 30923 16451 30929
rect 16393 30920 16405 30923
rect 16172 30892 16405 30920
rect 16172 30880 16178 30892
rect 16393 30889 16405 30892
rect 16439 30889 16451 30923
rect 16393 30883 16451 30889
rect 21082 30880 21088 30932
rect 21140 30920 21146 30932
rect 21729 30923 21787 30929
rect 21729 30920 21741 30923
rect 21140 30892 21741 30920
rect 21140 30880 21146 30892
rect 21729 30889 21741 30892
rect 21775 30889 21787 30923
rect 22554 30920 22560 30932
rect 22515 30892 22560 30920
rect 21729 30883 21787 30889
rect 22554 30880 22560 30892
rect 22612 30880 22618 30932
rect 23658 30880 23664 30932
rect 23716 30880 23722 30932
rect 28350 30880 28356 30932
rect 28408 30920 28414 30932
rect 28537 30923 28595 30929
rect 28537 30920 28549 30923
rect 28408 30892 28549 30920
rect 28408 30880 28414 30892
rect 28537 30889 28549 30892
rect 28583 30889 28595 30923
rect 28537 30883 28595 30889
rect 32214 30880 32220 30932
rect 32272 30920 32278 30932
rect 32861 30923 32919 30929
rect 32861 30920 32873 30923
rect 32272 30892 32873 30920
rect 32272 30880 32278 30892
rect 32861 30889 32873 30892
rect 32907 30889 32919 30923
rect 32861 30883 32919 30889
rect 12158 30852 12164 30864
rect 2792 30824 12164 30852
rect 1762 30676 1768 30728
rect 1820 30716 1826 30728
rect 2792 30725 2820 30824
rect 12158 30812 12164 30824
rect 12216 30812 12222 30864
rect 13262 30812 13268 30864
rect 13320 30852 13326 30864
rect 19518 30852 19524 30864
rect 13320 30824 19524 30852
rect 13320 30812 13326 30824
rect 19518 30812 19524 30824
rect 19576 30812 19582 30864
rect 21450 30852 21456 30864
rect 19628 30824 21456 30852
rect 9953 30787 10011 30793
rect 9953 30753 9965 30787
rect 9999 30784 10011 30787
rect 9999 30756 10916 30784
rect 9999 30753 10011 30756
rect 9953 30747 10011 30753
rect 2041 30719 2099 30725
rect 2041 30716 2053 30719
rect 1820 30688 2053 30716
rect 1820 30676 1826 30688
rect 2041 30685 2053 30688
rect 2087 30685 2099 30719
rect 2041 30679 2099 30685
rect 2777 30719 2835 30725
rect 2777 30685 2789 30719
rect 2823 30685 2835 30719
rect 2777 30679 2835 30685
rect 10410 30676 10416 30728
rect 10468 30716 10474 30728
rect 10643 30719 10701 30725
rect 10643 30716 10655 30719
rect 10468 30688 10655 30716
rect 10468 30676 10474 30688
rect 10643 30685 10655 30688
rect 10689 30685 10701 30719
rect 10778 30716 10784 30728
rect 10739 30688 10784 30716
rect 10643 30679 10701 30685
rect 10778 30676 10784 30688
rect 10836 30676 10842 30728
rect 10888 30725 10916 30756
rect 10980 30756 12204 30784
rect 10873 30719 10931 30725
rect 10873 30685 10885 30719
rect 10919 30685 10931 30719
rect 10873 30679 10931 30685
rect 9585 30651 9643 30657
rect 9585 30617 9597 30651
rect 9631 30648 9643 30651
rect 9674 30648 9680 30660
rect 9631 30620 9680 30648
rect 9631 30617 9643 30620
rect 9585 30611 9643 30617
rect 9674 30608 9680 30620
rect 9732 30608 9738 30660
rect 9769 30651 9827 30657
rect 9769 30617 9781 30651
rect 9815 30648 9827 30651
rect 10042 30648 10048 30660
rect 9815 30620 10048 30648
rect 9815 30617 9827 30620
rect 9769 30611 9827 30617
rect 10042 30608 10048 30620
rect 10100 30608 10106 30660
rect 10796 30648 10824 30676
rect 10980 30648 11008 30756
rect 11057 30719 11115 30725
rect 11057 30685 11069 30719
rect 11103 30685 11115 30719
rect 11057 30679 11115 30685
rect 10796 30620 11008 30648
rect 10870 30540 10876 30592
rect 10928 30580 10934 30592
rect 11072 30580 11100 30679
rect 11146 30676 11152 30728
rect 11204 30716 11210 30728
rect 12176 30725 12204 30756
rect 13354 30744 13360 30796
rect 13412 30784 13418 30796
rect 13412 30756 19564 30784
rect 13412 30744 13418 30756
rect 12069 30719 12127 30725
rect 12069 30716 12081 30719
rect 11204 30688 12081 30716
rect 11204 30676 11210 30688
rect 12069 30685 12081 30688
rect 12115 30685 12127 30719
rect 12069 30679 12127 30685
rect 12161 30719 12219 30725
rect 12161 30685 12173 30719
rect 12207 30685 12219 30719
rect 12161 30679 12219 30685
rect 12253 30719 12311 30725
rect 12253 30685 12265 30719
rect 12299 30685 12311 30719
rect 12434 30716 12440 30728
rect 12395 30688 12440 30716
rect 12253 30679 12311 30685
rect 12268 30648 12296 30679
rect 12434 30676 12440 30688
rect 12492 30676 12498 30728
rect 13262 30716 13268 30728
rect 13223 30688 13268 30716
rect 13262 30676 13268 30688
rect 13320 30676 13326 30728
rect 14090 30716 14096 30728
rect 14051 30688 14096 30716
rect 14090 30676 14096 30688
rect 14148 30676 14154 30728
rect 15470 30676 15476 30728
rect 15528 30716 15534 30728
rect 19536 30725 19564 30756
rect 19628 30725 19656 30824
rect 21450 30812 21456 30824
rect 21508 30812 21514 30864
rect 20717 30787 20775 30793
rect 20717 30784 20729 30787
rect 19720 30756 20729 30784
rect 19720 30725 19748 30756
rect 20717 30753 20729 30756
rect 20763 30753 20775 30787
rect 20717 30747 20775 30753
rect 23017 30787 23075 30793
rect 23017 30753 23029 30787
rect 23063 30784 23075 30787
rect 23106 30784 23112 30796
rect 23063 30756 23112 30784
rect 23063 30753 23075 30756
rect 23017 30747 23075 30753
rect 23106 30744 23112 30756
rect 23164 30744 23170 30796
rect 23676 30728 23704 30880
rect 27522 30812 27528 30864
rect 27580 30812 27586 30864
rect 27540 30784 27568 30812
rect 27540 30756 28396 30784
rect 16669 30719 16727 30725
rect 16669 30716 16681 30719
rect 15528 30688 16681 30716
rect 15528 30676 15534 30688
rect 16669 30685 16681 30688
rect 16715 30685 16727 30719
rect 16669 30679 16727 30685
rect 19521 30719 19579 30725
rect 19521 30685 19533 30719
rect 19567 30685 19579 30719
rect 19521 30679 19579 30685
rect 19613 30719 19671 30725
rect 19613 30685 19625 30719
rect 19659 30685 19671 30719
rect 19613 30679 19671 30685
rect 19705 30719 19763 30725
rect 19705 30685 19717 30719
rect 19751 30685 19763 30719
rect 19705 30679 19763 30685
rect 19889 30719 19947 30725
rect 19889 30685 19901 30719
rect 19935 30685 19947 30719
rect 20346 30716 20352 30728
rect 20307 30688 20352 30716
rect 19889 30679 19947 30685
rect 12618 30648 12624 30660
rect 12268 30620 12624 30648
rect 12618 30608 12624 30620
rect 12676 30608 12682 30660
rect 13357 30651 13415 30657
rect 13357 30617 13369 30651
rect 13403 30648 13415 30651
rect 14277 30651 14335 30657
rect 14277 30648 14289 30651
rect 13403 30620 14289 30648
rect 13403 30617 13415 30620
rect 13357 30611 13415 30617
rect 14277 30617 14289 30620
rect 14323 30617 14335 30651
rect 15930 30648 15936 30660
rect 15891 30620 15936 30648
rect 14277 30611 14335 30617
rect 15930 30608 15936 30620
rect 15988 30608 15994 30660
rect 16393 30651 16451 30657
rect 16393 30617 16405 30651
rect 16439 30648 16451 30651
rect 17402 30648 17408 30660
rect 16439 30620 17408 30648
rect 16439 30617 16451 30620
rect 16393 30611 16451 30617
rect 17402 30608 17408 30620
rect 17460 30608 17466 30660
rect 19426 30608 19432 30660
rect 19484 30648 19490 30660
rect 19904 30648 19932 30679
rect 20346 30676 20352 30688
rect 20404 30716 20410 30728
rect 21361 30719 21419 30725
rect 20404 30688 20668 30716
rect 20404 30676 20410 30688
rect 20530 30648 20536 30660
rect 19484 30620 19932 30648
rect 20491 30620 20536 30648
rect 19484 30608 19490 30620
rect 20530 30608 20536 30620
rect 20588 30608 20594 30660
rect 20640 30648 20668 30688
rect 21361 30685 21373 30719
rect 21407 30716 21419 30719
rect 22189 30719 22247 30725
rect 22189 30716 22201 30719
rect 21407 30688 22201 30716
rect 21407 30685 21419 30688
rect 21361 30679 21419 30685
rect 22189 30685 22201 30688
rect 22235 30716 22247 30719
rect 22646 30716 22652 30728
rect 22235 30688 22652 30716
rect 22235 30685 22247 30688
rect 22189 30679 22247 30685
rect 22646 30676 22652 30688
rect 22704 30676 22710 30728
rect 22738 30676 22744 30728
rect 22796 30716 22802 30728
rect 23293 30719 23351 30725
rect 23293 30716 23305 30719
rect 22796 30688 23305 30716
rect 22796 30676 22802 30688
rect 23293 30685 23305 30688
rect 23339 30685 23351 30719
rect 23293 30679 23351 30685
rect 23658 30676 23664 30728
rect 23716 30676 23722 30728
rect 26329 30719 26387 30725
rect 26329 30685 26341 30719
rect 26375 30716 26387 30719
rect 27062 30716 27068 30728
rect 26375 30688 27068 30716
rect 26375 30685 26387 30688
rect 26329 30679 26387 30685
rect 27062 30676 27068 30688
rect 27120 30716 27126 30728
rect 27522 30716 27528 30728
rect 27120 30688 27528 30716
rect 27120 30676 27126 30688
rect 27522 30676 27528 30688
rect 27580 30676 27586 30728
rect 28166 30716 28172 30728
rect 28127 30688 28172 30716
rect 28166 30676 28172 30688
rect 28224 30676 28230 30728
rect 28368 30725 28396 30756
rect 30834 30744 30840 30796
rect 30892 30784 30898 30796
rect 33413 30787 33471 30793
rect 33413 30784 33425 30787
rect 30892 30756 33425 30784
rect 30892 30744 30898 30756
rect 33413 30753 33425 30756
rect 33459 30753 33471 30787
rect 33413 30747 33471 30753
rect 28353 30719 28411 30725
rect 28353 30685 28365 30719
rect 28399 30685 28411 30719
rect 29730 30716 29736 30728
rect 29691 30688 29736 30716
rect 28353 30679 28411 30685
rect 29730 30676 29736 30688
rect 29788 30676 29794 30728
rect 29822 30676 29828 30728
rect 29880 30716 29886 30728
rect 29989 30719 30047 30725
rect 29989 30716 30001 30719
rect 29880 30688 30001 30716
rect 29880 30676 29886 30688
rect 29989 30685 30001 30688
rect 30035 30685 30047 30719
rect 29989 30679 30047 30685
rect 31938 30676 31944 30728
rect 31996 30716 32002 30728
rect 32217 30719 32275 30725
rect 32217 30716 32229 30719
rect 31996 30688 32229 30716
rect 31996 30676 32002 30688
rect 32217 30685 32229 30688
rect 32263 30685 32275 30719
rect 32217 30679 32275 30685
rect 33226 30676 33232 30728
rect 33284 30716 33290 30728
rect 33321 30719 33379 30725
rect 33321 30716 33333 30719
rect 33284 30688 33333 30716
rect 33284 30676 33290 30688
rect 33321 30685 33333 30688
rect 33367 30685 33379 30719
rect 33321 30679 33379 30685
rect 20714 30648 20720 30660
rect 20640 30620 20720 30648
rect 20714 30608 20720 30620
rect 20772 30608 20778 30660
rect 20806 30608 20812 30660
rect 20864 30648 20870 30660
rect 21266 30648 21272 30660
rect 20864 30620 21272 30648
rect 20864 30608 20870 30620
rect 21266 30608 21272 30620
rect 21324 30608 21330 30660
rect 21542 30648 21548 30660
rect 21503 30620 21548 30648
rect 21542 30608 21548 30620
rect 21600 30608 21606 30660
rect 22373 30651 22431 30657
rect 22373 30617 22385 30651
rect 22419 30648 22431 30651
rect 25038 30648 25044 30660
rect 22419 30620 25044 30648
rect 22419 30617 22431 30620
rect 22373 30611 22431 30617
rect 25038 30608 25044 30620
rect 25096 30608 25102 30660
rect 25774 30608 25780 30660
rect 25832 30648 25838 30660
rect 26574 30651 26632 30657
rect 26574 30648 26586 30651
rect 25832 30620 26586 30648
rect 25832 30608 25838 30620
rect 26574 30617 26586 30620
rect 26620 30617 26632 30651
rect 26574 30611 26632 30617
rect 32033 30651 32091 30657
rect 32033 30617 32045 30651
rect 32079 30617 32091 30651
rect 32033 30611 32091 30617
rect 32401 30651 32459 30657
rect 32401 30617 32413 30651
rect 32447 30648 32459 30651
rect 32950 30648 32956 30660
rect 32447 30620 32956 30648
rect 32447 30617 32459 30620
rect 32401 30611 32459 30617
rect 12434 30580 12440 30592
rect 10928 30552 12440 30580
rect 10928 30540 10934 30552
rect 12434 30540 12440 30552
rect 12492 30540 12498 30592
rect 16577 30583 16635 30589
rect 16577 30549 16589 30583
rect 16623 30580 16635 30583
rect 17586 30580 17592 30592
rect 16623 30552 17592 30580
rect 16623 30549 16635 30552
rect 16577 30543 16635 30549
rect 17586 30540 17592 30552
rect 17644 30540 17650 30592
rect 19245 30583 19303 30589
rect 19245 30549 19257 30583
rect 19291 30580 19303 30583
rect 19334 30580 19340 30592
rect 19291 30552 19340 30580
rect 19291 30549 19303 30552
rect 19245 30543 19303 30549
rect 19334 30540 19340 30552
rect 19392 30540 19398 30592
rect 20070 30540 20076 30592
rect 20128 30580 20134 30592
rect 23566 30580 23572 30592
rect 20128 30552 23572 30580
rect 20128 30540 20134 30552
rect 23566 30540 23572 30552
rect 23624 30540 23630 30592
rect 27154 30540 27160 30592
rect 27212 30580 27218 30592
rect 27430 30580 27436 30592
rect 27212 30552 27436 30580
rect 27212 30540 27218 30552
rect 27430 30540 27436 30552
rect 27488 30580 27494 30592
rect 27709 30583 27767 30589
rect 27709 30580 27721 30583
rect 27488 30552 27721 30580
rect 27488 30540 27494 30552
rect 27709 30549 27721 30552
rect 27755 30549 27767 30583
rect 27709 30543 27767 30549
rect 30006 30540 30012 30592
rect 30064 30580 30070 30592
rect 31113 30583 31171 30589
rect 31113 30580 31125 30583
rect 30064 30552 31125 30580
rect 30064 30540 30070 30552
rect 31113 30549 31125 30552
rect 31159 30549 31171 30583
rect 32048 30580 32076 30611
rect 32950 30608 32956 30620
rect 33008 30608 33014 30660
rect 33134 30580 33140 30592
rect 32048 30552 33140 30580
rect 31113 30543 31171 30549
rect 33134 30540 33140 30552
rect 33192 30540 33198 30592
rect 33229 30583 33287 30589
rect 33229 30549 33241 30583
rect 33275 30580 33287 30583
rect 33410 30580 33416 30592
rect 33275 30552 33416 30580
rect 33275 30549 33287 30552
rect 33229 30543 33287 30549
rect 33410 30540 33416 30552
rect 33468 30540 33474 30592
rect 1104 30490 48852 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 48852 30490
rect 1104 30416 48852 30438
rect 15930 30336 15936 30388
rect 15988 30376 15994 30388
rect 15988 30348 27476 30376
rect 15988 30336 15994 30348
rect 9674 30268 9680 30320
rect 9732 30308 9738 30320
rect 10413 30311 10471 30317
rect 10413 30308 10425 30311
rect 9732 30280 10425 30308
rect 9732 30268 9738 30280
rect 10413 30277 10425 30280
rect 10459 30308 10471 30311
rect 12250 30308 12256 30320
rect 10459 30280 12256 30308
rect 10459 30277 10471 30280
rect 10413 30271 10471 30277
rect 12250 30268 12256 30280
rect 12308 30268 12314 30320
rect 17126 30268 17132 30320
rect 17184 30308 17190 30320
rect 17865 30311 17923 30317
rect 17865 30308 17877 30311
rect 17184 30280 17877 30308
rect 17184 30268 17190 30280
rect 17865 30277 17877 30280
rect 17911 30277 17923 30311
rect 18414 30308 18420 30320
rect 18375 30280 18420 30308
rect 17865 30271 17923 30277
rect 18414 30268 18420 30280
rect 18472 30268 18478 30320
rect 19334 30317 19340 30320
rect 19328 30271 19340 30317
rect 19392 30308 19398 30320
rect 19392 30280 19428 30308
rect 19334 30268 19340 30271
rect 19392 30268 19398 30280
rect 23106 30268 23112 30320
rect 23164 30308 23170 30320
rect 23385 30311 23443 30317
rect 23385 30308 23397 30311
rect 23164 30280 23397 30308
rect 23164 30268 23170 30280
rect 23385 30277 23397 30280
rect 23431 30277 23443 30311
rect 27448 30308 27476 30348
rect 27522 30336 27528 30388
rect 27580 30376 27586 30388
rect 29549 30379 29607 30385
rect 29549 30376 29561 30379
rect 27580 30348 29561 30376
rect 27580 30336 27586 30348
rect 29549 30345 29561 30348
rect 29595 30376 29607 30379
rect 29730 30376 29736 30388
rect 29595 30348 29736 30376
rect 29595 30345 29607 30348
rect 29549 30339 29607 30345
rect 29730 30336 29736 30348
rect 29788 30336 29794 30388
rect 45462 30376 45468 30388
rect 29840 30348 45468 30376
rect 29454 30308 29460 30320
rect 27448 30280 27936 30308
rect 29415 30280 29460 30308
rect 23385 30271 23443 30277
rect 1762 30240 1768 30252
rect 1723 30212 1768 30240
rect 1762 30200 1768 30212
rect 1820 30200 1826 30252
rect 4798 30240 4804 30252
rect 4759 30212 4804 30240
rect 4798 30200 4804 30212
rect 4856 30200 4862 30252
rect 8748 30243 8806 30249
rect 8748 30209 8760 30243
rect 8794 30240 8806 30243
rect 10226 30240 10232 30252
rect 8794 30212 10232 30240
rect 8794 30209 8806 30212
rect 8748 30203 8806 30209
rect 10226 30200 10232 30212
rect 10284 30200 10290 30252
rect 10594 30240 10600 30252
rect 10555 30212 10600 30240
rect 10594 30200 10600 30212
rect 10652 30200 10658 30252
rect 10778 30200 10784 30252
rect 10836 30240 10842 30252
rect 16022 30240 16028 30252
rect 10836 30212 16028 30240
rect 10836 30200 10842 30212
rect 16022 30200 16028 30212
rect 16080 30240 16086 30252
rect 16298 30240 16304 30252
rect 16080 30212 16304 30240
rect 16080 30200 16086 30212
rect 16298 30200 16304 30212
rect 16356 30200 16362 30252
rect 17683 30243 17741 30249
rect 17683 30209 17695 30243
rect 17729 30209 17741 30243
rect 17683 30203 17741 30209
rect 1949 30175 2007 30181
rect 1949 30141 1961 30175
rect 1995 30172 2007 30175
rect 2130 30172 2136 30184
rect 1995 30144 2136 30172
rect 1995 30141 2007 30144
rect 1949 30135 2007 30141
rect 2130 30132 2136 30144
rect 2188 30132 2194 30184
rect 2774 30132 2780 30184
rect 2832 30172 2838 30184
rect 2832 30144 2877 30172
rect 2832 30132 2838 30144
rect 7742 30132 7748 30184
rect 7800 30172 7806 30184
rect 8478 30172 8484 30184
rect 7800 30144 8484 30172
rect 7800 30132 7806 30144
rect 8478 30132 8484 30144
rect 8536 30132 8542 30184
rect 17696 30172 17724 30203
rect 17770 30200 17776 30252
rect 17828 30240 17834 30252
rect 20993 30243 21051 30249
rect 17828 30212 20116 30240
rect 17828 30200 17834 30212
rect 19061 30175 19119 30181
rect 17696 30144 17954 30172
rect 4062 30064 4068 30116
rect 4120 30104 4126 30116
rect 4617 30107 4675 30113
rect 4617 30104 4629 30107
rect 4120 30076 4629 30104
rect 4120 30064 4126 30076
rect 4617 30073 4629 30076
rect 4663 30073 4675 30107
rect 4617 30067 4675 30073
rect 12434 30064 12440 30116
rect 12492 30104 12498 30116
rect 17770 30104 17776 30116
rect 12492 30076 17776 30104
rect 12492 30064 12498 30076
rect 17770 30064 17776 30076
rect 17828 30064 17834 30116
rect 17926 30104 17954 30144
rect 19061 30141 19073 30175
rect 19107 30141 19119 30175
rect 19061 30135 19119 30141
rect 18598 30104 18604 30116
rect 17926 30076 18604 30104
rect 18598 30064 18604 30076
rect 18656 30064 18662 30116
rect 9861 30039 9919 30045
rect 9861 30005 9873 30039
rect 9907 30036 9919 30039
rect 10594 30036 10600 30048
rect 9907 30008 10600 30036
rect 9907 30005 9919 30008
rect 9861 29999 9919 30005
rect 10594 29996 10600 30008
rect 10652 29996 10658 30048
rect 10686 29996 10692 30048
rect 10744 30036 10750 30048
rect 10781 30039 10839 30045
rect 10781 30036 10793 30039
rect 10744 30008 10793 30036
rect 10744 29996 10750 30008
rect 10781 30005 10793 30008
rect 10827 30005 10839 30039
rect 19076 30036 19104 30135
rect 20088 30104 20116 30212
rect 20993 30209 21005 30243
rect 21039 30240 21051 30243
rect 21358 30240 21364 30252
rect 21039 30212 21364 30240
rect 21039 30209 21051 30212
rect 20993 30203 21051 30209
rect 21358 30200 21364 30212
rect 21416 30200 21422 30252
rect 21821 30243 21879 30249
rect 21821 30209 21833 30243
rect 21867 30240 21879 30243
rect 23201 30243 23259 30249
rect 23201 30240 23213 30243
rect 21867 30212 23213 30240
rect 21867 30209 21879 30212
rect 21821 30203 21879 30209
rect 23201 30209 23213 30212
rect 23247 30240 23259 30243
rect 27338 30240 27344 30252
rect 23247 30212 27344 30240
rect 23247 30209 23259 30212
rect 23201 30203 23259 30209
rect 27338 30200 27344 30212
rect 27396 30200 27402 30252
rect 27614 30200 27620 30252
rect 27672 30240 27678 30252
rect 27781 30243 27839 30249
rect 27781 30240 27793 30243
rect 27672 30212 27793 30240
rect 27672 30200 27678 30212
rect 27781 30209 27793 30212
rect 27827 30209 27839 30243
rect 27908 30240 27936 30280
rect 29454 30268 29460 30280
rect 29512 30268 29518 30320
rect 29840 30240 29868 30348
rect 45462 30336 45468 30348
rect 45520 30336 45526 30388
rect 32493 30311 32551 30317
rect 32493 30277 32505 30311
rect 32539 30308 32551 30311
rect 33842 30311 33900 30317
rect 33842 30308 33854 30311
rect 32539 30280 33854 30308
rect 32539 30277 32551 30280
rect 32493 30271 32551 30277
rect 33842 30277 33854 30280
rect 33888 30277 33900 30311
rect 33842 30271 33900 30277
rect 27908 30212 29868 30240
rect 32769 30243 32827 30249
rect 27781 30203 27839 30209
rect 32769 30209 32781 30243
rect 32815 30209 32827 30243
rect 32769 30203 32827 30209
rect 32861 30243 32919 30249
rect 32861 30209 32873 30243
rect 32907 30209 32919 30243
rect 32861 30203 32919 30209
rect 21376 30172 21404 30200
rect 22097 30175 22155 30181
rect 22097 30172 22109 30175
rect 21376 30144 22109 30172
rect 22097 30141 22109 30144
rect 22143 30141 22155 30175
rect 27522 30172 27528 30184
rect 27483 30144 27528 30172
rect 22097 30135 22155 30141
rect 27522 30132 27528 30144
rect 27580 30132 27586 30184
rect 32784 30172 32812 30203
rect 31726 30144 32812 30172
rect 20441 30107 20499 30113
rect 20088 30076 20208 30104
rect 20070 30036 20076 30048
rect 19076 30008 20076 30036
rect 10781 29999 10839 30005
rect 20070 29996 20076 30008
rect 20128 29996 20134 30048
rect 20180 30036 20208 30076
rect 20441 30073 20453 30107
rect 20487 30104 20499 30107
rect 20530 30104 20536 30116
rect 20487 30076 20536 30104
rect 20487 30073 20499 30076
rect 20441 30067 20499 30073
rect 20530 30064 20536 30076
rect 20588 30104 20594 30116
rect 31726 30104 31754 30144
rect 32876 30116 32904 30203
rect 32950 30200 32956 30252
rect 33008 30240 33014 30252
rect 33137 30243 33195 30249
rect 33008 30212 33053 30240
rect 33008 30200 33014 30212
rect 33137 30209 33149 30243
rect 33183 30240 33195 30243
rect 33502 30240 33508 30252
rect 33183 30212 33508 30240
rect 33183 30209 33195 30212
rect 33137 30203 33195 30209
rect 33502 30200 33508 30212
rect 33560 30200 33566 30252
rect 47946 30240 47952 30252
rect 47907 30212 47952 30240
rect 47946 30200 47952 30212
rect 48004 30200 48010 30252
rect 33042 30132 33048 30184
rect 33100 30172 33106 30184
rect 33594 30172 33600 30184
rect 33100 30144 33600 30172
rect 33100 30132 33106 30144
rect 33594 30132 33600 30144
rect 33652 30132 33658 30184
rect 20588 30076 26924 30104
rect 20588 30064 20594 30076
rect 20622 30036 20628 30048
rect 20180 30008 20628 30036
rect 20622 29996 20628 30008
rect 20680 30036 20686 30048
rect 21177 30039 21235 30045
rect 21177 30036 21189 30039
rect 20680 30008 21189 30036
rect 20680 29996 20686 30008
rect 21177 30005 21189 30008
rect 21223 30005 21235 30039
rect 21177 29999 21235 30005
rect 22002 29996 22008 30048
rect 22060 30036 22066 30048
rect 25590 30036 25596 30048
rect 22060 30008 25596 30036
rect 22060 29996 22066 30008
rect 25590 29996 25596 30008
rect 25648 29996 25654 30048
rect 26896 30036 26924 30076
rect 28460 30076 31754 30104
rect 28460 30036 28488 30076
rect 32398 30064 32404 30116
rect 32456 30104 32462 30116
rect 32858 30104 32864 30116
rect 32456 30076 32864 30104
rect 32456 30064 32462 30076
rect 32858 30064 32864 30076
rect 32916 30064 32922 30116
rect 26896 30008 28488 30036
rect 28718 29996 28724 30048
rect 28776 30036 28782 30048
rect 28905 30039 28963 30045
rect 28905 30036 28917 30039
rect 28776 30008 28917 30036
rect 28776 29996 28782 30008
rect 28905 30005 28917 30008
rect 28951 30005 28963 30039
rect 28905 29999 28963 30005
rect 34606 29996 34612 30048
rect 34664 30036 34670 30048
rect 34977 30039 35035 30045
rect 34977 30036 34989 30039
rect 34664 30008 34989 30036
rect 34664 29996 34670 30008
rect 34977 30005 34989 30008
rect 35023 30005 35035 30039
rect 48038 30036 48044 30048
rect 47999 30008 48044 30036
rect 34977 29999 35035 30005
rect 48038 29996 48044 30008
rect 48096 29996 48102 30048
rect 1104 29946 48852 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 48852 29946
rect 1104 29872 48852 29894
rect 2130 29832 2136 29844
rect 2091 29804 2136 29832
rect 2130 29792 2136 29804
rect 2188 29792 2194 29844
rect 10226 29832 10232 29844
rect 10187 29804 10232 29832
rect 10226 29792 10232 29804
rect 10284 29792 10290 29844
rect 10502 29792 10508 29844
rect 10560 29832 10566 29844
rect 12253 29835 12311 29841
rect 12253 29832 12265 29835
rect 10560 29804 12265 29832
rect 10560 29792 10566 29804
rect 12253 29801 12265 29804
rect 12299 29801 12311 29835
rect 20346 29832 20352 29844
rect 12253 29795 12311 29801
rect 12406 29804 20352 29832
rect 2682 29724 2688 29776
rect 2740 29764 2746 29776
rect 12406 29764 12434 29804
rect 20346 29792 20352 29804
rect 20404 29792 20410 29844
rect 20898 29792 20904 29844
rect 20956 29832 20962 29844
rect 32398 29832 32404 29844
rect 20956 29804 32404 29832
rect 20956 29792 20962 29804
rect 32398 29792 32404 29804
rect 32456 29792 32462 29844
rect 33134 29792 33140 29844
rect 33192 29832 33198 29844
rect 33413 29835 33471 29841
rect 33413 29832 33425 29835
rect 33192 29804 33425 29832
rect 33192 29792 33198 29804
rect 33413 29801 33425 29804
rect 33459 29801 33471 29835
rect 33413 29795 33471 29801
rect 2740 29736 12434 29764
rect 2740 29724 2746 29736
rect 13722 29724 13728 29776
rect 13780 29764 13786 29776
rect 48038 29764 48044 29776
rect 13780 29736 22784 29764
rect 13780 29724 13786 29736
rect 10778 29696 10784 29708
rect 10612 29668 10784 29696
rect 1581 29631 1639 29637
rect 1581 29597 1593 29631
rect 1627 29628 1639 29631
rect 1762 29628 1768 29640
rect 1627 29600 1768 29628
rect 1627 29597 1639 29600
rect 1581 29591 1639 29597
rect 1762 29588 1768 29600
rect 1820 29588 1826 29640
rect 2041 29631 2099 29637
rect 2041 29597 2053 29631
rect 2087 29628 2099 29631
rect 2685 29631 2743 29637
rect 2685 29628 2697 29631
rect 2087 29600 2697 29628
rect 2087 29597 2099 29600
rect 2041 29591 2099 29597
rect 2685 29597 2697 29600
rect 2731 29628 2743 29631
rect 9122 29628 9128 29640
rect 2731 29600 7236 29628
rect 9083 29600 9128 29628
rect 2731 29597 2743 29600
rect 2685 29591 2743 29597
rect 7208 29560 7236 29600
rect 9122 29588 9128 29600
rect 9180 29588 9186 29640
rect 10502 29628 10508 29640
rect 10463 29600 10508 29628
rect 10502 29588 10508 29600
rect 10560 29588 10566 29640
rect 10612 29637 10640 29668
rect 10778 29656 10784 29668
rect 10836 29656 10842 29708
rect 12434 29656 12440 29708
rect 12492 29696 12498 29708
rect 16298 29696 16304 29708
rect 12492 29668 12537 29696
rect 16259 29668 16304 29696
rect 12492 29656 12498 29668
rect 16298 29656 16304 29668
rect 16356 29656 16362 29708
rect 17218 29656 17224 29708
rect 17276 29696 17282 29708
rect 22002 29696 22008 29708
rect 17276 29668 22008 29696
rect 17276 29656 17282 29668
rect 22002 29656 22008 29668
rect 22060 29656 22066 29708
rect 10597 29631 10655 29637
rect 10597 29597 10609 29631
rect 10643 29597 10655 29631
rect 10597 29591 10655 29597
rect 10686 29588 10692 29640
rect 10744 29628 10750 29640
rect 10744 29600 10789 29628
rect 10744 29588 10750 29600
rect 10870 29588 10876 29640
rect 10928 29628 10934 29640
rect 12529 29631 12587 29637
rect 10928 29600 10973 29628
rect 10928 29588 10934 29600
rect 12529 29597 12541 29631
rect 12575 29597 12587 29631
rect 14366 29628 14372 29640
rect 14327 29600 14372 29628
rect 12529 29591 12587 29597
rect 11698 29560 11704 29572
rect 7208 29532 11704 29560
rect 11698 29520 11704 29532
rect 11756 29520 11762 29572
rect 12250 29560 12256 29572
rect 12211 29532 12256 29560
rect 12250 29520 12256 29532
rect 12308 29520 12314 29572
rect 12544 29560 12572 29591
rect 14366 29588 14372 29600
rect 14424 29588 14430 29640
rect 14645 29631 14703 29637
rect 14645 29597 14657 29631
rect 14691 29628 14703 29631
rect 15378 29628 15384 29640
rect 14691 29600 15384 29628
rect 14691 29597 14703 29600
rect 14645 29591 14703 29597
rect 15378 29588 15384 29600
rect 15436 29588 15442 29640
rect 15841 29631 15899 29637
rect 15841 29597 15853 29631
rect 15887 29597 15899 29631
rect 15841 29591 15899 29597
rect 12406 29532 12572 29560
rect 14384 29560 14412 29588
rect 15856 29560 15884 29591
rect 16022 29588 16028 29640
rect 16080 29628 16086 29640
rect 16577 29631 16635 29637
rect 16577 29628 16589 29631
rect 16080 29600 16589 29628
rect 16080 29588 16086 29600
rect 16577 29597 16589 29600
rect 16623 29628 16635 29631
rect 17770 29628 17776 29640
rect 16623 29600 17776 29628
rect 16623 29597 16635 29600
rect 16577 29591 16635 29597
rect 17770 29588 17776 29600
rect 17828 29588 17834 29640
rect 18598 29588 18604 29640
rect 18656 29628 18662 29640
rect 20073 29631 20131 29637
rect 20073 29628 20085 29631
rect 18656 29600 20085 29628
rect 18656 29588 18662 29600
rect 20073 29597 20085 29600
rect 20119 29597 20131 29631
rect 20714 29628 20720 29640
rect 20675 29600 20720 29628
rect 20073 29591 20131 29597
rect 20714 29588 20720 29600
rect 20772 29588 20778 29640
rect 20898 29628 20904 29640
rect 20859 29600 20904 29628
rect 20898 29588 20904 29600
rect 20956 29588 20962 29640
rect 14384 29532 15884 29560
rect 17957 29563 18015 29569
rect 1946 29452 1952 29504
rect 2004 29492 2010 29504
rect 2777 29495 2835 29501
rect 2777 29492 2789 29495
rect 2004 29464 2789 29492
rect 2004 29452 2010 29464
rect 2777 29461 2789 29464
rect 2823 29461 2835 29495
rect 8938 29492 8944 29504
rect 8899 29464 8944 29492
rect 2777 29455 2835 29461
rect 8938 29452 8944 29464
rect 8996 29452 9002 29504
rect 10226 29452 10232 29504
rect 10284 29492 10290 29504
rect 10410 29492 10416 29504
rect 10284 29464 10416 29492
rect 10284 29452 10290 29464
rect 10410 29452 10416 29464
rect 10468 29492 10474 29504
rect 12406 29492 12434 29532
rect 17957 29529 17969 29563
rect 18003 29529 18015 29563
rect 17957 29523 18015 29529
rect 18141 29563 18199 29569
rect 18141 29529 18153 29563
rect 18187 29560 18199 29563
rect 19334 29560 19340 29572
rect 18187 29532 19340 29560
rect 18187 29529 18199 29532
rect 18141 29523 18199 29529
rect 10468 29464 12434 29492
rect 12713 29495 12771 29501
rect 10468 29452 10474 29464
rect 12713 29461 12725 29495
rect 12759 29492 12771 29495
rect 13630 29492 13636 29504
rect 12759 29464 13636 29492
rect 12759 29461 12771 29464
rect 12713 29455 12771 29461
rect 13630 29452 13636 29464
rect 13688 29452 13694 29504
rect 14185 29495 14243 29501
rect 14185 29461 14197 29495
rect 14231 29492 14243 29495
rect 14366 29492 14372 29504
rect 14231 29464 14372 29492
rect 14231 29461 14243 29464
rect 14185 29455 14243 29461
rect 14366 29452 14372 29464
rect 14424 29452 14430 29504
rect 14550 29492 14556 29504
rect 14511 29464 14556 29492
rect 14550 29452 14556 29464
rect 14608 29452 14614 29504
rect 15657 29495 15715 29501
rect 15657 29461 15669 29495
rect 15703 29492 15715 29495
rect 16758 29492 16764 29504
rect 15703 29464 16764 29492
rect 15703 29461 15715 29464
rect 15657 29455 15715 29461
rect 16758 29452 16764 29464
rect 16816 29492 16822 29504
rect 17972 29492 18000 29523
rect 19334 29520 19340 29532
rect 19392 29520 19398 29572
rect 20732 29560 20760 29588
rect 22756 29560 22784 29736
rect 24688 29736 48044 29764
rect 23017 29699 23075 29705
rect 23017 29665 23029 29699
rect 23063 29696 23075 29699
rect 23106 29696 23112 29708
rect 23063 29668 23112 29696
rect 23063 29665 23075 29668
rect 23017 29659 23075 29665
rect 23106 29656 23112 29668
rect 23164 29656 23170 29708
rect 23293 29631 23351 29637
rect 23293 29597 23305 29631
rect 23339 29628 23351 29631
rect 23474 29628 23480 29640
rect 23339 29600 23480 29628
rect 23339 29597 23351 29600
rect 23293 29591 23351 29597
rect 23474 29588 23480 29600
rect 23532 29588 23538 29640
rect 24688 29637 24716 29736
rect 48038 29724 48044 29736
rect 48096 29724 48102 29776
rect 24946 29696 24952 29708
rect 24780 29668 24952 29696
rect 24780 29637 24808 29668
rect 24946 29656 24952 29668
rect 25004 29656 25010 29708
rect 27246 29656 27252 29708
rect 27304 29696 27310 29708
rect 27525 29699 27583 29705
rect 27525 29696 27537 29699
rect 27304 29668 27537 29696
rect 27304 29656 27310 29668
rect 27525 29665 27537 29668
rect 27571 29665 27583 29699
rect 27525 29659 27583 29665
rect 32674 29656 32680 29708
rect 32732 29696 32738 29708
rect 32732 29668 32904 29696
rect 32732 29656 32738 29668
rect 24673 29631 24731 29637
rect 24673 29597 24685 29631
rect 24719 29597 24731 29631
rect 24673 29591 24731 29597
rect 24765 29631 24823 29637
rect 24765 29597 24777 29631
rect 24811 29597 24823 29631
rect 24765 29591 24823 29597
rect 24854 29588 24860 29640
rect 24912 29628 24918 29640
rect 25041 29631 25099 29637
rect 24912 29600 24957 29628
rect 24912 29588 24918 29600
rect 25041 29597 25053 29631
rect 25087 29628 25099 29631
rect 25130 29628 25136 29640
rect 25087 29600 25136 29628
rect 25087 29597 25099 29600
rect 25041 29591 25099 29597
rect 25130 29588 25136 29600
rect 25188 29588 25194 29640
rect 25590 29628 25596 29640
rect 25551 29600 25596 29628
rect 25590 29588 25596 29600
rect 25648 29588 25654 29640
rect 27801 29631 27859 29637
rect 27801 29597 27813 29631
rect 27847 29628 27859 29631
rect 28166 29628 28172 29640
rect 27847 29600 28172 29628
rect 27847 29597 27859 29600
rect 27801 29591 27859 29597
rect 28166 29588 28172 29600
rect 28224 29628 28230 29640
rect 28902 29628 28908 29640
rect 28224 29600 28908 29628
rect 28224 29588 28230 29600
rect 28902 29588 28908 29600
rect 28960 29628 28966 29640
rect 31389 29631 31447 29637
rect 31389 29628 31401 29631
rect 28960 29600 31401 29628
rect 28960 29588 28966 29600
rect 31389 29597 31401 29600
rect 31435 29628 31447 29631
rect 32769 29631 32827 29637
rect 32769 29628 32781 29631
rect 31435 29600 32781 29628
rect 31435 29597 31447 29600
rect 31389 29591 31447 29597
rect 32769 29597 32781 29600
rect 32815 29597 32827 29631
rect 32876 29628 32904 29668
rect 33778 29656 33784 29708
rect 33836 29696 33842 29708
rect 33873 29699 33931 29705
rect 33873 29696 33885 29699
rect 33836 29668 33885 29696
rect 33836 29656 33842 29668
rect 33873 29665 33885 29668
rect 33919 29665 33931 29699
rect 33873 29659 33931 29665
rect 33962 29656 33968 29708
rect 34020 29696 34026 29708
rect 38010 29696 38016 29708
rect 34020 29668 34065 29696
rect 37971 29668 38016 29696
rect 34020 29656 34026 29668
rect 38010 29656 38016 29668
rect 38068 29656 38074 29708
rect 36173 29631 36231 29637
rect 36173 29628 36185 29631
rect 32876 29600 36185 29628
rect 32769 29591 32827 29597
rect 36173 29597 36185 29600
rect 36219 29597 36231 29631
rect 36173 29591 36231 29597
rect 28350 29560 28356 29572
rect 20732 29532 22094 29560
rect 22756 29532 28356 29560
rect 18322 29492 18328 29504
rect 16816 29464 18000 29492
rect 18283 29464 18328 29492
rect 16816 29452 16822 29464
rect 18322 29452 18328 29464
rect 18380 29452 18386 29504
rect 20070 29452 20076 29504
rect 20128 29492 20134 29504
rect 20165 29495 20223 29501
rect 20165 29492 20177 29495
rect 20128 29464 20177 29492
rect 20128 29452 20134 29464
rect 20165 29461 20177 29464
rect 20211 29461 20223 29495
rect 20165 29455 20223 29461
rect 20806 29452 20812 29504
rect 20864 29492 20870 29504
rect 21085 29495 21143 29501
rect 21085 29492 21097 29495
rect 20864 29464 21097 29492
rect 20864 29452 20870 29464
rect 21085 29461 21097 29464
rect 21131 29461 21143 29495
rect 22066 29492 22094 29532
rect 28350 29520 28356 29532
rect 28408 29520 28414 29572
rect 31202 29560 31208 29572
rect 31163 29532 31208 29560
rect 31202 29520 31208 29532
rect 31260 29520 31266 29572
rect 32585 29563 32643 29569
rect 32585 29529 32597 29563
rect 32631 29560 32643 29563
rect 33318 29560 33324 29572
rect 32631 29532 33324 29560
rect 32631 29529 32643 29532
rect 32585 29523 32643 29529
rect 33318 29520 33324 29532
rect 33376 29520 33382 29572
rect 36357 29563 36415 29569
rect 36357 29529 36369 29563
rect 36403 29560 36415 29563
rect 36446 29560 36452 29572
rect 36403 29532 36452 29560
rect 36403 29529 36415 29532
rect 36357 29523 36415 29529
rect 36446 29520 36452 29532
rect 36504 29520 36510 29572
rect 22922 29492 22928 29504
rect 22066 29464 22928 29492
rect 21085 29455 21143 29461
rect 22922 29452 22928 29464
rect 22980 29452 22986 29504
rect 24394 29492 24400 29504
rect 24355 29464 24400 29492
rect 24394 29452 24400 29464
rect 24452 29452 24458 29504
rect 24578 29452 24584 29504
rect 24636 29492 24642 29504
rect 24762 29492 24768 29504
rect 24636 29464 24768 29492
rect 24636 29452 24642 29464
rect 24762 29452 24768 29464
rect 24820 29452 24826 29504
rect 25038 29452 25044 29504
rect 25096 29492 25102 29504
rect 25685 29495 25743 29501
rect 25685 29492 25697 29495
rect 25096 29464 25697 29492
rect 25096 29452 25102 29464
rect 25685 29461 25697 29464
rect 25731 29461 25743 29495
rect 25685 29455 25743 29461
rect 31478 29452 31484 29504
rect 31536 29492 31542 29504
rect 31573 29495 31631 29501
rect 31573 29492 31585 29495
rect 31536 29464 31585 29492
rect 31536 29452 31542 29464
rect 31573 29461 31585 29464
rect 31619 29461 31631 29495
rect 31573 29455 31631 29461
rect 32953 29495 33011 29501
rect 32953 29461 32965 29495
rect 32999 29492 33011 29495
rect 33042 29492 33048 29504
rect 32999 29464 33048 29492
rect 32999 29461 33011 29464
rect 32953 29455 33011 29461
rect 33042 29452 33048 29464
rect 33100 29452 33106 29504
rect 33781 29495 33839 29501
rect 33781 29461 33793 29495
rect 33827 29492 33839 29495
rect 34606 29492 34612 29504
rect 33827 29464 34612 29492
rect 33827 29461 33839 29464
rect 33781 29455 33839 29461
rect 34606 29452 34612 29464
rect 34664 29452 34670 29504
rect 1104 29402 48852 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 48852 29402
rect 1104 29328 48852 29350
rect 9217 29291 9275 29297
rect 9217 29257 9229 29291
rect 9263 29288 9275 29291
rect 10226 29288 10232 29300
rect 9263 29260 10232 29288
rect 9263 29257 9275 29260
rect 9217 29251 9275 29257
rect 1946 29220 1952 29232
rect 1907 29192 1952 29220
rect 1946 29180 1952 29192
rect 2004 29180 2010 29232
rect 8104 29223 8162 29229
rect 8104 29189 8116 29223
rect 8150 29220 8162 29223
rect 8938 29220 8944 29232
rect 8150 29192 8944 29220
rect 8150 29189 8162 29192
rect 8104 29183 8162 29189
rect 8938 29180 8944 29192
rect 8996 29180 9002 29232
rect 9692 29229 9720 29260
rect 10226 29248 10232 29260
rect 10284 29248 10290 29300
rect 13722 29288 13728 29300
rect 13683 29260 13728 29288
rect 13722 29248 13728 29260
rect 13780 29248 13786 29300
rect 18049 29291 18107 29297
rect 18049 29257 18061 29291
rect 18095 29288 18107 29291
rect 18138 29288 18144 29300
rect 18095 29260 18144 29288
rect 18095 29257 18107 29260
rect 18049 29251 18107 29257
rect 18138 29248 18144 29260
rect 18196 29248 18202 29300
rect 19334 29248 19340 29300
rect 19392 29288 19398 29300
rect 19889 29291 19947 29297
rect 19889 29288 19901 29291
rect 19392 29260 19901 29288
rect 19392 29248 19398 29260
rect 19889 29257 19901 29260
rect 19935 29257 19947 29291
rect 19889 29251 19947 29257
rect 24029 29291 24087 29297
rect 24029 29257 24041 29291
rect 24075 29288 24087 29291
rect 24854 29288 24860 29300
rect 24075 29260 24860 29288
rect 24075 29257 24087 29260
rect 24029 29251 24087 29257
rect 24854 29248 24860 29260
rect 24912 29248 24918 29300
rect 25869 29291 25927 29297
rect 25869 29257 25881 29291
rect 25915 29288 25927 29291
rect 25915 29260 28212 29288
rect 25915 29257 25927 29260
rect 25869 29251 25927 29257
rect 9677 29223 9735 29229
rect 9677 29189 9689 29223
rect 9723 29189 9735 29223
rect 9677 29183 9735 29189
rect 9858 29180 9864 29232
rect 9916 29229 9922 29232
rect 9916 29223 9935 29229
rect 9923 29189 9935 29223
rect 15470 29220 15476 29232
rect 15431 29192 15476 29220
rect 9916 29183 9935 29189
rect 9916 29180 9922 29183
rect 15470 29180 15476 29192
rect 15528 29180 15534 29232
rect 16574 29220 16580 29232
rect 15948 29192 16580 29220
rect 1762 29152 1768 29164
rect 1723 29124 1768 29152
rect 1762 29112 1768 29124
rect 1820 29112 1826 29164
rect 4062 29112 4068 29164
rect 4120 29152 4126 29164
rect 11514 29152 11520 29164
rect 4120 29124 9720 29152
rect 11475 29124 11520 29152
rect 4120 29112 4126 29124
rect 9692 29096 9720 29124
rect 11514 29112 11520 29124
rect 11572 29112 11578 29164
rect 11606 29112 11612 29164
rect 11664 29152 11670 29164
rect 11773 29155 11831 29161
rect 11773 29152 11785 29155
rect 11664 29124 11785 29152
rect 11664 29112 11670 29124
rect 11773 29121 11785 29124
rect 11819 29121 11831 29155
rect 11773 29115 11831 29121
rect 12894 29112 12900 29164
rect 12952 29152 12958 29164
rect 13449 29155 13507 29161
rect 13449 29152 13461 29155
rect 12952 29124 13461 29152
rect 12952 29112 12958 29124
rect 13449 29121 13461 29124
rect 13495 29121 13507 29155
rect 13630 29152 13636 29164
rect 13591 29124 13636 29152
rect 13449 29115 13507 29121
rect 13630 29112 13636 29124
rect 13688 29112 13694 29164
rect 14366 29152 14372 29164
rect 14327 29124 14372 29152
rect 14366 29112 14372 29124
rect 14424 29112 14430 29164
rect 15746 29152 15752 29164
rect 15707 29124 15752 29152
rect 15746 29112 15752 29124
rect 15804 29112 15810 29164
rect 15948 29161 15976 29192
rect 16574 29180 16580 29192
rect 16632 29180 16638 29232
rect 20070 29220 20076 29232
rect 16684 29192 20076 29220
rect 16684 29161 16712 29192
rect 16942 29161 16948 29164
rect 15841 29155 15899 29161
rect 15841 29121 15853 29155
rect 15887 29121 15899 29155
rect 15841 29115 15899 29121
rect 15933 29155 15991 29161
rect 15933 29121 15945 29155
rect 15979 29121 15991 29155
rect 15933 29115 15991 29121
rect 16117 29155 16175 29161
rect 16117 29121 16129 29155
rect 16163 29121 16175 29155
rect 16117 29115 16175 29121
rect 16669 29155 16727 29161
rect 16669 29121 16681 29155
rect 16715 29121 16727 29155
rect 16936 29152 16948 29161
rect 16903 29124 16948 29152
rect 16669 29115 16727 29121
rect 16936 29115 16948 29124
rect 3326 29084 3332 29096
rect 3287 29056 3332 29084
rect 3326 29044 3332 29056
rect 3384 29044 3390 29096
rect 7742 29044 7748 29096
rect 7800 29084 7806 29096
rect 7837 29087 7895 29093
rect 7837 29084 7849 29087
rect 7800 29056 7849 29084
rect 7800 29044 7806 29056
rect 7837 29053 7849 29056
rect 7883 29053 7895 29087
rect 7837 29047 7895 29053
rect 9674 29044 9680 29096
rect 9732 29044 9738 29096
rect 15856 29084 15884 29115
rect 16022 29084 16028 29096
rect 15856 29056 16028 29084
rect 16022 29044 16028 29056
rect 16080 29044 16086 29096
rect 8846 28976 8852 29028
rect 8904 29016 8910 29028
rect 10045 29019 10103 29025
rect 10045 29016 10057 29019
rect 8904 28988 10057 29016
rect 8904 28976 8910 28988
rect 10045 28985 10057 28988
rect 10091 28985 10103 29019
rect 10045 28979 10103 28985
rect 1394 28908 1400 28960
rect 1452 28948 1458 28960
rect 4249 28951 4307 28957
rect 4249 28948 4261 28951
rect 1452 28920 4261 28948
rect 1452 28908 1458 28920
rect 4249 28917 4261 28920
rect 4295 28917 4307 28951
rect 4249 28911 4307 28917
rect 9766 28908 9772 28960
rect 9824 28948 9830 28960
rect 9861 28951 9919 28957
rect 9861 28948 9873 28951
rect 9824 28920 9873 28948
rect 9824 28908 9830 28920
rect 9861 28917 9873 28920
rect 9907 28948 9919 28951
rect 10502 28948 10508 28960
rect 9907 28920 10508 28948
rect 9907 28917 9919 28920
rect 9861 28911 9919 28917
rect 10502 28908 10508 28920
rect 10560 28908 10566 28960
rect 12526 28908 12532 28960
rect 12584 28948 12590 28960
rect 12897 28951 12955 28957
rect 12897 28948 12909 28951
rect 12584 28920 12909 28948
rect 12584 28908 12590 28920
rect 12897 28917 12909 28920
rect 12943 28917 12955 28951
rect 12897 28911 12955 28917
rect 13354 28908 13360 28960
rect 13412 28948 13418 28960
rect 14461 28951 14519 28957
rect 14461 28948 14473 28951
rect 13412 28920 14473 28948
rect 13412 28908 13418 28920
rect 14461 28917 14473 28920
rect 14507 28917 14519 28951
rect 14461 28911 14519 28917
rect 15654 28908 15660 28960
rect 15712 28948 15718 28960
rect 16022 28948 16028 28960
rect 15712 28920 16028 28948
rect 15712 28908 15718 28920
rect 16022 28908 16028 28920
rect 16080 28908 16086 28960
rect 16132 28948 16160 29115
rect 16942 29112 16948 29115
rect 17000 29112 17006 29164
rect 18524 29161 18552 29192
rect 20070 29180 20076 29192
rect 20128 29180 20134 29232
rect 24394 29180 24400 29232
rect 24452 29220 24458 29232
rect 24734 29223 24792 29229
rect 24734 29220 24746 29223
rect 24452 29192 24746 29220
rect 24452 29180 24458 29192
rect 24734 29189 24746 29192
rect 24780 29189 24792 29223
rect 24734 29183 24792 29189
rect 18509 29155 18567 29161
rect 18509 29121 18521 29155
rect 18555 29121 18567 29155
rect 18509 29115 18567 29121
rect 18598 29112 18604 29164
rect 18656 29152 18662 29164
rect 18765 29155 18823 29161
rect 18765 29152 18777 29155
rect 18656 29124 18777 29152
rect 18656 29112 18662 29124
rect 18765 29121 18777 29124
rect 18811 29121 18823 29155
rect 18765 29115 18823 29121
rect 20346 29112 20352 29164
rect 20404 29152 20410 29164
rect 20579 29155 20637 29161
rect 20579 29152 20591 29155
rect 20404 29124 20591 29152
rect 20404 29112 20410 29124
rect 20579 29121 20591 29124
rect 20625 29121 20637 29155
rect 20579 29115 20637 29121
rect 20717 29155 20775 29161
rect 20717 29121 20729 29155
rect 20763 29121 20775 29155
rect 20717 29115 20775 29121
rect 20732 29084 20760 29115
rect 20806 29112 20812 29164
rect 20864 29152 20870 29164
rect 20864 29124 20909 29152
rect 20864 29112 20870 29124
rect 20990 29112 20996 29164
rect 21048 29152 21054 29164
rect 21048 29124 21093 29152
rect 21048 29112 21054 29124
rect 22002 29112 22008 29164
rect 22060 29161 22066 29164
rect 22060 29155 22109 29161
rect 22183 29155 22189 29167
rect 22060 29121 22063 29155
rect 22097 29121 22109 29155
rect 22144 29127 22189 29155
rect 22060 29115 22109 29121
rect 22183 29115 22189 29127
rect 22241 29115 22247 29167
rect 22060 29112 22066 29115
rect 22278 29112 22284 29164
rect 22336 29161 22342 29164
rect 22336 29152 22344 29161
rect 22465 29155 22523 29161
rect 22336 29124 22381 29152
rect 22336 29115 22344 29124
rect 22465 29121 22477 29155
rect 22511 29152 22523 29155
rect 22554 29152 22560 29164
rect 22511 29124 22560 29152
rect 22511 29121 22523 29124
rect 22465 29115 22523 29121
rect 22336 29112 22342 29115
rect 22554 29112 22560 29124
rect 22612 29112 22618 29164
rect 22922 29112 22928 29164
rect 22980 29152 22986 29164
rect 23661 29155 23719 29161
rect 23661 29152 23673 29155
rect 22980 29124 23673 29152
rect 22980 29112 22986 29124
rect 23661 29121 23673 29124
rect 23707 29121 23719 29155
rect 23661 29115 23719 29121
rect 23845 29155 23903 29161
rect 23845 29121 23857 29155
rect 23891 29152 23903 29155
rect 25884 29152 25912 29251
rect 27525 29223 27583 29229
rect 27525 29189 27537 29223
rect 27571 29220 27583 29223
rect 27614 29220 27620 29232
rect 27571 29192 27620 29220
rect 27571 29189 27583 29192
rect 27525 29183 27583 29189
rect 27614 29180 27620 29192
rect 27672 29220 27678 29232
rect 28074 29220 28080 29232
rect 27672 29192 28080 29220
rect 27672 29180 27678 29192
rect 28074 29180 28080 29192
rect 28132 29180 28138 29232
rect 28184 29220 28212 29260
rect 28350 29248 28356 29300
rect 28408 29288 28414 29300
rect 32674 29288 32680 29300
rect 28408 29260 32680 29288
rect 28408 29248 28414 29260
rect 32674 29248 32680 29260
rect 32732 29248 32738 29300
rect 36446 29288 36452 29300
rect 36407 29260 36452 29288
rect 36446 29248 36452 29260
rect 36504 29248 36510 29300
rect 47302 29248 47308 29300
rect 47360 29288 47366 29300
rect 47486 29288 47492 29300
rect 47360 29260 47492 29288
rect 47360 29248 47366 29260
rect 47486 29248 47492 29260
rect 47544 29248 47550 29300
rect 28184 29192 28488 29220
rect 27338 29152 27344 29164
rect 23891 29124 25912 29152
rect 27299 29124 27344 29152
rect 23891 29121 23903 29124
rect 23845 29115 23903 29121
rect 27338 29112 27344 29124
rect 27396 29112 27402 29164
rect 27982 29152 27988 29164
rect 27943 29124 27988 29152
rect 27982 29112 27988 29124
rect 28040 29112 28046 29164
rect 28167 29155 28225 29161
rect 28167 29121 28179 29155
rect 28213 29121 28225 29155
rect 28460 29152 28488 29192
rect 30190 29180 30196 29232
rect 30248 29220 30254 29232
rect 32490 29220 32496 29232
rect 30248 29192 31248 29220
rect 32451 29192 32496 29220
rect 30248 29180 30254 29192
rect 31220 29161 31248 29192
rect 32490 29180 32496 29192
rect 32548 29180 32554 29232
rect 33042 29180 33048 29232
rect 33100 29180 33106 29232
rect 31021 29155 31079 29161
rect 31021 29152 31033 29155
rect 28460 29124 31033 29152
rect 28167 29115 28225 29121
rect 31021 29121 31033 29124
rect 31067 29121 31079 29155
rect 31021 29115 31079 29121
rect 31113 29155 31171 29161
rect 31113 29121 31125 29155
rect 31159 29121 31171 29155
rect 31113 29115 31171 29121
rect 31205 29155 31263 29161
rect 31205 29121 31217 29155
rect 31251 29121 31263 29155
rect 31205 29115 31263 29121
rect 31389 29155 31447 29161
rect 31389 29121 31401 29155
rect 31435 29152 31447 29155
rect 31754 29152 31760 29164
rect 31435 29124 31760 29152
rect 31435 29121 31447 29124
rect 31389 29115 31447 29121
rect 24486 29084 24492 29096
rect 20732 29056 21306 29084
rect 24447 29056 24492 29084
rect 21174 29016 21180 29028
rect 19444 28988 21180 29016
rect 17310 28948 17316 28960
rect 16132 28920 17316 28948
rect 17310 28908 17316 28920
rect 17368 28948 17374 28960
rect 18046 28948 18052 28960
rect 17368 28920 18052 28948
rect 17368 28908 17374 28920
rect 18046 28908 18052 28920
rect 18104 28948 18110 28960
rect 19444 28948 19472 28988
rect 21174 28976 21180 28988
rect 21232 28976 21238 29028
rect 20346 28948 20352 28960
rect 18104 28920 19472 28948
rect 20307 28920 20352 28948
rect 18104 28908 18110 28920
rect 20346 28908 20352 28920
rect 20404 28908 20410 28960
rect 21278 28948 21306 29056
rect 24486 29044 24492 29056
rect 24544 29044 24550 29096
rect 28184 29028 28212 29115
rect 29457 29087 29515 29093
rect 29457 29084 29469 29087
rect 28460 29056 29469 29084
rect 21821 29019 21879 29025
rect 21821 28985 21833 29019
rect 21867 29016 21879 29019
rect 22094 29016 22100 29028
rect 21867 28988 22100 29016
rect 21867 28985 21879 28988
rect 21821 28979 21879 28985
rect 22094 28976 22100 28988
rect 22152 28976 22158 29028
rect 28166 28976 28172 29028
rect 28224 28976 28230 29028
rect 28350 29016 28356 29028
rect 28311 28988 28356 29016
rect 28350 28976 28356 28988
rect 28408 28976 28414 29028
rect 21450 28948 21456 28960
rect 21278 28920 21456 28948
rect 21450 28908 21456 28920
rect 21508 28948 21514 28960
rect 24854 28948 24860 28960
rect 21508 28920 24860 28948
rect 21508 28908 21514 28920
rect 24854 28908 24860 28920
rect 24912 28908 24918 28960
rect 28074 28908 28080 28960
rect 28132 28948 28138 28960
rect 28460 28948 28488 29056
rect 29457 29053 29469 29056
rect 29503 29053 29515 29087
rect 29457 29047 29515 29053
rect 29733 29087 29791 29093
rect 29733 29053 29745 29087
rect 29779 29084 29791 29087
rect 29779 29056 31064 29084
rect 29779 29053 29791 29056
rect 29733 29047 29791 29053
rect 30742 28948 30748 28960
rect 28132 28920 28488 28948
rect 30703 28920 30748 28948
rect 28132 28908 28138 28920
rect 30742 28908 30748 28920
rect 30800 28908 30806 28960
rect 31036 28948 31064 29056
rect 31128 29028 31156 29115
rect 31110 28976 31116 29028
rect 31168 28976 31174 29028
rect 31404 29016 31432 29115
rect 31754 29112 31760 29124
rect 31812 29112 31818 29164
rect 32398 29112 32404 29164
rect 32456 29152 32462 29164
rect 32723 29155 32781 29161
rect 32723 29152 32735 29155
rect 32456 29124 32735 29152
rect 32456 29112 32462 29124
rect 32723 29121 32735 29124
rect 32769 29121 32781 29155
rect 32858 29152 32864 29164
rect 32819 29124 32864 29152
rect 32723 29115 32781 29121
rect 32858 29112 32864 29124
rect 32916 29112 32922 29164
rect 32953 29158 33011 29164
rect 32953 29124 32965 29158
rect 32999 29152 33011 29158
rect 33060 29152 33088 29180
rect 32999 29124 33088 29152
rect 33131 29155 33189 29161
rect 32953 29118 33011 29124
rect 33131 29121 33143 29155
rect 33177 29150 33189 29155
rect 33502 29152 33508 29164
rect 33244 29150 33508 29152
rect 33177 29124 33508 29150
rect 33177 29122 33272 29124
rect 33177 29121 33189 29122
rect 33131 29115 33189 29121
rect 33502 29112 33508 29124
rect 33560 29112 33566 29164
rect 33594 29112 33600 29164
rect 33652 29152 33658 29164
rect 33689 29155 33747 29161
rect 33689 29152 33701 29155
rect 33652 29124 33701 29152
rect 33652 29112 33658 29124
rect 33689 29121 33701 29124
rect 33735 29121 33747 29155
rect 33689 29115 33747 29121
rect 33778 29112 33784 29164
rect 33836 29152 33842 29164
rect 33945 29155 34003 29161
rect 33945 29152 33957 29155
rect 33836 29124 33957 29152
rect 33836 29112 33842 29124
rect 33945 29121 33957 29124
rect 33991 29121 34003 29155
rect 36354 29152 36360 29164
rect 36315 29124 36360 29152
rect 33945 29115 34003 29121
rect 36354 29112 36360 29124
rect 36412 29112 36418 29164
rect 46290 29112 46296 29164
rect 46348 29152 46354 29164
rect 47581 29155 47639 29161
rect 47581 29152 47593 29155
rect 46348 29124 47593 29152
rect 46348 29112 46354 29124
rect 47581 29121 47593 29124
rect 47627 29121 47639 29155
rect 47581 29115 47639 29121
rect 32490 29044 32496 29096
rect 32548 29084 32554 29096
rect 33612 29084 33640 29112
rect 32548 29056 33640 29084
rect 32548 29044 32554 29056
rect 47486 29044 47492 29096
rect 47544 29084 47550 29096
rect 47762 29084 47768 29096
rect 47544 29056 47768 29084
rect 47544 29044 47550 29056
rect 47762 29044 47768 29056
rect 47820 29044 47826 29096
rect 31220 28988 31432 29016
rect 35069 29019 35127 29025
rect 31220 28948 31248 28988
rect 35069 28985 35081 29019
rect 35115 29016 35127 29019
rect 35526 29016 35532 29028
rect 35115 28988 35532 29016
rect 35115 28985 35127 28988
rect 35069 28979 35127 28985
rect 35526 28976 35532 28988
rect 35584 28976 35590 29028
rect 47670 28948 47676 28960
rect 31036 28920 31248 28948
rect 47631 28920 47676 28948
rect 47670 28908 47676 28920
rect 47728 28908 47734 28960
rect 1104 28858 48852 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 48852 28858
rect 1104 28784 48852 28806
rect 8205 28747 8263 28753
rect 8205 28713 8217 28747
rect 8251 28744 8263 28747
rect 8294 28744 8300 28756
rect 8251 28716 8300 28744
rect 8251 28713 8263 28716
rect 8205 28707 8263 28713
rect 8294 28704 8300 28716
rect 8352 28704 8358 28756
rect 8389 28747 8447 28753
rect 8389 28713 8401 28747
rect 8435 28744 8447 28747
rect 9122 28744 9128 28756
rect 8435 28716 9128 28744
rect 8435 28713 8447 28716
rect 8389 28707 8447 28713
rect 9122 28704 9128 28716
rect 9180 28704 9186 28756
rect 11333 28747 11391 28753
rect 11333 28713 11345 28747
rect 11379 28744 11391 28747
rect 11606 28744 11612 28756
rect 11379 28716 11612 28744
rect 11379 28713 11391 28716
rect 11333 28707 11391 28713
rect 11606 28704 11612 28716
rect 11664 28704 11670 28756
rect 15654 28744 15660 28756
rect 15567 28716 15660 28744
rect 15654 28704 15660 28716
rect 15712 28744 15718 28756
rect 17405 28747 17463 28753
rect 15712 28716 16160 28744
rect 15712 28704 15718 28716
rect 7837 28679 7895 28685
rect 7837 28645 7849 28679
rect 7883 28676 7895 28679
rect 8846 28676 8852 28688
rect 7883 28648 8852 28676
rect 7883 28645 7895 28648
rect 7837 28639 7895 28645
rect 8846 28636 8852 28648
rect 8904 28636 8910 28688
rect 1394 28608 1400 28620
rect 1355 28580 1400 28608
rect 1394 28568 1400 28580
rect 1452 28568 1458 28620
rect 2774 28568 2780 28620
rect 2832 28608 2838 28620
rect 9585 28611 9643 28617
rect 2832 28580 2877 28608
rect 2832 28568 2838 28580
rect 9585 28577 9597 28611
rect 9631 28577 9643 28611
rect 9585 28571 9643 28577
rect 1581 28475 1639 28481
rect 1581 28441 1593 28475
rect 1627 28472 1639 28475
rect 2314 28472 2320 28484
rect 1627 28444 2320 28472
rect 1627 28441 1639 28444
rect 1581 28435 1639 28441
rect 2314 28432 2320 28444
rect 2372 28432 2378 28484
rect 8205 28475 8263 28481
rect 8205 28441 8217 28475
rect 8251 28472 8263 28475
rect 8251 28444 9444 28472
rect 8251 28441 8263 28444
rect 8205 28435 8263 28441
rect 9416 28413 9444 28444
rect 9401 28407 9459 28413
rect 9401 28373 9413 28407
rect 9447 28373 9459 28407
rect 9600 28404 9628 28571
rect 9766 28568 9772 28620
rect 9824 28608 9830 28620
rect 12161 28611 12219 28617
rect 9824 28580 9869 28608
rect 9824 28568 9830 28580
rect 12161 28577 12173 28611
rect 12207 28608 12219 28611
rect 13265 28611 13323 28617
rect 13265 28608 13277 28611
rect 12207 28580 13277 28608
rect 12207 28577 12219 28580
rect 12161 28571 12219 28577
rect 13265 28577 13277 28580
rect 13311 28608 13323 28611
rect 13354 28608 13360 28620
rect 13311 28580 13360 28608
rect 13311 28577 13323 28580
rect 13265 28571 13323 28577
rect 13354 28568 13360 28580
rect 13412 28568 13418 28620
rect 13541 28611 13599 28617
rect 13541 28577 13553 28611
rect 13587 28608 13599 28611
rect 13998 28608 14004 28620
rect 13587 28580 14004 28608
rect 13587 28577 13599 28580
rect 13541 28571 13599 28577
rect 13998 28568 14004 28580
rect 14056 28568 14062 28620
rect 16132 28617 16160 28716
rect 17405 28713 17417 28747
rect 17451 28744 17463 28747
rect 18598 28744 18604 28756
rect 17451 28716 18604 28744
rect 17451 28713 17463 28716
rect 17405 28707 17463 28713
rect 18598 28704 18604 28716
rect 18656 28704 18662 28756
rect 20898 28704 20904 28756
rect 20956 28744 20962 28756
rect 21361 28747 21419 28753
rect 21361 28744 21373 28747
rect 20956 28716 21373 28744
rect 20956 28704 20962 28716
rect 21361 28713 21373 28716
rect 21407 28713 21419 28747
rect 21361 28707 21419 28713
rect 27982 28704 27988 28756
rect 28040 28744 28046 28756
rect 28261 28747 28319 28753
rect 28261 28744 28273 28747
rect 28040 28716 28273 28744
rect 28040 28704 28046 28716
rect 28261 28713 28273 28716
rect 28307 28713 28319 28747
rect 28261 28707 28319 28713
rect 31202 28704 31208 28756
rect 31260 28744 31266 28756
rect 31481 28747 31539 28753
rect 31481 28744 31493 28747
rect 31260 28716 31493 28744
rect 31260 28704 31266 28716
rect 31481 28713 31493 28716
rect 31527 28713 31539 28747
rect 31481 28707 31539 28713
rect 33318 28704 33324 28756
rect 33376 28744 33382 28756
rect 33413 28747 33471 28753
rect 33413 28744 33425 28747
rect 33376 28716 33425 28744
rect 33376 28704 33382 28716
rect 33413 28713 33425 28716
rect 33459 28713 33471 28747
rect 33413 28707 33471 28713
rect 17770 28636 17776 28688
rect 17828 28636 17834 28688
rect 30484 28648 32168 28676
rect 16117 28611 16175 28617
rect 16117 28577 16129 28611
rect 16163 28577 16175 28611
rect 16117 28571 16175 28577
rect 9677 28543 9735 28549
rect 9677 28509 9689 28543
rect 9723 28509 9735 28543
rect 9677 28503 9735 28509
rect 9861 28543 9919 28549
rect 9861 28509 9873 28543
rect 9907 28540 9919 28543
rect 10226 28540 10232 28552
rect 9907 28512 10232 28540
rect 9907 28509 9919 28512
rect 9861 28503 9919 28509
rect 9692 28472 9720 28503
rect 10226 28500 10232 28512
rect 10284 28500 10290 28552
rect 11514 28540 11520 28552
rect 11475 28512 11520 28540
rect 11514 28500 11520 28512
rect 11572 28500 11578 28552
rect 12250 28540 12256 28552
rect 12211 28512 12256 28540
rect 12250 28500 12256 28512
rect 12308 28500 12314 28552
rect 12345 28543 12403 28549
rect 12345 28509 12357 28543
rect 12391 28509 12403 28543
rect 12345 28503 12403 28509
rect 12437 28543 12495 28549
rect 12437 28509 12449 28543
rect 12483 28540 12495 28543
rect 12526 28540 12532 28552
rect 12483 28512 12532 28540
rect 12483 28509 12495 28512
rect 12437 28503 12495 28509
rect 10962 28472 10968 28484
rect 9692 28444 10968 28472
rect 10962 28432 10968 28444
rect 11020 28432 11026 28484
rect 12360 28472 12388 28503
rect 12526 28500 12532 28512
rect 12584 28500 12590 28552
rect 13173 28543 13231 28549
rect 13173 28509 13185 28543
rect 13219 28509 13231 28543
rect 14274 28540 14280 28552
rect 14235 28512 14280 28540
rect 13173 28503 13231 28509
rect 12710 28472 12716 28484
rect 12360 28444 12716 28472
rect 12452 28416 12480 28444
rect 12710 28432 12716 28444
rect 12768 28432 12774 28484
rect 12986 28432 12992 28484
rect 13044 28472 13050 28484
rect 13188 28472 13216 28503
rect 14274 28500 14280 28512
rect 14332 28500 14338 28552
rect 15746 28540 15752 28552
rect 14384 28512 15752 28540
rect 14384 28472 14412 28512
rect 15746 28500 15752 28512
rect 15804 28540 15810 28552
rect 17788 28549 17816 28636
rect 18322 28608 18328 28620
rect 17880 28580 18328 28608
rect 17880 28549 17908 28580
rect 18322 28568 18328 28580
rect 18380 28568 18386 28620
rect 21818 28608 21824 28620
rect 21779 28580 21824 28608
rect 21818 28568 21824 28580
rect 21876 28568 21882 28620
rect 24486 28568 24492 28620
rect 24544 28608 24550 28620
rect 24673 28611 24731 28617
rect 24673 28608 24685 28611
rect 24544 28580 24685 28608
rect 24544 28568 24550 28580
rect 24673 28577 24685 28580
rect 24719 28577 24731 28611
rect 28718 28608 28724 28620
rect 28679 28580 28724 28608
rect 24673 28571 24731 28577
rect 28718 28568 28724 28580
rect 28776 28568 28782 28620
rect 30484 28617 30512 28648
rect 28905 28611 28963 28617
rect 28905 28577 28917 28611
rect 28951 28608 28963 28611
rect 30469 28611 30527 28617
rect 30469 28608 30481 28611
rect 28951 28580 30481 28608
rect 28951 28577 28963 28580
rect 28905 28571 28963 28577
rect 30469 28577 30481 28580
rect 30515 28577 30527 28611
rect 30469 28571 30527 28577
rect 31386 28568 31392 28620
rect 31444 28608 31450 28620
rect 32140 28617 32168 28648
rect 31941 28611 31999 28617
rect 31941 28608 31953 28611
rect 31444 28580 31953 28608
rect 31444 28568 31450 28580
rect 31941 28577 31953 28580
rect 31987 28577 31999 28611
rect 31941 28571 31999 28577
rect 32125 28611 32183 28617
rect 32125 28577 32137 28611
rect 32171 28608 32183 28611
rect 32953 28611 33011 28617
rect 32953 28608 32965 28611
rect 32171 28580 32965 28608
rect 32171 28577 32183 28580
rect 32125 28571 32183 28577
rect 32953 28577 32965 28580
rect 32999 28608 33011 28611
rect 33962 28608 33968 28620
rect 32999 28580 33968 28608
rect 32999 28577 33011 28580
rect 32953 28571 33011 28577
rect 33962 28568 33968 28580
rect 34020 28568 34026 28620
rect 46477 28611 46535 28617
rect 46477 28577 46489 28611
rect 46523 28608 46535 28611
rect 47670 28608 47676 28620
rect 46523 28580 47676 28608
rect 46523 28577 46535 28580
rect 46477 28571 46535 28577
rect 47670 28568 47676 28580
rect 47728 28568 47734 28620
rect 48130 28608 48136 28620
rect 48091 28580 48136 28608
rect 48130 28568 48136 28580
rect 48188 28568 48194 28620
rect 16393 28543 16451 28549
rect 16393 28540 16405 28543
rect 15804 28512 16405 28540
rect 15804 28500 15810 28512
rect 16393 28509 16405 28512
rect 16439 28509 16451 28543
rect 17661 28543 17719 28549
rect 17661 28540 17673 28543
rect 16393 28503 16451 28509
rect 17650 28509 17673 28540
rect 17707 28509 17719 28543
rect 17650 28503 17719 28509
rect 17770 28543 17828 28549
rect 17770 28509 17782 28543
rect 17816 28509 17828 28543
rect 17770 28503 17828 28509
rect 17870 28543 17928 28549
rect 17870 28509 17882 28543
rect 17916 28509 17928 28543
rect 18046 28540 18052 28552
rect 18007 28512 18052 28540
rect 17870 28503 17928 28509
rect 13044 28444 14412 28472
rect 14544 28475 14602 28481
rect 13044 28432 13050 28444
rect 14544 28441 14556 28475
rect 14590 28472 14602 28475
rect 14642 28472 14648 28484
rect 14590 28444 14648 28472
rect 14590 28441 14602 28444
rect 14544 28435 14602 28441
rect 14642 28432 14648 28444
rect 14700 28432 14706 28484
rect 14734 28432 14740 28484
rect 14792 28472 14798 28484
rect 17650 28472 17678 28503
rect 18046 28500 18052 28512
rect 18104 28500 18110 28552
rect 19981 28543 20039 28549
rect 19981 28509 19993 28543
rect 20027 28540 20039 28543
rect 20070 28540 20076 28552
rect 20027 28512 20076 28540
rect 20027 28509 20039 28512
rect 19981 28503 20039 28509
rect 20070 28500 20076 28512
rect 20128 28540 20134 28552
rect 21836 28540 21864 28568
rect 22094 28549 22100 28552
rect 20128 28512 21864 28540
rect 20128 28500 20134 28512
rect 22088 28503 22100 28549
rect 22152 28540 22158 28552
rect 27341 28543 27399 28549
rect 22152 28512 22188 28540
rect 22094 28500 22100 28503
rect 22152 28500 22158 28512
rect 27341 28509 27353 28543
rect 27387 28540 27399 28543
rect 27614 28540 27620 28552
rect 27387 28512 27620 28540
rect 27387 28509 27399 28512
rect 27341 28503 27399 28509
rect 27614 28500 27620 28512
rect 27672 28500 27678 28552
rect 28810 28500 28816 28552
rect 28868 28540 28874 28552
rect 30285 28543 30343 28549
rect 30285 28540 30297 28543
rect 28868 28512 30297 28540
rect 28868 28500 28874 28512
rect 30285 28509 30297 28512
rect 30331 28509 30343 28543
rect 30285 28503 30343 28509
rect 31849 28543 31907 28549
rect 31849 28509 31861 28543
rect 31895 28540 31907 28543
rect 33778 28540 33784 28552
rect 31895 28512 33784 28540
rect 31895 28509 31907 28512
rect 31849 28503 31907 28509
rect 33778 28500 33784 28512
rect 33836 28500 33842 28552
rect 33873 28543 33931 28549
rect 33873 28509 33885 28543
rect 33919 28540 33931 28543
rect 34422 28540 34428 28552
rect 33919 28512 34428 28540
rect 33919 28509 33931 28512
rect 33873 28503 33931 28509
rect 34422 28500 34428 28512
rect 34480 28500 34486 28552
rect 46293 28543 46351 28549
rect 46293 28509 46305 28543
rect 46339 28509 46351 28543
rect 46293 28503 46351 28509
rect 14792 28444 17678 28472
rect 20248 28475 20306 28481
rect 14792 28432 14798 28444
rect 20248 28441 20260 28475
rect 20294 28472 20306 28475
rect 20346 28472 20352 28484
rect 20294 28444 20352 28472
rect 20294 28441 20306 28444
rect 20248 28435 20306 28441
rect 20346 28432 20352 28444
rect 20404 28432 20410 28484
rect 24578 28432 24584 28484
rect 24636 28472 24642 28484
rect 24918 28475 24976 28481
rect 24918 28472 24930 28475
rect 24636 28444 24930 28472
rect 24636 28432 24642 28444
rect 24918 28441 24930 28444
rect 24964 28441 24976 28475
rect 24918 28435 24976 28441
rect 32582 28432 32588 28484
rect 32640 28472 32646 28484
rect 32769 28475 32827 28481
rect 32769 28472 32781 28475
rect 32640 28444 32781 28472
rect 32640 28432 32646 28444
rect 32769 28441 32781 28444
rect 32815 28441 32827 28475
rect 46308 28472 46336 28503
rect 47670 28472 47676 28484
rect 46308 28444 47676 28472
rect 32769 28435 32827 28441
rect 47670 28432 47676 28444
rect 47728 28432 47734 28484
rect 9950 28404 9956 28416
rect 9600 28376 9956 28404
rect 9401 28367 9459 28373
rect 9950 28364 9956 28376
rect 10008 28364 10014 28416
rect 11974 28404 11980 28416
rect 11935 28376 11980 28404
rect 11974 28364 11980 28376
rect 12032 28364 12038 28416
rect 12434 28364 12440 28416
rect 12492 28364 12498 28416
rect 23201 28407 23259 28413
rect 23201 28373 23213 28407
rect 23247 28404 23259 28407
rect 23474 28404 23480 28416
rect 23247 28376 23480 28404
rect 23247 28373 23259 28376
rect 23201 28367 23259 28373
rect 23474 28364 23480 28376
rect 23532 28364 23538 28416
rect 26050 28404 26056 28416
rect 26011 28376 26056 28404
rect 26050 28364 26056 28376
rect 26108 28364 26114 28416
rect 27430 28404 27436 28416
rect 27391 28376 27436 28404
rect 27430 28364 27436 28376
rect 27488 28364 27494 28416
rect 28626 28404 28632 28416
rect 28587 28376 28632 28404
rect 28626 28364 28632 28376
rect 28684 28364 28690 28416
rect 29822 28404 29828 28416
rect 29783 28376 29828 28404
rect 29822 28364 29828 28376
rect 29880 28364 29886 28416
rect 30193 28407 30251 28413
rect 30193 28373 30205 28407
rect 30239 28404 30251 28407
rect 31570 28404 31576 28416
rect 30239 28376 31576 28404
rect 30239 28373 30251 28376
rect 30193 28367 30251 28373
rect 31570 28364 31576 28376
rect 31628 28364 31634 28416
rect 33781 28407 33839 28413
rect 33781 28373 33793 28407
rect 33827 28404 33839 28407
rect 35526 28404 35532 28416
rect 33827 28376 35532 28404
rect 33827 28373 33839 28376
rect 33781 28367 33839 28373
rect 35526 28364 35532 28376
rect 35584 28364 35590 28416
rect 1104 28314 48852 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 48852 28314
rect 1104 28240 48852 28262
rect 2314 28200 2320 28212
rect 2275 28172 2320 28200
rect 2314 28160 2320 28172
rect 2372 28160 2378 28212
rect 8294 28160 8300 28212
rect 8352 28200 8358 28212
rect 8352 28172 11468 28200
rect 8352 28160 8358 28172
rect 8389 28135 8447 28141
rect 8389 28101 8401 28135
rect 8435 28132 8447 28135
rect 11440 28132 11468 28172
rect 11514 28160 11520 28212
rect 11572 28200 11578 28212
rect 12161 28203 12219 28209
rect 12161 28200 12173 28203
rect 11572 28172 12173 28200
rect 11572 28160 11578 28172
rect 12161 28169 12173 28172
rect 12207 28169 12219 28203
rect 12161 28163 12219 28169
rect 12250 28160 12256 28212
rect 12308 28200 12314 28212
rect 12986 28200 12992 28212
rect 12308 28172 12992 28200
rect 12308 28160 12314 28172
rect 12986 28160 12992 28172
rect 13044 28160 13050 28212
rect 13081 28203 13139 28209
rect 13081 28169 13093 28203
rect 13127 28200 13139 28203
rect 14366 28200 14372 28212
rect 13127 28172 14372 28200
rect 13127 28169 13139 28172
rect 13081 28163 13139 28169
rect 14366 28160 14372 28172
rect 14424 28160 14430 28212
rect 14642 28200 14648 28212
rect 14603 28172 14648 28200
rect 14642 28160 14648 28172
rect 14700 28160 14706 28212
rect 16574 28160 16580 28212
rect 16632 28200 16638 28212
rect 17037 28203 17095 28209
rect 17037 28200 17049 28203
rect 16632 28172 17049 28200
rect 16632 28160 16638 28172
rect 17037 28169 17049 28172
rect 17083 28169 17095 28203
rect 17037 28163 17095 28169
rect 22278 28160 22284 28212
rect 22336 28200 22342 28212
rect 23293 28203 23351 28209
rect 23293 28200 23305 28203
rect 22336 28172 23305 28200
rect 22336 28160 22342 28172
rect 23293 28169 23305 28172
rect 23339 28169 23351 28203
rect 23293 28163 23351 28169
rect 24489 28203 24547 28209
rect 24489 28169 24501 28203
rect 24535 28200 24547 28203
rect 24578 28200 24584 28212
rect 24535 28172 24584 28200
rect 24535 28169 24547 28172
rect 24489 28163 24547 28169
rect 24578 28160 24584 28172
rect 24636 28160 24642 28212
rect 33778 28160 33784 28212
rect 33836 28200 33842 28212
rect 33873 28203 33931 28209
rect 33873 28200 33885 28203
rect 33836 28172 33885 28200
rect 33836 28160 33842 28172
rect 33873 28169 33885 28172
rect 33919 28169 33931 28203
rect 33873 28163 33931 28169
rect 11882 28132 11888 28144
rect 8435 28104 9904 28132
rect 11440 28104 11888 28132
rect 8435 28101 8447 28104
rect 8389 28095 8447 28101
rect 9876 28076 9904 28104
rect 11882 28092 11888 28104
rect 11940 28132 11946 28144
rect 11977 28135 12035 28141
rect 11977 28132 11989 28135
rect 11940 28104 11989 28132
rect 11940 28092 11946 28104
rect 11977 28101 11989 28104
rect 12023 28132 12035 28135
rect 14090 28132 14096 28144
rect 12023 28104 14096 28132
rect 12023 28101 12035 28104
rect 11977 28095 12035 28101
rect 2225 28067 2283 28073
rect 2225 28033 2237 28067
rect 2271 28064 2283 28067
rect 3510 28064 3516 28076
rect 2271 28036 3516 28064
rect 2271 28033 2283 28036
rect 2225 28027 2283 28033
rect 3510 28024 3516 28036
rect 3568 28024 3574 28076
rect 7929 28067 7987 28073
rect 7929 28033 7941 28067
rect 7975 28064 7987 28067
rect 8294 28064 8300 28076
rect 7975 28036 8300 28064
rect 7975 28033 7987 28036
rect 7929 28027 7987 28033
rect 8294 28024 8300 28036
rect 8352 28024 8358 28076
rect 8573 28067 8631 28073
rect 8573 28033 8585 28067
rect 8619 28064 8631 28067
rect 9493 28067 9551 28073
rect 8619 28036 9260 28064
rect 8619 28033 8631 28036
rect 8573 28027 8631 28033
rect 9232 28005 9260 28036
rect 9493 28033 9505 28067
rect 9539 28064 9551 28067
rect 9766 28064 9772 28076
rect 9539 28036 9772 28064
rect 9539 28033 9551 28036
rect 9493 28027 9551 28033
rect 9766 28024 9772 28036
rect 9824 28024 9830 28076
rect 9858 28024 9864 28076
rect 9916 28064 9922 28076
rect 10505 28067 10563 28073
rect 10505 28064 10517 28067
rect 9916 28036 10517 28064
rect 9916 28024 9922 28036
rect 10505 28033 10517 28036
rect 10551 28033 10563 28067
rect 10505 28027 10563 28033
rect 10689 28067 10747 28073
rect 10689 28033 10701 28067
rect 10735 28033 10747 28067
rect 10689 28027 10747 28033
rect 9217 27999 9275 28005
rect 9217 27965 9229 27999
rect 9263 27996 9275 27999
rect 9306 27996 9312 28008
rect 9263 27968 9312 27996
rect 9263 27965 9275 27968
rect 9217 27959 9275 27965
rect 9306 27956 9312 27968
rect 9364 27956 9370 28008
rect 9784 27996 9812 28024
rect 10704 27996 10732 28027
rect 12710 28024 12716 28076
rect 12768 28064 12774 28076
rect 12897 28067 12955 28073
rect 12897 28064 12909 28067
rect 12768 28036 12909 28064
rect 12768 28024 12774 28036
rect 12897 28033 12909 28036
rect 12943 28064 12955 28067
rect 12986 28064 12992 28076
rect 12943 28036 12992 28064
rect 12943 28033 12955 28036
rect 12897 28027 12955 28033
rect 12986 28024 12992 28036
rect 13044 28024 13050 28076
rect 13832 28073 13860 28104
rect 14090 28092 14096 28104
rect 14148 28092 14154 28144
rect 16669 28135 16727 28141
rect 16669 28101 16681 28135
rect 16715 28132 16727 28135
rect 16758 28132 16764 28144
rect 16715 28104 16764 28132
rect 16715 28101 16727 28104
rect 16669 28095 16727 28101
rect 16758 28092 16764 28104
rect 16816 28092 16822 28144
rect 16853 28135 16911 28141
rect 16853 28101 16865 28135
rect 16899 28132 16911 28135
rect 18138 28132 18144 28144
rect 16899 28104 18144 28132
rect 16899 28101 16911 28104
rect 16853 28095 16911 28101
rect 18138 28092 18144 28104
rect 18196 28092 18202 28144
rect 20990 28092 20996 28144
rect 21048 28132 21054 28144
rect 22554 28132 22560 28144
rect 21048 28104 22560 28132
rect 21048 28092 21054 28104
rect 13817 28067 13875 28073
rect 13817 28033 13829 28067
rect 13863 28033 13875 28067
rect 13998 28064 14004 28076
rect 13959 28036 14004 28064
rect 13817 28027 13875 28033
rect 13998 28024 14004 28036
rect 14056 28024 14062 28076
rect 14185 28067 14243 28073
rect 14185 28033 14197 28067
rect 14231 28064 14243 28067
rect 14829 28067 14887 28073
rect 14829 28064 14841 28067
rect 14231 28036 14841 28064
rect 14231 28033 14243 28036
rect 14185 28027 14243 28033
rect 14829 28033 14841 28036
rect 14875 28033 14887 28067
rect 14829 28027 14887 28033
rect 22051 28067 22109 28073
rect 22051 28033 22063 28067
rect 22097 28033 22109 28067
rect 22186 28064 22192 28076
rect 22147 28036 22192 28064
rect 22051 28027 22109 28033
rect 9784 27968 10732 27996
rect 11609 27999 11667 28005
rect 11609 27965 11621 27999
rect 11655 27996 11667 27999
rect 12158 27996 12164 28008
rect 11655 27968 12164 27996
rect 11655 27965 11667 27968
rect 11609 27959 11667 27965
rect 12158 27956 12164 27968
rect 12216 27996 12222 28008
rect 13265 27999 13323 28005
rect 13265 27996 13277 27999
rect 12216 27968 13277 27996
rect 12216 27956 12222 27968
rect 13265 27965 13277 27968
rect 13311 27965 13323 27999
rect 22066 27996 22094 28027
rect 22186 28024 22192 28036
rect 22244 28024 22250 28076
rect 22278 28024 22284 28076
rect 22336 28064 22342 28076
rect 22480 28073 22508 28104
rect 22554 28092 22560 28104
rect 22612 28132 22618 28144
rect 32490 28132 32496 28144
rect 22612 28104 25176 28132
rect 22612 28092 22618 28104
rect 25148 28076 25176 28104
rect 30208 28104 32496 28132
rect 22465 28067 22523 28073
rect 22336 28036 22381 28064
rect 22336 28024 22342 28036
rect 22465 28033 22477 28067
rect 22511 28033 22523 28067
rect 22922 28064 22928 28076
rect 22883 28036 22928 28064
rect 22465 28027 22523 28033
rect 22922 28024 22928 28036
rect 22980 28024 22986 28076
rect 23109 28067 23167 28073
rect 23109 28033 23121 28067
rect 23155 28064 23167 28067
rect 23474 28064 23480 28076
rect 23155 28036 23480 28064
rect 23155 28033 23167 28036
rect 23109 28027 23167 28033
rect 23474 28024 23480 28036
rect 23532 28024 23538 28076
rect 24394 28024 24400 28076
rect 24452 28064 24458 28076
rect 24719 28067 24777 28073
rect 24719 28064 24731 28067
rect 24452 28036 24731 28064
rect 24452 28024 24458 28036
rect 24719 28033 24731 28036
rect 24765 28033 24777 28067
rect 24854 28064 24860 28076
rect 24815 28036 24860 28064
rect 24719 28027 24777 28033
rect 24854 28024 24860 28036
rect 24912 28024 24918 28076
rect 24946 28024 24952 28076
rect 25004 28064 25010 28076
rect 25004 28036 25049 28064
rect 25004 28024 25010 28036
rect 25130 28024 25136 28076
rect 25188 28064 25194 28076
rect 25188 28036 25233 28064
rect 25188 28024 25194 28036
rect 27614 28024 27620 28076
rect 27672 28064 27678 28076
rect 30208 28073 30236 28104
rect 32490 28092 32496 28104
rect 32548 28092 32554 28144
rect 27965 28067 28023 28073
rect 27965 28064 27977 28067
rect 27672 28036 27977 28064
rect 27672 28024 27678 28036
rect 27965 28033 27977 28036
rect 28011 28033 28023 28067
rect 27965 28027 28023 28033
rect 30193 28067 30251 28073
rect 30193 28033 30205 28067
rect 30239 28033 30251 28067
rect 30193 28027 30251 28033
rect 30460 28067 30518 28073
rect 30460 28033 30472 28067
rect 30506 28064 30518 28067
rect 30742 28064 30748 28076
rect 30506 28036 30748 28064
rect 30506 28033 30518 28036
rect 30460 28027 30518 28033
rect 30742 28024 30748 28036
rect 30800 28024 30806 28076
rect 31938 28024 31944 28076
rect 31996 28064 32002 28076
rect 32749 28067 32807 28073
rect 32749 28064 32761 28067
rect 31996 28036 32761 28064
rect 31996 28024 32002 28036
rect 32749 28033 32761 28036
rect 32795 28033 32807 28067
rect 47946 28064 47952 28076
rect 47907 28036 47952 28064
rect 32749 28027 32807 28033
rect 47946 28024 47952 28036
rect 48004 28024 48010 28076
rect 22830 27996 22836 28008
rect 22066 27968 22836 27996
rect 13265 27959 13323 27965
rect 22830 27956 22836 27968
rect 22888 27956 22894 28008
rect 27522 27956 27528 28008
rect 27580 27996 27586 28008
rect 27709 27999 27767 28005
rect 27709 27996 27721 27999
rect 27580 27968 27721 27996
rect 27580 27956 27586 27968
rect 27709 27965 27721 27968
rect 27755 27965 27767 27999
rect 32490 27996 32496 28008
rect 32451 27968 32496 27996
rect 27709 27959 27767 27965
rect 12526 27888 12532 27940
rect 12584 27928 12590 27940
rect 12713 27931 12771 27937
rect 12713 27928 12725 27931
rect 12584 27900 12725 27928
rect 12584 27888 12590 27900
rect 12713 27897 12725 27900
rect 12759 27897 12771 27931
rect 12713 27891 12771 27897
rect 20254 27888 20260 27940
rect 20312 27928 20318 27940
rect 25774 27928 25780 27940
rect 20312 27900 25780 27928
rect 20312 27888 20318 27900
rect 25774 27888 25780 27900
rect 25832 27888 25838 27940
rect 7282 27820 7288 27872
rect 7340 27860 7346 27872
rect 7745 27863 7803 27869
rect 7745 27860 7757 27863
rect 7340 27832 7757 27860
rect 7340 27820 7346 27832
rect 7745 27829 7757 27832
rect 7791 27829 7803 27863
rect 8754 27860 8760 27872
rect 8715 27832 8760 27860
rect 7745 27823 7803 27829
rect 8754 27820 8760 27832
rect 8812 27820 8818 27872
rect 9674 27820 9680 27872
rect 9732 27860 9738 27872
rect 10597 27863 10655 27869
rect 10597 27860 10609 27863
rect 9732 27832 10609 27860
rect 9732 27820 9738 27832
rect 10597 27829 10609 27832
rect 10643 27829 10655 27863
rect 11974 27860 11980 27872
rect 11935 27832 11980 27860
rect 10597 27823 10655 27829
rect 11974 27820 11980 27832
rect 12032 27820 12038 27872
rect 21821 27863 21879 27869
rect 21821 27829 21833 27863
rect 21867 27860 21879 27863
rect 22094 27860 22100 27872
rect 21867 27832 22100 27860
rect 21867 27829 21879 27832
rect 21821 27823 21879 27829
rect 22094 27820 22100 27832
rect 22152 27820 22158 27872
rect 27724 27860 27752 27959
rect 32490 27956 32496 27968
rect 32548 27956 32554 28008
rect 31128 27900 31754 27928
rect 27890 27860 27896 27872
rect 27724 27832 27896 27860
rect 27890 27820 27896 27832
rect 27948 27820 27954 27872
rect 28626 27820 28632 27872
rect 28684 27860 28690 27872
rect 29089 27863 29147 27869
rect 29089 27860 29101 27863
rect 28684 27832 29101 27860
rect 28684 27820 28690 27832
rect 29089 27829 29101 27832
rect 29135 27860 29147 27863
rect 31128 27860 31156 27900
rect 31570 27860 31576 27872
rect 29135 27832 31156 27860
rect 31531 27832 31576 27860
rect 29135 27829 29147 27832
rect 29089 27823 29147 27829
rect 31570 27820 31576 27832
rect 31628 27820 31634 27872
rect 31726 27860 31754 27900
rect 32398 27860 32404 27872
rect 31726 27832 32404 27860
rect 32398 27820 32404 27832
rect 32456 27820 32462 27872
rect 32508 27860 32536 27956
rect 32766 27860 32772 27872
rect 32508 27832 32772 27860
rect 32766 27820 32772 27832
rect 32824 27820 32830 27872
rect 44174 27820 44180 27872
rect 44232 27860 44238 27872
rect 48041 27863 48099 27869
rect 48041 27860 48053 27863
rect 44232 27832 48053 27860
rect 44232 27820 44238 27832
rect 48041 27829 48053 27832
rect 48087 27829 48099 27863
rect 48041 27823 48099 27829
rect 1104 27770 48852 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 48852 27770
rect 1104 27696 48852 27718
rect 9858 27656 9864 27668
rect 9819 27628 9864 27656
rect 9858 27616 9864 27628
rect 9916 27616 9922 27668
rect 12710 27656 12716 27668
rect 12671 27628 12716 27656
rect 12710 27616 12716 27628
rect 12768 27616 12774 27668
rect 24946 27656 24952 27668
rect 24907 27628 24952 27656
rect 24946 27616 24952 27628
rect 25004 27616 25010 27668
rect 27172 27628 27844 27656
rect 10962 27548 10968 27600
rect 11020 27588 11026 27600
rect 12894 27588 12900 27600
rect 11020 27560 12434 27588
rect 12855 27560 12900 27588
rect 11020 27548 11026 27560
rect 9030 27480 9036 27532
rect 9088 27520 9094 27532
rect 9088 27492 11100 27520
rect 9088 27480 9094 27492
rect 1394 27412 1400 27464
rect 1452 27452 1458 27464
rect 1581 27455 1639 27461
rect 1581 27452 1593 27455
rect 1452 27424 1593 27452
rect 1452 27412 1458 27424
rect 1581 27421 1593 27424
rect 1627 27421 1639 27455
rect 2038 27452 2044 27464
rect 1999 27424 2044 27452
rect 1581 27415 1639 27421
rect 2038 27412 2044 27424
rect 2096 27452 2102 27464
rect 2314 27452 2320 27464
rect 2096 27424 2320 27452
rect 2096 27412 2102 27424
rect 2314 27412 2320 27424
rect 2372 27412 2378 27464
rect 2869 27455 2927 27461
rect 2869 27452 2881 27455
rect 2746 27424 2881 27452
rect 1762 27344 1768 27396
rect 1820 27384 1826 27396
rect 2746 27384 2774 27424
rect 2869 27421 2881 27424
rect 2915 27421 2927 27455
rect 2869 27415 2927 27421
rect 7009 27455 7067 27461
rect 7009 27421 7021 27455
rect 7055 27452 7067 27455
rect 7742 27452 7748 27464
rect 7055 27424 7748 27452
rect 7055 27421 7067 27424
rect 7009 27415 7067 27421
rect 7742 27412 7748 27424
rect 7800 27412 7806 27464
rect 9585 27455 9643 27461
rect 9585 27421 9597 27455
rect 9631 27421 9643 27455
rect 9585 27415 9643 27421
rect 9677 27455 9735 27461
rect 9677 27421 9689 27455
rect 9723 27452 9735 27455
rect 9950 27452 9956 27464
rect 9723 27424 9956 27452
rect 9723 27421 9735 27424
rect 9677 27415 9735 27421
rect 7282 27393 7288 27396
rect 7276 27384 7288 27393
rect 1820 27356 2774 27384
rect 7243 27356 7288 27384
rect 1820 27344 1826 27356
rect 7276 27347 7288 27356
rect 7282 27344 7288 27347
rect 7340 27344 7346 27396
rect 9600 27384 9628 27415
rect 9950 27412 9956 27424
rect 10008 27452 10014 27464
rect 10321 27455 10379 27461
rect 10321 27452 10333 27455
rect 10008 27424 10333 27452
rect 10008 27412 10014 27424
rect 10321 27421 10333 27424
rect 10367 27452 10379 27455
rect 10870 27452 10876 27464
rect 10367 27424 10876 27452
rect 10367 27421 10379 27424
rect 10321 27415 10379 27421
rect 10870 27412 10876 27424
rect 10928 27412 10934 27464
rect 10410 27384 10416 27396
rect 9600 27356 10416 27384
rect 10410 27344 10416 27356
rect 10468 27384 10474 27396
rect 10505 27387 10563 27393
rect 10505 27384 10517 27387
rect 10468 27356 10517 27384
rect 10468 27344 10474 27356
rect 10505 27353 10517 27356
rect 10551 27384 10563 27387
rect 10962 27384 10968 27396
rect 10551 27356 10968 27384
rect 10551 27353 10563 27356
rect 10505 27347 10563 27353
rect 10962 27344 10968 27356
rect 11020 27344 11026 27396
rect 1946 27276 1952 27328
rect 2004 27316 2010 27328
rect 2133 27319 2191 27325
rect 2133 27316 2145 27319
rect 2004 27288 2145 27316
rect 2004 27276 2010 27288
rect 2133 27285 2145 27288
rect 2179 27285 2191 27319
rect 2133 27279 2191 27285
rect 8389 27319 8447 27325
rect 8389 27285 8401 27319
rect 8435 27316 8447 27319
rect 9306 27316 9312 27328
rect 8435 27288 9312 27316
rect 8435 27285 8447 27288
rect 8389 27279 8447 27285
rect 9306 27276 9312 27288
rect 9364 27276 9370 27328
rect 10686 27316 10692 27328
rect 10647 27288 10692 27316
rect 10686 27276 10692 27288
rect 10744 27276 10750 27328
rect 11072 27316 11100 27492
rect 12406 27452 12434 27560
rect 12894 27548 12900 27560
rect 12952 27548 12958 27600
rect 14274 27548 14280 27600
rect 14332 27588 14338 27600
rect 17126 27588 17132 27600
rect 14332 27560 17132 27588
rect 14332 27548 14338 27560
rect 17126 27548 17132 27560
rect 17184 27548 17190 27600
rect 26050 27548 26056 27600
rect 26108 27588 26114 27600
rect 27172 27588 27200 27628
rect 26108 27560 27200 27588
rect 27249 27591 27307 27597
rect 26108 27548 26114 27560
rect 27249 27557 27261 27591
rect 27295 27588 27307 27591
rect 27614 27588 27620 27600
rect 27295 27560 27620 27588
rect 27295 27557 27307 27560
rect 27249 27551 27307 27557
rect 27614 27548 27620 27560
rect 27672 27548 27678 27600
rect 27706 27548 27712 27600
rect 27764 27548 27770 27600
rect 27816 27588 27844 27628
rect 30190 27588 30196 27600
rect 27816 27560 29960 27588
rect 30151 27560 30196 27588
rect 12526 27480 12532 27532
rect 12584 27520 12590 27532
rect 17586 27520 17592 27532
rect 12584 27492 17592 27520
rect 12584 27480 12590 27492
rect 17586 27480 17592 27492
rect 17644 27480 17650 27532
rect 21818 27480 21824 27532
rect 21876 27520 21882 27532
rect 22005 27523 22063 27529
rect 22005 27520 22017 27523
rect 21876 27492 22017 27520
rect 21876 27480 21882 27492
rect 22005 27489 22017 27492
rect 22051 27489 22063 27523
rect 22005 27483 22063 27489
rect 12713 27455 12771 27461
rect 12713 27452 12725 27455
rect 12406 27424 12725 27452
rect 12713 27421 12725 27424
rect 12759 27421 12771 27455
rect 12713 27415 12771 27421
rect 16758 27412 16764 27464
rect 16816 27452 16822 27464
rect 17862 27452 17868 27464
rect 16816 27424 17868 27452
rect 16816 27412 16822 27424
rect 17862 27412 17868 27424
rect 17920 27452 17926 27464
rect 17957 27455 18015 27461
rect 17957 27452 17969 27455
rect 17920 27424 17969 27452
rect 17920 27412 17926 27424
rect 17957 27421 17969 27424
rect 18003 27421 18015 27455
rect 17957 27415 18015 27421
rect 20162 27412 20168 27464
rect 20220 27452 20226 27464
rect 20257 27455 20315 27461
rect 20257 27452 20269 27455
rect 20220 27424 20269 27452
rect 20220 27412 20226 27424
rect 20257 27421 20269 27424
rect 20303 27421 20315 27455
rect 22020 27452 22048 27483
rect 23474 27480 23480 27532
rect 23532 27520 23538 27532
rect 27724 27520 27752 27548
rect 28350 27520 28356 27532
rect 23532 27492 27568 27520
rect 23532 27480 23538 27492
rect 24486 27452 24492 27464
rect 22020 27424 24492 27452
rect 20257 27415 20315 27421
rect 24486 27412 24492 27424
rect 24544 27412 24550 27464
rect 27540 27461 27568 27492
rect 27629 27492 27752 27520
rect 27816 27492 28356 27520
rect 27629 27461 27657 27492
rect 27525 27455 27583 27461
rect 27525 27421 27537 27455
rect 27571 27421 27583 27455
rect 27525 27415 27583 27421
rect 27614 27455 27672 27461
rect 27614 27421 27626 27455
rect 27660 27421 27672 27455
rect 27614 27415 27672 27421
rect 27730 27455 27788 27461
rect 27730 27421 27742 27455
rect 27776 27452 27788 27455
rect 27816 27452 27844 27492
rect 28350 27480 28356 27492
rect 28408 27480 28414 27532
rect 27776 27424 27844 27452
rect 27893 27455 27951 27461
rect 27776 27421 27788 27424
rect 27730 27415 27788 27421
rect 27893 27421 27905 27455
rect 27939 27452 27951 27455
rect 27982 27452 27988 27464
rect 27939 27424 27988 27452
rect 27939 27421 27951 27424
rect 27893 27415 27951 27421
rect 27982 27412 27988 27424
rect 28040 27412 28046 27464
rect 29822 27452 29828 27464
rect 29783 27424 29828 27452
rect 29822 27412 29828 27424
rect 29880 27412 29886 27464
rect 29932 27452 29960 27560
rect 30190 27548 30196 27560
rect 30248 27548 30254 27600
rect 30929 27591 30987 27597
rect 30929 27557 30941 27591
rect 30975 27588 30987 27591
rect 31938 27588 31944 27600
rect 30975 27560 31944 27588
rect 30975 27557 30987 27560
rect 30929 27551 30987 27557
rect 31938 27548 31944 27560
rect 31996 27548 32002 27600
rect 47670 27588 47676 27600
rect 47631 27560 47676 27588
rect 47670 27548 47676 27560
rect 47728 27548 47734 27600
rect 31159 27455 31217 27461
rect 31159 27452 31171 27455
rect 29932 27424 31171 27452
rect 31159 27421 31171 27424
rect 31205 27421 31217 27455
rect 31159 27415 31217 27421
rect 31297 27455 31355 27461
rect 31297 27421 31309 27455
rect 31343 27421 31355 27455
rect 31297 27415 31355 27421
rect 31389 27455 31447 27461
rect 31389 27421 31401 27455
rect 31435 27452 31447 27455
rect 31478 27452 31484 27464
rect 31435 27424 31484 27452
rect 31435 27421 31447 27424
rect 31389 27415 31447 27421
rect 12437 27387 12495 27393
rect 12437 27353 12449 27387
rect 12483 27384 12495 27387
rect 12618 27384 12624 27396
rect 12483 27356 12624 27384
rect 12483 27353 12495 27356
rect 12437 27347 12495 27353
rect 12618 27344 12624 27356
rect 12676 27384 12682 27396
rect 14734 27384 14740 27396
rect 12676 27356 14740 27384
rect 12676 27344 12682 27356
rect 14734 27344 14740 27356
rect 14792 27344 14798 27396
rect 18141 27387 18199 27393
rect 18141 27353 18153 27387
rect 18187 27384 18199 27387
rect 19426 27384 19432 27396
rect 18187 27356 19432 27384
rect 18187 27353 18199 27356
rect 18141 27347 18199 27353
rect 19426 27344 19432 27356
rect 19484 27344 19490 27396
rect 19518 27344 19524 27396
rect 19576 27384 19582 27396
rect 20806 27384 20812 27396
rect 19576 27356 20812 27384
rect 19576 27344 19582 27356
rect 20806 27344 20812 27356
rect 20864 27344 20870 27396
rect 22094 27344 22100 27396
rect 22152 27384 22158 27396
rect 22250 27387 22308 27393
rect 22250 27384 22262 27387
rect 22152 27356 22262 27384
rect 22152 27344 22158 27356
rect 22250 27353 22262 27356
rect 22296 27353 22308 27387
rect 22250 27347 22308 27353
rect 22922 27344 22928 27396
rect 22980 27384 22986 27396
rect 24581 27387 24639 27393
rect 24581 27384 24593 27387
rect 22980 27356 24593 27384
rect 22980 27344 22986 27356
rect 24581 27353 24593 27356
rect 24627 27353 24639 27387
rect 24581 27347 24639 27353
rect 24765 27387 24823 27393
rect 24765 27353 24777 27387
rect 24811 27384 24823 27387
rect 26050 27384 26056 27396
rect 24811 27356 26056 27384
rect 24811 27353 24823 27356
rect 24765 27347 24823 27353
rect 26050 27344 26056 27356
rect 26108 27344 26114 27396
rect 28902 27344 28908 27396
rect 28960 27384 28966 27396
rect 30009 27387 30067 27393
rect 30009 27384 30021 27387
rect 28960 27356 30021 27384
rect 28960 27344 28966 27356
rect 30009 27353 30021 27356
rect 30055 27353 30067 27387
rect 31312 27384 31340 27415
rect 31478 27412 31484 27424
rect 31536 27412 31542 27464
rect 31573 27455 31631 27461
rect 31573 27421 31585 27455
rect 31619 27452 31631 27455
rect 31754 27452 31760 27464
rect 31619 27424 31760 27452
rect 31619 27421 31631 27424
rect 31573 27415 31631 27421
rect 31754 27412 31760 27424
rect 31812 27412 31818 27464
rect 32125 27455 32183 27461
rect 32125 27421 32137 27455
rect 32171 27452 32183 27455
rect 32306 27452 32312 27464
rect 32171 27424 32312 27452
rect 32171 27421 32183 27424
rect 32125 27415 32183 27421
rect 32306 27412 32312 27424
rect 32364 27412 32370 27464
rect 30009 27347 30067 27353
rect 31128 27356 31340 27384
rect 31128 27328 31156 27356
rect 12802 27316 12808 27328
rect 11072 27288 12808 27316
rect 12802 27276 12808 27288
rect 12860 27276 12866 27328
rect 17034 27276 17040 27328
rect 17092 27316 17098 27328
rect 17770 27316 17776 27328
rect 17092 27288 17776 27316
rect 17092 27276 17098 27288
rect 17770 27276 17776 27288
rect 17828 27276 17834 27328
rect 18230 27276 18236 27328
rect 18288 27316 18294 27328
rect 18325 27319 18383 27325
rect 18325 27316 18337 27319
rect 18288 27288 18337 27316
rect 18288 27276 18294 27288
rect 18325 27285 18337 27288
rect 18371 27285 18383 27319
rect 18325 27279 18383 27285
rect 23385 27319 23443 27325
rect 23385 27285 23397 27319
rect 23431 27316 23443 27319
rect 23474 27316 23480 27328
rect 23431 27288 23480 27316
rect 23431 27285 23443 27288
rect 23385 27279 23443 27285
rect 23474 27276 23480 27288
rect 23532 27276 23538 27328
rect 31110 27276 31116 27328
rect 31168 27276 31174 27328
rect 32217 27319 32275 27325
rect 32217 27285 32229 27319
rect 32263 27316 32275 27319
rect 32858 27316 32864 27328
rect 32263 27288 32864 27316
rect 32263 27285 32275 27288
rect 32217 27279 32275 27285
rect 32858 27276 32864 27288
rect 32916 27276 32922 27328
rect 1104 27226 48852 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 48852 27226
rect 1104 27152 48852 27174
rect 8507 27115 8565 27121
rect 8507 27081 8519 27115
rect 8553 27112 8565 27115
rect 8754 27112 8760 27124
rect 8553 27084 8760 27112
rect 8553 27081 8565 27084
rect 8507 27075 8565 27081
rect 8754 27072 8760 27084
rect 8812 27072 8818 27124
rect 11882 27072 11888 27124
rect 11940 27112 11946 27124
rect 12069 27115 12127 27121
rect 12069 27112 12081 27115
rect 11940 27084 12081 27112
rect 11940 27072 11946 27084
rect 12069 27081 12081 27084
rect 12115 27081 12127 27115
rect 12069 27075 12127 27081
rect 12802 27072 12808 27124
rect 12860 27112 12866 27124
rect 12860 27084 22094 27112
rect 12860 27072 12866 27084
rect 1946 27044 1952 27056
rect 1907 27016 1952 27044
rect 1946 27004 1952 27016
rect 2004 27004 2010 27056
rect 8297 27047 8355 27053
rect 8297 27013 8309 27047
rect 8343 27044 8355 27047
rect 8386 27044 8392 27056
rect 8343 27016 8392 27044
rect 8343 27013 8355 27016
rect 8297 27007 8355 27013
rect 8386 27004 8392 27016
rect 8444 27004 8450 27056
rect 9493 27047 9551 27053
rect 9493 27013 9505 27047
rect 9539 27044 9551 27047
rect 10318 27044 10324 27056
rect 9539 27016 10324 27044
rect 9539 27013 9551 27016
rect 9493 27007 9551 27013
rect 10318 27004 10324 27016
rect 10376 27044 10382 27056
rect 11974 27044 11980 27056
rect 10376 27016 11980 27044
rect 10376 27004 10382 27016
rect 11974 27004 11980 27016
rect 12032 27004 12038 27056
rect 12986 27004 12992 27056
rect 13044 27044 13050 27056
rect 13044 27016 15608 27044
rect 13044 27004 13050 27016
rect 1762 26976 1768 26988
rect 1723 26948 1768 26976
rect 1762 26936 1768 26948
rect 1820 26936 1826 26988
rect 9125 26979 9183 26985
rect 9125 26945 9137 26979
rect 9171 26976 9183 26979
rect 9858 26976 9864 26988
rect 9171 26948 9864 26976
rect 9171 26945 9183 26948
rect 9125 26939 9183 26945
rect 9858 26936 9864 26948
rect 9916 26936 9922 26988
rect 10410 26976 10416 26988
rect 10371 26948 10416 26976
rect 10410 26936 10416 26948
rect 10468 26936 10474 26988
rect 14016 26985 14044 27016
rect 14001 26979 14059 26985
rect 14001 26945 14013 26979
rect 14047 26945 14059 26979
rect 14001 26939 14059 26945
rect 14090 26979 14148 26985
rect 14090 26945 14102 26979
rect 14136 26945 14148 26979
rect 14090 26939 14148 26945
rect 2774 26868 2780 26920
rect 2832 26908 2838 26920
rect 9674 26908 9680 26920
rect 2832 26880 2877 26908
rect 9416 26880 9680 26908
rect 2832 26868 2838 26880
rect 8294 26800 8300 26852
rect 8352 26840 8358 26852
rect 8665 26843 8723 26849
rect 8665 26840 8677 26843
rect 8352 26812 8677 26840
rect 8352 26800 8358 26812
rect 8665 26809 8677 26812
rect 8711 26809 8723 26843
rect 8665 26803 8723 26809
rect 8481 26775 8539 26781
rect 8481 26741 8493 26775
rect 8527 26772 8539 26775
rect 9416 26772 9444 26880
rect 9674 26868 9680 26880
rect 9732 26868 9738 26920
rect 10134 26908 10140 26920
rect 10095 26880 10140 26908
rect 10134 26868 10140 26880
rect 10192 26868 10198 26920
rect 10686 26840 10692 26852
rect 9508 26812 10692 26840
rect 9508 26781 9536 26812
rect 10686 26800 10692 26812
rect 10744 26800 10750 26852
rect 13354 26800 13360 26852
rect 13412 26840 13418 26852
rect 14108 26840 14136 26939
rect 14182 26936 14188 26988
rect 14240 26976 14246 26988
rect 14366 26976 14372 26988
rect 14240 26948 14285 26976
rect 14327 26948 14372 26976
rect 14240 26936 14246 26948
rect 14366 26936 14372 26948
rect 14424 26936 14430 26988
rect 15580 26985 15608 27016
rect 17770 27004 17776 27056
rect 17828 27044 17834 27056
rect 19061 27047 19119 27053
rect 17828 27016 18181 27044
rect 17828 27004 17834 27016
rect 15565 26979 15623 26985
rect 15565 26945 15577 26979
rect 15611 26976 15623 26979
rect 16899 26979 16957 26985
rect 16899 26976 16911 26979
rect 15611 26948 16911 26976
rect 15611 26945 15623 26948
rect 15565 26939 15623 26945
rect 16899 26945 16911 26948
rect 16945 26945 16957 26979
rect 16899 26939 16957 26945
rect 17014 26936 17020 26988
rect 17072 26985 17078 26988
rect 17072 26979 17092 26985
rect 17080 26945 17092 26979
rect 17072 26939 17092 26945
rect 17150 26979 17208 26985
rect 17150 26945 17162 26979
rect 17196 26976 17208 26979
rect 17196 26948 17264 26976
rect 17196 26945 17208 26948
rect 17150 26939 17208 26945
rect 17072 26936 17078 26939
rect 15289 26911 15347 26917
rect 15289 26877 15301 26911
rect 15335 26908 15347 26911
rect 15470 26908 15476 26920
rect 15335 26880 15476 26908
rect 15335 26877 15347 26880
rect 15289 26871 15347 26877
rect 15470 26868 15476 26880
rect 15528 26868 15534 26920
rect 17236 26852 17264 26948
rect 17310 26936 17316 26988
rect 17368 26976 17374 26988
rect 17368 26948 17413 26976
rect 17368 26936 17374 26948
rect 17586 26936 17592 26988
rect 17644 26976 17650 26988
rect 18153 26985 18181 27016
rect 19061 27013 19073 27047
rect 19107 27044 19119 27047
rect 20530 27044 20536 27056
rect 19107 27016 20536 27044
rect 19107 27013 19119 27016
rect 19061 27007 19119 27013
rect 20530 27004 20536 27016
rect 20588 27004 20594 27056
rect 18049 26979 18107 26985
rect 17893 26976 18061 26979
rect 17644 26951 18061 26976
rect 17644 26948 17921 26951
rect 17972 26948 18021 26951
rect 17644 26936 17650 26948
rect 18049 26945 18061 26951
rect 18095 26945 18107 26979
rect 18049 26939 18107 26945
rect 18141 26979 18199 26985
rect 18141 26945 18153 26979
rect 18187 26945 18199 26979
rect 18141 26939 18199 26945
rect 18230 26936 18236 26988
rect 18288 26976 18294 26988
rect 18417 26979 18475 26985
rect 18288 26948 18333 26976
rect 18288 26936 18294 26948
rect 18417 26945 18429 26979
rect 18463 26976 18475 26979
rect 18506 26976 18512 26988
rect 18463 26948 18512 26976
rect 18463 26945 18475 26948
rect 18417 26939 18475 26945
rect 18506 26936 18512 26948
rect 18564 26936 18570 26988
rect 18877 26979 18935 26985
rect 18877 26945 18889 26979
rect 18923 26945 18935 26979
rect 18877 26939 18935 26945
rect 13412 26812 14136 26840
rect 13412 26800 13418 26812
rect 17218 26800 17224 26852
rect 17276 26800 17282 26852
rect 17328 26840 17356 26936
rect 17862 26868 17868 26920
rect 17920 26908 17926 26920
rect 18892 26908 18920 26939
rect 20162 26936 20168 26988
rect 20220 26976 20226 26988
rect 20257 26979 20315 26985
rect 20257 26976 20269 26979
rect 20220 26948 20269 26976
rect 20220 26936 20226 26948
rect 20257 26945 20269 26948
rect 20303 26945 20315 26979
rect 20257 26939 20315 26945
rect 17920 26880 18920 26908
rect 20533 26911 20591 26917
rect 17920 26868 17926 26880
rect 20533 26877 20545 26911
rect 20579 26877 20591 26911
rect 20533 26871 20591 26877
rect 18506 26840 18512 26852
rect 17328 26812 18512 26840
rect 18506 26800 18512 26812
rect 18564 26800 18570 26852
rect 20254 26800 20260 26852
rect 20312 26840 20318 26852
rect 20548 26840 20576 26871
rect 20312 26812 20576 26840
rect 22066 26840 22094 27084
rect 22278 27072 22284 27124
rect 22336 27112 22342 27124
rect 23385 27115 23443 27121
rect 23385 27112 23397 27115
rect 22336 27084 23397 27112
rect 22336 27072 22342 27084
rect 23385 27081 23397 27084
rect 23431 27081 23443 27115
rect 23385 27075 23443 27081
rect 23934 27072 23940 27124
rect 23992 27112 23998 27124
rect 24210 27112 24216 27124
rect 23992 27084 24216 27112
rect 23992 27072 23998 27084
rect 24210 27072 24216 27084
rect 24268 27072 24274 27124
rect 25038 27112 25044 27124
rect 24964 27084 25044 27112
rect 25038 27072 25044 27084
rect 25096 27112 25102 27124
rect 27706 27112 27712 27124
rect 25096 27084 27712 27112
rect 25096 27072 25102 27084
rect 27706 27072 27712 27084
rect 27764 27112 27770 27124
rect 31110 27112 31116 27124
rect 27764 27084 31116 27112
rect 27764 27072 27770 27084
rect 31110 27072 31116 27084
rect 31168 27072 31174 27124
rect 23017 27047 23075 27053
rect 23017 27013 23029 27047
rect 23063 27044 23075 27047
rect 24118 27044 24124 27056
rect 23063 27016 24124 27044
rect 23063 27013 23075 27016
rect 23017 27007 23075 27013
rect 24118 27004 24124 27016
rect 24176 27004 24182 27056
rect 23201 26979 23259 26985
rect 23201 26945 23213 26979
rect 23247 26945 23259 26979
rect 23201 26939 23259 26945
rect 23216 26908 23244 26939
rect 23842 26936 23848 26988
rect 23900 26976 23906 26988
rect 24210 26976 24216 26988
rect 23900 26948 24216 26976
rect 23900 26936 23906 26948
rect 24210 26936 24216 26948
rect 24268 26936 24274 26988
rect 24762 26936 24768 26988
rect 24820 26976 24826 26988
rect 25069 26985 25097 27072
rect 26421 27047 26479 27053
rect 26421 27044 26433 27047
rect 25240 27016 26433 27044
rect 25154 26985 25212 26991
rect 24949 26979 25007 26985
rect 24949 26976 24961 26979
rect 24820 26948 24961 26976
rect 24820 26936 24826 26948
rect 24949 26945 24961 26948
rect 24995 26945 25007 26979
rect 24949 26939 25007 26945
rect 25041 26979 25099 26985
rect 25041 26945 25053 26979
rect 25087 26945 25099 26979
rect 25154 26951 25166 26985
rect 25200 26982 25212 26985
rect 25240 26982 25268 27016
rect 26421 27013 26433 27016
rect 26467 27013 26479 27047
rect 26421 27007 26479 27013
rect 27724 26991 27752 27072
rect 28629 27047 28687 27053
rect 28629 27013 28641 27047
rect 28675 27044 28687 27047
rect 28902 27044 28908 27056
rect 28675 27016 28908 27044
rect 28675 27013 28687 27016
rect 28629 27007 28687 27013
rect 28902 27004 28908 27016
rect 28960 27004 28966 27056
rect 32398 27004 32404 27056
rect 32456 27044 32462 27056
rect 34885 27047 34943 27053
rect 32456 27016 32996 27044
rect 32456 27004 32462 27016
rect 25200 26954 25268 26982
rect 25317 26982 25375 26985
rect 25317 26979 25452 26982
rect 25200 26951 25212 26954
rect 25154 26945 25212 26951
rect 25317 26945 25329 26979
rect 25363 26976 25452 26979
rect 25590 26976 25596 26988
rect 25363 26954 25596 26976
rect 25363 26945 25375 26954
rect 25424 26948 25596 26954
rect 25041 26939 25099 26945
rect 25317 26939 25375 26945
rect 25590 26936 25596 26948
rect 25648 26936 25654 26988
rect 26050 26976 26056 26988
rect 26011 26948 26056 26976
rect 26050 26936 26056 26948
rect 26108 26936 26114 26988
rect 26237 26979 26295 26985
rect 26237 26945 26249 26979
rect 26283 26976 26295 26979
rect 26510 26976 26516 26988
rect 26283 26948 26516 26976
rect 26283 26945 26295 26948
rect 26237 26939 26295 26945
rect 26510 26936 26516 26948
rect 26568 26936 26574 26988
rect 27706 26985 27764 26991
rect 27617 26979 27675 26985
rect 27617 26976 27629 26979
rect 26620 26948 27629 26976
rect 23474 26908 23480 26920
rect 23216 26880 23480 26908
rect 23474 26868 23480 26880
rect 23532 26908 23538 26920
rect 26620 26908 26648 26948
rect 27617 26945 27629 26948
rect 27663 26945 27675 26979
rect 27706 26951 27718 26985
rect 27752 26951 27764 26985
rect 27706 26945 27764 26951
rect 27801 26979 27859 26985
rect 27801 26945 27813 26979
rect 27847 26945 27859 26979
rect 27982 26976 27988 26988
rect 27943 26948 27988 26976
rect 27617 26939 27675 26945
rect 27801 26939 27859 26945
rect 23532 26880 26648 26908
rect 27816 26908 27844 26939
rect 27982 26936 27988 26948
rect 28040 26936 28046 26988
rect 28445 26979 28503 26985
rect 28445 26945 28457 26979
rect 28491 26976 28503 26979
rect 28534 26976 28540 26988
rect 28491 26948 28540 26976
rect 28491 26945 28503 26948
rect 28445 26939 28503 26945
rect 28534 26936 28540 26948
rect 28592 26936 28598 26988
rect 31202 26976 31208 26988
rect 31163 26948 31208 26976
rect 31202 26936 31208 26948
rect 31260 26936 31266 26988
rect 32858 26976 32864 26988
rect 32819 26948 32864 26976
rect 32858 26936 32864 26948
rect 32916 26936 32922 26988
rect 32968 26985 32996 27016
rect 34885 27013 34897 27047
rect 34931 27044 34943 27047
rect 36446 27044 36452 27056
rect 34931 27016 36452 27044
rect 34931 27013 34943 27016
rect 34885 27007 34943 27013
rect 36446 27004 36452 27016
rect 36504 27004 36510 27056
rect 32953 26979 33011 26985
rect 32953 26945 32965 26979
rect 32999 26945 33011 26979
rect 32953 26939 33011 26945
rect 33045 26979 33103 26985
rect 33045 26945 33057 26979
rect 33091 26945 33103 26979
rect 33226 26976 33232 26988
rect 33187 26948 33232 26976
rect 33045 26939 33103 26945
rect 28813 26911 28871 26917
rect 28813 26908 28825 26911
rect 27816 26880 28825 26908
rect 23532 26868 23538 26880
rect 28813 26877 28825 26880
rect 28859 26877 28871 26911
rect 31754 26908 31760 26920
rect 28813 26871 28871 26877
rect 31726 26868 31760 26908
rect 31812 26868 31818 26920
rect 33060 26908 33088 26939
rect 33226 26936 33232 26948
rect 33284 26936 33290 26988
rect 35069 26979 35127 26985
rect 35069 26945 35081 26979
rect 35115 26976 35127 26979
rect 35710 26976 35716 26988
rect 35115 26948 35716 26976
rect 35115 26945 35127 26948
rect 35069 26939 35127 26945
rect 35710 26936 35716 26948
rect 35768 26936 35774 26988
rect 35342 26908 35348 26920
rect 33060 26880 35348 26908
rect 35342 26868 35348 26880
rect 35400 26868 35406 26920
rect 31726 26840 31754 26868
rect 22066 26812 31754 26840
rect 20312 26800 20318 26812
rect 8527 26744 9444 26772
rect 9493 26775 9551 26781
rect 8527 26741 8539 26744
rect 8481 26735 8539 26741
rect 9493 26741 9505 26775
rect 9539 26741 9551 26775
rect 9674 26772 9680 26784
rect 9635 26744 9680 26772
rect 9493 26735 9551 26741
rect 9674 26732 9680 26744
rect 9732 26732 9738 26784
rect 13725 26775 13783 26781
rect 13725 26741 13737 26775
rect 13771 26772 13783 26775
rect 14458 26772 14464 26784
rect 13771 26744 14464 26772
rect 13771 26741 13783 26744
rect 13725 26735 13783 26741
rect 14458 26732 14464 26744
rect 14516 26732 14522 26784
rect 16666 26772 16672 26784
rect 16627 26744 16672 26772
rect 16666 26732 16672 26744
rect 16724 26732 16730 26784
rect 17773 26775 17831 26781
rect 17773 26741 17785 26775
rect 17819 26772 17831 26775
rect 18230 26772 18236 26784
rect 17819 26744 18236 26772
rect 17819 26741 17831 26744
rect 17773 26735 17831 26741
rect 18230 26732 18236 26744
rect 18288 26732 18294 26784
rect 18322 26732 18328 26784
rect 18380 26772 18386 26784
rect 19245 26775 19303 26781
rect 19245 26772 19257 26775
rect 18380 26744 19257 26772
rect 18380 26732 18386 26744
rect 19245 26741 19257 26744
rect 19291 26741 19303 26775
rect 24670 26772 24676 26784
rect 24631 26744 24676 26772
rect 19245 26735 19303 26741
rect 24670 26732 24676 26744
rect 24728 26732 24734 26784
rect 25038 26732 25044 26784
rect 25096 26772 25102 26784
rect 25590 26772 25596 26784
rect 25096 26744 25596 26772
rect 25096 26732 25102 26744
rect 25590 26732 25596 26744
rect 25648 26732 25654 26784
rect 27341 26775 27399 26781
rect 27341 26741 27353 26775
rect 27387 26772 27399 26775
rect 27982 26772 27988 26784
rect 27387 26744 27988 26772
rect 27387 26741 27399 26744
rect 27341 26735 27399 26741
rect 27982 26732 27988 26744
rect 28040 26732 28046 26784
rect 30558 26732 30564 26784
rect 30616 26772 30622 26784
rect 31297 26775 31355 26781
rect 31297 26772 31309 26775
rect 30616 26744 31309 26772
rect 30616 26732 30622 26744
rect 31297 26741 31309 26744
rect 31343 26741 31355 26775
rect 31297 26735 31355 26741
rect 32585 26775 32643 26781
rect 32585 26741 32597 26775
rect 32631 26772 32643 26775
rect 32858 26772 32864 26784
rect 32631 26744 32864 26772
rect 32631 26741 32643 26744
rect 32585 26735 32643 26741
rect 32858 26732 32864 26744
rect 32916 26732 32922 26784
rect 35253 26775 35311 26781
rect 35253 26741 35265 26775
rect 35299 26772 35311 26775
rect 35618 26772 35624 26784
rect 35299 26744 35624 26772
rect 35299 26741 35311 26744
rect 35253 26735 35311 26741
rect 35618 26732 35624 26744
rect 35676 26732 35682 26784
rect 1104 26682 48852 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 48852 26682
rect 1104 26608 48852 26630
rect 11422 26568 11428 26580
rect 11383 26540 11428 26568
rect 11422 26528 11428 26540
rect 11480 26528 11486 26580
rect 13449 26571 13507 26577
rect 13449 26537 13461 26571
rect 13495 26568 13507 26571
rect 14366 26568 14372 26580
rect 13495 26540 14372 26568
rect 13495 26537 13507 26540
rect 13449 26531 13507 26537
rect 14366 26528 14372 26540
rect 14424 26528 14430 26580
rect 17126 26568 17132 26580
rect 16776 26540 17132 26568
rect 1302 26460 1308 26512
rect 1360 26500 1366 26512
rect 1578 26500 1584 26512
rect 1360 26472 1584 26500
rect 1360 26460 1366 26472
rect 1578 26460 1584 26472
rect 1636 26460 1642 26512
rect 10134 26460 10140 26512
rect 10192 26500 10198 26512
rect 10321 26503 10379 26509
rect 10321 26500 10333 26503
rect 10192 26472 10333 26500
rect 10192 26460 10198 26472
rect 10321 26469 10333 26472
rect 10367 26500 10379 26503
rect 10778 26500 10784 26512
rect 10367 26472 10784 26500
rect 10367 26469 10379 26472
rect 10321 26463 10379 26469
rect 10778 26460 10784 26472
rect 10836 26460 10842 26512
rect 10870 26460 10876 26512
rect 10928 26500 10934 26512
rect 11609 26503 11667 26509
rect 11609 26500 11621 26503
rect 10928 26472 11621 26500
rect 10928 26460 10934 26472
rect 11609 26469 11621 26472
rect 11655 26469 11667 26503
rect 11609 26463 11667 26469
rect 1394 26432 1400 26444
rect 1355 26404 1400 26432
rect 1394 26392 1400 26404
rect 1452 26392 1458 26444
rect 2774 26392 2780 26444
rect 2832 26432 2838 26444
rect 16776 26441 16804 26540
rect 17126 26528 17132 26540
rect 17184 26528 17190 26580
rect 26050 26528 26056 26580
rect 26108 26568 26114 26580
rect 26697 26571 26755 26577
rect 26697 26568 26709 26571
rect 26108 26540 26709 26568
rect 26108 26528 26114 26540
rect 26697 26537 26709 26540
rect 26743 26537 26755 26571
rect 26697 26531 26755 26537
rect 28534 26528 28540 26580
rect 28592 26568 28598 26580
rect 29549 26571 29607 26577
rect 29549 26568 29561 26571
rect 28592 26540 29561 26568
rect 28592 26528 28598 26540
rect 29549 26537 29561 26540
rect 29595 26537 29607 26571
rect 29549 26531 29607 26537
rect 31202 26528 31208 26580
rect 31260 26568 31266 26580
rect 31757 26571 31815 26577
rect 31757 26568 31769 26571
rect 31260 26540 31769 26568
rect 31260 26528 31266 26540
rect 31757 26537 31769 26540
rect 31803 26568 31815 26571
rect 37274 26568 37280 26580
rect 31803 26540 37280 26568
rect 31803 26537 31815 26540
rect 31757 26531 31815 26537
rect 37274 26528 37280 26540
rect 37332 26528 37338 26580
rect 20530 26460 20536 26512
rect 20588 26500 20594 26512
rect 20625 26503 20683 26509
rect 20625 26500 20637 26503
rect 20588 26472 20637 26500
rect 20588 26460 20594 26472
rect 20625 26469 20637 26472
rect 20671 26469 20683 26503
rect 28994 26500 29000 26512
rect 20625 26463 20683 26469
rect 27356 26472 29000 26500
rect 16761 26435 16819 26441
rect 2832 26404 2877 26432
rect 2832 26392 2838 26404
rect 16761 26401 16773 26435
rect 16807 26401 16819 26435
rect 16761 26395 16819 26401
rect 24486 26392 24492 26444
rect 24544 26432 24550 26444
rect 24857 26435 24915 26441
rect 24857 26432 24869 26435
rect 24544 26404 24869 26432
rect 24544 26392 24550 26404
rect 24857 26401 24869 26404
rect 24903 26401 24915 26435
rect 27154 26432 27160 26444
rect 27115 26404 27160 26432
rect 24857 26395 24915 26401
rect 27154 26392 27160 26404
rect 27212 26392 27218 26444
rect 27356 26441 27384 26472
rect 28994 26460 29000 26472
rect 29052 26500 29058 26512
rect 34149 26503 34207 26509
rect 29052 26472 30144 26500
rect 29052 26460 29058 26472
rect 27341 26435 27399 26441
rect 27341 26401 27353 26435
rect 27387 26401 27399 26435
rect 30006 26432 30012 26444
rect 29967 26404 30012 26432
rect 27341 26395 27399 26401
rect 30006 26392 30012 26404
rect 30064 26392 30070 26444
rect 30116 26441 30144 26472
rect 34149 26469 34161 26503
rect 34195 26469 34207 26503
rect 34149 26463 34207 26469
rect 30101 26435 30159 26441
rect 30101 26401 30113 26435
rect 30147 26432 30159 26435
rect 30147 26404 30972 26432
rect 30147 26401 30159 26404
rect 30101 26395 30159 26401
rect 7742 26324 7748 26376
rect 7800 26364 7806 26376
rect 8941 26367 8999 26373
rect 8941 26364 8953 26367
rect 7800 26336 8953 26364
rect 7800 26324 7806 26336
rect 8941 26333 8953 26336
rect 8987 26333 8999 26367
rect 12158 26364 12164 26376
rect 12119 26336 12164 26364
rect 8941 26327 8999 26333
rect 12158 26324 12164 26336
rect 12216 26324 12222 26376
rect 12526 26324 12532 26376
rect 12584 26324 12590 26376
rect 13354 26364 13360 26376
rect 13315 26336 13360 26364
rect 13354 26324 13360 26336
rect 13412 26324 13418 26376
rect 13541 26367 13599 26373
rect 13541 26333 13553 26367
rect 13587 26333 13599 26367
rect 13541 26327 13599 26333
rect 14185 26367 14243 26373
rect 14185 26333 14197 26367
rect 14231 26364 14243 26367
rect 14274 26364 14280 26376
rect 14231 26336 14280 26364
rect 14231 26333 14243 26336
rect 14185 26327 14243 26333
rect 1578 26296 1584 26308
rect 1539 26268 1584 26296
rect 1578 26256 1584 26268
rect 1636 26256 1642 26308
rect 9214 26305 9220 26308
rect 9208 26259 9220 26305
rect 9272 26296 9278 26308
rect 11241 26299 11299 26305
rect 9272 26268 9308 26296
rect 9214 26256 9220 26259
rect 9272 26256 9278 26268
rect 11241 26265 11253 26299
rect 11287 26265 11299 26299
rect 11241 26259 11299 26265
rect 11457 26299 11515 26305
rect 11457 26265 11469 26299
rect 11503 26296 11515 26299
rect 11790 26296 11796 26308
rect 11503 26268 11796 26296
rect 11503 26265 11515 26268
rect 11457 26259 11515 26265
rect 10962 26188 10968 26240
rect 11020 26228 11026 26240
rect 11256 26228 11284 26259
rect 11790 26256 11796 26268
rect 11848 26296 11854 26308
rect 12176 26296 12204 26324
rect 11848 26268 12204 26296
rect 12345 26299 12403 26305
rect 11848 26256 11854 26268
rect 12345 26265 12357 26299
rect 12391 26296 12403 26299
rect 12544 26296 12572 26324
rect 13170 26296 13176 26308
rect 12391 26268 13176 26296
rect 12391 26265 12403 26268
rect 12345 26259 12403 26265
rect 13170 26256 13176 26268
rect 13228 26256 13234 26308
rect 13556 26296 13584 26327
rect 14274 26324 14280 26336
rect 14332 26324 14338 26376
rect 14458 26373 14464 26376
rect 14452 26364 14464 26373
rect 14419 26336 14464 26364
rect 14452 26327 14464 26336
rect 14458 26324 14464 26327
rect 14516 26324 14522 26376
rect 16666 26324 16672 26376
rect 16724 26364 16730 26376
rect 17017 26367 17075 26373
rect 17017 26364 17029 26367
rect 16724 26336 17029 26364
rect 16724 26324 16730 26336
rect 17017 26333 17029 26336
rect 17063 26333 17075 26367
rect 17017 26327 17075 26333
rect 19245 26367 19303 26373
rect 19245 26333 19257 26367
rect 19291 26364 19303 26367
rect 20070 26364 20076 26376
rect 19291 26336 20076 26364
rect 19291 26333 19303 26336
rect 19245 26327 19303 26333
rect 20070 26324 20076 26336
rect 20128 26324 20134 26376
rect 24670 26324 24676 26376
rect 24728 26364 24734 26376
rect 30944 26373 30972 26404
rect 33962 26392 33968 26444
rect 34020 26432 34026 26444
rect 34164 26432 34192 26463
rect 37001 26435 37059 26441
rect 37001 26432 37013 26435
rect 34020 26404 37013 26432
rect 34020 26392 34026 26404
rect 37001 26401 37013 26404
rect 37047 26401 37059 26435
rect 37001 26395 37059 26401
rect 25113 26367 25171 26373
rect 25113 26364 25125 26367
rect 24728 26336 25125 26364
rect 24728 26324 24734 26336
rect 25113 26333 25125 26336
rect 25159 26333 25171 26367
rect 25113 26327 25171 26333
rect 30929 26367 30987 26373
rect 30929 26333 30941 26367
rect 30975 26333 30987 26367
rect 30929 26327 30987 26333
rect 31386 26324 31392 26376
rect 31444 26364 31450 26376
rect 31573 26367 31631 26373
rect 31573 26364 31585 26367
rect 31444 26336 31585 26364
rect 31444 26324 31450 26336
rect 31573 26333 31585 26336
rect 31619 26333 31631 26367
rect 32766 26364 32772 26376
rect 32727 26336 32772 26364
rect 31573 26327 31631 26333
rect 32766 26324 32772 26336
rect 32824 26324 32830 26376
rect 32858 26324 32864 26376
rect 32916 26364 32922 26376
rect 33025 26367 33083 26373
rect 33025 26364 33037 26367
rect 32916 26336 33037 26364
rect 32916 26324 32922 26336
rect 33025 26333 33037 26336
rect 33071 26333 33083 26367
rect 33025 26327 33083 26333
rect 34698 26324 34704 26376
rect 34756 26364 34762 26376
rect 34977 26367 35035 26373
rect 34977 26364 34989 26367
rect 34756 26336 34989 26364
rect 34756 26324 34762 26336
rect 34977 26333 34989 26336
rect 35023 26333 35035 26367
rect 34977 26327 35035 26333
rect 35069 26367 35127 26373
rect 35069 26333 35081 26367
rect 35115 26333 35127 26367
rect 35069 26327 35127 26333
rect 35161 26367 35219 26373
rect 35161 26333 35173 26367
rect 35207 26364 35219 26367
rect 35250 26364 35256 26376
rect 35207 26336 35256 26364
rect 35207 26333 35219 26336
rect 35161 26327 35219 26333
rect 15286 26296 15292 26308
rect 13556 26268 15292 26296
rect 15286 26256 15292 26268
rect 15344 26256 15350 26308
rect 17954 26256 17960 26308
rect 18012 26296 18018 26308
rect 19490 26299 19548 26305
rect 19490 26296 19502 26299
rect 18012 26268 19502 26296
rect 18012 26256 18018 26268
rect 19490 26265 19502 26268
rect 19536 26265 19548 26299
rect 31110 26296 31116 26308
rect 31071 26268 31116 26296
rect 19490 26259 19548 26265
rect 31110 26256 31116 26268
rect 31168 26256 31174 26308
rect 33778 26256 33784 26308
rect 33836 26296 33842 26308
rect 35084 26296 35112 26327
rect 35250 26324 35256 26336
rect 35308 26324 35314 26376
rect 35345 26367 35403 26373
rect 35345 26333 35357 26367
rect 35391 26364 35403 26367
rect 35618 26364 35624 26376
rect 35391 26336 35624 26364
rect 35391 26333 35403 26336
rect 35345 26327 35403 26333
rect 35618 26324 35624 26336
rect 35676 26324 35682 26376
rect 33836 26268 35112 26296
rect 37185 26299 37243 26305
rect 33836 26256 33842 26268
rect 37185 26265 37197 26299
rect 37231 26296 37243 26299
rect 37366 26296 37372 26308
rect 37231 26268 37372 26296
rect 37231 26265 37243 26268
rect 37185 26259 37243 26265
rect 37366 26256 37372 26268
rect 37424 26256 37430 26308
rect 38841 26299 38899 26305
rect 38841 26265 38853 26299
rect 38887 26296 38899 26299
rect 46014 26296 46020 26308
rect 38887 26268 46020 26296
rect 38887 26265 38899 26268
rect 38841 26259 38899 26265
rect 46014 26256 46020 26268
rect 46072 26256 46078 26308
rect 47946 26296 47952 26308
rect 47907 26268 47952 26296
rect 47946 26256 47952 26268
rect 48004 26256 48010 26308
rect 48130 26296 48136 26308
rect 48091 26268 48136 26296
rect 48130 26256 48136 26268
rect 48188 26256 48194 26308
rect 12250 26228 12256 26240
rect 11020 26200 12256 26228
rect 11020 26188 11026 26200
rect 12250 26188 12256 26200
rect 12308 26188 12314 26240
rect 12526 26228 12532 26240
rect 12487 26200 12532 26228
rect 12526 26188 12532 26200
rect 12584 26188 12590 26240
rect 15562 26228 15568 26240
rect 15523 26200 15568 26228
rect 15562 26188 15568 26200
rect 15620 26188 15626 26240
rect 18046 26188 18052 26240
rect 18104 26228 18110 26240
rect 18141 26231 18199 26237
rect 18141 26228 18153 26231
rect 18104 26200 18153 26228
rect 18104 26188 18110 26200
rect 18141 26197 18153 26200
rect 18187 26228 18199 26231
rect 18782 26228 18788 26240
rect 18187 26200 18788 26228
rect 18187 26197 18199 26200
rect 18141 26191 18199 26197
rect 18782 26188 18788 26200
rect 18840 26188 18846 26240
rect 22278 26188 22284 26240
rect 22336 26228 22342 26240
rect 23934 26228 23940 26240
rect 22336 26200 23940 26228
rect 22336 26188 22342 26200
rect 23934 26188 23940 26200
rect 23992 26188 23998 26240
rect 26234 26228 26240 26240
rect 26147 26200 26240 26228
rect 26234 26188 26240 26200
rect 26292 26228 26298 26240
rect 27065 26231 27123 26237
rect 27065 26228 27077 26231
rect 26292 26200 27077 26228
rect 26292 26188 26298 26200
rect 27065 26197 27077 26200
rect 27111 26197 27123 26231
rect 27065 26191 27123 26197
rect 29270 26188 29276 26240
rect 29328 26228 29334 26240
rect 29917 26231 29975 26237
rect 29917 26228 29929 26231
rect 29328 26200 29929 26228
rect 29328 26188 29334 26200
rect 29917 26197 29929 26200
rect 29963 26197 29975 26231
rect 34698 26228 34704 26240
rect 34659 26200 34704 26228
rect 29917 26191 29975 26197
rect 34698 26188 34704 26200
rect 34756 26188 34762 26240
rect 36538 26188 36544 26240
rect 36596 26228 36602 26240
rect 46566 26228 46572 26240
rect 36596 26200 46572 26228
rect 36596 26188 36602 26200
rect 46566 26188 46572 26200
rect 46624 26188 46630 26240
rect 1104 26138 48852 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 48852 26138
rect 1104 26064 48852 26086
rect 1578 25984 1584 26036
rect 1636 26024 1642 26036
rect 2225 26027 2283 26033
rect 2225 26024 2237 26027
rect 1636 25996 2237 26024
rect 1636 25984 1642 25996
rect 2225 25993 2237 25996
rect 2271 25993 2283 26027
rect 2225 25987 2283 25993
rect 9125 26027 9183 26033
rect 9125 25993 9137 26027
rect 9171 26024 9183 26027
rect 9214 26024 9220 26036
rect 9171 25996 9220 26024
rect 9171 25993 9183 25996
rect 9125 25987 9183 25993
rect 9214 25984 9220 25996
rect 9272 25984 9278 26036
rect 10318 26024 10324 26036
rect 10279 25996 10324 26024
rect 10318 25984 10324 25996
rect 10376 25984 10382 26036
rect 12250 25984 12256 26036
rect 12308 26024 12314 26036
rect 12710 26024 12716 26036
rect 12308 25996 12716 26024
rect 12308 25984 12314 25996
rect 12710 25984 12716 25996
rect 12768 26024 12774 26036
rect 13722 26024 13728 26036
rect 12768 25996 13728 26024
rect 12768 25984 12774 25996
rect 13722 25984 13728 25996
rect 13780 25984 13786 26036
rect 15286 26024 15292 26036
rect 15247 25996 15292 26024
rect 15286 25984 15292 25996
rect 15344 25984 15350 26036
rect 17218 25984 17224 26036
rect 17276 26024 17282 26036
rect 17589 26027 17647 26033
rect 17589 26024 17601 26027
rect 17276 25996 17601 26024
rect 17276 25984 17282 25996
rect 17589 25993 17601 25996
rect 17635 25993 17647 26027
rect 17589 25987 17647 25993
rect 19426 25984 19432 26036
rect 19484 26024 19490 26036
rect 19521 26027 19579 26033
rect 19521 26024 19533 26027
rect 19484 25996 19533 26024
rect 19484 25984 19490 25996
rect 19521 25993 19533 25996
rect 19567 25993 19579 26027
rect 19521 25987 19579 25993
rect 20162 25984 20168 26036
rect 20220 26024 20226 26036
rect 20257 26027 20315 26033
rect 20257 26024 20269 26027
rect 20220 25996 20269 26024
rect 20220 25984 20226 25996
rect 20257 25993 20269 25996
rect 20303 25993 20315 26027
rect 20257 25987 20315 25993
rect 21818 25984 21824 26036
rect 21876 26024 21882 26036
rect 25866 26024 25872 26036
rect 21876 25996 25872 26024
rect 21876 25984 21882 25996
rect 25866 25984 25872 25996
rect 25924 25984 25930 26036
rect 27341 26027 27399 26033
rect 27341 25993 27353 26027
rect 27387 26024 27399 26027
rect 28258 26024 28264 26036
rect 27387 25996 28264 26024
rect 27387 25993 27399 25996
rect 27341 25987 27399 25993
rect 28258 25984 28264 25996
rect 28316 25984 28322 26036
rect 29270 26024 29276 26036
rect 29231 25996 29276 26024
rect 29270 25984 29276 25996
rect 29328 25984 29334 26036
rect 32950 26024 32956 26036
rect 29380 25996 32956 26024
rect 11974 25916 11980 25968
rect 12032 25956 12038 25968
rect 12069 25959 12127 25965
rect 12069 25956 12081 25959
rect 12032 25928 12081 25956
rect 12032 25916 12038 25928
rect 12069 25925 12081 25928
rect 12115 25925 12127 25959
rect 12069 25919 12127 25925
rect 12434 25916 12440 25968
rect 12492 25956 12498 25968
rect 22278 25956 22284 25968
rect 12492 25928 22284 25956
rect 12492 25916 12498 25928
rect 22278 25916 22284 25928
rect 22336 25916 22342 25968
rect 24486 25956 24492 25968
rect 23492 25928 24492 25956
rect 23492 25900 23520 25928
rect 24486 25916 24492 25928
rect 24544 25916 24550 25968
rect 28626 25956 28632 25968
rect 25608 25928 28632 25956
rect 1394 25888 1400 25900
rect 1355 25860 1400 25888
rect 1394 25848 1400 25860
rect 1452 25848 1458 25900
rect 1762 25848 1768 25900
rect 1820 25888 1826 25900
rect 2133 25891 2191 25897
rect 2133 25888 2145 25891
rect 1820 25860 2145 25888
rect 1820 25848 1826 25860
rect 2133 25857 2145 25860
rect 2179 25888 2191 25891
rect 7098 25888 7104 25900
rect 2179 25860 2774 25888
rect 7059 25860 7104 25888
rect 2179 25857 2191 25860
rect 2133 25851 2191 25857
rect 2746 25820 2774 25860
rect 7098 25848 7104 25860
rect 7156 25848 7162 25900
rect 9309 25891 9367 25897
rect 9309 25857 9321 25891
rect 9355 25888 9367 25891
rect 9674 25888 9680 25900
rect 9355 25860 9680 25888
rect 9355 25857 9367 25860
rect 9309 25851 9367 25857
rect 9674 25848 9680 25860
rect 9732 25848 9738 25900
rect 9953 25891 10011 25897
rect 9953 25857 9965 25891
rect 9999 25888 10011 25891
rect 10870 25888 10876 25900
rect 9999 25860 10876 25888
rect 9999 25857 10011 25860
rect 9953 25851 10011 25857
rect 10870 25848 10876 25860
rect 10928 25848 10934 25900
rect 12802 25888 12808 25900
rect 12715 25860 12808 25888
rect 12802 25848 12808 25860
rect 12860 25888 12866 25900
rect 14090 25888 14096 25900
rect 12860 25860 14096 25888
rect 12860 25848 12866 25860
rect 14090 25848 14096 25860
rect 14148 25848 14154 25900
rect 14921 25891 14979 25897
rect 14921 25857 14933 25891
rect 14967 25888 14979 25891
rect 15562 25888 15568 25900
rect 14967 25860 15568 25888
rect 14967 25857 14979 25860
rect 14921 25851 14979 25857
rect 15562 25848 15568 25860
rect 15620 25848 15626 25900
rect 15746 25888 15752 25900
rect 15707 25860 15752 25888
rect 15746 25848 15752 25860
rect 15804 25848 15810 25900
rect 16758 25848 16764 25900
rect 16816 25888 16822 25900
rect 17221 25891 17279 25897
rect 17221 25888 17233 25891
rect 16816 25860 17233 25888
rect 16816 25848 16822 25860
rect 17221 25857 17233 25860
rect 17267 25857 17279 25891
rect 17221 25851 17279 25857
rect 17405 25891 17463 25897
rect 17405 25857 17417 25891
rect 17451 25888 17463 25891
rect 18046 25888 18052 25900
rect 17451 25860 18052 25888
rect 17451 25857 17463 25860
rect 17405 25851 17463 25857
rect 18046 25848 18052 25860
rect 18104 25848 18110 25900
rect 18230 25848 18236 25900
rect 18288 25888 18294 25900
rect 18397 25891 18455 25897
rect 18397 25888 18409 25891
rect 18288 25860 18409 25888
rect 18288 25848 18294 25860
rect 18397 25857 18409 25860
rect 18443 25857 18455 25891
rect 20073 25891 20131 25897
rect 20073 25888 20085 25891
rect 18397 25851 18455 25857
rect 19904 25860 20085 25888
rect 12434 25820 12440 25832
rect 2746 25792 12440 25820
rect 12434 25780 12440 25792
rect 12492 25780 12498 25832
rect 14826 25780 14832 25832
rect 14884 25820 14890 25832
rect 15013 25823 15071 25829
rect 15013 25820 15025 25823
rect 14884 25792 15025 25820
rect 14884 25780 14890 25792
rect 15013 25789 15025 25792
rect 15059 25820 15071 25823
rect 15654 25820 15660 25832
rect 15059 25792 15660 25820
rect 15059 25789 15071 25792
rect 15013 25783 15071 25789
rect 15654 25780 15660 25792
rect 15712 25780 15718 25832
rect 17126 25780 17132 25832
rect 17184 25820 17190 25832
rect 18141 25823 18199 25829
rect 18141 25820 18153 25823
rect 17184 25792 18153 25820
rect 17184 25780 17190 25792
rect 18141 25789 18153 25792
rect 18187 25789 18199 25823
rect 18141 25783 18199 25789
rect 11698 25752 11704 25764
rect 11659 25724 11704 25752
rect 11698 25712 11704 25724
rect 11756 25712 11762 25764
rect 12526 25752 12532 25764
rect 12084 25724 12532 25752
rect 1578 25684 1584 25696
rect 1539 25656 1584 25684
rect 1578 25644 1584 25656
rect 1636 25644 1642 25696
rect 6730 25644 6736 25696
rect 6788 25684 6794 25696
rect 7193 25687 7251 25693
rect 7193 25684 7205 25687
rect 6788 25656 7205 25684
rect 6788 25644 6794 25656
rect 7193 25653 7205 25656
rect 7239 25653 7251 25687
rect 10318 25684 10324 25696
rect 10279 25656 10324 25684
rect 7193 25647 7251 25653
rect 10318 25644 10324 25656
rect 10376 25644 10382 25696
rect 10502 25684 10508 25696
rect 10463 25656 10508 25684
rect 10502 25644 10508 25656
rect 10560 25644 10566 25696
rect 12084 25693 12112 25724
rect 12526 25712 12532 25724
rect 12584 25712 12590 25764
rect 19904 25752 19932 25860
rect 20073 25857 20085 25860
rect 20119 25857 20131 25891
rect 20073 25851 20131 25857
rect 20809 25891 20867 25897
rect 20809 25857 20821 25891
rect 20855 25857 20867 25891
rect 20809 25851 20867 25857
rect 19978 25780 19984 25832
rect 20036 25820 20042 25832
rect 20438 25820 20444 25832
rect 20036 25792 20444 25820
rect 20036 25780 20042 25792
rect 20438 25780 20444 25792
rect 20496 25820 20502 25832
rect 20824 25820 20852 25851
rect 22462 25848 22468 25900
rect 22520 25888 22526 25900
rect 23474 25888 23480 25900
rect 22520 25860 22565 25888
rect 23387 25860 23480 25888
rect 22520 25848 22526 25860
rect 23474 25848 23480 25860
rect 23532 25848 23538 25900
rect 25608 25897 25636 25928
rect 28626 25916 28632 25928
rect 28684 25956 28690 25968
rect 29380 25956 29408 25996
rect 32950 25984 32956 25996
rect 33008 25984 33014 26036
rect 33226 25984 33232 26036
rect 33284 26024 33290 26036
rect 34333 26027 34391 26033
rect 34333 26024 34345 26027
rect 33284 25996 34345 26024
rect 33284 25984 33290 25996
rect 34333 25993 34345 25996
rect 34379 25993 34391 26027
rect 36538 26024 36544 26036
rect 34333 25987 34391 25993
rect 34440 25996 36544 26024
rect 28684 25928 29408 25956
rect 28684 25916 28690 25928
rect 29546 25916 29552 25968
rect 29604 25956 29610 25968
rect 33962 25956 33968 25968
rect 29604 25928 33088 25956
rect 33923 25928 33968 25956
rect 29604 25916 29610 25928
rect 33060 25900 33088 25928
rect 33962 25916 33968 25928
rect 34020 25916 34026 25968
rect 34440 25956 34468 25996
rect 36538 25984 36544 25996
rect 36596 25984 36602 26036
rect 37366 26024 37372 26036
rect 37327 25996 37372 26024
rect 37366 25984 37372 25996
rect 37424 25984 37430 26036
rect 34072 25928 34468 25956
rect 23744 25891 23802 25897
rect 23744 25857 23756 25891
rect 23790 25888 23802 25891
rect 25593 25891 25651 25897
rect 23790 25860 25360 25888
rect 23790 25857 23802 25860
rect 23744 25851 23802 25857
rect 25332 25829 25360 25860
rect 25593 25857 25605 25891
rect 25639 25857 25651 25891
rect 25593 25851 25651 25857
rect 25685 25891 25743 25897
rect 25685 25857 25697 25891
rect 25731 25857 25743 25891
rect 25685 25851 25743 25857
rect 25777 25891 25835 25897
rect 25777 25857 25789 25891
rect 25823 25888 25835 25891
rect 25866 25888 25872 25900
rect 25823 25860 25872 25888
rect 25823 25857 25835 25860
rect 25777 25851 25835 25857
rect 20496 25792 20852 25820
rect 25317 25823 25375 25829
rect 20496 25780 20502 25792
rect 25317 25789 25329 25823
rect 25363 25789 25375 25823
rect 25700 25820 25728 25851
rect 25866 25848 25872 25860
rect 25924 25848 25930 25900
rect 25961 25891 26019 25897
rect 25961 25857 25973 25891
rect 26007 25888 26019 25891
rect 26050 25888 26056 25900
rect 26007 25860 26056 25888
rect 26007 25857 26019 25860
rect 25961 25851 26019 25857
rect 26050 25848 26056 25860
rect 26108 25848 26114 25900
rect 26878 25848 26884 25900
rect 26936 25888 26942 25900
rect 27157 25891 27215 25897
rect 27157 25888 27169 25891
rect 26936 25860 27169 25888
rect 26936 25848 26942 25860
rect 27157 25857 27169 25860
rect 27203 25857 27215 25891
rect 27157 25851 27215 25857
rect 27982 25848 27988 25900
rect 28040 25888 28046 25900
rect 28149 25891 28207 25897
rect 28149 25888 28161 25891
rect 28040 25860 28161 25888
rect 28040 25848 28046 25860
rect 28149 25857 28161 25860
rect 28195 25857 28207 25891
rect 28149 25851 28207 25857
rect 30745 25891 30803 25897
rect 30745 25857 30757 25891
rect 30791 25888 30803 25891
rect 31386 25888 31392 25900
rect 30791 25860 31392 25888
rect 30791 25857 30803 25860
rect 30745 25851 30803 25857
rect 31386 25848 31392 25860
rect 31444 25888 31450 25900
rect 32125 25891 32183 25897
rect 32125 25888 32137 25891
rect 31444 25860 32137 25888
rect 31444 25848 31450 25860
rect 32125 25857 32137 25860
rect 32171 25857 32183 25891
rect 33042 25888 33048 25900
rect 33003 25860 33048 25888
rect 32125 25851 32183 25857
rect 33042 25848 33048 25860
rect 33100 25848 33106 25900
rect 33336 25888 33456 25894
rect 34072 25888 34100 25928
rect 34698 25916 34704 25968
rect 34756 25956 34762 25968
rect 35406 25959 35464 25965
rect 35406 25956 35418 25959
rect 34756 25928 35418 25956
rect 34756 25916 34762 25928
rect 35406 25925 35418 25928
rect 35452 25925 35464 25959
rect 35406 25919 35464 25925
rect 33244 25866 34100 25888
rect 33244 25860 33364 25866
rect 33428 25860 34100 25866
rect 34149 25891 34207 25897
rect 26234 25820 26240 25832
rect 25700 25792 26240 25820
rect 25317 25783 25375 25789
rect 26234 25780 26240 25792
rect 26292 25780 26298 25832
rect 27890 25820 27896 25832
rect 27851 25792 27896 25820
rect 27890 25780 27896 25792
rect 27948 25780 27954 25832
rect 30926 25820 30932 25832
rect 30887 25792 30932 25820
rect 30926 25780 30932 25792
rect 30984 25820 30990 25832
rect 33244 25820 33272 25860
rect 34149 25857 34161 25891
rect 34195 25857 34207 25891
rect 37274 25888 37280 25900
rect 37235 25860 37280 25888
rect 34149 25851 34207 25857
rect 30984 25792 33272 25820
rect 30984 25780 30990 25792
rect 20162 25752 20168 25764
rect 19904 25724 20168 25752
rect 20162 25712 20168 25724
rect 20220 25752 20226 25764
rect 27706 25752 27712 25764
rect 20220 25724 22600 25752
rect 20220 25712 20226 25724
rect 12069 25687 12127 25693
rect 12069 25653 12081 25687
rect 12115 25653 12127 25687
rect 12069 25647 12127 25653
rect 12253 25687 12311 25693
rect 12253 25653 12265 25687
rect 12299 25684 12311 25687
rect 12618 25684 12624 25696
rect 12299 25656 12624 25684
rect 12299 25653 12311 25656
rect 12253 25647 12311 25653
rect 12618 25644 12624 25656
rect 12676 25644 12682 25696
rect 12989 25687 13047 25693
rect 12989 25653 13001 25687
rect 13035 25684 13047 25687
rect 13170 25684 13176 25696
rect 13035 25656 13176 25684
rect 13035 25653 13047 25656
rect 12989 25647 13047 25653
rect 13170 25644 13176 25656
rect 13228 25644 13234 25696
rect 14274 25644 14280 25696
rect 14332 25684 14338 25696
rect 14550 25684 14556 25696
rect 14332 25656 14556 25684
rect 14332 25644 14338 25656
rect 14550 25644 14556 25656
rect 14608 25684 14614 25696
rect 15841 25687 15899 25693
rect 15841 25684 15853 25687
rect 14608 25656 15853 25684
rect 14608 25644 14614 25656
rect 15841 25653 15853 25656
rect 15887 25653 15899 25687
rect 15841 25647 15899 25653
rect 20346 25644 20352 25696
rect 20404 25684 20410 25696
rect 22572 25693 22600 25724
rect 24412 25724 27712 25752
rect 20901 25687 20959 25693
rect 20901 25684 20913 25687
rect 20404 25656 20913 25684
rect 20404 25644 20410 25656
rect 20901 25653 20913 25656
rect 20947 25653 20959 25687
rect 20901 25647 20959 25653
rect 22557 25687 22615 25693
rect 22557 25653 22569 25687
rect 22603 25684 22615 25687
rect 24412 25684 24440 25724
rect 27706 25712 27712 25724
rect 27764 25712 27770 25764
rect 31110 25712 31116 25764
rect 31168 25752 31174 25764
rect 34164 25752 34192 25851
rect 37274 25848 37280 25860
rect 37332 25848 37338 25900
rect 34698 25780 34704 25832
rect 34756 25820 34762 25832
rect 35161 25823 35219 25829
rect 35161 25820 35173 25823
rect 34756 25792 35173 25820
rect 34756 25780 34762 25792
rect 35161 25789 35173 25792
rect 35207 25789 35219 25823
rect 35161 25783 35219 25789
rect 31168 25724 34192 25752
rect 31168 25712 31174 25724
rect 36446 25712 36452 25764
rect 36504 25752 36510 25764
rect 36541 25755 36599 25761
rect 36541 25752 36553 25755
rect 36504 25724 36553 25752
rect 36504 25712 36510 25724
rect 36541 25721 36553 25724
rect 36587 25721 36599 25755
rect 36541 25715 36599 25721
rect 37366 25712 37372 25764
rect 37424 25752 37430 25764
rect 45646 25752 45652 25764
rect 37424 25724 45652 25752
rect 37424 25712 37430 25724
rect 45646 25712 45652 25724
rect 45704 25712 45710 25764
rect 24854 25684 24860 25696
rect 22603 25656 24440 25684
rect 24815 25656 24860 25684
rect 22603 25653 22615 25656
rect 22557 25647 22615 25653
rect 24854 25644 24860 25656
rect 24912 25644 24918 25696
rect 27614 25644 27620 25696
rect 27672 25684 27678 25696
rect 28810 25684 28816 25696
rect 27672 25656 28816 25684
rect 27672 25644 27678 25656
rect 28810 25644 28816 25656
rect 28868 25684 28874 25696
rect 32582 25684 32588 25696
rect 28868 25656 32588 25684
rect 28868 25644 28874 25656
rect 32582 25644 32588 25656
rect 32640 25644 32646 25696
rect 33042 25644 33048 25696
rect 33100 25684 33106 25696
rect 37384 25684 37412 25712
rect 33100 25656 37412 25684
rect 33100 25644 33106 25656
rect 1104 25594 48852 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 48852 25594
rect 1104 25520 48852 25542
rect 7098 25440 7104 25492
rect 7156 25480 7162 25492
rect 7156 25452 9628 25480
rect 7156 25440 7162 25452
rect 9600 25412 9628 25452
rect 10318 25440 10324 25492
rect 10376 25480 10382 25492
rect 11057 25483 11115 25489
rect 11057 25480 11069 25483
rect 10376 25452 11069 25480
rect 10376 25440 10382 25452
rect 11057 25449 11069 25452
rect 11103 25449 11115 25483
rect 11057 25443 11115 25449
rect 11974 25440 11980 25492
rect 12032 25480 12038 25492
rect 12713 25483 12771 25489
rect 12713 25480 12725 25483
rect 12032 25452 12725 25480
rect 12032 25440 12038 25452
rect 12713 25449 12725 25452
rect 12759 25449 12771 25483
rect 12713 25443 12771 25449
rect 12894 25440 12900 25492
rect 12952 25480 12958 25492
rect 17034 25480 17040 25492
rect 12952 25452 17040 25480
rect 12952 25440 12958 25452
rect 17034 25440 17040 25452
rect 17092 25440 17098 25492
rect 24765 25483 24823 25489
rect 17144 25452 24716 25480
rect 17144 25412 17172 25452
rect 24688 25412 24716 25452
rect 24765 25449 24777 25483
rect 24811 25480 24823 25483
rect 26050 25480 26056 25492
rect 24811 25452 26056 25480
rect 24811 25449 24823 25452
rect 24765 25443 24823 25449
rect 26050 25440 26056 25452
rect 26108 25440 26114 25492
rect 27525 25483 27583 25489
rect 27525 25449 27537 25483
rect 27571 25480 27583 25483
rect 27614 25480 27620 25492
rect 27571 25452 27620 25480
rect 27571 25449 27583 25452
rect 27525 25443 27583 25449
rect 27614 25440 27620 25452
rect 27672 25440 27678 25492
rect 27706 25440 27712 25492
rect 27764 25480 27770 25492
rect 30006 25480 30012 25492
rect 27764 25452 30012 25480
rect 27764 25440 27770 25452
rect 30006 25440 30012 25452
rect 30064 25440 30070 25492
rect 30926 25412 30932 25424
rect 6564 25384 9536 25412
rect 9600 25384 17172 25412
rect 17236 25384 22094 25412
rect 24688 25384 30932 25412
rect 6564 25353 6592 25384
rect 6549 25347 6607 25353
rect 6549 25313 6561 25347
rect 6595 25313 6607 25347
rect 6730 25344 6736 25356
rect 6691 25316 6736 25344
rect 6549 25307 6607 25313
rect 6730 25304 6736 25316
rect 6788 25304 6794 25356
rect 8110 25344 8116 25356
rect 8071 25316 8116 25344
rect 8110 25304 8116 25316
rect 8168 25304 8174 25356
rect 9508 25344 9536 25384
rect 17236 25344 17264 25384
rect 9508 25316 17264 25344
rect 17865 25347 17923 25353
rect 17865 25313 17877 25347
rect 17911 25344 17923 25347
rect 17954 25344 17960 25356
rect 17911 25316 17960 25344
rect 17911 25313 17923 25316
rect 17865 25307 17923 25313
rect 17954 25304 17960 25316
rect 18012 25304 18018 25356
rect 19426 25304 19432 25356
rect 19484 25344 19490 25356
rect 20165 25347 20223 25353
rect 20165 25344 20177 25347
rect 19484 25316 20177 25344
rect 19484 25304 19490 25316
rect 20165 25313 20177 25316
rect 20211 25313 20223 25347
rect 20346 25344 20352 25356
rect 20307 25316 20352 25344
rect 20165 25307 20223 25313
rect 20346 25304 20352 25316
rect 20404 25304 20410 25356
rect 21542 25344 21548 25356
rect 21503 25316 21548 25344
rect 21542 25304 21548 25316
rect 21600 25304 21606 25356
rect 9125 25279 9183 25285
rect 9125 25245 9137 25279
rect 9171 25276 9183 25279
rect 10502 25276 10508 25288
rect 9171 25248 10508 25276
rect 9171 25245 9183 25248
rect 9125 25239 9183 25245
rect 10502 25236 10508 25248
rect 10560 25236 10566 25288
rect 10873 25279 10931 25285
rect 10873 25245 10885 25279
rect 10919 25276 10931 25279
rect 10962 25276 10968 25288
rect 10919 25248 10968 25276
rect 10919 25245 10931 25248
rect 10873 25239 10931 25245
rect 10962 25236 10968 25248
rect 11020 25236 11026 25288
rect 11422 25236 11428 25288
rect 11480 25276 11486 25288
rect 11609 25279 11667 25285
rect 11609 25276 11621 25279
rect 11480 25248 11621 25276
rect 11480 25236 11486 25248
rect 11609 25245 11621 25248
rect 11655 25245 11667 25279
rect 11609 25239 11667 25245
rect 11701 25279 11759 25285
rect 11701 25245 11713 25279
rect 11747 25276 11759 25279
rect 11790 25276 11796 25288
rect 11747 25248 11796 25276
rect 11747 25245 11759 25248
rect 11701 25239 11759 25245
rect 10689 25211 10747 25217
rect 10689 25177 10701 25211
rect 10735 25177 10747 25211
rect 11624 25208 11652 25239
rect 11790 25236 11796 25248
rect 11848 25236 11854 25288
rect 12713 25279 12771 25285
rect 12713 25245 12725 25279
rect 12759 25276 12771 25279
rect 12894 25276 12900 25288
rect 12759 25248 12900 25276
rect 12759 25245 12771 25248
rect 12713 25239 12771 25245
rect 12894 25236 12900 25248
rect 12952 25236 12958 25288
rect 12989 25279 13047 25285
rect 12989 25245 13001 25279
rect 13035 25276 13047 25279
rect 13354 25276 13360 25288
rect 13035 25248 13360 25276
rect 13035 25245 13047 25248
rect 12989 25239 13047 25245
rect 13354 25236 13360 25248
rect 13412 25236 13418 25288
rect 14090 25276 14096 25288
rect 14051 25248 14096 25276
rect 14090 25236 14096 25248
rect 14148 25236 14154 25288
rect 14274 25276 14280 25288
rect 14235 25248 14280 25276
rect 14274 25236 14280 25248
rect 14332 25236 14338 25288
rect 18095 25279 18153 25285
rect 18095 25276 18107 25279
rect 14384 25248 18107 25276
rect 12802 25208 12808 25220
rect 11624 25180 12808 25208
rect 10689 25171 10747 25177
rect 8938 25140 8944 25152
rect 8899 25112 8944 25140
rect 8938 25100 8944 25112
rect 8996 25100 9002 25152
rect 10704 25140 10732 25171
rect 12802 25168 12808 25180
rect 12860 25168 12866 25220
rect 13722 25168 13728 25220
rect 13780 25208 13786 25220
rect 14384 25208 14412 25248
rect 18095 25245 18107 25248
rect 18141 25245 18153 25279
rect 18095 25239 18153 25245
rect 18233 25279 18291 25285
rect 18233 25245 18245 25279
rect 18279 25245 18291 25279
rect 18233 25239 18291 25245
rect 13780 25180 14412 25208
rect 13780 25168 13786 25180
rect 17770 25168 17776 25220
rect 17828 25208 17834 25220
rect 18248 25208 18276 25239
rect 18322 25236 18328 25288
rect 18380 25276 18386 25288
rect 18509 25279 18567 25285
rect 18380 25248 18425 25276
rect 18380 25236 18386 25248
rect 18509 25245 18521 25279
rect 18555 25245 18567 25279
rect 22066 25276 22094 25384
rect 30926 25372 30932 25384
rect 30984 25372 30990 25424
rect 34606 25372 34612 25424
rect 34664 25412 34670 25424
rect 34882 25412 34888 25424
rect 34664 25384 34888 25412
rect 34664 25372 34670 25384
rect 34882 25372 34888 25384
rect 34940 25372 34946 25424
rect 22462 25304 22468 25356
rect 22520 25344 22526 25356
rect 23842 25344 23848 25356
rect 22520 25316 23848 25344
rect 22520 25304 22526 25316
rect 23842 25304 23848 25316
rect 23900 25344 23906 25356
rect 25866 25344 25872 25356
rect 23900 25316 25872 25344
rect 23900 25304 23906 25316
rect 25866 25304 25872 25316
rect 25924 25304 25930 25356
rect 29270 25344 29276 25356
rect 28736 25316 29276 25344
rect 24397 25279 24455 25285
rect 24397 25276 24409 25279
rect 22066 25248 24409 25276
rect 18509 25239 18567 25245
rect 24397 25245 24409 25248
rect 24443 25276 24455 25279
rect 24854 25276 24860 25288
rect 24443 25248 24860 25276
rect 24443 25245 24455 25248
rect 24397 25239 24455 25245
rect 17828 25180 18276 25208
rect 18524 25208 18552 25239
rect 24854 25236 24860 25248
rect 24912 25236 24918 25288
rect 26878 25236 26884 25288
rect 26936 25276 26942 25288
rect 27341 25279 27399 25285
rect 27341 25276 27353 25279
rect 26936 25248 27353 25276
rect 26936 25236 26942 25248
rect 27341 25245 27353 25248
rect 27387 25245 27399 25279
rect 28350 25276 28356 25288
rect 27341 25239 27399 25245
rect 27632 25248 28356 25276
rect 20622 25208 20628 25220
rect 18524 25180 20628 25208
rect 17828 25168 17834 25180
rect 20622 25168 20628 25180
rect 20680 25208 20686 25220
rect 21818 25208 21824 25220
rect 20680 25180 21824 25208
rect 20680 25168 20686 25180
rect 21818 25168 21824 25180
rect 21876 25168 21882 25220
rect 24486 25168 24492 25220
rect 24544 25208 24550 25220
rect 24581 25211 24639 25217
rect 24581 25208 24593 25211
rect 24544 25180 24593 25208
rect 24544 25168 24550 25180
rect 24581 25177 24593 25180
rect 24627 25208 24639 25211
rect 27632 25208 27660 25248
rect 28350 25236 28356 25248
rect 28408 25236 28414 25288
rect 28626 25285 28632 25288
rect 28609 25279 28632 25285
rect 28609 25245 28621 25279
rect 28609 25239 28632 25245
rect 28626 25236 28632 25239
rect 28684 25236 28690 25288
rect 28736 25285 28764 25316
rect 29270 25304 29276 25316
rect 29328 25304 29334 25356
rect 30558 25344 30564 25356
rect 30519 25316 30564 25344
rect 30558 25304 30564 25316
rect 30616 25304 30622 25356
rect 31754 25304 31760 25356
rect 31812 25344 31818 25356
rect 35526 25344 35532 25356
rect 31812 25316 31857 25344
rect 35084 25316 35532 25344
rect 31812 25304 31818 25316
rect 28721 25279 28779 25285
rect 28721 25245 28733 25279
rect 28767 25245 28779 25279
rect 28721 25239 28779 25245
rect 28813 25279 28871 25285
rect 28813 25245 28825 25279
rect 28859 25245 28871 25279
rect 28813 25239 28871 25245
rect 28997 25279 29055 25285
rect 28997 25245 29009 25279
rect 29043 25276 29055 25279
rect 29917 25279 29975 25285
rect 29917 25276 29929 25279
rect 29043 25248 29929 25276
rect 29043 25245 29055 25248
rect 28997 25239 29055 25245
rect 29917 25245 29929 25248
rect 29963 25245 29975 25279
rect 30374 25276 30380 25288
rect 30335 25248 30380 25276
rect 29917 25239 29975 25245
rect 24627 25180 27660 25208
rect 28828 25208 28856 25239
rect 30374 25236 30380 25248
rect 30432 25236 30438 25288
rect 32677 25279 32735 25285
rect 32677 25245 32689 25279
rect 32723 25276 32735 25279
rect 32766 25276 32772 25288
rect 32723 25248 32772 25276
rect 32723 25245 32735 25248
rect 32677 25239 32735 25245
rect 32766 25236 32772 25248
rect 32824 25276 32830 25288
rect 34698 25276 34704 25288
rect 32824 25248 34704 25276
rect 32824 25236 32830 25248
rect 34698 25236 34704 25248
rect 34756 25236 34762 25288
rect 34790 25236 34796 25288
rect 34848 25276 34854 25288
rect 35084 25285 35112 25316
rect 35526 25304 35532 25316
rect 35584 25304 35590 25356
rect 36446 25304 36452 25356
rect 36504 25344 36510 25356
rect 37369 25347 37427 25353
rect 37369 25344 37381 25347
rect 36504 25316 37381 25344
rect 36504 25304 36510 25316
rect 37369 25313 37381 25316
rect 37415 25313 37427 25347
rect 37369 25307 37427 25313
rect 34977 25279 35035 25285
rect 34977 25276 34989 25279
rect 34848 25248 34989 25276
rect 34848 25236 34854 25248
rect 34977 25245 34989 25248
rect 35023 25245 35035 25279
rect 34977 25239 35035 25245
rect 35069 25279 35127 25285
rect 35069 25245 35081 25279
rect 35115 25245 35127 25279
rect 35069 25239 35127 25245
rect 35158 25236 35164 25288
rect 35216 25276 35222 25288
rect 35345 25279 35403 25285
rect 35216 25248 35261 25276
rect 35216 25236 35222 25248
rect 35345 25245 35357 25279
rect 35391 25276 35403 25279
rect 35894 25276 35900 25288
rect 35391 25248 35900 25276
rect 35391 25245 35403 25248
rect 35345 25239 35403 25245
rect 35894 25236 35900 25248
rect 35952 25236 35958 25288
rect 36725 25279 36783 25285
rect 36725 25245 36737 25279
rect 36771 25276 36783 25279
rect 37274 25276 37280 25288
rect 36771 25248 37280 25276
rect 36771 25245 36783 25248
rect 36725 25239 36783 25245
rect 37274 25236 37280 25248
rect 37332 25236 37338 25288
rect 47854 25276 47860 25288
rect 47815 25248 47860 25276
rect 47854 25236 47860 25248
rect 47912 25236 47918 25288
rect 29362 25208 29368 25220
rect 28828 25180 29368 25208
rect 24627 25177 24639 25180
rect 24581 25171 24639 25177
rect 29362 25168 29368 25180
rect 29420 25168 29426 25220
rect 29549 25211 29607 25217
rect 29549 25177 29561 25211
rect 29595 25177 29607 25211
rect 29549 25171 29607 25177
rect 11698 25140 11704 25152
rect 10704 25112 11704 25140
rect 11698 25100 11704 25112
rect 11756 25140 11762 25152
rect 11885 25143 11943 25149
rect 11885 25140 11897 25143
rect 11756 25112 11897 25140
rect 11756 25100 11762 25112
rect 11885 25109 11897 25112
rect 11931 25109 11943 25143
rect 12894 25140 12900 25152
rect 12855 25112 12900 25140
rect 11885 25103 11943 25109
rect 12894 25100 12900 25112
rect 12952 25100 12958 25152
rect 13814 25100 13820 25152
rect 13872 25140 13878 25152
rect 14461 25143 14519 25149
rect 14461 25140 14473 25143
rect 13872 25112 14473 25140
rect 13872 25100 13878 25112
rect 14461 25109 14473 25112
rect 14507 25109 14519 25143
rect 14461 25103 14519 25109
rect 17034 25100 17040 25152
rect 17092 25140 17098 25152
rect 21634 25140 21640 25152
rect 17092 25112 21640 25140
rect 17092 25100 17098 25112
rect 21634 25100 21640 25112
rect 21692 25140 21698 25152
rect 27154 25140 27160 25152
rect 21692 25112 27160 25140
rect 21692 25100 21698 25112
rect 27154 25100 27160 25112
rect 27212 25140 27218 25152
rect 27338 25140 27344 25152
rect 27212 25112 27344 25140
rect 27212 25100 27218 25112
rect 27338 25100 27344 25112
rect 27396 25100 27402 25152
rect 28353 25143 28411 25149
rect 28353 25109 28365 25143
rect 28399 25140 28411 25143
rect 29454 25140 29460 25152
rect 28399 25112 29460 25140
rect 28399 25109 28411 25112
rect 28353 25103 28411 25109
rect 29454 25100 29460 25112
rect 29512 25100 29518 25152
rect 29564 25140 29592 25171
rect 29638 25168 29644 25220
rect 29696 25208 29702 25220
rect 29733 25211 29791 25217
rect 29733 25208 29745 25211
rect 29696 25180 29745 25208
rect 29696 25168 29702 25180
rect 29733 25177 29745 25180
rect 29779 25208 29791 25211
rect 31110 25208 31116 25220
rect 29779 25180 31116 25208
rect 29779 25177 29791 25180
rect 29733 25171 29791 25177
rect 31110 25168 31116 25180
rect 31168 25168 31174 25220
rect 32944 25211 33002 25217
rect 32944 25177 32956 25211
rect 32990 25208 33002 25211
rect 33318 25208 33324 25220
rect 32990 25180 33324 25208
rect 32990 25177 33002 25180
rect 32944 25171 33002 25177
rect 33318 25168 33324 25180
rect 33376 25168 33382 25220
rect 34606 25168 34612 25220
rect 34664 25208 34670 25220
rect 34808 25208 34836 25236
rect 34664 25180 34836 25208
rect 36817 25211 36875 25217
rect 34664 25168 34670 25180
rect 36817 25177 36829 25211
rect 36863 25208 36875 25211
rect 37553 25211 37611 25217
rect 37553 25208 37565 25211
rect 36863 25180 37565 25208
rect 36863 25177 36875 25180
rect 36817 25171 36875 25177
rect 37553 25177 37565 25180
rect 37599 25177 37611 25211
rect 37553 25171 37611 25177
rect 39209 25211 39267 25217
rect 39209 25177 39221 25211
rect 39255 25208 39267 25211
rect 48498 25208 48504 25220
rect 39255 25180 48504 25208
rect 39255 25177 39267 25180
rect 39209 25171 39267 25177
rect 48498 25168 48504 25180
rect 48556 25168 48562 25220
rect 30374 25140 30380 25152
rect 29564 25112 30380 25140
rect 30374 25100 30380 25112
rect 30432 25100 30438 25152
rect 34057 25143 34115 25149
rect 34057 25109 34069 25143
rect 34103 25140 34115 25143
rect 34514 25140 34520 25152
rect 34103 25112 34520 25140
rect 34103 25109 34115 25112
rect 34057 25103 34115 25109
rect 34514 25100 34520 25112
rect 34572 25100 34578 25152
rect 34701 25143 34759 25149
rect 34701 25109 34713 25143
rect 34747 25140 34759 25143
rect 35618 25140 35624 25152
rect 34747 25112 35624 25140
rect 34747 25109 34759 25112
rect 34701 25103 34759 25109
rect 35618 25100 35624 25112
rect 35676 25100 35682 25152
rect 39942 25100 39948 25152
rect 40000 25140 40006 25152
rect 48041 25143 48099 25149
rect 48041 25140 48053 25143
rect 40000 25112 48053 25140
rect 40000 25100 40006 25112
rect 48041 25109 48053 25112
rect 48087 25109 48099 25143
rect 48041 25103 48099 25109
rect 1104 25050 48852 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 48852 25050
rect 1104 24976 48852 24998
rect 9398 24896 9404 24948
rect 9456 24936 9462 24948
rect 29546 24936 29552 24948
rect 9456 24908 29552 24936
rect 9456 24896 9462 24908
rect 29546 24896 29552 24908
rect 29604 24896 29610 24948
rect 30374 24896 30380 24948
rect 30432 24936 30438 24948
rect 30745 24939 30803 24945
rect 30745 24936 30757 24939
rect 30432 24908 30757 24936
rect 30432 24896 30438 24908
rect 30745 24905 30757 24908
rect 30791 24905 30803 24939
rect 31386 24936 31392 24948
rect 31347 24908 31392 24936
rect 30745 24899 30803 24905
rect 31386 24896 31392 24908
rect 31444 24936 31450 24948
rect 31444 24908 31754 24936
rect 31444 24896 31450 24908
rect 14826 24868 14832 24880
rect 14787 24840 14832 24868
rect 14826 24828 14832 24840
rect 14884 24828 14890 24880
rect 22094 24877 22100 24880
rect 22088 24831 22100 24877
rect 22152 24868 22158 24880
rect 22152 24840 22188 24868
rect 27080 24840 27292 24868
rect 22094 24828 22100 24831
rect 22152 24828 22158 24840
rect 7742 24800 7748 24812
rect 7703 24772 7748 24800
rect 7742 24760 7748 24772
rect 7800 24760 7806 24812
rect 8012 24803 8070 24809
rect 8012 24769 8024 24803
rect 8058 24800 8070 24803
rect 8938 24800 8944 24812
rect 8058 24772 8944 24800
rect 8058 24769 8070 24772
rect 8012 24763 8070 24769
rect 8938 24760 8944 24772
rect 8996 24760 9002 24812
rect 10137 24803 10195 24809
rect 10137 24769 10149 24803
rect 10183 24769 10195 24803
rect 10137 24763 10195 24769
rect 10321 24803 10379 24809
rect 10321 24769 10333 24803
rect 10367 24800 10379 24803
rect 10778 24800 10784 24812
rect 10367 24772 10784 24800
rect 10367 24769 10379 24772
rect 10321 24763 10379 24769
rect 10152 24732 10180 24763
rect 10778 24760 10784 24772
rect 10836 24760 10842 24812
rect 14182 24760 14188 24812
rect 14240 24800 14246 24812
rect 14921 24803 14979 24809
rect 14921 24800 14933 24803
rect 14240 24772 14933 24800
rect 14240 24760 14246 24772
rect 14921 24769 14933 24772
rect 14967 24769 14979 24803
rect 14921 24763 14979 24769
rect 15010 24760 15016 24812
rect 15068 24800 15074 24812
rect 15068 24772 15884 24800
rect 15068 24760 15074 24772
rect 10594 24732 10600 24744
rect 10152 24704 10600 24732
rect 10594 24692 10600 24704
rect 10652 24692 10658 24744
rect 14461 24735 14519 24741
rect 14461 24701 14473 24735
rect 14507 24732 14519 24735
rect 15746 24732 15752 24744
rect 14507 24704 15752 24732
rect 14507 24701 14519 24704
rect 14461 24695 14519 24701
rect 15746 24692 15752 24704
rect 15804 24692 15810 24744
rect 15856 24732 15884 24772
rect 21560 24772 23152 24800
rect 21560 24732 21588 24772
rect 21818 24732 21824 24744
rect 15856 24704 21588 24732
rect 21779 24704 21824 24732
rect 21818 24692 21824 24704
rect 21876 24692 21882 24744
rect 23124 24732 23152 24772
rect 25866 24760 25872 24812
rect 25924 24800 25930 24812
rect 26053 24803 26111 24809
rect 26053 24800 26065 24803
rect 25924 24772 26065 24800
rect 25924 24760 25930 24772
rect 26053 24769 26065 24772
rect 26099 24769 26111 24803
rect 26878 24800 26884 24812
rect 26053 24763 26111 24769
rect 26160 24772 26884 24800
rect 26160 24732 26188 24772
rect 26878 24760 26884 24772
rect 26936 24760 26942 24812
rect 26973 24803 27031 24809
rect 26973 24769 26985 24803
rect 27019 24800 27031 24803
rect 27080 24800 27108 24840
rect 27019 24772 27108 24800
rect 27157 24803 27215 24809
rect 27019 24769 27031 24772
rect 26973 24763 27031 24769
rect 27157 24769 27169 24803
rect 27203 24769 27215 24803
rect 27157 24763 27215 24769
rect 23124 24704 26188 24732
rect 11790 24624 11796 24676
rect 11848 24664 11854 24676
rect 20622 24664 20628 24676
rect 11848 24636 20628 24664
rect 11848 24624 11854 24636
rect 20622 24624 20628 24636
rect 20680 24624 20686 24676
rect 23124 24664 23152 24704
rect 26234 24692 26240 24744
rect 26292 24732 26298 24744
rect 27172 24732 27200 24763
rect 26292 24704 27200 24732
rect 27264 24732 27292 24840
rect 27706 24828 27712 24880
rect 27764 24868 27770 24880
rect 27801 24871 27859 24877
rect 27801 24868 27813 24871
rect 27764 24840 27813 24868
rect 27764 24828 27770 24840
rect 27801 24837 27813 24840
rect 27847 24837 27859 24871
rect 28001 24871 28059 24877
rect 28001 24868 28013 24871
rect 27801 24831 27859 24837
rect 28000 24837 28013 24868
rect 28047 24837 28059 24871
rect 28000 24831 28059 24837
rect 27338 24760 27344 24812
rect 27396 24800 27402 24812
rect 28000 24800 28028 24831
rect 28258 24828 28264 24880
rect 28316 24868 28322 24880
rect 31726 24868 31754 24908
rect 33778 24896 33784 24948
rect 33836 24936 33842 24948
rect 35158 24936 35164 24948
rect 33836 24908 35164 24936
rect 33836 24896 33842 24908
rect 35158 24896 35164 24908
rect 35216 24896 35222 24948
rect 35618 24877 35624 24880
rect 32493 24871 32551 24877
rect 32493 24868 32505 24871
rect 28316 24840 28764 24868
rect 31726 24840 32505 24868
rect 28316 24828 28322 24840
rect 28626 24800 28632 24812
rect 27396 24772 27441 24800
rect 28000 24772 28632 24800
rect 27396 24760 27402 24772
rect 28626 24760 28632 24772
rect 28684 24760 28690 24812
rect 28736 24809 28764 24840
rect 32493 24837 32505 24840
rect 32539 24837 32551 24871
rect 35612 24868 35624 24877
rect 35579 24840 35624 24868
rect 32493 24831 32551 24837
rect 35612 24831 35624 24840
rect 35618 24828 35624 24831
rect 35676 24828 35682 24880
rect 28721 24803 28779 24809
rect 28721 24769 28733 24803
rect 28767 24769 28779 24803
rect 28721 24763 28779 24769
rect 28905 24803 28963 24809
rect 28905 24769 28917 24803
rect 28951 24800 28963 24803
rect 28994 24800 29000 24812
rect 28951 24772 29000 24800
rect 28951 24769 28963 24772
rect 28905 24763 28963 24769
rect 28994 24760 29000 24772
rect 29052 24760 29058 24812
rect 29454 24760 29460 24812
rect 29512 24800 29518 24812
rect 29621 24803 29679 24809
rect 29621 24800 29633 24803
rect 29512 24772 29633 24800
rect 29512 24760 29518 24772
rect 29621 24769 29633 24772
rect 29667 24769 29679 24803
rect 29621 24763 29679 24769
rect 30006 24760 30012 24812
rect 30064 24800 30070 24812
rect 31205 24803 31263 24809
rect 31205 24800 31217 24803
rect 30064 24772 31217 24800
rect 30064 24760 30070 24772
rect 31205 24769 31217 24772
rect 31251 24769 31263 24803
rect 31205 24763 31263 24769
rect 31726 24772 36400 24800
rect 27798 24732 27804 24744
rect 27264 24704 27804 24732
rect 26292 24692 26298 24704
rect 23201 24667 23259 24673
rect 23201 24664 23213 24667
rect 23124 24636 23213 24664
rect 23201 24633 23213 24636
rect 23247 24633 23259 24667
rect 23201 24627 23259 24633
rect 24394 24624 24400 24676
rect 24452 24664 24458 24676
rect 24452 24636 26280 24664
rect 24452 24624 24458 24636
rect 9122 24596 9128 24608
rect 9083 24568 9128 24596
rect 9122 24556 9128 24568
rect 9180 24556 9186 24608
rect 10226 24596 10232 24608
rect 10187 24568 10232 24596
rect 10226 24556 10232 24568
rect 10284 24556 10290 24608
rect 10318 24556 10324 24608
rect 10376 24596 10382 24608
rect 11882 24596 11888 24608
rect 10376 24568 11888 24596
rect 10376 24556 10382 24568
rect 11882 24556 11888 24568
rect 11940 24556 11946 24608
rect 14090 24556 14096 24608
rect 14148 24596 14154 24608
rect 14645 24599 14703 24605
rect 14645 24596 14657 24599
rect 14148 24568 14657 24596
rect 14148 24556 14154 24568
rect 14645 24565 14657 24568
rect 14691 24565 14703 24599
rect 26050 24596 26056 24608
rect 26011 24568 26056 24596
rect 14645 24559 14703 24565
rect 26050 24556 26056 24568
rect 26108 24556 26114 24608
rect 26252 24596 26280 24636
rect 26326 24624 26332 24676
rect 26384 24664 26390 24676
rect 27264 24664 27292 24704
rect 27798 24692 27804 24704
rect 27856 24692 27862 24744
rect 27890 24692 27896 24744
rect 27948 24732 27954 24744
rect 29365 24735 29423 24741
rect 29365 24732 29377 24735
rect 27948 24704 29377 24732
rect 27948 24692 27954 24704
rect 29365 24701 29377 24704
rect 29411 24701 29423 24735
rect 29365 24695 29423 24701
rect 30374 24692 30380 24744
rect 30432 24732 30438 24744
rect 31726 24732 31754 24772
rect 34238 24732 34244 24744
rect 30432 24704 31754 24732
rect 34199 24704 34244 24732
rect 30432 24692 30438 24704
rect 34238 24692 34244 24704
rect 34296 24692 34302 24744
rect 34698 24692 34704 24744
rect 34756 24732 34762 24744
rect 35345 24735 35403 24741
rect 35345 24732 35357 24735
rect 34756 24704 35357 24732
rect 34756 24692 34762 24704
rect 35345 24701 35357 24704
rect 35391 24701 35403 24735
rect 36372 24732 36400 24772
rect 37274 24760 37280 24812
rect 37332 24800 37338 24812
rect 37461 24803 37519 24809
rect 37461 24800 37473 24803
rect 37332 24772 37473 24800
rect 37332 24760 37338 24772
rect 37461 24769 37473 24772
rect 37507 24800 37519 24803
rect 38105 24803 38163 24809
rect 38105 24800 38117 24803
rect 37507 24772 38117 24800
rect 37507 24769 37519 24772
rect 37461 24763 37519 24769
rect 38105 24769 38117 24772
rect 38151 24769 38163 24803
rect 47302 24800 47308 24812
rect 38105 24763 38163 24769
rect 41386 24772 47308 24800
rect 41386 24732 41414 24772
rect 47302 24760 47308 24772
rect 47360 24760 47366 24812
rect 47578 24800 47584 24812
rect 47539 24772 47584 24800
rect 47578 24760 47584 24772
rect 47636 24760 47642 24812
rect 36372 24704 41414 24732
rect 35345 24695 35403 24701
rect 28902 24664 28908 24676
rect 26384 24636 27292 24664
rect 27724 24636 28908 24664
rect 26384 24624 26390 24636
rect 27724 24596 27752 24636
rect 28902 24624 28908 24636
rect 28960 24624 28966 24676
rect 47596 24664 47624 24760
rect 30300 24636 31340 24664
rect 26252 24568 27752 24596
rect 27798 24556 27804 24608
rect 27856 24596 27862 24608
rect 27985 24599 28043 24605
rect 27985 24596 27997 24599
rect 27856 24568 27997 24596
rect 27856 24556 27862 24568
rect 27985 24565 27997 24568
rect 28031 24565 28043 24599
rect 27985 24559 28043 24565
rect 28074 24556 28080 24608
rect 28132 24596 28138 24608
rect 28169 24599 28227 24605
rect 28169 24596 28181 24599
rect 28132 24568 28181 24596
rect 28132 24556 28138 24568
rect 28169 24565 28181 24568
rect 28215 24565 28227 24599
rect 28169 24559 28227 24565
rect 28534 24556 28540 24608
rect 28592 24596 28598 24608
rect 30300 24596 30328 24636
rect 28592 24568 30328 24596
rect 31312 24596 31340 24636
rect 36280 24636 47624 24664
rect 33042 24596 33048 24608
rect 31312 24568 33048 24596
rect 28592 24556 28598 24568
rect 33042 24556 33048 24568
rect 33100 24556 33106 24608
rect 33226 24556 33232 24608
rect 33284 24596 33290 24608
rect 36280 24596 36308 24636
rect 36722 24596 36728 24608
rect 33284 24568 36308 24596
rect 36683 24568 36728 24596
rect 33284 24556 33290 24568
rect 36722 24556 36728 24568
rect 36780 24556 36786 24608
rect 37553 24599 37611 24605
rect 37553 24565 37565 24599
rect 37599 24596 37611 24599
rect 37642 24596 37648 24608
rect 37599 24568 37648 24596
rect 37599 24565 37611 24568
rect 37553 24559 37611 24565
rect 37642 24556 37648 24568
rect 37700 24556 37706 24608
rect 38194 24596 38200 24608
rect 38155 24568 38200 24596
rect 38194 24556 38200 24568
rect 38252 24556 38258 24608
rect 46290 24556 46296 24608
rect 46348 24596 46354 24608
rect 47029 24599 47087 24605
rect 47029 24596 47041 24599
rect 46348 24568 47041 24596
rect 46348 24556 46354 24568
rect 47029 24565 47041 24568
rect 47075 24565 47087 24599
rect 47670 24596 47676 24608
rect 47631 24568 47676 24596
rect 47029 24559 47087 24565
rect 47670 24556 47676 24568
rect 47728 24556 47734 24608
rect 1104 24506 48852 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 48852 24506
rect 1104 24432 48852 24454
rect 9861 24395 9919 24401
rect 9861 24361 9873 24395
rect 9907 24392 9919 24395
rect 12713 24395 12771 24401
rect 9907 24364 12434 24392
rect 9907 24361 9919 24364
rect 9861 24355 9919 24361
rect 9306 24324 9312 24336
rect 9267 24296 9312 24324
rect 9306 24284 9312 24296
rect 9364 24284 9370 24336
rect 9401 24327 9459 24333
rect 9401 24293 9413 24327
rect 9447 24324 9459 24327
rect 9447 24296 11100 24324
rect 9447 24293 9459 24296
rect 9401 24287 9459 24293
rect 10226 24256 10232 24268
rect 10187 24228 10232 24256
rect 10226 24216 10232 24228
rect 10284 24216 10290 24268
rect 10502 24216 10508 24268
rect 10560 24256 10566 24268
rect 10962 24256 10968 24268
rect 10560 24228 10968 24256
rect 10560 24216 10566 24228
rect 10962 24216 10968 24228
rect 11020 24216 11026 24268
rect 11072 24256 11100 24296
rect 11146 24284 11152 24336
rect 11204 24324 11210 24336
rect 11204 24296 11249 24324
rect 11204 24284 11210 24296
rect 11238 24256 11244 24268
rect 11072 24228 11244 24256
rect 11238 24216 11244 24228
rect 11296 24216 11302 24268
rect 11790 24256 11796 24268
rect 11751 24228 11796 24256
rect 11790 24216 11796 24228
rect 11848 24216 11854 24268
rect 12406 24256 12434 24364
rect 12713 24361 12725 24395
rect 12759 24392 12771 24395
rect 12894 24392 12900 24404
rect 12759 24364 12900 24392
rect 12759 24361 12771 24364
rect 12713 24355 12771 24361
rect 12894 24352 12900 24364
rect 12952 24352 12958 24404
rect 22738 24352 22744 24404
rect 22796 24392 22802 24404
rect 23382 24392 23388 24404
rect 22796 24364 23388 24392
rect 22796 24352 22802 24364
rect 23382 24352 23388 24364
rect 23440 24352 23446 24404
rect 25976 24364 27660 24392
rect 13081 24259 13139 24265
rect 13081 24256 13093 24259
rect 12406 24228 13093 24256
rect 13081 24225 13093 24228
rect 13127 24225 13139 24259
rect 13081 24219 13139 24225
rect 13173 24259 13231 24265
rect 13173 24225 13185 24259
rect 13219 24256 13231 24259
rect 13814 24256 13820 24268
rect 13219 24228 13820 24256
rect 13219 24225 13231 24228
rect 13173 24219 13231 24225
rect 13814 24216 13820 24228
rect 13872 24216 13878 24268
rect 14182 24216 14188 24268
rect 14240 24256 14246 24268
rect 14461 24259 14519 24265
rect 14461 24256 14473 24259
rect 14240 24228 14473 24256
rect 14240 24216 14246 24228
rect 14461 24225 14473 24228
rect 14507 24225 14519 24259
rect 25976 24256 26004 24364
rect 26326 24324 26332 24336
rect 14461 24219 14519 24225
rect 18340 24228 26004 24256
rect 26068 24296 26332 24324
rect 8846 24148 8852 24200
rect 8904 24188 8910 24200
rect 10045 24191 10103 24197
rect 10045 24188 10057 24191
rect 8904 24160 10057 24188
rect 8904 24148 8910 24160
rect 10045 24157 10057 24160
rect 10091 24157 10103 24191
rect 10045 24151 10103 24157
rect 10134 24148 10140 24200
rect 10192 24188 10198 24200
rect 10192 24160 10237 24188
rect 10192 24148 10198 24160
rect 10318 24148 10324 24200
rect 10376 24188 10382 24200
rect 10870 24188 10876 24200
rect 10376 24160 10876 24188
rect 10376 24148 10382 24160
rect 10870 24148 10876 24160
rect 10928 24148 10934 24200
rect 11882 24188 11888 24200
rect 11843 24160 11888 24188
rect 11882 24148 11888 24160
rect 11940 24148 11946 24200
rect 12894 24188 12900 24200
rect 12855 24160 12900 24188
rect 12894 24148 12900 24160
rect 12952 24148 12958 24200
rect 12989 24191 13047 24197
rect 12989 24157 13001 24191
rect 13035 24188 13047 24191
rect 13906 24188 13912 24200
rect 13035 24160 13912 24188
rect 13035 24157 13047 24160
rect 12989 24151 13047 24157
rect 13906 24148 13912 24160
rect 13964 24148 13970 24200
rect 14090 24188 14096 24200
rect 14051 24160 14096 24188
rect 14090 24148 14096 24160
rect 14148 24148 14154 24200
rect 14277 24191 14335 24197
rect 14277 24157 14289 24191
rect 14323 24157 14335 24191
rect 14277 24151 14335 24157
rect 14369 24191 14427 24197
rect 14369 24157 14381 24191
rect 14415 24157 14427 24191
rect 14369 24151 14427 24157
rect 14645 24191 14703 24197
rect 14645 24157 14657 24191
rect 14691 24188 14703 24191
rect 14826 24188 14832 24200
rect 14691 24160 14832 24188
rect 14691 24157 14703 24160
rect 14645 24151 14703 24157
rect 1854 24120 1860 24132
rect 1815 24092 1860 24120
rect 1854 24080 1860 24092
rect 1912 24080 1918 24132
rect 2041 24123 2099 24129
rect 2041 24089 2053 24123
rect 2087 24120 2099 24123
rect 2682 24120 2688 24132
rect 2087 24092 2688 24120
rect 2087 24089 2099 24092
rect 2041 24083 2099 24089
rect 2682 24080 2688 24092
rect 2740 24080 2746 24132
rect 8941 24123 8999 24129
rect 8941 24089 8953 24123
rect 8987 24089 8999 24123
rect 8941 24083 8999 24089
rect 8956 24052 8984 24083
rect 9122 24080 9128 24132
rect 9180 24120 9186 24132
rect 10962 24120 10968 24132
rect 9180 24092 10968 24120
rect 9180 24080 9186 24092
rect 10962 24080 10968 24092
rect 11020 24080 11026 24132
rect 11422 24080 11428 24132
rect 11480 24120 11486 24132
rect 14292 24120 14320 24151
rect 11480 24092 14320 24120
rect 11480 24080 11486 24092
rect 9398 24052 9404 24064
rect 8956 24024 9404 24052
rect 9398 24012 9404 24024
rect 9456 24052 9462 24064
rect 11698 24052 11704 24064
rect 9456 24024 11704 24052
rect 9456 24012 9462 24024
rect 11698 24012 11704 24024
rect 11756 24012 11762 24064
rect 11882 24012 11888 24064
rect 11940 24052 11946 24064
rect 12253 24055 12311 24061
rect 12253 24052 12265 24055
rect 11940 24024 12265 24052
rect 11940 24012 11946 24024
rect 12253 24021 12265 24024
rect 12299 24052 12311 24055
rect 14384 24052 14412 24151
rect 14826 24148 14832 24160
rect 14884 24148 14890 24200
rect 15286 24148 15292 24200
rect 15344 24188 15350 24200
rect 15473 24191 15531 24197
rect 15344 24160 15389 24188
rect 15344 24148 15350 24160
rect 15473 24157 15485 24191
rect 15519 24157 15531 24191
rect 15473 24151 15531 24157
rect 16025 24191 16083 24197
rect 16025 24157 16037 24191
rect 16071 24188 16083 24191
rect 17310 24188 17316 24200
rect 16071 24160 17316 24188
rect 16071 24157 16083 24160
rect 16025 24151 16083 24157
rect 14918 24080 14924 24132
rect 14976 24120 14982 24132
rect 15488 24120 15516 24151
rect 17310 24148 17316 24160
rect 17368 24148 17374 24200
rect 18340 24197 18368 24228
rect 17773 24191 17831 24197
rect 17773 24157 17785 24191
rect 17819 24188 17831 24191
rect 18325 24191 18383 24197
rect 18325 24188 18337 24191
rect 17819 24160 18337 24188
rect 17819 24157 17831 24160
rect 17773 24151 17831 24157
rect 18325 24157 18337 24160
rect 18371 24157 18383 24191
rect 18325 24151 18383 24157
rect 18417 24191 18475 24197
rect 18417 24157 18429 24191
rect 18463 24157 18475 24191
rect 18417 24151 18475 24157
rect 18509 24191 18567 24197
rect 18509 24157 18521 24191
rect 18555 24157 18567 24191
rect 18690 24188 18696 24200
rect 18651 24160 18696 24188
rect 18509 24151 18567 24157
rect 14976 24092 15516 24120
rect 16292 24123 16350 24129
rect 14976 24080 14982 24092
rect 16292 24089 16304 24123
rect 16338 24120 16350 24123
rect 16666 24120 16672 24132
rect 16338 24092 16672 24120
rect 16338 24089 16350 24092
rect 16292 24083 16350 24089
rect 16666 24080 16672 24092
rect 16724 24080 16730 24132
rect 18230 24080 18236 24132
rect 18288 24120 18294 24132
rect 18432 24120 18460 24151
rect 18288 24092 18460 24120
rect 18524 24120 18552 24151
rect 18690 24148 18696 24160
rect 18748 24148 18754 24200
rect 19978 24148 19984 24200
rect 20036 24188 20042 24200
rect 20254 24188 20260 24200
rect 20036 24160 20260 24188
rect 20036 24148 20042 24160
rect 20254 24148 20260 24160
rect 20312 24188 20318 24200
rect 24397 24191 24455 24197
rect 20312 24160 24348 24188
rect 20312 24148 20318 24160
rect 19426 24120 19432 24132
rect 18524 24092 19432 24120
rect 18288 24080 18294 24092
rect 19426 24080 19432 24092
rect 19484 24080 19490 24132
rect 20346 24080 20352 24132
rect 20404 24120 20410 24132
rect 20441 24123 20499 24129
rect 20441 24120 20453 24123
rect 20404 24092 20453 24120
rect 20404 24080 20410 24092
rect 20441 24089 20453 24092
rect 20487 24089 20499 24123
rect 20622 24120 20628 24132
rect 20583 24092 20628 24120
rect 20441 24083 20499 24089
rect 20622 24080 20628 24092
rect 20680 24080 20686 24132
rect 22094 24080 22100 24132
rect 22152 24120 22158 24132
rect 24320 24120 24348 24160
rect 24397 24157 24409 24191
rect 24443 24188 24455 24191
rect 24762 24188 24768 24200
rect 24443 24160 24768 24188
rect 24443 24157 24455 24160
rect 24397 24151 24455 24157
rect 24762 24148 24768 24160
rect 24820 24148 24826 24200
rect 26068 24197 26096 24296
rect 26326 24284 26332 24296
rect 26384 24284 26390 24336
rect 27632 24324 27660 24364
rect 29362 24352 29368 24404
rect 29420 24392 29426 24404
rect 30098 24392 30104 24404
rect 29420 24364 30104 24392
rect 29420 24352 29426 24364
rect 30098 24352 30104 24364
rect 30156 24352 30162 24404
rect 30650 24352 30656 24404
rect 30708 24392 30714 24404
rect 31846 24392 31852 24404
rect 30708 24364 31852 24392
rect 30708 24352 30714 24364
rect 31846 24352 31852 24364
rect 31904 24392 31910 24404
rect 32401 24395 32459 24401
rect 32401 24392 32413 24395
rect 31904 24364 32413 24392
rect 31904 24352 31910 24364
rect 32401 24361 32413 24364
rect 32447 24361 32459 24395
rect 33318 24392 33324 24404
rect 33279 24364 33324 24392
rect 32401 24355 32459 24361
rect 33318 24352 33324 24364
rect 33376 24352 33382 24404
rect 33502 24352 33508 24404
rect 33560 24392 33566 24404
rect 34238 24392 34244 24404
rect 33560 24364 34244 24392
rect 33560 24352 33566 24364
rect 34238 24352 34244 24364
rect 34296 24392 34302 24404
rect 35526 24392 35532 24404
rect 34296 24364 35532 24392
rect 34296 24352 34302 24364
rect 35526 24352 35532 24364
rect 35584 24352 35590 24404
rect 35894 24392 35900 24404
rect 35855 24364 35900 24392
rect 35894 24352 35900 24364
rect 35952 24352 35958 24404
rect 48038 24392 48044 24404
rect 36280 24364 48044 24392
rect 36280 24324 36308 24364
rect 48038 24352 48044 24364
rect 48096 24352 48102 24404
rect 27632 24296 36308 24324
rect 36446 24284 36452 24336
rect 36504 24324 36510 24336
rect 45002 24324 45008 24336
rect 36504 24296 45008 24324
rect 36504 24284 36510 24296
rect 45002 24284 45008 24296
rect 45060 24284 45066 24336
rect 28000 24228 28849 24256
rect 26053 24191 26111 24197
rect 26053 24157 26065 24191
rect 26099 24157 26111 24191
rect 26053 24151 26111 24157
rect 26142 24148 26148 24200
rect 26200 24188 26206 24200
rect 26237 24191 26295 24197
rect 26237 24188 26249 24191
rect 26200 24160 26249 24188
rect 26200 24148 26206 24160
rect 26237 24157 26249 24160
rect 26283 24157 26295 24191
rect 26237 24151 26295 24157
rect 26697 24191 26755 24197
rect 26697 24157 26709 24191
rect 26743 24188 26755 24191
rect 27890 24188 27896 24200
rect 26743 24160 27896 24188
rect 26743 24157 26755 24160
rect 26697 24151 26755 24157
rect 27890 24148 27896 24160
rect 27948 24148 27954 24200
rect 26964 24123 27022 24129
rect 22152 24092 22197 24120
rect 24320 24092 26924 24120
rect 22152 24080 22158 24092
rect 14826 24052 14832 24064
rect 12299 24024 14412 24052
rect 14787 24024 14832 24052
rect 12299 24021 12311 24024
rect 12253 24015 12311 24021
rect 14826 24012 14832 24024
rect 14884 24012 14890 24064
rect 15473 24055 15531 24061
rect 15473 24021 15485 24055
rect 15519 24052 15531 24055
rect 15562 24052 15568 24064
rect 15519 24024 15568 24052
rect 15519 24021 15531 24024
rect 15473 24015 15531 24021
rect 15562 24012 15568 24024
rect 15620 24012 15626 24064
rect 17402 24052 17408 24064
rect 17363 24024 17408 24052
rect 17402 24012 17408 24024
rect 17460 24012 17466 24064
rect 18046 24052 18052 24064
rect 18007 24024 18052 24052
rect 18046 24012 18052 24024
rect 18104 24012 18110 24064
rect 20809 24055 20867 24061
rect 20809 24021 20821 24055
rect 20855 24052 20867 24055
rect 21174 24052 21180 24064
rect 20855 24024 21180 24052
rect 20855 24021 20867 24024
rect 20809 24015 20867 24021
rect 21174 24012 21180 24024
rect 21232 24012 21238 24064
rect 24489 24055 24547 24061
rect 24489 24021 24501 24055
rect 24535 24052 24547 24055
rect 24854 24052 24860 24064
rect 24535 24024 24860 24052
rect 24535 24021 24547 24024
rect 24489 24015 24547 24021
rect 24854 24012 24860 24024
rect 24912 24012 24918 24064
rect 25498 24012 25504 24064
rect 25556 24052 25562 24064
rect 26050 24052 26056 24064
rect 25556 24024 26056 24052
rect 25556 24012 25562 24024
rect 26050 24012 26056 24024
rect 26108 24012 26114 24064
rect 26145 24055 26203 24061
rect 26145 24021 26157 24055
rect 26191 24052 26203 24055
rect 26786 24052 26792 24064
rect 26191 24024 26792 24052
rect 26191 24021 26203 24024
rect 26145 24015 26203 24021
rect 26786 24012 26792 24024
rect 26844 24012 26850 24064
rect 26896 24052 26924 24092
rect 26964 24089 26976 24123
rect 27010 24120 27022 24123
rect 27062 24120 27068 24132
rect 27010 24092 27068 24120
rect 27010 24089 27022 24092
rect 26964 24083 27022 24089
rect 27062 24080 27068 24092
rect 27120 24080 27126 24132
rect 28000 24120 28028 24228
rect 28537 24191 28595 24197
rect 28537 24188 28549 24191
rect 27172 24092 28028 24120
rect 28092 24160 28549 24188
rect 27172 24052 27200 24092
rect 26896 24024 27200 24052
rect 27522 24012 27528 24064
rect 27580 24052 27586 24064
rect 28092 24061 28120 24160
rect 28537 24157 28549 24160
rect 28583 24157 28595 24191
rect 28718 24188 28724 24200
rect 28679 24160 28724 24188
rect 28537 24151 28595 24157
rect 28718 24148 28724 24160
rect 28776 24148 28782 24200
rect 28821 24188 28849 24228
rect 28902 24216 28908 24268
rect 28960 24256 28966 24268
rect 31294 24256 31300 24268
rect 28960 24228 31300 24256
rect 28960 24216 28966 24228
rect 31294 24216 31300 24228
rect 31352 24216 31358 24268
rect 31570 24216 31576 24268
rect 31628 24256 31634 24268
rect 37642 24256 37648 24268
rect 31628 24228 33732 24256
rect 37603 24228 37648 24256
rect 31628 24216 31634 24228
rect 28821 24160 31754 24188
rect 28902 24080 28908 24132
rect 28960 24120 28966 24132
rect 30009 24123 30067 24129
rect 30009 24120 30021 24123
rect 28960 24092 30021 24120
rect 28960 24080 28966 24092
rect 30009 24089 30021 24092
rect 30055 24089 30067 24123
rect 30009 24083 30067 24089
rect 31113 24123 31171 24129
rect 31113 24089 31125 24123
rect 31159 24120 31171 24123
rect 31386 24120 31392 24132
rect 31159 24092 31392 24120
rect 31159 24089 31171 24092
rect 31113 24083 31171 24089
rect 31386 24080 31392 24092
rect 31444 24080 31450 24132
rect 31726 24120 31754 24160
rect 32858 24148 32864 24200
rect 32916 24188 32922 24200
rect 33704 24197 33732 24228
rect 37642 24216 37648 24228
rect 37700 24216 37706 24268
rect 46290 24256 46296 24268
rect 46251 24228 46296 24256
rect 46290 24216 46296 24228
rect 46348 24216 46354 24268
rect 46477 24259 46535 24265
rect 46477 24225 46489 24259
rect 46523 24256 46535 24259
rect 47670 24256 47676 24268
rect 46523 24228 47676 24256
rect 46523 24225 46535 24228
rect 46477 24219 46535 24225
rect 47670 24216 47676 24228
rect 47728 24216 47734 24268
rect 48130 24256 48136 24268
rect 48091 24228 48136 24256
rect 48130 24216 48136 24228
rect 48188 24216 48194 24268
rect 33597 24191 33655 24197
rect 33597 24188 33609 24191
rect 32916 24160 33609 24188
rect 32916 24148 32922 24160
rect 33597 24157 33609 24160
rect 33643 24157 33655 24191
rect 33597 24151 33655 24157
rect 33689 24191 33747 24197
rect 33689 24157 33701 24191
rect 33735 24157 33747 24191
rect 33689 24151 33747 24157
rect 33778 24148 33784 24200
rect 33836 24188 33842 24200
rect 33965 24191 34023 24197
rect 33836 24160 33929 24188
rect 33836 24148 33842 24160
rect 33965 24157 33977 24191
rect 34011 24188 34023 24191
rect 35069 24191 35127 24197
rect 35069 24188 35081 24191
rect 34011 24160 35081 24188
rect 34011 24157 34023 24160
rect 33965 24151 34023 24157
rect 35069 24157 35081 24160
rect 35115 24157 35127 24191
rect 35069 24151 35127 24157
rect 35529 24191 35587 24197
rect 35529 24157 35541 24191
rect 35575 24188 35587 24191
rect 36722 24188 36728 24200
rect 35575 24160 36728 24188
rect 35575 24157 35587 24160
rect 35529 24151 35587 24157
rect 36722 24148 36728 24160
rect 36780 24148 36786 24200
rect 37461 24191 37519 24197
rect 37461 24157 37473 24191
rect 37507 24157 37519 24191
rect 37461 24151 37519 24157
rect 33226 24120 33232 24132
rect 31726 24092 33232 24120
rect 33226 24080 33232 24092
rect 33284 24080 33290 24132
rect 28077 24055 28135 24061
rect 28077 24052 28089 24055
rect 27580 24024 28089 24052
rect 27580 24012 27586 24024
rect 28077 24021 28089 24024
rect 28123 24021 28135 24055
rect 28626 24052 28632 24064
rect 28587 24024 28632 24052
rect 28077 24015 28135 24021
rect 28626 24012 28632 24024
rect 28684 24012 28690 24064
rect 30098 24012 30104 24064
rect 30156 24052 30162 24064
rect 33796 24052 33824 24148
rect 34514 24080 34520 24132
rect 34572 24120 34578 24132
rect 34701 24123 34759 24129
rect 34701 24120 34713 24123
rect 34572 24092 34713 24120
rect 34572 24080 34578 24092
rect 34701 24089 34713 24092
rect 34747 24089 34759 24123
rect 34882 24120 34888 24132
rect 34843 24092 34888 24120
rect 34701 24083 34759 24089
rect 30156 24024 33824 24052
rect 34716 24052 34744 24083
rect 34882 24080 34888 24092
rect 34940 24120 34946 24132
rect 35710 24120 35716 24132
rect 34940 24092 35716 24120
rect 34940 24080 34946 24092
rect 35710 24080 35716 24092
rect 35768 24120 35774 24132
rect 35986 24120 35992 24132
rect 35768 24092 35992 24120
rect 35768 24080 35774 24092
rect 35986 24080 35992 24092
rect 36044 24080 36050 24132
rect 37476 24052 37504 24151
rect 39298 24120 39304 24132
rect 39259 24092 39304 24120
rect 39298 24080 39304 24092
rect 39356 24080 39362 24132
rect 34716 24024 37504 24052
rect 30156 24012 30162 24024
rect 1104 23962 48852 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 48852 23962
rect 1104 23888 48852 23910
rect 8846 23848 8852 23860
rect 8807 23820 8852 23848
rect 8846 23808 8852 23820
rect 8904 23808 8910 23860
rect 10965 23851 11023 23857
rect 10965 23817 10977 23851
rect 11011 23848 11023 23851
rect 12894 23848 12900 23860
rect 11011 23820 12900 23848
rect 11011 23817 11023 23820
rect 10965 23811 11023 23817
rect 12894 23808 12900 23820
rect 12952 23808 12958 23860
rect 13814 23808 13820 23860
rect 13872 23848 13878 23860
rect 14001 23851 14059 23857
rect 14001 23848 14013 23851
rect 13872 23820 14013 23848
rect 13872 23808 13878 23820
rect 14001 23817 14013 23820
rect 14047 23817 14059 23851
rect 14001 23811 14059 23817
rect 14826 23808 14832 23860
rect 14884 23848 14890 23860
rect 15765 23851 15823 23857
rect 15765 23848 15777 23851
rect 14884 23820 15777 23848
rect 14884 23808 14890 23820
rect 15765 23817 15777 23820
rect 15811 23817 15823 23851
rect 16666 23848 16672 23860
rect 16627 23820 16672 23848
rect 15765 23811 15823 23817
rect 16666 23808 16672 23820
rect 16724 23808 16730 23860
rect 18230 23848 18236 23860
rect 17144 23820 18236 23848
rect 1486 23740 1492 23792
rect 1544 23780 1550 23792
rect 14274 23780 14280 23792
rect 1544 23752 12434 23780
rect 1544 23740 1550 23752
rect 8389 23715 8447 23721
rect 8389 23681 8401 23715
rect 8435 23712 8447 23715
rect 9214 23712 9220 23724
rect 8435 23684 9220 23712
rect 8435 23681 8447 23684
rect 8389 23675 8447 23681
rect 9214 23672 9220 23684
rect 9272 23672 9278 23724
rect 9309 23715 9367 23721
rect 9309 23681 9321 23715
rect 9355 23712 9367 23715
rect 9398 23712 9404 23724
rect 9355 23684 9404 23712
rect 9355 23681 9367 23684
rect 9309 23675 9367 23681
rect 9324 23576 9352 23675
rect 9398 23672 9404 23684
rect 9456 23672 9462 23724
rect 10229 23715 10287 23721
rect 10229 23681 10241 23715
rect 10275 23712 10287 23715
rect 10275 23684 10364 23712
rect 10275 23681 10287 23684
rect 10229 23675 10287 23681
rect 8680 23548 9352 23576
rect 10336 23576 10364 23684
rect 10410 23672 10416 23724
rect 10468 23712 10474 23724
rect 10594 23712 10600 23724
rect 10468 23684 10513 23712
rect 10555 23684 10600 23712
rect 10468 23672 10474 23684
rect 10594 23672 10600 23684
rect 10652 23672 10658 23724
rect 10778 23712 10784 23724
rect 10739 23684 10784 23712
rect 10778 23672 10784 23684
rect 10836 23672 10842 23724
rect 10870 23672 10876 23724
rect 10928 23712 10934 23724
rect 11517 23715 11575 23721
rect 11517 23712 11529 23715
rect 10928 23684 11529 23712
rect 10928 23672 10934 23684
rect 11517 23681 11529 23684
rect 11563 23681 11575 23715
rect 11698 23712 11704 23724
rect 11659 23684 11704 23712
rect 11517 23675 11575 23681
rect 11698 23672 11704 23684
rect 11756 23672 11762 23724
rect 11793 23715 11851 23721
rect 11793 23681 11805 23715
rect 11839 23681 11851 23715
rect 11900 23711 12020 23712
rect 11793 23675 11851 23681
rect 11890 23705 12020 23711
rect 10502 23644 10508 23656
rect 10463 23616 10508 23644
rect 10502 23604 10508 23616
rect 10560 23604 10566 23656
rect 10962 23604 10968 23656
rect 11020 23644 11026 23656
rect 11808 23644 11836 23675
rect 11890 23671 11902 23705
rect 11936 23684 12020 23705
rect 11936 23671 11948 23684
rect 11890 23665 11948 23671
rect 11020 23616 11836 23644
rect 11020 23604 11026 23616
rect 11517 23579 11575 23585
rect 11517 23576 11529 23579
rect 10336 23548 11529 23576
rect 2038 23508 2044 23520
rect 1999 23480 2044 23508
rect 2038 23468 2044 23480
rect 2096 23468 2102 23520
rect 8680 23517 8708 23548
rect 11517 23545 11529 23548
rect 11563 23545 11575 23579
rect 11517 23539 11575 23545
rect 8665 23511 8723 23517
rect 8665 23477 8677 23511
rect 8711 23477 8723 23511
rect 8665 23471 8723 23477
rect 9306 23468 9312 23520
rect 9364 23508 9370 23520
rect 9401 23511 9459 23517
rect 9401 23508 9413 23511
rect 9364 23480 9413 23508
rect 9364 23468 9370 23480
rect 9401 23477 9413 23480
rect 9447 23477 9459 23511
rect 9401 23471 9459 23477
rect 9769 23511 9827 23517
rect 9769 23477 9781 23511
rect 9815 23508 9827 23511
rect 10134 23508 10140 23520
rect 9815 23480 10140 23508
rect 9815 23477 9827 23480
rect 9769 23471 9827 23477
rect 10134 23468 10140 23480
rect 10192 23508 10198 23520
rect 10318 23508 10324 23520
rect 10192 23480 10324 23508
rect 10192 23468 10198 23480
rect 10318 23468 10324 23480
rect 10376 23468 10382 23520
rect 10410 23468 10416 23520
rect 10468 23508 10474 23520
rect 11992 23508 12020 23684
rect 12406 23644 12434 23752
rect 13832 23752 14280 23780
rect 12618 23712 12624 23724
rect 12579 23684 12624 23712
rect 12618 23672 12624 23684
rect 12676 23672 12682 23724
rect 13832 23721 13860 23752
rect 14274 23740 14280 23752
rect 14332 23740 14338 23792
rect 14642 23740 14648 23792
rect 14700 23780 14706 23792
rect 14918 23780 14924 23792
rect 14700 23752 14924 23780
rect 14700 23740 14706 23752
rect 14918 23740 14924 23752
rect 14976 23740 14982 23792
rect 15562 23780 15568 23792
rect 15523 23752 15568 23780
rect 15562 23740 15568 23752
rect 15620 23740 15626 23792
rect 17144 23780 17172 23820
rect 18230 23808 18236 23820
rect 18288 23808 18294 23860
rect 20254 23808 20260 23860
rect 20312 23848 20318 23860
rect 20806 23848 20812 23860
rect 20312 23820 20812 23848
rect 20312 23808 20318 23820
rect 20806 23808 20812 23820
rect 20864 23808 20870 23860
rect 27798 23848 27804 23860
rect 20916 23820 27614 23848
rect 27759 23820 27804 23848
rect 17052 23752 17172 23780
rect 13817 23715 13875 23721
rect 13817 23681 13829 23715
rect 13863 23681 13875 23715
rect 13817 23675 13875 23681
rect 14090 23672 14096 23724
rect 14148 23712 14154 23724
rect 14737 23715 14795 23721
rect 14148 23684 14193 23712
rect 14148 23672 14154 23684
rect 14737 23681 14749 23715
rect 14783 23712 14795 23715
rect 15286 23712 15292 23724
rect 14783 23684 15292 23712
rect 14783 23681 14795 23684
rect 14737 23675 14795 23681
rect 15286 23672 15292 23684
rect 15344 23672 15350 23724
rect 17052 23721 17080 23752
rect 18046 23740 18052 23792
rect 18104 23780 18110 23792
rect 18478 23783 18536 23789
rect 18478 23780 18490 23783
rect 18104 23752 18490 23780
rect 18104 23740 18110 23752
rect 18478 23749 18490 23752
rect 18524 23749 18536 23783
rect 18690 23780 18696 23792
rect 18478 23743 18536 23749
rect 18616 23752 18696 23780
rect 16945 23715 17003 23721
rect 16945 23681 16957 23715
rect 16991 23681 17003 23715
rect 16945 23675 17003 23681
rect 17037 23715 17095 23721
rect 17037 23681 17049 23715
rect 17083 23681 17095 23715
rect 17037 23675 17095 23681
rect 16960 23644 16988 23675
rect 17126 23672 17132 23724
rect 17184 23712 17190 23724
rect 17313 23715 17371 23721
rect 17184 23684 17229 23712
rect 17184 23672 17190 23684
rect 17313 23681 17325 23715
rect 17359 23712 17371 23715
rect 18138 23712 18144 23724
rect 17359 23684 18144 23712
rect 17359 23681 17371 23684
rect 17313 23675 17371 23681
rect 18138 23672 18144 23684
rect 18196 23712 18202 23724
rect 18616 23712 18644 23752
rect 18690 23740 18696 23752
rect 18748 23740 18754 23792
rect 20916 23721 20944 23820
rect 23474 23780 23480 23792
rect 22066 23752 23480 23780
rect 18196 23684 18644 23712
rect 20901 23715 20959 23721
rect 18196 23672 18202 23684
rect 20901 23681 20913 23715
rect 20947 23681 20959 23715
rect 20901 23675 20959 23681
rect 20993 23715 21051 23721
rect 20993 23681 21005 23715
rect 21039 23681 21051 23715
rect 20993 23675 21051 23681
rect 21090 23718 21148 23724
rect 21090 23684 21102 23718
rect 21136 23684 21148 23718
rect 21090 23678 21148 23684
rect 12406 23616 16988 23644
rect 17862 23604 17868 23656
rect 17920 23644 17926 23656
rect 18233 23647 18291 23653
rect 18233 23644 18245 23647
rect 17920 23616 18245 23644
rect 17920 23604 17926 23616
rect 18233 23613 18245 23616
rect 18279 23613 18291 23647
rect 18233 23607 18291 23613
rect 17310 23536 17316 23588
rect 17368 23576 17374 23588
rect 17880 23576 17908 23604
rect 17368 23548 17908 23576
rect 17368 23536 17374 23548
rect 20898 23536 20904 23588
rect 20956 23576 20962 23588
rect 21008 23576 21036 23675
rect 21102 23644 21130 23678
rect 21266 23672 21272 23724
rect 21324 23712 21330 23724
rect 21324 23684 21369 23712
rect 21324 23672 21330 23684
rect 21818 23672 21824 23724
rect 21876 23712 21882 23724
rect 22066 23712 22094 23752
rect 22480 23721 22508 23752
rect 23474 23740 23480 23752
rect 23532 23740 23538 23792
rect 24305 23783 24363 23789
rect 24305 23749 24317 23783
rect 24351 23749 24363 23783
rect 24854 23780 24860 23792
rect 24305 23743 24363 23749
rect 24679 23752 24860 23780
rect 21876 23684 22094 23712
rect 22465 23715 22523 23721
rect 21876 23672 21882 23684
rect 22465 23681 22477 23715
rect 22511 23712 22523 23715
rect 22732 23715 22790 23721
rect 22511 23684 22545 23712
rect 22511 23681 22523 23684
rect 22465 23675 22523 23681
rect 22732 23681 22744 23715
rect 22778 23712 22790 23715
rect 24320 23712 24348 23743
rect 22778 23684 24348 23712
rect 22778 23681 22790 23684
rect 22732 23675 22790 23681
rect 24486 23672 24492 23724
rect 24544 23712 24550 23724
rect 24679 23721 24707 23752
rect 24854 23740 24860 23752
rect 24912 23740 24918 23792
rect 25409 23783 25467 23789
rect 25409 23749 25421 23783
rect 25455 23780 25467 23783
rect 25498 23780 25504 23792
rect 25455 23752 25504 23780
rect 25455 23749 25467 23752
rect 25409 23743 25467 23749
rect 25498 23740 25504 23752
rect 25556 23740 25562 23792
rect 27586 23780 27614 23820
rect 27798 23808 27804 23820
rect 27856 23808 27862 23860
rect 27890 23808 27896 23860
rect 27948 23848 27954 23860
rect 28902 23848 28908 23860
rect 27948 23820 28908 23848
rect 27948 23808 27954 23820
rect 28902 23808 28908 23820
rect 28960 23808 28966 23860
rect 29638 23848 29644 23860
rect 29599 23820 29644 23848
rect 29638 23808 29644 23820
rect 29696 23808 29702 23860
rect 31570 23808 31576 23860
rect 31628 23848 31634 23860
rect 48041 23851 48099 23857
rect 48041 23848 48053 23851
rect 31628 23820 48053 23848
rect 31628 23808 31634 23820
rect 48041 23817 48053 23820
rect 48087 23817 48099 23851
rect 48041 23811 48099 23817
rect 33778 23780 33784 23792
rect 27586 23752 33784 23780
rect 33778 23740 33784 23752
rect 33836 23740 33842 23792
rect 35342 23740 35348 23792
rect 35400 23780 35406 23792
rect 47486 23780 47492 23792
rect 35400 23752 47492 23780
rect 35400 23740 35406 23752
rect 47486 23740 47492 23752
rect 47544 23740 47550 23792
rect 47946 23780 47952 23792
rect 47907 23752 47952 23780
rect 47946 23740 47952 23752
rect 48004 23740 48010 23792
rect 34906 23724 34964 23727
rect 24581 23715 24639 23721
rect 24581 23712 24593 23715
rect 24544 23684 24593 23712
rect 24544 23672 24550 23684
rect 24581 23681 24593 23684
rect 24627 23681 24639 23715
rect 24581 23675 24639 23681
rect 24670 23715 24728 23721
rect 24670 23681 24682 23715
rect 24716 23681 24728 23715
rect 24670 23675 24728 23681
rect 24765 23715 24823 23721
rect 24765 23681 24777 23715
rect 24811 23681 24823 23715
rect 24765 23675 24823 23681
rect 24949 23715 25007 23721
rect 24949 23681 24961 23715
rect 24995 23712 25007 23715
rect 25038 23712 25044 23724
rect 24995 23684 25044 23712
rect 24995 23681 25007 23684
rect 24949 23675 25007 23681
rect 21174 23644 21180 23656
rect 21102 23616 21180 23644
rect 21174 23604 21180 23616
rect 21232 23604 21238 23656
rect 24118 23604 24124 23656
rect 24176 23644 24182 23656
rect 24780 23644 24808 23675
rect 25038 23672 25044 23684
rect 25096 23672 25102 23724
rect 25590 23712 25596 23724
rect 25551 23684 25596 23712
rect 25590 23672 25596 23684
rect 25648 23672 25654 23724
rect 27433 23715 27491 23721
rect 27433 23681 27445 23715
rect 27479 23712 27491 23715
rect 27522 23712 27528 23724
rect 27479 23684 27528 23712
rect 27479 23681 27491 23684
rect 27433 23675 27491 23681
rect 27522 23672 27528 23684
rect 27580 23672 27586 23724
rect 27617 23715 27675 23721
rect 27617 23681 27629 23715
rect 27663 23712 27675 23715
rect 28994 23712 29000 23724
rect 27663 23684 29000 23712
rect 27663 23681 27675 23684
rect 27617 23675 27675 23681
rect 28994 23672 29000 23684
rect 29052 23712 29058 23724
rect 29825 23715 29883 23721
rect 29825 23712 29837 23715
rect 29052 23684 29837 23712
rect 29052 23672 29058 23684
rect 29825 23681 29837 23684
rect 29871 23681 29883 23715
rect 29825 23675 29883 23681
rect 30006 23672 30012 23724
rect 30064 23712 30070 23724
rect 30101 23715 30159 23721
rect 30101 23712 30113 23715
rect 30064 23684 30113 23712
rect 30064 23672 30070 23684
rect 30101 23681 30113 23684
rect 30147 23681 30159 23715
rect 30101 23675 30159 23681
rect 30650 23672 30656 23724
rect 30708 23712 30714 23724
rect 31021 23715 31079 23721
rect 31021 23712 31033 23715
rect 30708 23684 31033 23712
rect 30708 23672 30714 23684
rect 31021 23681 31033 23684
rect 31067 23681 31079 23715
rect 31021 23675 31079 23681
rect 31297 23715 31355 23721
rect 31297 23681 31309 23715
rect 31343 23712 31355 23715
rect 31662 23712 31668 23724
rect 31343 23684 31668 23712
rect 31343 23681 31355 23684
rect 31297 23675 31355 23681
rect 31662 23672 31668 23684
rect 31720 23672 31726 23724
rect 32122 23712 32128 23724
rect 32083 23684 32128 23712
rect 32122 23672 32128 23684
rect 32180 23672 32186 23724
rect 32214 23672 32220 23724
rect 32272 23712 32278 23724
rect 33042 23712 33048 23724
rect 32272 23684 33048 23712
rect 32272 23672 32278 23684
rect 33042 23672 33048 23684
rect 33100 23712 33106 23724
rect 33321 23715 33379 23721
rect 33321 23712 33333 23715
rect 33100 23684 33333 23712
rect 33100 23672 33106 23684
rect 33321 23681 33333 23684
rect 33367 23712 33379 23715
rect 34514 23712 34520 23724
rect 33367 23684 34520 23712
rect 33367 23681 33379 23684
rect 33321 23675 33379 23681
rect 34514 23672 34520 23684
rect 34572 23672 34578 23724
rect 34606 23672 34612 23724
rect 34664 23712 34670 23724
rect 34906 23721 34949 23724
rect 34701 23715 34759 23721
rect 34701 23712 34713 23715
rect 34664 23684 34713 23712
rect 34664 23672 34670 23684
rect 34701 23681 34713 23684
rect 34747 23681 34759 23715
rect 34806 23715 34864 23721
rect 34806 23708 34818 23715
rect 34701 23675 34759 23681
rect 34790 23656 34796 23708
rect 34852 23681 34864 23715
rect 34906 23687 34918 23721
rect 34906 23681 34949 23687
rect 34848 23675 34864 23681
rect 34848 23656 34854 23675
rect 34943 23672 34949 23681
rect 35001 23672 35007 23724
rect 35069 23716 35127 23721
rect 35069 23715 35265 23716
rect 35069 23681 35081 23715
rect 35115 23712 35265 23715
rect 35529 23715 35587 23721
rect 35618 23715 35624 23724
rect 35115 23688 35449 23712
rect 35115 23681 35127 23688
rect 35237 23684 35449 23688
rect 35069 23675 35127 23681
rect 24176 23616 24808 23644
rect 24176 23604 24182 23616
rect 25498 23604 25504 23656
rect 25556 23644 25562 23656
rect 28626 23644 28632 23656
rect 25556 23616 28632 23644
rect 25556 23604 25562 23616
rect 28626 23604 28632 23616
rect 28684 23604 28690 23656
rect 30374 23644 30380 23656
rect 28736 23616 30380 23644
rect 20956 23548 21036 23576
rect 20956 23536 20962 23548
rect 23566 23536 23572 23588
rect 23624 23576 23630 23588
rect 23845 23579 23903 23585
rect 23845 23576 23857 23579
rect 23624 23548 23857 23576
rect 23624 23536 23630 23548
rect 23845 23545 23857 23548
rect 23891 23576 23903 23579
rect 24486 23576 24492 23588
rect 23891 23548 24492 23576
rect 23891 23545 23903 23548
rect 23845 23539 23903 23545
rect 24486 23536 24492 23548
rect 24544 23536 24550 23588
rect 27706 23536 27712 23588
rect 27764 23576 27770 23588
rect 28258 23576 28264 23588
rect 27764 23548 28264 23576
rect 27764 23536 27770 23548
rect 28258 23536 28264 23548
rect 28316 23536 28322 23588
rect 10468 23480 12020 23508
rect 10468 23468 10474 23480
rect 12434 23468 12440 23520
rect 12492 23508 12498 23520
rect 13633 23511 13691 23517
rect 12492 23480 12537 23508
rect 12492 23468 12498 23480
rect 13633 23477 13645 23511
rect 13679 23508 13691 23511
rect 14366 23508 14372 23520
rect 13679 23480 14372 23508
rect 13679 23477 13691 23480
rect 13633 23471 13691 23477
rect 14366 23468 14372 23480
rect 14424 23468 14430 23520
rect 15105 23511 15163 23517
rect 15105 23477 15117 23511
rect 15151 23508 15163 23511
rect 15749 23511 15807 23517
rect 15749 23508 15761 23511
rect 15151 23480 15761 23508
rect 15151 23477 15163 23480
rect 15105 23471 15163 23477
rect 15749 23477 15761 23480
rect 15795 23477 15807 23511
rect 15930 23508 15936 23520
rect 15891 23480 15936 23508
rect 15749 23471 15807 23477
rect 15930 23468 15936 23480
rect 15988 23468 15994 23520
rect 19518 23468 19524 23520
rect 19576 23508 19582 23520
rect 19613 23511 19671 23517
rect 19613 23508 19625 23511
rect 19576 23480 19625 23508
rect 19576 23468 19582 23480
rect 19613 23477 19625 23480
rect 19659 23477 19671 23511
rect 19613 23471 19671 23477
rect 20625 23511 20683 23517
rect 20625 23477 20637 23511
rect 20671 23508 20683 23511
rect 20714 23508 20720 23520
rect 20671 23480 20720 23508
rect 20671 23477 20683 23480
rect 20625 23471 20683 23477
rect 20714 23468 20720 23480
rect 20772 23468 20778 23520
rect 24762 23468 24768 23520
rect 24820 23508 24826 23520
rect 25777 23511 25835 23517
rect 25777 23508 25789 23511
rect 24820 23480 25789 23508
rect 24820 23468 24826 23480
rect 25777 23477 25789 23480
rect 25823 23477 25835 23511
rect 25777 23471 25835 23477
rect 25866 23468 25872 23520
rect 25924 23508 25930 23520
rect 28736 23508 28764 23616
rect 30374 23604 30380 23616
rect 30432 23604 30438 23656
rect 30466 23604 30472 23656
rect 30524 23644 30530 23656
rect 30742 23644 30748 23656
rect 30524 23616 30748 23644
rect 30524 23604 30530 23616
rect 30742 23604 30748 23616
rect 30800 23604 30806 23656
rect 31205 23647 31263 23653
rect 31205 23613 31217 23647
rect 31251 23644 31263 23647
rect 32582 23644 32588 23656
rect 31251 23616 32588 23644
rect 31251 23613 31263 23616
rect 31205 23607 31263 23613
rect 32582 23604 32588 23616
rect 32640 23604 32646 23656
rect 35421 23644 35449 23684
rect 35529 23681 35541 23715
rect 35575 23687 35624 23715
rect 35575 23681 35587 23687
rect 35529 23675 35587 23681
rect 35618 23672 35624 23687
rect 35676 23672 35682 23724
rect 35721 23715 35779 23721
rect 35721 23681 35733 23715
rect 35767 23712 35779 23715
rect 35986 23712 35992 23724
rect 35767 23684 35992 23712
rect 35767 23681 35779 23684
rect 35721 23675 35779 23681
rect 35986 23672 35992 23684
rect 36044 23672 36050 23724
rect 36722 23672 36728 23724
rect 36780 23712 36786 23724
rect 37369 23715 37427 23721
rect 37369 23712 37381 23715
rect 36780 23684 37381 23712
rect 36780 23672 36786 23684
rect 37369 23681 37381 23684
rect 37415 23681 37427 23715
rect 37369 23675 37427 23681
rect 37553 23647 37611 23653
rect 35421 23616 35940 23644
rect 29914 23536 29920 23588
rect 29972 23576 29978 23588
rect 31481 23579 31539 23585
rect 31481 23576 31493 23579
rect 29972 23548 31493 23576
rect 29972 23536 29978 23548
rect 31481 23545 31493 23548
rect 31527 23545 31539 23579
rect 31481 23539 31539 23545
rect 33778 23536 33784 23588
rect 33836 23576 33842 23588
rect 35342 23576 35348 23588
rect 33836 23548 35348 23576
rect 33836 23536 33842 23548
rect 35342 23536 35348 23548
rect 35400 23536 35406 23588
rect 35912 23585 35940 23616
rect 37553 23613 37565 23647
rect 37599 23644 37611 23647
rect 38194 23644 38200 23656
rect 37599 23616 38200 23644
rect 37599 23613 37611 23616
rect 37553 23607 37611 23613
rect 38194 23604 38200 23616
rect 38252 23604 38258 23656
rect 39209 23647 39267 23653
rect 39209 23613 39221 23647
rect 39255 23644 39267 23647
rect 43438 23644 43444 23656
rect 39255 23616 43444 23644
rect 39255 23613 39267 23616
rect 39209 23607 39267 23613
rect 43438 23604 43444 23616
rect 43496 23604 43502 23656
rect 35897 23579 35955 23585
rect 35897 23545 35909 23579
rect 35943 23545 35955 23579
rect 35897 23539 35955 23545
rect 36078 23536 36084 23588
rect 36136 23576 36142 23588
rect 46658 23576 46664 23588
rect 36136 23548 46664 23576
rect 36136 23536 36142 23548
rect 46658 23536 46664 23548
rect 46716 23536 46722 23588
rect 25924 23480 28764 23508
rect 30285 23511 30343 23517
rect 25924 23468 25930 23480
rect 30285 23477 30297 23511
rect 30331 23508 30343 23511
rect 30558 23508 30564 23520
rect 30331 23480 30564 23508
rect 30331 23477 30343 23480
rect 30285 23471 30343 23477
rect 30558 23468 30564 23480
rect 30616 23468 30622 23520
rect 30742 23468 30748 23520
rect 30800 23508 30806 23520
rect 31018 23508 31024 23520
rect 30800 23480 31024 23508
rect 30800 23468 30806 23480
rect 31018 23468 31024 23480
rect 31076 23468 31082 23520
rect 34425 23511 34483 23517
rect 34425 23477 34437 23511
rect 34471 23508 34483 23511
rect 34790 23508 34796 23520
rect 34471 23480 34796 23508
rect 34471 23477 34483 23480
rect 34425 23471 34483 23477
rect 34790 23468 34796 23480
rect 34848 23468 34854 23520
rect 35526 23468 35532 23520
rect 35584 23508 35590 23520
rect 45554 23508 45560 23520
rect 35584 23480 45560 23508
rect 35584 23468 35590 23480
rect 45554 23468 45560 23480
rect 45612 23468 45618 23520
rect 1104 23418 48852 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 48852 23418
rect 1104 23344 48852 23366
rect 1578 23264 1584 23316
rect 1636 23304 1642 23316
rect 1636 23276 25544 23304
rect 1636 23264 1642 23276
rect 10597 23239 10655 23245
rect 10597 23205 10609 23239
rect 10643 23236 10655 23239
rect 11698 23236 11704 23248
rect 10643 23208 11704 23236
rect 10643 23205 10655 23208
rect 10597 23199 10655 23205
rect 11698 23196 11704 23208
rect 11756 23196 11762 23248
rect 13357 23239 13415 23245
rect 13357 23205 13369 23239
rect 13403 23205 13415 23239
rect 16853 23239 16911 23245
rect 13357 23199 13415 23205
rect 14568 23208 16804 23236
rect 1397 23171 1455 23177
rect 1397 23137 1409 23171
rect 1443 23168 1455 23171
rect 2038 23168 2044 23180
rect 1443 23140 2044 23168
rect 1443 23137 1455 23140
rect 1397 23131 1455 23137
rect 2038 23128 2044 23140
rect 2096 23128 2102 23180
rect 2774 23128 2780 23180
rect 2832 23168 2838 23180
rect 10318 23168 10324 23180
rect 2832 23140 2877 23168
rect 10279 23140 10324 23168
rect 2832 23128 2838 23140
rect 10318 23128 10324 23140
rect 10376 23128 10382 23180
rect 10413 23171 10471 23177
rect 10413 23137 10425 23171
rect 10459 23168 10471 23171
rect 11882 23168 11888 23180
rect 10459 23140 11888 23168
rect 10459 23137 10471 23140
rect 10413 23131 10471 23137
rect 11882 23128 11888 23140
rect 11940 23128 11946 23180
rect 13262 23128 13268 23180
rect 13320 23168 13326 23180
rect 13372 23168 13400 23199
rect 14093 23171 14151 23177
rect 14093 23168 14105 23171
rect 13320 23140 14105 23168
rect 13320 23128 13326 23140
rect 14093 23137 14105 23140
rect 14139 23137 14151 23171
rect 14568 23168 14596 23208
rect 15654 23168 15660 23180
rect 14093 23131 14151 23137
rect 14200 23140 14596 23168
rect 15615 23140 15660 23168
rect 9953 23103 10011 23109
rect 9953 23069 9965 23103
rect 9999 23100 10011 23103
rect 10778 23100 10784 23112
rect 9999 23072 10784 23100
rect 9999 23069 10011 23072
rect 9953 23063 10011 23069
rect 10778 23060 10784 23072
rect 10836 23060 10842 23112
rect 11977 23103 12035 23109
rect 11977 23069 11989 23103
rect 12023 23100 12035 23103
rect 12986 23100 12992 23112
rect 12023 23072 12992 23100
rect 12023 23069 12035 23072
rect 11977 23063 12035 23069
rect 12986 23060 12992 23072
rect 13044 23060 13050 23112
rect 13078 23060 13084 23112
rect 13136 23100 13142 23112
rect 14200 23100 14228 23140
rect 15654 23128 15660 23140
rect 15712 23128 15718 23180
rect 16574 23128 16580 23180
rect 16632 23168 16638 23180
rect 16632 23140 16712 23168
rect 16632 23128 16638 23140
rect 13136 23072 14228 23100
rect 13136 23060 13142 23072
rect 14274 23060 14280 23112
rect 14332 23100 14338 23112
rect 14369 23103 14427 23109
rect 14369 23100 14381 23103
rect 14332 23072 14381 23100
rect 14332 23060 14338 23072
rect 14369 23069 14381 23072
rect 14415 23069 14427 23103
rect 14369 23063 14427 23069
rect 14734 23060 14740 23112
rect 14792 23100 14798 23112
rect 16684 23109 16712 23140
rect 15565 23103 15623 23109
rect 15565 23100 15577 23103
rect 14792 23072 15577 23100
rect 14792 23060 14798 23072
rect 15565 23069 15577 23072
rect 15611 23069 15623 23103
rect 15565 23063 15623 23069
rect 16669 23103 16727 23109
rect 16669 23069 16681 23103
rect 16715 23069 16727 23103
rect 16669 23063 16727 23069
rect 1581 23035 1639 23041
rect 1581 23001 1593 23035
rect 1627 23032 1639 23035
rect 2590 23032 2596 23044
rect 1627 23004 2596 23032
rect 1627 23001 1639 23004
rect 1581 22995 1639 23001
rect 2590 22992 2596 23004
rect 2648 22992 2654 23044
rect 12244 23035 12302 23041
rect 12244 23001 12256 23035
rect 12290 23032 12302 23035
rect 12434 23032 12440 23044
rect 12290 23004 12440 23032
rect 12290 23001 12302 23004
rect 12244 22995 12302 23001
rect 12434 22992 12440 23004
rect 12492 22992 12498 23044
rect 16485 23035 16543 23041
rect 14384 23004 16068 23032
rect 6914 22924 6920 22976
rect 6972 22964 6978 22976
rect 14384 22964 14412 23004
rect 6972 22936 14412 22964
rect 6972 22924 6978 22936
rect 14458 22924 14464 22976
rect 14516 22964 14522 22976
rect 15933 22967 15991 22973
rect 15933 22964 15945 22967
rect 14516 22936 15945 22964
rect 14516 22924 14522 22936
rect 15933 22933 15945 22936
rect 15979 22933 15991 22967
rect 16040 22964 16068 23004
rect 16485 23001 16497 23035
rect 16531 23032 16543 23035
rect 16574 23032 16580 23044
rect 16531 23004 16580 23032
rect 16531 23001 16543 23004
rect 16485 22995 16543 23001
rect 16574 22992 16580 23004
rect 16632 22992 16638 23044
rect 16776 23032 16804 23208
rect 16853 23205 16865 23239
rect 16899 23236 16911 23239
rect 17126 23236 17132 23248
rect 16899 23208 17132 23236
rect 16899 23205 16911 23208
rect 16853 23199 16911 23205
rect 17126 23196 17132 23208
rect 17184 23196 17190 23248
rect 19426 23196 19432 23248
rect 19484 23236 19490 23248
rect 19613 23239 19671 23245
rect 19613 23236 19625 23239
rect 19484 23208 19625 23236
rect 19484 23196 19490 23208
rect 19613 23205 19625 23208
rect 19659 23205 19671 23239
rect 25516 23236 25544 23276
rect 25590 23264 25596 23316
rect 25648 23304 25654 23316
rect 25777 23307 25835 23313
rect 25777 23304 25789 23307
rect 25648 23276 25789 23304
rect 25648 23264 25654 23276
rect 25777 23273 25789 23276
rect 25823 23304 25835 23307
rect 25866 23304 25872 23316
rect 25823 23276 25872 23304
rect 25823 23273 25835 23276
rect 25777 23267 25835 23273
rect 25866 23264 25872 23276
rect 25924 23264 25930 23316
rect 27062 23264 27068 23316
rect 27120 23304 27126 23316
rect 27433 23307 27491 23313
rect 27433 23304 27445 23307
rect 27120 23276 27445 23304
rect 27120 23264 27126 23276
rect 27433 23273 27445 23276
rect 27479 23273 27491 23307
rect 27433 23267 27491 23273
rect 29917 23307 29975 23313
rect 29917 23273 29929 23307
rect 29963 23304 29975 23307
rect 31110 23304 31116 23316
rect 29963 23276 31116 23304
rect 29963 23273 29975 23276
rect 29917 23267 29975 23273
rect 31110 23264 31116 23276
rect 31168 23264 31174 23316
rect 44174 23304 44180 23316
rect 31726 23276 44180 23304
rect 29362 23236 29368 23248
rect 25516 23208 29368 23236
rect 19613 23199 19671 23205
rect 29362 23196 29368 23208
rect 29420 23196 29426 23248
rect 29454 23196 29460 23248
rect 29512 23236 29518 23248
rect 31726 23236 31754 23276
rect 44174 23264 44180 23276
rect 44232 23264 44238 23316
rect 29512 23208 31754 23236
rect 29512 23196 29518 23208
rect 32950 23196 32956 23248
rect 33008 23236 33014 23248
rect 33686 23236 33692 23248
rect 33008 23208 33692 23236
rect 33008 23196 33014 23208
rect 33686 23196 33692 23208
rect 33744 23196 33750 23248
rect 17218 23128 17224 23180
rect 17276 23168 17282 23180
rect 17276 23140 17448 23168
rect 17276 23128 17282 23140
rect 16850 23060 16856 23112
rect 16908 23100 16914 23112
rect 17310 23100 17316 23112
rect 16908 23072 17316 23100
rect 16908 23060 16914 23072
rect 17310 23060 17316 23072
rect 17368 23060 17374 23112
rect 17420 23100 17448 23140
rect 23474 23128 23480 23180
rect 23532 23168 23538 23180
rect 24397 23171 24455 23177
rect 24397 23168 24409 23171
rect 23532 23140 24409 23168
rect 23532 23128 23538 23140
rect 24397 23137 24409 23140
rect 24443 23137 24455 23171
rect 29638 23168 29644 23180
rect 24397 23131 24455 23137
rect 26620 23140 29644 23168
rect 17569 23103 17627 23109
rect 17569 23100 17581 23103
rect 17420 23072 17581 23100
rect 17569 23069 17581 23072
rect 17615 23069 17627 23103
rect 17569 23063 17627 23069
rect 17862 23060 17868 23112
rect 17920 23100 17926 23112
rect 20441 23103 20499 23109
rect 20441 23100 20453 23103
rect 17920 23072 20453 23100
rect 17920 23060 17926 23072
rect 20441 23069 20453 23072
rect 20487 23100 20499 23103
rect 22281 23103 22339 23109
rect 22281 23100 22293 23103
rect 20487 23072 22293 23100
rect 20487 23069 20499 23072
rect 20441 23063 20499 23069
rect 22281 23069 22293 23072
rect 22327 23100 22339 23103
rect 22370 23100 22376 23112
rect 22327 23072 22376 23100
rect 22327 23069 22339 23072
rect 22281 23063 22339 23069
rect 22370 23060 22376 23072
rect 22428 23060 22434 23112
rect 23934 23060 23940 23112
rect 23992 23100 23998 23112
rect 26620 23100 26648 23140
rect 29638 23128 29644 23140
rect 29696 23168 29702 23180
rect 29733 23171 29791 23177
rect 29733 23168 29745 23171
rect 29696 23140 29745 23168
rect 29696 23128 29702 23140
rect 29733 23137 29745 23140
rect 29779 23137 29791 23171
rect 33962 23168 33968 23180
rect 29733 23131 29791 23137
rect 29840 23140 33968 23168
rect 26786 23100 26792 23112
rect 23992 23072 26648 23100
rect 26747 23072 26792 23100
rect 23992 23060 23998 23072
rect 26786 23060 26792 23072
rect 26844 23060 26850 23112
rect 26973 23103 27031 23109
rect 26973 23069 26985 23103
rect 27019 23100 27031 23103
rect 27062 23100 27068 23112
rect 27019 23072 27068 23100
rect 27019 23069 27031 23072
rect 26973 23063 27031 23069
rect 27062 23060 27068 23072
rect 27120 23100 27126 23112
rect 27430 23100 27436 23112
rect 27120 23072 27436 23100
rect 27120 23060 27126 23072
rect 27430 23060 27436 23072
rect 27488 23060 27494 23112
rect 27617 23103 27675 23109
rect 27617 23069 27629 23103
rect 27663 23100 27675 23103
rect 28074 23100 28080 23112
rect 27663 23072 28080 23100
rect 27663 23069 27675 23072
rect 27617 23063 27675 23069
rect 28074 23060 28080 23072
rect 28132 23060 28138 23112
rect 28537 23103 28595 23109
rect 28537 23069 28549 23103
rect 28583 23100 28595 23103
rect 28626 23100 28632 23112
rect 28583 23072 28632 23100
rect 28583 23069 28595 23072
rect 28537 23063 28595 23069
rect 28626 23060 28632 23072
rect 28684 23100 28690 23112
rect 29840 23100 29868 23140
rect 33962 23128 33968 23140
rect 34020 23128 34026 23180
rect 34698 23168 34704 23180
rect 34659 23140 34704 23168
rect 34698 23128 34704 23140
rect 34756 23128 34762 23180
rect 28684 23072 29868 23100
rect 29917 23103 29975 23109
rect 28684 23060 28690 23072
rect 29917 23069 29929 23103
rect 29963 23069 29975 23103
rect 29917 23063 29975 23069
rect 19150 23032 19156 23044
rect 16776 23004 19156 23032
rect 19150 22992 19156 23004
rect 19208 22992 19214 23044
rect 19245 23035 19303 23041
rect 19245 23001 19257 23035
rect 19291 23032 19303 23035
rect 19334 23032 19340 23044
rect 19291 23004 19340 23032
rect 19291 23001 19303 23004
rect 19245 22995 19303 23001
rect 19334 22992 19340 23004
rect 19392 22992 19398 23044
rect 19426 22992 19432 23044
rect 19484 23032 19490 23044
rect 20714 23041 20720 23044
rect 20708 23032 20720 23041
rect 19484 23004 19529 23032
rect 20675 23004 20720 23032
rect 19484 22992 19490 23004
rect 20708 22995 20720 23004
rect 20714 22992 20720 22995
rect 20772 22992 20778 23044
rect 20806 22992 20812 23044
rect 20864 23032 20870 23044
rect 22526 23035 22584 23041
rect 22526 23032 22538 23035
rect 20864 23004 22538 23032
rect 20864 22992 20870 23004
rect 22526 23001 22538 23004
rect 22572 23001 22584 23035
rect 22526 22995 22584 23001
rect 24664 23035 24722 23041
rect 24664 23001 24676 23035
rect 24710 23032 24722 23035
rect 24946 23032 24952 23044
rect 24710 23004 24952 23032
rect 24710 23001 24722 23004
rect 24664 22995 24722 23001
rect 24946 22992 24952 23004
rect 25004 22992 25010 23044
rect 27890 22992 27896 23044
rect 27948 23032 27954 23044
rect 28169 23035 28227 23041
rect 28169 23032 28181 23035
rect 27948 23004 28181 23032
rect 27948 22992 27954 23004
rect 28169 23001 28181 23004
rect 28215 23001 28227 23035
rect 28169 22995 28227 23001
rect 29362 22992 29368 23044
rect 29420 23032 29426 23044
rect 29641 23035 29699 23041
rect 29641 23032 29653 23035
rect 29420 23004 29653 23032
rect 29420 22992 29426 23004
rect 29641 23001 29653 23004
rect 29687 23001 29699 23035
rect 29641 22995 29699 23001
rect 29932 23032 29960 23063
rect 30558 23060 30564 23112
rect 30616 23100 30622 23112
rect 30653 23103 30711 23109
rect 30653 23100 30665 23103
rect 30616 23072 30665 23100
rect 30616 23060 30622 23072
rect 30653 23069 30665 23072
rect 30699 23100 30711 23103
rect 31757 23103 31815 23109
rect 31757 23100 31769 23103
rect 30699 23072 31769 23100
rect 30699 23069 30711 23072
rect 30653 23063 30711 23069
rect 31757 23069 31769 23072
rect 31803 23100 31815 23103
rect 32122 23100 32128 23112
rect 31803 23072 32128 23100
rect 31803 23069 31815 23072
rect 31757 23063 31815 23069
rect 32122 23060 32128 23072
rect 32180 23060 32186 23112
rect 32306 23060 32312 23112
rect 32364 23100 32370 23112
rect 33042 23100 33048 23112
rect 32364 23072 33048 23100
rect 32364 23060 32370 23072
rect 33042 23060 33048 23072
rect 33100 23100 33106 23112
rect 33321 23103 33379 23109
rect 33321 23100 33333 23103
rect 33100 23072 33333 23100
rect 33100 23060 33106 23072
rect 33321 23069 33333 23072
rect 33367 23069 33379 23103
rect 38286 23100 38292 23112
rect 33321 23063 33379 23069
rect 34440 23072 38292 23100
rect 29932 23004 30420 23032
rect 17954 22964 17960 22976
rect 16040 22936 17960 22964
rect 15933 22927 15991 22933
rect 17954 22924 17960 22936
rect 18012 22924 18018 22976
rect 18046 22924 18052 22976
rect 18104 22964 18110 22976
rect 18693 22967 18751 22973
rect 18693 22964 18705 22967
rect 18104 22936 18705 22964
rect 18104 22924 18110 22936
rect 18693 22933 18705 22936
rect 18739 22933 18751 22967
rect 18693 22927 18751 22933
rect 20622 22924 20628 22976
rect 20680 22964 20686 22976
rect 21821 22967 21879 22973
rect 21821 22964 21833 22967
rect 20680 22936 21833 22964
rect 20680 22924 20686 22936
rect 21821 22933 21833 22936
rect 21867 22933 21879 22967
rect 23658 22964 23664 22976
rect 23619 22936 23664 22964
rect 21821 22927 21879 22933
rect 23658 22924 23664 22936
rect 23716 22924 23722 22976
rect 25774 22924 25780 22976
rect 25832 22964 25838 22976
rect 29932 22964 29960 23004
rect 25832 22936 29960 22964
rect 30101 22967 30159 22973
rect 25832 22924 25838 22936
rect 30101 22933 30113 22967
rect 30147 22964 30159 22967
rect 30282 22964 30288 22976
rect 30147 22936 30288 22964
rect 30147 22933 30159 22936
rect 30101 22927 30159 22933
rect 30282 22924 30288 22936
rect 30340 22924 30346 22976
rect 30392 22964 30420 23004
rect 30466 22992 30472 23044
rect 30524 23032 30530 23044
rect 31021 23035 31079 23041
rect 31021 23032 31033 23035
rect 30524 23004 31033 23032
rect 30524 22992 30530 23004
rect 31021 23001 31033 23004
rect 31067 23001 31079 23035
rect 31021 22995 31079 23001
rect 30926 22964 30932 22976
rect 30392 22936 30932 22964
rect 30926 22924 30932 22936
rect 30984 22924 30990 22976
rect 31036 22964 31064 22995
rect 31110 22992 31116 23044
rect 31168 23032 31174 23044
rect 34440 23032 34468 23072
rect 38286 23060 38292 23072
rect 38344 23060 38350 23112
rect 48130 23100 48136 23112
rect 48091 23072 48136 23100
rect 48130 23060 48136 23072
rect 48188 23060 48194 23112
rect 31168 23004 34468 23032
rect 31168 22992 31174 23004
rect 34514 22992 34520 23044
rect 34572 23032 34578 23044
rect 34946 23035 35004 23041
rect 34946 23032 34958 23035
rect 34572 23004 34958 23032
rect 34572 22992 34578 23004
rect 34946 23001 34958 23004
rect 34992 23001 35004 23035
rect 34946 22995 35004 23001
rect 35820 23004 41414 23032
rect 32950 22964 32956 22976
rect 31036 22936 32956 22964
rect 32950 22924 32956 22936
rect 33008 22924 33014 22976
rect 33042 22924 33048 22976
rect 33100 22964 33106 22976
rect 35820 22964 35848 23004
rect 33100 22936 35848 22964
rect 33100 22924 33106 22936
rect 35894 22924 35900 22976
rect 35952 22964 35958 22976
rect 36081 22967 36139 22973
rect 36081 22964 36093 22967
rect 35952 22936 36093 22964
rect 35952 22924 35958 22936
rect 36081 22933 36093 22936
rect 36127 22933 36139 22967
rect 41386 22964 41414 23004
rect 46106 22964 46112 22976
rect 41386 22936 46112 22964
rect 36081 22927 36139 22933
rect 46106 22924 46112 22936
rect 46164 22924 46170 22976
rect 47578 22924 47584 22976
rect 47636 22964 47642 22976
rect 47949 22967 48007 22973
rect 47949 22964 47961 22967
rect 47636 22936 47961 22964
rect 47636 22924 47642 22936
rect 47949 22933 47961 22936
rect 47995 22933 48007 22967
rect 47949 22927 48007 22933
rect 1104 22874 48852 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 48852 22874
rect 1104 22800 48852 22822
rect 2590 22760 2596 22772
rect 2551 22732 2596 22760
rect 2590 22720 2596 22732
rect 2648 22720 2654 22772
rect 10594 22720 10600 22772
rect 10652 22760 10658 22772
rect 10965 22763 11023 22769
rect 10965 22760 10977 22763
rect 10652 22732 10977 22760
rect 10652 22720 10658 22732
rect 10965 22729 10977 22732
rect 11011 22729 11023 22763
rect 10965 22723 11023 22729
rect 13814 22720 13820 22772
rect 13872 22760 13878 22772
rect 14274 22760 14280 22772
rect 13872 22732 14280 22760
rect 13872 22720 13878 22732
rect 14274 22720 14280 22732
rect 14332 22720 14338 22772
rect 14458 22760 14464 22772
rect 14419 22732 14464 22760
rect 14458 22720 14464 22732
rect 14516 22720 14522 22772
rect 17218 22720 17224 22772
rect 17276 22760 17282 22772
rect 17865 22763 17923 22769
rect 17865 22760 17877 22763
rect 17276 22732 17877 22760
rect 17276 22720 17282 22732
rect 17865 22729 17877 22732
rect 17911 22729 17923 22763
rect 17865 22723 17923 22729
rect 17954 22720 17960 22772
rect 18012 22760 18018 22772
rect 23934 22760 23940 22772
rect 18012 22732 23940 22760
rect 18012 22720 18018 22732
rect 23934 22720 23940 22732
rect 23992 22720 23998 22772
rect 24029 22763 24087 22769
rect 24029 22729 24041 22763
rect 24075 22760 24087 22763
rect 24118 22760 24124 22772
rect 24075 22732 24124 22760
rect 24075 22729 24087 22732
rect 24029 22723 24087 22729
rect 24118 22720 24124 22732
rect 24176 22720 24182 22772
rect 25222 22760 25228 22772
rect 24780 22732 25228 22760
rect 24780 22704 24808 22732
rect 25222 22720 25228 22732
rect 25280 22720 25286 22772
rect 26694 22720 26700 22772
rect 26752 22760 26758 22772
rect 30834 22760 30840 22772
rect 26752 22732 30840 22760
rect 26752 22720 26758 22732
rect 30834 22720 30840 22732
rect 30892 22720 30898 22772
rect 33134 22720 33140 22772
rect 33192 22760 33198 22772
rect 36354 22760 36360 22772
rect 33192 22732 36360 22760
rect 33192 22720 33198 22732
rect 36354 22720 36360 22732
rect 36412 22720 36418 22772
rect 2041 22695 2099 22701
rect 2041 22661 2053 22695
rect 2087 22692 2099 22695
rect 13078 22692 13084 22704
rect 2087 22664 13084 22692
rect 2087 22661 2099 22664
rect 2041 22655 2099 22661
rect 13078 22652 13084 22664
rect 13136 22652 13142 22704
rect 13262 22692 13268 22704
rect 13223 22664 13268 22692
rect 13262 22652 13268 22664
rect 13320 22652 13326 22704
rect 13481 22695 13539 22701
rect 13481 22661 13493 22695
rect 13527 22692 13539 22695
rect 14090 22692 14096 22704
rect 13527 22664 14096 22692
rect 13527 22661 13539 22664
rect 13481 22655 13539 22661
rect 1854 22624 1860 22636
rect 1815 22596 1860 22624
rect 1854 22584 1860 22596
rect 1912 22584 1918 22636
rect 2498 22624 2504 22636
rect 2459 22596 2504 22624
rect 2498 22584 2504 22596
rect 2556 22584 2562 22636
rect 9490 22584 9496 22636
rect 9548 22624 9554 22636
rect 9861 22627 9919 22633
rect 9861 22624 9873 22627
rect 9548 22596 9873 22624
rect 9548 22584 9554 22596
rect 9861 22593 9873 22596
rect 9907 22624 9919 22627
rect 10689 22627 10747 22633
rect 10689 22624 10701 22627
rect 9907 22596 10701 22624
rect 9907 22593 9919 22596
rect 9861 22587 9919 22593
rect 10689 22593 10701 22596
rect 10735 22624 10747 22627
rect 10778 22624 10784 22636
rect 10735 22596 10784 22624
rect 10735 22593 10747 22596
rect 10689 22587 10747 22593
rect 10778 22584 10784 22596
rect 10836 22584 10842 22636
rect 14016 22624 14044 22664
rect 14090 22652 14096 22664
rect 14148 22652 14154 22704
rect 14366 22692 14372 22704
rect 14327 22664 14372 22692
rect 14366 22652 14372 22664
rect 14424 22652 14430 22704
rect 14578 22695 14636 22701
rect 14578 22661 14590 22695
rect 14624 22692 14636 22695
rect 15930 22692 15936 22704
rect 14624 22664 15936 22692
rect 14624 22661 14636 22664
rect 14578 22655 14636 22661
rect 15930 22652 15936 22664
rect 15988 22652 15994 22704
rect 20625 22695 20683 22701
rect 18110 22664 19334 22692
rect 14458 22624 14464 22636
rect 14016 22596 14464 22624
rect 14458 22584 14464 22596
rect 14516 22584 14522 22636
rect 18110 22633 18138 22664
rect 17589 22627 17647 22633
rect 17589 22593 17601 22627
rect 17635 22624 17647 22627
rect 18095 22627 18153 22633
rect 18095 22624 18107 22627
rect 17635 22596 18107 22624
rect 17635 22593 17647 22596
rect 17589 22587 17647 22593
rect 18095 22593 18107 22596
rect 18141 22593 18153 22627
rect 18230 22624 18236 22636
rect 18191 22596 18236 22624
rect 18095 22587 18153 22593
rect 18230 22584 18236 22596
rect 18288 22584 18294 22636
rect 18322 22584 18328 22636
rect 18380 22624 18386 22636
rect 18509 22627 18567 22633
rect 18380 22596 18425 22624
rect 18380 22584 18386 22596
rect 18509 22593 18521 22627
rect 18555 22593 18567 22627
rect 19306 22624 19334 22664
rect 20625 22661 20637 22695
rect 20671 22692 20683 22695
rect 20714 22692 20720 22704
rect 20671 22664 20720 22692
rect 20671 22661 20683 22664
rect 20625 22655 20683 22661
rect 20714 22652 20720 22664
rect 20772 22652 20778 22704
rect 20896 22664 24164 22692
rect 19886 22624 19892 22636
rect 19306 22596 19892 22624
rect 18509 22587 18567 22593
rect 9950 22556 9956 22568
rect 10008 22567 10014 22568
rect 9863 22528 9956 22556
rect 9950 22516 9956 22528
rect 10008 22556 10088 22567
rect 10229 22559 10287 22565
rect 10008 22539 10180 22556
rect 10008 22516 10014 22539
rect 10060 22528 10180 22539
rect 10152 22488 10180 22528
rect 10229 22525 10241 22559
rect 10275 22556 10287 22559
rect 10410 22556 10416 22568
rect 10275 22528 10416 22556
rect 10275 22525 10287 22528
rect 10229 22519 10287 22525
rect 10410 22516 10416 22528
rect 10468 22516 10474 22568
rect 10962 22556 10968 22568
rect 10875 22528 10968 22556
rect 10962 22516 10968 22528
rect 11020 22556 11026 22568
rect 13722 22556 13728 22568
rect 11020 22528 13728 22556
rect 11020 22516 11026 22528
rect 13722 22516 13728 22528
rect 13780 22516 13786 22568
rect 14016 22565 14143 22567
rect 14016 22559 14158 22565
rect 14016 22556 14112 22559
rect 13924 22539 14112 22556
rect 13924 22528 14044 22539
rect 10781 22491 10839 22497
rect 10781 22488 10793 22491
rect 10152 22460 10793 22488
rect 10781 22457 10793 22460
rect 10827 22457 10839 22491
rect 10781 22451 10839 22457
rect 13633 22491 13691 22497
rect 13633 22457 13645 22491
rect 13679 22488 13691 22491
rect 13924 22488 13952 22528
rect 14100 22525 14112 22539
rect 14146 22525 14158 22559
rect 18524 22556 18552 22587
rect 19886 22584 19892 22596
rect 19944 22584 19950 22636
rect 20896 22633 20924 22664
rect 20896 22627 20959 22633
rect 20896 22599 20913 22627
rect 20901 22593 20913 22599
rect 20947 22593 20959 22627
rect 20901 22587 20959 22593
rect 20993 22627 21051 22633
rect 20993 22593 21005 22627
rect 21039 22593 21051 22627
rect 20993 22587 21051 22593
rect 14100 22519 14158 22525
rect 18340 22528 18552 22556
rect 13679 22460 13952 22488
rect 13679 22457 13691 22460
rect 13633 22451 13691 22457
rect 9766 22380 9772 22432
rect 9824 22420 9830 22432
rect 10410 22420 10416 22432
rect 9824 22392 10416 22420
rect 9824 22380 9830 22392
rect 10410 22380 10416 22392
rect 10468 22380 10474 22432
rect 10796 22420 10824 22451
rect 14274 22448 14280 22500
rect 14332 22488 14338 22500
rect 14826 22488 14832 22500
rect 14332 22460 14832 22488
rect 14332 22448 14338 22460
rect 14826 22448 14832 22460
rect 14884 22448 14890 22500
rect 14918 22448 14924 22500
rect 14976 22488 14982 22500
rect 17954 22488 17960 22500
rect 14976 22460 17960 22488
rect 14976 22448 14982 22460
rect 17954 22448 17960 22460
rect 18012 22448 18018 22500
rect 18138 22448 18144 22500
rect 18196 22488 18202 22500
rect 18340 22488 18368 22528
rect 20070 22516 20076 22568
rect 20128 22556 20134 22568
rect 21008 22556 21036 22587
rect 21082 22584 21088 22636
rect 21140 22633 21146 22636
rect 21140 22624 21148 22633
rect 21140 22596 21185 22624
rect 21140 22587 21148 22596
rect 21140 22584 21146 22587
rect 21266 22584 21272 22636
rect 21324 22624 21330 22636
rect 21324 22596 21369 22624
rect 21324 22584 21330 22596
rect 20128 22528 21036 22556
rect 20128 22516 20134 22528
rect 20916 22500 20944 22528
rect 18196 22460 18368 22488
rect 18196 22448 18202 22460
rect 18414 22448 18420 22500
rect 18472 22488 18478 22500
rect 19426 22488 19432 22500
rect 18472 22460 19432 22488
rect 18472 22448 18478 22460
rect 19426 22448 19432 22460
rect 19484 22448 19490 22500
rect 20898 22448 20904 22500
rect 20956 22448 20962 22500
rect 13449 22423 13507 22429
rect 13449 22420 13461 22423
rect 10796 22392 13461 22420
rect 13449 22389 13461 22392
rect 13495 22420 13507 22423
rect 13814 22420 13820 22432
rect 13495 22392 13820 22420
rect 13495 22389 13507 22392
rect 13449 22383 13507 22389
rect 13814 22380 13820 22392
rect 13872 22380 13878 22432
rect 13906 22380 13912 22432
rect 13964 22420 13970 22432
rect 14737 22423 14795 22429
rect 14737 22420 14749 22423
rect 13964 22392 14749 22420
rect 13964 22380 13970 22392
rect 14737 22389 14749 22392
rect 14783 22389 14795 22423
rect 14737 22383 14795 22389
rect 16022 22380 16028 22432
rect 16080 22420 16086 22432
rect 20806 22420 20812 22432
rect 16080 22392 20812 22420
rect 16080 22380 16086 22392
rect 20806 22380 20812 22392
rect 20864 22380 20870 22432
rect 24136 22420 24164 22664
rect 24762 22652 24768 22704
rect 24820 22652 24826 22704
rect 25133 22695 25191 22701
rect 25133 22661 25145 22695
rect 25179 22692 25191 22695
rect 25777 22695 25835 22701
rect 25777 22692 25789 22695
rect 25179 22664 25789 22692
rect 25179 22661 25191 22664
rect 25133 22655 25191 22661
rect 25777 22661 25789 22664
rect 25823 22661 25835 22695
rect 25777 22655 25835 22661
rect 26142 22652 26148 22704
rect 26200 22692 26206 22704
rect 30742 22692 30748 22704
rect 26200 22664 30748 22692
rect 26200 22652 26206 22664
rect 30742 22652 30748 22664
rect 30800 22652 30806 22704
rect 31021 22695 31079 22701
rect 31021 22661 31033 22695
rect 31067 22692 31079 22695
rect 31110 22692 31116 22704
rect 31067 22664 31116 22692
rect 31067 22661 31079 22664
rect 31021 22655 31079 22661
rect 31110 22652 31116 22664
rect 31168 22652 31174 22704
rect 31220 22664 32812 22692
rect 24213 22627 24271 22633
rect 24213 22593 24225 22627
rect 24259 22593 24271 22627
rect 24394 22624 24400 22636
rect 24355 22596 24400 22624
rect 24213 22587 24271 22593
rect 24228 22556 24256 22587
rect 24394 22584 24400 22596
rect 24452 22584 24458 22636
rect 24489 22627 24547 22633
rect 24489 22593 24501 22627
rect 24535 22624 24547 22627
rect 24780 22624 24808 22652
rect 24535 22596 24808 22624
rect 24949 22627 25007 22633
rect 24535 22593 24547 22596
rect 24489 22587 24547 22593
rect 24949 22593 24961 22627
rect 24995 22593 25007 22627
rect 25222 22624 25228 22636
rect 25183 22596 25228 22624
rect 24949 22587 25007 22593
rect 24762 22556 24768 22568
rect 24228 22528 24768 22556
rect 24762 22516 24768 22528
rect 24820 22516 24826 22568
rect 24964 22556 24992 22587
rect 25222 22584 25228 22596
rect 25280 22584 25286 22636
rect 25498 22584 25504 22636
rect 25556 22624 25562 22636
rect 25685 22627 25743 22633
rect 25685 22624 25697 22627
rect 25556 22596 25697 22624
rect 25556 22584 25562 22596
rect 25685 22593 25697 22596
rect 25731 22593 25743 22627
rect 25866 22624 25872 22636
rect 25827 22596 25872 22624
rect 25685 22587 25743 22593
rect 25866 22584 25872 22596
rect 25924 22584 25930 22636
rect 29454 22624 29460 22636
rect 29415 22596 29460 22624
rect 29454 22584 29460 22596
rect 29512 22584 29518 22636
rect 29638 22584 29644 22636
rect 29696 22624 29702 22636
rect 29733 22627 29791 22633
rect 29733 22624 29745 22627
rect 29696 22596 29745 22624
rect 29696 22584 29702 22596
rect 29733 22593 29745 22596
rect 29779 22593 29791 22627
rect 29733 22587 29791 22593
rect 30834 22584 30840 22636
rect 30892 22624 30898 22636
rect 31220 22624 31248 22664
rect 30892 22596 31248 22624
rect 31337 22627 31395 22633
rect 30892 22584 30898 22596
rect 31337 22593 31349 22627
rect 31383 22624 31395 22627
rect 31478 22624 31484 22636
rect 31383 22596 31484 22624
rect 31383 22593 31395 22596
rect 31337 22587 31395 22593
rect 31478 22584 31484 22596
rect 31536 22584 31542 22636
rect 32122 22584 32128 22636
rect 32180 22624 32186 22636
rect 32784 22633 32812 22664
rect 33594 22652 33600 22704
rect 33652 22692 33658 22704
rect 47118 22692 47124 22704
rect 33652 22664 47124 22692
rect 33652 22652 33658 22664
rect 47118 22652 47124 22664
rect 47176 22652 47182 22704
rect 47394 22652 47400 22704
rect 47452 22692 47458 22704
rect 47452 22664 47808 22692
rect 47452 22652 47458 22664
rect 32217 22627 32275 22633
rect 32217 22624 32229 22627
rect 32180 22596 32229 22624
rect 32180 22584 32186 22596
rect 32217 22593 32229 22596
rect 32263 22593 32275 22627
rect 32217 22587 32275 22593
rect 32769 22627 32827 22633
rect 32769 22593 32781 22627
rect 32815 22624 32827 22627
rect 33134 22624 33140 22636
rect 32815 22596 33140 22624
rect 32815 22593 32827 22596
rect 32769 22587 32827 22593
rect 33134 22584 33140 22596
rect 33192 22584 33198 22636
rect 35710 22624 35716 22636
rect 35671 22596 35716 22624
rect 35710 22584 35716 22596
rect 35768 22584 35774 22636
rect 35894 22624 35900 22636
rect 35855 22596 35900 22624
rect 35894 22584 35900 22596
rect 35952 22624 35958 22636
rect 36078 22624 36084 22636
rect 35952 22596 36084 22624
rect 35952 22584 35958 22596
rect 36078 22584 36084 22596
rect 36136 22584 36142 22636
rect 47578 22624 47584 22636
rect 47539 22596 47584 22624
rect 47578 22584 47584 22596
rect 47636 22584 47642 22636
rect 47780 22633 47808 22664
rect 47765 22627 47823 22633
rect 47765 22593 47777 22627
rect 47811 22593 47823 22627
rect 47765 22587 47823 22593
rect 25130 22556 25136 22568
rect 24964 22528 25136 22556
rect 25130 22516 25136 22528
rect 25188 22516 25194 22568
rect 29546 22556 29552 22568
rect 29507 22528 29552 22556
rect 29546 22516 29552 22528
rect 29604 22516 29610 22568
rect 31205 22559 31263 22565
rect 31205 22525 31217 22559
rect 31251 22556 31263 22559
rect 31570 22556 31576 22568
rect 31251 22528 31576 22556
rect 31251 22525 31263 22528
rect 31205 22519 31263 22525
rect 31570 22516 31576 22528
rect 31628 22516 31634 22568
rect 33413 22559 33471 22565
rect 33413 22525 33425 22559
rect 33459 22525 33471 22559
rect 33594 22556 33600 22568
rect 33555 22528 33600 22556
rect 33413 22519 33471 22525
rect 24946 22488 24952 22500
rect 24907 22460 24952 22488
rect 24946 22448 24952 22460
rect 25004 22448 25010 22500
rect 25222 22448 25228 22500
rect 25280 22488 25286 22500
rect 25280 22460 31202 22488
rect 25280 22448 25286 22460
rect 26142 22420 26148 22432
rect 24136 22392 26148 22420
rect 26142 22380 26148 22392
rect 26200 22380 26206 22432
rect 29362 22380 29368 22432
rect 29420 22420 29426 22432
rect 29457 22423 29515 22429
rect 29457 22420 29469 22423
rect 29420 22392 29469 22420
rect 29420 22380 29426 22392
rect 29457 22389 29469 22392
rect 29503 22389 29515 22423
rect 29457 22383 29515 22389
rect 29917 22423 29975 22429
rect 29917 22389 29929 22423
rect 29963 22420 29975 22423
rect 31021 22423 31079 22429
rect 31021 22420 31033 22423
rect 29963 22392 31033 22420
rect 29963 22389 29975 22392
rect 29917 22383 29975 22389
rect 31021 22389 31033 22392
rect 31067 22389 31079 22423
rect 31174 22420 31202 22460
rect 31386 22448 31392 22500
rect 31444 22488 31450 22500
rect 31481 22491 31539 22497
rect 31481 22488 31493 22491
rect 31444 22460 31493 22488
rect 31444 22448 31450 22460
rect 31481 22457 31493 22460
rect 31527 22457 31539 22491
rect 31481 22451 31539 22457
rect 33428 22420 33456 22519
rect 33594 22516 33600 22528
rect 33652 22516 33658 22568
rect 35253 22559 35311 22565
rect 35253 22525 35265 22559
rect 35299 22556 35311 22559
rect 42058 22556 42064 22568
rect 35299 22528 42064 22556
rect 35299 22525 35311 22528
rect 35253 22519 35311 22525
rect 42058 22516 42064 22528
rect 42116 22516 42122 22568
rect 35618 22448 35624 22500
rect 35676 22488 35682 22500
rect 36262 22488 36268 22500
rect 35676 22460 36268 22488
rect 35676 22448 35682 22460
rect 36262 22448 36268 22460
rect 36320 22448 36326 22500
rect 31174 22392 33456 22420
rect 31021 22383 31079 22389
rect 34606 22380 34612 22432
rect 34664 22420 34670 22432
rect 36081 22423 36139 22429
rect 36081 22420 36093 22423
rect 34664 22392 36093 22420
rect 34664 22380 34670 22392
rect 36081 22389 36093 22392
rect 36127 22389 36139 22423
rect 47670 22420 47676 22432
rect 47631 22392 47676 22420
rect 36081 22383 36139 22389
rect 47670 22380 47676 22392
rect 47728 22380 47734 22432
rect 1104 22330 48852 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 48852 22330
rect 1104 22256 48852 22278
rect 4798 22176 4804 22228
rect 4856 22216 4862 22228
rect 18141 22219 18199 22225
rect 4856 22188 17264 22216
rect 4856 22176 4862 22188
rect 9490 22108 9496 22160
rect 9548 22148 9554 22160
rect 10045 22151 10103 22157
rect 10045 22148 10057 22151
rect 9548 22120 10057 22148
rect 9548 22108 9554 22120
rect 10045 22117 10057 22120
rect 10091 22117 10103 22151
rect 10045 22111 10103 22117
rect 14277 22151 14335 22157
rect 14277 22117 14289 22151
rect 14323 22148 14335 22151
rect 15286 22148 15292 22160
rect 14323 22120 15292 22148
rect 14323 22117 14335 22120
rect 14277 22111 14335 22117
rect 15286 22108 15292 22120
rect 15344 22108 15350 22160
rect 17236 22148 17264 22188
rect 18141 22185 18153 22219
rect 18187 22216 18199 22219
rect 18322 22216 18328 22228
rect 18187 22188 18328 22216
rect 18187 22185 18199 22188
rect 18141 22179 18199 22185
rect 18322 22176 18328 22188
rect 18380 22176 18386 22228
rect 20901 22219 20959 22225
rect 18432 22188 20208 22216
rect 18432 22148 18460 22188
rect 17236 22120 18460 22148
rect 18506 22108 18512 22160
rect 18564 22148 18570 22160
rect 20070 22148 20076 22160
rect 18564 22120 20076 22148
rect 18564 22108 18570 22120
rect 20070 22108 20076 22120
rect 20128 22108 20134 22160
rect 20180 22148 20208 22188
rect 20901 22185 20913 22219
rect 20947 22216 20959 22219
rect 21082 22216 21088 22228
rect 20947 22188 21088 22216
rect 20947 22185 20959 22188
rect 20901 22179 20959 22185
rect 21082 22176 21088 22188
rect 21140 22176 21146 22228
rect 28813 22219 28871 22225
rect 28813 22185 28825 22219
rect 28859 22216 28871 22219
rect 29454 22216 29460 22228
rect 28859 22188 29460 22216
rect 28859 22185 28871 22188
rect 28813 22179 28871 22185
rect 29454 22176 29460 22188
rect 29512 22176 29518 22228
rect 29730 22216 29736 22228
rect 29691 22188 29736 22216
rect 29730 22176 29736 22188
rect 29788 22176 29794 22228
rect 29840 22188 30049 22216
rect 26694 22148 26700 22160
rect 20180 22120 26700 22148
rect 26694 22108 26700 22120
rect 26752 22108 26758 22160
rect 26878 22108 26884 22160
rect 26936 22148 26942 22160
rect 29840 22148 29868 22188
rect 26936 22120 29868 22148
rect 30021 22148 30049 22188
rect 30190 22176 30196 22228
rect 30248 22216 30254 22228
rect 30834 22216 30840 22228
rect 30248 22188 30293 22216
rect 30795 22188 30840 22216
rect 30248 22176 30254 22188
rect 30834 22176 30840 22188
rect 30892 22176 30898 22228
rect 31297 22219 31355 22225
rect 31297 22185 31309 22219
rect 31343 22216 31355 22219
rect 31478 22216 31484 22228
rect 31343 22188 31484 22216
rect 31343 22185 31355 22188
rect 31297 22179 31355 22185
rect 31478 22176 31484 22188
rect 31536 22176 31542 22228
rect 46934 22216 46940 22228
rect 33336 22188 46940 22216
rect 33336 22148 33364 22188
rect 46934 22176 46940 22188
rect 46992 22176 46998 22228
rect 47854 22216 47860 22228
rect 47815 22188 47860 22216
rect 47854 22176 47860 22188
rect 47912 22176 47918 22228
rect 30021 22120 33364 22148
rect 33428 22120 33916 22148
rect 26936 22108 26942 22120
rect 7834 22040 7840 22092
rect 7892 22080 7898 22092
rect 14461 22083 14519 22089
rect 7892 22052 14412 22080
rect 7892 22040 7898 22052
rect 6825 22015 6883 22021
rect 6825 21981 6837 22015
rect 6871 22012 6883 22015
rect 8018 22012 8024 22024
rect 6871 21984 8024 22012
rect 6871 21981 6883 21984
rect 6825 21975 6883 21981
rect 8018 21972 8024 21984
rect 8076 21972 8082 22024
rect 9950 22012 9956 22024
rect 9911 21984 9956 22012
rect 9950 21972 9956 21984
rect 10008 21972 10014 22024
rect 14090 21972 14096 22024
rect 14148 22012 14154 22024
rect 14185 22015 14243 22021
rect 14185 22012 14197 22015
rect 14148 21984 14197 22012
rect 14148 21972 14154 21984
rect 14185 21981 14197 21984
rect 14231 21981 14243 22015
rect 14384 22012 14412 22052
rect 14461 22049 14473 22083
rect 14507 22080 14519 22083
rect 14550 22080 14556 22092
rect 14507 22052 14556 22080
rect 14507 22049 14519 22052
rect 14461 22043 14519 22049
rect 14550 22040 14556 22052
rect 14608 22040 14614 22092
rect 17218 22040 17224 22092
rect 17276 22080 17282 22092
rect 25593 22083 25651 22089
rect 17276 22052 25452 22080
rect 17276 22040 17282 22052
rect 14384 21984 14596 22012
rect 14185 21975 14243 21981
rect 7092 21947 7150 21953
rect 7092 21913 7104 21947
rect 7138 21944 7150 21947
rect 7138 21916 10088 21944
rect 7138 21913 7150 21916
rect 7092 21907 7150 21913
rect 2314 21836 2320 21888
rect 2372 21876 2378 21888
rect 7190 21876 7196 21888
rect 2372 21848 7196 21876
rect 2372 21836 2378 21848
rect 7190 21836 7196 21848
rect 7248 21836 7254 21888
rect 7282 21836 7288 21888
rect 7340 21876 7346 21888
rect 8205 21879 8263 21885
rect 8205 21876 8217 21879
rect 7340 21848 8217 21876
rect 7340 21836 7346 21848
rect 8205 21845 8217 21848
rect 8251 21845 8263 21879
rect 9950 21876 9956 21888
rect 9911 21848 9956 21876
rect 8205 21839 8263 21845
rect 9950 21836 9956 21848
rect 10008 21836 10014 21888
rect 10060 21876 10088 21916
rect 10134 21904 10140 21956
rect 10192 21944 10198 21956
rect 10229 21947 10287 21953
rect 10229 21944 10241 21947
rect 10192 21916 10241 21944
rect 10192 21904 10198 21916
rect 10229 21913 10241 21916
rect 10275 21944 10287 21947
rect 10962 21944 10968 21956
rect 10275 21916 10968 21944
rect 10275 21913 10287 21916
rect 10229 21907 10287 21913
rect 10962 21904 10968 21916
rect 11020 21904 11026 21956
rect 14458 21944 14464 21956
rect 14419 21916 14464 21944
rect 14458 21904 14464 21916
rect 14516 21904 14522 21956
rect 14568 21944 14596 21984
rect 16666 21972 16672 22024
rect 16724 22012 16730 22024
rect 17773 22015 17831 22021
rect 17773 22012 17785 22015
rect 16724 21984 17785 22012
rect 16724 21972 16730 21984
rect 17773 21981 17785 21984
rect 17819 21981 17831 22015
rect 17954 22012 17960 22024
rect 17915 21984 17960 22012
rect 17773 21975 17831 21981
rect 17586 21944 17592 21956
rect 14568 21916 17592 21944
rect 17586 21904 17592 21916
rect 17644 21904 17650 21956
rect 17788 21944 17816 21975
rect 17954 21972 17960 21984
rect 18012 21972 18018 22024
rect 19426 21972 19432 22024
rect 19484 22012 19490 22024
rect 19889 22015 19947 22021
rect 19889 22012 19901 22015
rect 19484 21984 19901 22012
rect 19484 21972 19490 21984
rect 19889 21981 19901 21984
rect 19935 22012 19947 22015
rect 20622 22012 20628 22024
rect 19935 21984 20628 22012
rect 19935 21981 19947 21984
rect 19889 21975 19947 21981
rect 20622 21972 20628 21984
rect 20680 21972 20686 22024
rect 20990 21972 20996 22024
rect 21048 22012 21054 22024
rect 24854 22012 24860 22024
rect 21048 21984 24860 22012
rect 21048 21972 21054 21984
rect 24854 21972 24860 21984
rect 24912 21972 24918 22024
rect 25130 22012 25136 22024
rect 25091 21984 25136 22012
rect 25130 21972 25136 21984
rect 25188 21972 25194 22024
rect 19334 21944 19340 21956
rect 17788 21916 19340 21944
rect 19334 21904 19340 21916
rect 19392 21904 19398 21956
rect 20346 21904 20352 21956
rect 20404 21944 20410 21956
rect 20533 21947 20591 21953
rect 20533 21944 20545 21947
rect 20404 21916 20545 21944
rect 20404 21904 20410 21916
rect 20533 21913 20545 21916
rect 20579 21913 20591 21947
rect 20533 21907 20591 21913
rect 20717 21947 20775 21953
rect 20717 21913 20729 21947
rect 20763 21944 20775 21947
rect 22186 21944 22192 21956
rect 20763 21916 22192 21944
rect 20763 21913 20775 21916
rect 20717 21907 20775 21913
rect 22186 21904 22192 21916
rect 22244 21904 22250 21956
rect 22278 21904 22284 21956
rect 22336 21944 22342 21956
rect 25314 21944 25320 21956
rect 22336 21916 25320 21944
rect 22336 21904 22342 21916
rect 25314 21904 25320 21916
rect 25372 21904 25378 21956
rect 25225 21879 25283 21885
rect 25225 21876 25237 21879
rect 10060 21848 25237 21876
rect 25225 21845 25237 21848
rect 25271 21845 25283 21879
rect 25424 21876 25452 22052
rect 25593 22049 25605 22083
rect 25639 22080 25651 22083
rect 26326 22080 26332 22092
rect 25639 22052 26332 22080
rect 25639 22049 25651 22052
rect 25593 22043 25651 22049
rect 26326 22040 26332 22052
rect 26384 22040 26390 22092
rect 28534 22040 28540 22092
rect 28592 22080 28598 22092
rect 28629 22083 28687 22089
rect 28629 22080 28641 22083
rect 28592 22052 28641 22080
rect 28592 22040 28598 22052
rect 28629 22049 28641 22052
rect 28675 22049 28687 22083
rect 28629 22043 28687 22049
rect 28718 22040 28724 22092
rect 28776 22080 28782 22092
rect 29638 22080 29644 22092
rect 28776 22052 29644 22080
rect 28776 22040 28782 22052
rect 29638 22040 29644 22052
rect 29696 22040 29702 22092
rect 29825 22083 29883 22089
rect 29825 22049 29837 22083
rect 29871 22049 29883 22083
rect 30926 22080 30932 22092
rect 30887 22052 30932 22080
rect 29825 22046 29883 22049
rect 29825 22043 29960 22046
rect 25498 21972 25504 22024
rect 25556 22012 25562 22024
rect 26234 22012 26240 22024
rect 25556 21984 25601 22012
rect 26195 21984 26240 22012
rect 25556 21972 25562 21984
rect 26234 21972 26240 21984
rect 26292 21972 26298 22024
rect 26418 22012 26424 22024
rect 26379 21984 26424 22012
rect 26418 21972 26424 21984
rect 26476 21972 26482 22024
rect 26881 22015 26939 22021
rect 26881 21981 26893 22015
rect 26927 22012 26939 22015
rect 27798 22012 27804 22024
rect 26927 21984 27804 22012
rect 26927 21981 26939 21984
rect 26881 21975 26939 21981
rect 26234 21876 26240 21888
rect 25424 21848 26240 21876
rect 25225 21839 25283 21845
rect 26234 21836 26240 21848
rect 26292 21836 26298 21888
rect 26418 21876 26424 21888
rect 26379 21848 26424 21876
rect 26418 21836 26424 21848
rect 26476 21836 26482 21888
rect 26510 21836 26516 21888
rect 26568 21876 26574 21888
rect 26896 21876 26924 21975
rect 27798 21972 27804 21984
rect 27856 22012 27862 22024
rect 28810 22012 28816 22024
rect 27856 21984 28120 22012
rect 28771 21984 28816 22012
rect 27856 21972 27862 21984
rect 26568 21848 26924 21876
rect 26973 21879 27031 21885
rect 26568 21836 26574 21848
rect 26973 21845 26985 21879
rect 27019 21876 27031 21879
rect 27246 21876 27252 21888
rect 27019 21848 27252 21876
rect 27019 21845 27031 21848
rect 26973 21839 27031 21845
rect 27246 21836 27252 21848
rect 27304 21836 27310 21888
rect 28092 21876 28120 21984
rect 28810 21972 28816 21984
rect 28868 21972 28874 22024
rect 29730 22012 29736 22024
rect 28920 21984 29736 22012
rect 28258 21904 28264 21956
rect 28316 21944 28322 21956
rect 28537 21947 28595 21953
rect 28537 21944 28549 21947
rect 28316 21916 28549 21944
rect 28316 21904 28322 21916
rect 28537 21913 28549 21916
rect 28583 21913 28595 21947
rect 28537 21907 28595 21913
rect 28920 21876 28948 21984
rect 29730 21972 29736 21984
rect 29788 21972 29794 22024
rect 29840 22018 29960 22043
rect 30926 22040 30932 22052
rect 30984 22040 30990 22092
rect 32858 22040 32864 22092
rect 32916 22080 32922 22092
rect 33428 22080 33456 22120
rect 32916 22052 33456 22080
rect 32916 22040 32922 22052
rect 29178 21944 29184 21956
rect 29012 21916 29184 21944
rect 29012 21885 29040 21916
rect 29178 21904 29184 21916
rect 29236 21904 29242 21956
rect 29454 21904 29460 21956
rect 29512 21944 29518 21956
rect 29549 21947 29607 21953
rect 29549 21944 29561 21947
rect 29512 21916 29561 21944
rect 29512 21904 29518 21916
rect 29549 21913 29561 21916
rect 29595 21913 29607 21947
rect 29932 21944 29960 22018
rect 30006 21972 30012 22024
rect 30064 22012 30070 22024
rect 31113 22015 31171 22021
rect 30064 21984 30109 22012
rect 30064 21972 30070 21984
rect 31113 21981 31125 22015
rect 31159 22012 31171 22015
rect 31386 22012 31392 22024
rect 31159 21984 31392 22012
rect 31159 21981 31171 21984
rect 31113 21975 31171 21981
rect 31386 21972 31392 21984
rect 31444 21972 31450 22024
rect 31941 22015 31999 22021
rect 31941 21981 31953 22015
rect 31987 22012 31999 22015
rect 32122 22012 32128 22024
rect 31987 21984 32128 22012
rect 31987 21981 31999 21984
rect 31941 21975 31999 21981
rect 32122 21972 32128 21984
rect 32180 21972 32186 22024
rect 33410 21972 33416 22024
rect 33468 22012 33474 22024
rect 33888 22021 33916 22120
rect 36262 22108 36268 22160
rect 36320 22148 36326 22160
rect 36357 22151 36415 22157
rect 36357 22148 36369 22151
rect 36320 22120 36369 22148
rect 36320 22108 36326 22120
rect 36357 22117 36369 22120
rect 36403 22117 36415 22151
rect 47872 22148 47900 22176
rect 36357 22111 36415 22117
rect 47136 22120 47900 22148
rect 47136 22080 47164 22120
rect 47394 22080 47400 22092
rect 36004 22052 47164 22080
rect 47355 22052 47400 22080
rect 33781 22015 33839 22021
rect 33781 22012 33793 22015
rect 33468 21984 33793 22012
rect 33468 21972 33474 21984
rect 33781 21981 33793 21984
rect 33827 21981 33839 22015
rect 33781 21975 33839 21981
rect 33873 22015 33931 22021
rect 33873 21981 33885 22015
rect 33919 21981 33931 22015
rect 33873 21975 33931 21981
rect 33962 21972 33968 22024
rect 34020 22012 34026 22024
rect 34149 22015 34207 22021
rect 34020 21984 34065 22012
rect 34020 21972 34026 21984
rect 34149 21981 34161 22015
rect 34195 22012 34207 22015
rect 34606 22012 34612 22024
rect 34195 21984 34612 22012
rect 34195 21981 34207 21984
rect 34149 21975 34207 21981
rect 34606 21972 34612 21984
rect 34664 21972 34670 22024
rect 34698 21972 34704 22024
rect 34756 22012 34762 22024
rect 34977 22015 35035 22021
rect 34977 22012 34989 22015
rect 34756 21984 34989 22012
rect 34756 21972 34762 21984
rect 34977 21981 34989 21984
rect 35023 21981 35035 22015
rect 34977 21975 35035 21981
rect 30837 21947 30895 21953
rect 29932 21916 30604 21944
rect 29549 21907 29607 21913
rect 28092 21848 28948 21876
rect 28997 21879 29055 21885
rect 28997 21845 29009 21879
rect 29043 21845 29055 21879
rect 28997 21839 29055 21845
rect 29086 21836 29092 21888
rect 29144 21876 29150 21888
rect 29914 21876 29920 21888
rect 29144 21848 29920 21876
rect 29144 21836 29150 21848
rect 29914 21836 29920 21848
rect 29972 21836 29978 21888
rect 30576 21885 30604 21916
rect 30837 21913 30849 21947
rect 30883 21944 30895 21947
rect 31202 21944 31208 21956
rect 30883 21916 31208 21944
rect 30883 21913 30895 21916
rect 30837 21907 30895 21913
rect 31202 21904 31208 21916
rect 31260 21904 31266 21956
rect 31294 21904 31300 21956
rect 31352 21944 31358 21956
rect 32585 21947 32643 21953
rect 32585 21944 32597 21947
rect 31352 21916 32597 21944
rect 31352 21904 31358 21916
rect 32585 21913 32597 21916
rect 32631 21944 32643 21947
rect 32674 21944 32680 21956
rect 32631 21916 32680 21944
rect 32631 21913 32643 21916
rect 32585 21907 32643 21913
rect 32674 21904 32680 21916
rect 32732 21904 32738 21956
rect 33505 21947 33563 21953
rect 33505 21913 33517 21947
rect 33551 21944 33563 21947
rect 34514 21944 34520 21956
rect 33551 21916 34520 21944
rect 33551 21913 33563 21916
rect 33505 21907 33563 21913
rect 34514 21904 34520 21916
rect 34572 21904 34578 21956
rect 34790 21904 34796 21956
rect 34848 21944 34854 21956
rect 35222 21947 35280 21953
rect 35222 21944 35234 21947
rect 34848 21916 35234 21944
rect 34848 21904 34854 21916
rect 35222 21913 35234 21916
rect 35268 21913 35280 21947
rect 35222 21907 35280 21913
rect 30561 21879 30619 21885
rect 30561 21845 30573 21879
rect 30607 21876 30619 21879
rect 36004 21876 36032 22052
rect 47394 22040 47400 22052
rect 47452 22040 47458 22092
rect 36262 21972 36268 22024
rect 36320 22012 36326 22024
rect 36909 22015 36967 22021
rect 36909 22012 36921 22015
rect 36320 21984 36921 22012
rect 36320 21972 36326 21984
rect 36909 21981 36921 21984
rect 36955 21981 36967 22015
rect 36909 21975 36967 21981
rect 47489 22015 47547 22021
rect 47489 21981 47501 22015
rect 47535 22012 47547 22015
rect 47578 22012 47584 22024
rect 47535 21984 47584 22012
rect 47535 21981 47547 21984
rect 47489 21975 47547 21981
rect 47578 21972 47584 21984
rect 47636 21972 47642 22024
rect 47854 22012 47860 22024
rect 47815 21984 47860 22012
rect 47854 21972 47860 21984
rect 47912 21972 47918 22024
rect 37093 21947 37151 21953
rect 37093 21913 37105 21947
rect 37139 21944 37151 21947
rect 37366 21944 37372 21956
rect 37139 21916 37372 21944
rect 37139 21913 37151 21916
rect 37093 21907 37151 21913
rect 37366 21904 37372 21916
rect 37424 21904 37430 21956
rect 38749 21947 38807 21953
rect 38749 21913 38761 21947
rect 38795 21944 38807 21947
rect 40770 21944 40776 21956
rect 38795 21916 40776 21944
rect 38795 21913 38807 21916
rect 38749 21907 38807 21913
rect 40770 21904 40776 21916
rect 40828 21904 40834 21956
rect 30607 21848 36032 21876
rect 30607 21845 30619 21848
rect 30561 21839 30619 21845
rect 36170 21836 36176 21888
rect 36228 21876 36234 21888
rect 48041 21879 48099 21885
rect 48041 21876 48053 21879
rect 36228 21848 48053 21876
rect 36228 21836 36234 21848
rect 48041 21845 48053 21848
rect 48087 21845 48099 21879
rect 48041 21839 48099 21845
rect 1104 21786 48852 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 48852 21786
rect 1104 21712 48852 21734
rect 2682 21632 2688 21684
rect 2740 21672 2746 21684
rect 14550 21672 14556 21684
rect 2740 21644 14556 21672
rect 2740 21632 2746 21644
rect 14550 21632 14556 21644
rect 14608 21632 14614 21684
rect 14645 21675 14703 21681
rect 14645 21641 14657 21675
rect 14691 21672 14703 21675
rect 14826 21672 14832 21684
rect 14691 21644 14832 21672
rect 14691 21641 14703 21644
rect 14645 21635 14703 21641
rect 14826 21632 14832 21644
rect 14884 21632 14890 21684
rect 15654 21632 15660 21684
rect 15712 21672 15718 21684
rect 15749 21675 15807 21681
rect 15749 21672 15761 21675
rect 15712 21644 15761 21672
rect 15712 21632 15718 21644
rect 15749 21641 15761 21644
rect 15795 21641 15807 21675
rect 15749 21635 15807 21641
rect 19334 21632 19340 21684
rect 19392 21672 19398 21684
rect 19521 21675 19579 21681
rect 19521 21672 19533 21675
rect 19392 21644 19533 21672
rect 19392 21632 19398 21644
rect 19521 21641 19533 21644
rect 19567 21672 19579 21675
rect 20346 21672 20352 21684
rect 19567 21644 20352 21672
rect 19567 21641 19579 21644
rect 19521 21635 19579 21641
rect 20346 21632 20352 21644
rect 20404 21632 20410 21684
rect 20622 21632 20628 21684
rect 20680 21672 20686 21684
rect 25041 21675 25099 21681
rect 20680 21644 24808 21672
rect 20680 21632 20686 21644
rect 2406 21564 2412 21616
rect 2464 21604 2470 21616
rect 7098 21604 7104 21616
rect 2464 21576 7104 21604
rect 2464 21564 2470 21576
rect 7098 21564 7104 21576
rect 7156 21564 7162 21616
rect 7190 21564 7196 21616
rect 7248 21604 7254 21616
rect 17218 21604 17224 21616
rect 7248 21576 17224 21604
rect 7248 21564 7254 21576
rect 17218 21564 17224 21576
rect 17276 21564 17282 21616
rect 17402 21564 17408 21616
rect 17460 21604 17466 21616
rect 22278 21604 22284 21616
rect 17460 21576 22284 21604
rect 17460 21564 17466 21576
rect 22278 21564 22284 21576
rect 22336 21564 22342 21616
rect 22370 21564 22376 21616
rect 22428 21604 22434 21616
rect 22916 21607 22974 21613
rect 22428 21576 22692 21604
rect 22428 21564 22434 21576
rect 2222 21496 2228 21548
rect 2280 21496 2286 21548
rect 7282 21536 7288 21548
rect 7243 21508 7288 21536
rect 7282 21496 7288 21508
rect 7340 21496 7346 21548
rect 9950 21496 9956 21548
rect 10008 21536 10014 21548
rect 10226 21536 10232 21548
rect 10008 21508 10232 21536
rect 10008 21496 10014 21508
rect 10226 21496 10232 21508
rect 10284 21496 10290 21548
rect 13814 21496 13820 21548
rect 13872 21536 13878 21548
rect 14182 21536 14188 21548
rect 13872 21508 14188 21536
rect 13872 21496 13878 21508
rect 14182 21496 14188 21508
rect 14240 21496 14246 21548
rect 14458 21536 14464 21548
rect 14419 21508 14464 21536
rect 14458 21496 14464 21508
rect 14516 21496 14522 21548
rect 15378 21536 15384 21548
rect 15291 21508 15384 21536
rect 15378 21496 15384 21508
rect 15436 21536 15442 21548
rect 16482 21536 16488 21548
rect 15436 21508 16488 21536
rect 15436 21496 15442 21508
rect 16482 21496 16488 21508
rect 16540 21496 16546 21548
rect 19705 21539 19763 21545
rect 19705 21505 19717 21539
rect 19751 21505 19763 21539
rect 20162 21536 20168 21548
rect 20123 21508 20168 21536
rect 19705 21499 19763 21505
rect 2240 21332 2268 21496
rect 7466 21468 7472 21480
rect 7427 21440 7472 21468
rect 7466 21428 7472 21440
rect 7524 21428 7530 21480
rect 7745 21471 7803 21477
rect 7745 21468 7757 21471
rect 7576 21440 7757 21468
rect 3418 21360 3424 21412
rect 3476 21400 3482 21412
rect 7576 21400 7604 21440
rect 7745 21437 7757 21440
rect 7791 21437 7803 21471
rect 7745 21431 7803 21437
rect 11517 21471 11575 21477
rect 11517 21437 11529 21471
rect 11563 21437 11575 21471
rect 11517 21431 11575 21437
rect 11701 21471 11759 21477
rect 11701 21437 11713 21471
rect 11747 21468 11759 21471
rect 12158 21468 12164 21480
rect 11747 21440 12164 21468
rect 11747 21437 11759 21440
rect 11701 21431 11759 21437
rect 3476 21372 7604 21400
rect 3476 21360 3482 21372
rect 11532 21332 11560 21431
rect 12158 21428 12164 21440
rect 12216 21428 12222 21480
rect 13078 21468 13084 21480
rect 13039 21440 13084 21468
rect 13078 21428 13084 21440
rect 13136 21428 13142 21480
rect 14369 21471 14427 21477
rect 14369 21437 14381 21471
rect 14415 21468 14427 21471
rect 14642 21468 14648 21480
rect 14415 21440 14648 21468
rect 14415 21437 14427 21440
rect 14369 21431 14427 21437
rect 14642 21428 14648 21440
rect 14700 21428 14706 21480
rect 15286 21468 15292 21480
rect 15247 21440 15292 21468
rect 15286 21428 15292 21440
rect 15344 21428 15350 21480
rect 19720 21468 19748 21499
rect 20162 21496 20168 21508
rect 20220 21496 20226 21548
rect 21087 21539 21145 21545
rect 21087 21505 21099 21539
rect 21133 21505 21145 21539
rect 21087 21499 21145 21505
rect 20806 21468 20812 21480
rect 19720 21440 20812 21468
rect 20806 21428 20812 21440
rect 20864 21428 20870 21480
rect 21100 21468 21128 21499
rect 21266 21496 21272 21548
rect 21324 21536 21330 21548
rect 21821 21539 21879 21545
rect 21821 21536 21833 21539
rect 21324 21508 21833 21536
rect 21324 21496 21330 21508
rect 21821 21505 21833 21508
rect 21867 21505 21879 21539
rect 21821 21499 21879 21505
rect 22005 21539 22063 21545
rect 22005 21505 22017 21539
rect 22051 21536 22063 21539
rect 22554 21536 22560 21548
rect 22051 21508 22560 21536
rect 22051 21505 22063 21508
rect 22005 21499 22063 21505
rect 22554 21496 22560 21508
rect 22612 21496 22618 21548
rect 22664 21545 22692 21576
rect 22916 21573 22928 21607
rect 22962 21604 22974 21607
rect 23106 21604 23112 21616
rect 22962 21576 23112 21604
rect 22962 21573 22974 21576
rect 22916 21567 22974 21573
rect 23106 21564 23112 21576
rect 23164 21564 23170 21616
rect 22649 21539 22707 21545
rect 22649 21505 22661 21539
rect 22695 21505 22707 21539
rect 22649 21499 22707 21505
rect 22756 21508 24716 21536
rect 22370 21468 22376 21480
rect 21100 21440 22376 21468
rect 22370 21428 22376 21440
rect 22428 21428 22434 21480
rect 22756 21468 22784 21508
rect 22572 21440 22784 21468
rect 11606 21360 11612 21412
rect 11664 21400 11670 21412
rect 22572 21400 22600 21440
rect 24688 21400 24716 21508
rect 24780 21468 24808 21644
rect 25041 21641 25053 21675
rect 25087 21672 25099 21675
rect 25222 21672 25228 21684
rect 25087 21644 25228 21672
rect 25087 21641 25099 21644
rect 25041 21635 25099 21641
rect 25222 21632 25228 21644
rect 25280 21632 25286 21684
rect 25961 21675 26019 21681
rect 25961 21641 25973 21675
rect 26007 21672 26019 21675
rect 26050 21672 26056 21684
rect 26007 21644 26056 21672
rect 26007 21641 26019 21644
rect 25961 21635 26019 21641
rect 26050 21632 26056 21644
rect 26108 21632 26114 21684
rect 26234 21632 26240 21684
rect 26292 21672 26298 21684
rect 29822 21672 29828 21684
rect 26292 21644 29684 21672
rect 29783 21644 29828 21672
rect 26292 21632 26298 21644
rect 24854 21564 24860 21616
rect 24912 21604 24918 21616
rect 26329 21607 26387 21613
rect 26329 21604 26341 21607
rect 24912 21576 26341 21604
rect 24912 21564 24918 21576
rect 26329 21573 26341 21576
rect 26375 21573 26387 21607
rect 26329 21567 26387 21573
rect 26418 21564 26424 21616
rect 26476 21604 26482 21616
rect 26878 21604 26884 21616
rect 26476 21576 26884 21604
rect 26476 21564 26482 21576
rect 26878 21564 26884 21576
rect 26936 21604 26942 21616
rect 26973 21607 27031 21613
rect 26973 21604 26985 21607
rect 26936 21576 26985 21604
rect 26936 21564 26942 21576
rect 26973 21573 26985 21576
rect 27019 21573 27031 21607
rect 26973 21567 27031 21573
rect 27080 21576 28396 21604
rect 24946 21536 24952 21548
rect 24907 21508 24952 21536
rect 24946 21496 24952 21508
rect 25004 21496 25010 21548
rect 26050 21536 26056 21548
rect 26011 21508 26056 21536
rect 26050 21496 26056 21508
rect 26108 21496 26114 21548
rect 26142 21496 26148 21548
rect 26200 21536 26206 21548
rect 27080 21536 27108 21576
rect 27246 21536 27252 21548
rect 26200 21508 26245 21536
rect 26344 21508 27108 21536
rect 27207 21508 27252 21536
rect 26200 21496 26206 21508
rect 26344 21480 26372 21508
rect 27246 21496 27252 21508
rect 27304 21496 27310 21548
rect 28166 21496 28172 21548
rect 28224 21536 28230 21548
rect 28261 21539 28319 21545
rect 28261 21536 28273 21539
rect 28224 21508 28273 21536
rect 28224 21496 28230 21508
rect 28261 21505 28273 21508
rect 28307 21505 28319 21539
rect 28368 21536 28396 21576
rect 28442 21564 28448 21616
rect 28500 21604 28506 21616
rect 28718 21604 28724 21616
rect 28500 21576 28724 21604
rect 28500 21564 28506 21576
rect 28718 21564 28724 21576
rect 28776 21604 28782 21616
rect 29656 21604 29684 21644
rect 29822 21632 29828 21644
rect 29880 21632 29886 21684
rect 31294 21672 31300 21684
rect 29932 21644 31300 21672
rect 29932 21604 29960 21644
rect 31294 21632 31300 21644
rect 31352 21632 31358 21684
rect 31570 21672 31576 21684
rect 31531 21644 31576 21672
rect 31570 21632 31576 21644
rect 31628 21632 31634 21684
rect 31938 21632 31944 21684
rect 31996 21672 32002 21684
rect 32306 21672 32312 21684
rect 31996 21644 32312 21672
rect 31996 21632 32002 21644
rect 32306 21632 32312 21644
rect 32364 21632 32370 21684
rect 32582 21672 32588 21684
rect 32543 21644 32588 21672
rect 32582 21632 32588 21644
rect 32640 21632 32646 21684
rect 33137 21675 33195 21681
rect 33137 21641 33149 21675
rect 33183 21672 33195 21675
rect 33594 21672 33600 21684
rect 33183 21644 33600 21672
rect 33183 21641 33195 21644
rect 33137 21635 33195 21641
rect 33594 21632 33600 21644
rect 33652 21632 33658 21684
rect 36262 21632 36268 21684
rect 36320 21672 36326 21684
rect 36357 21675 36415 21681
rect 36357 21672 36369 21675
rect 36320 21644 36369 21672
rect 36320 21632 36326 21644
rect 36357 21641 36369 21644
rect 36403 21641 36415 21675
rect 37366 21672 37372 21684
rect 37327 21644 37372 21672
rect 36357 21635 36415 21641
rect 37366 21632 37372 21644
rect 37424 21632 37430 21684
rect 47854 21672 47860 21684
rect 45526 21644 47860 21672
rect 28776 21576 29500 21604
rect 29656 21576 29960 21604
rect 28776 21564 28782 21576
rect 28368 21508 28488 21536
rect 28261 21499 28319 21505
rect 25777 21471 25835 21477
rect 25777 21468 25789 21471
rect 24780 21440 25789 21468
rect 25777 21437 25789 21440
rect 25823 21468 25835 21471
rect 26326 21468 26332 21480
rect 25823 21440 26332 21468
rect 25823 21437 25835 21440
rect 25777 21431 25835 21437
rect 26326 21428 26332 21440
rect 26384 21428 26390 21480
rect 26418 21428 26424 21480
rect 26476 21468 26482 21480
rect 27157 21471 27215 21477
rect 27157 21468 27169 21471
rect 26476 21440 27169 21468
rect 26476 21428 26482 21440
rect 27157 21437 27169 21440
rect 27203 21468 27215 21471
rect 27338 21468 27344 21480
rect 27203 21440 27344 21468
rect 27203 21437 27215 21440
rect 27157 21431 27215 21437
rect 27338 21428 27344 21440
rect 27396 21468 27402 21480
rect 27614 21468 27620 21480
rect 27396 21440 27620 21468
rect 27396 21428 27402 21440
rect 27614 21428 27620 21440
rect 27672 21428 27678 21480
rect 28353 21471 28411 21477
rect 28353 21437 28365 21471
rect 28399 21437 28411 21471
rect 28460 21468 28488 21508
rect 28534 21496 28540 21548
rect 28592 21536 28598 21548
rect 29362 21536 29368 21548
rect 28592 21508 28637 21536
rect 29323 21508 29368 21536
rect 28592 21496 28598 21508
rect 29362 21496 29368 21508
rect 29420 21496 29426 21548
rect 29472 21536 29500 21576
rect 30006 21564 30012 21616
rect 30064 21604 30070 21616
rect 45526 21604 45554 21644
rect 47854 21632 47860 21644
rect 47912 21632 47918 21684
rect 47946 21604 47952 21616
rect 30064 21576 45554 21604
rect 47907 21576 47952 21604
rect 30064 21564 30070 21576
rect 47946 21564 47952 21576
rect 48004 21564 48010 21616
rect 29641 21539 29699 21545
rect 29641 21536 29653 21539
rect 29472 21508 29653 21536
rect 29641 21505 29653 21508
rect 29687 21505 29699 21539
rect 29641 21499 29699 21505
rect 30742 21496 30748 21548
rect 30800 21536 30806 21548
rect 31113 21539 31171 21545
rect 31113 21536 31125 21539
rect 30800 21508 31125 21536
rect 30800 21496 30806 21508
rect 31113 21505 31125 21508
rect 31159 21505 31171 21539
rect 31113 21499 31171 21505
rect 31389 21539 31447 21545
rect 31389 21505 31401 21539
rect 31435 21536 31447 21539
rect 31938 21536 31944 21548
rect 31435 21508 31944 21536
rect 31435 21505 31447 21508
rect 31389 21499 31447 21505
rect 31938 21496 31944 21508
rect 31996 21496 32002 21548
rect 32125 21539 32183 21545
rect 32125 21505 32137 21539
rect 32171 21505 32183 21539
rect 32125 21499 32183 21505
rect 32401 21539 32459 21545
rect 32401 21505 32413 21539
rect 32447 21536 32459 21539
rect 32490 21536 32496 21548
rect 32447 21508 32496 21536
rect 32447 21505 32459 21508
rect 32401 21499 32459 21505
rect 29454 21468 29460 21480
rect 28460 21440 29460 21468
rect 28353 21431 28411 21437
rect 26970 21400 26976 21412
rect 11664 21372 22600 21400
rect 23584 21372 24164 21400
rect 24688 21372 26976 21400
rect 11664 21360 11670 21372
rect 12250 21332 12256 21344
rect 2240 21304 12256 21332
rect 12250 21292 12256 21304
rect 12308 21292 12314 21344
rect 14090 21292 14096 21344
rect 14148 21332 14154 21344
rect 14461 21335 14519 21341
rect 14461 21332 14473 21335
rect 14148 21304 14473 21332
rect 14148 21292 14154 21304
rect 14461 21301 14473 21304
rect 14507 21332 14519 21335
rect 15378 21332 15384 21344
rect 14507 21304 15384 21332
rect 14507 21301 14519 21304
rect 14461 21295 14519 21301
rect 15378 21292 15384 21304
rect 15436 21292 15442 21344
rect 16758 21292 16764 21344
rect 16816 21332 16822 21344
rect 18230 21332 18236 21344
rect 16816 21304 18236 21332
rect 16816 21292 16822 21304
rect 18230 21292 18236 21304
rect 18288 21292 18294 21344
rect 20346 21332 20352 21344
rect 20307 21304 20352 21332
rect 20346 21292 20352 21304
rect 20404 21292 20410 21344
rect 20714 21292 20720 21344
rect 20772 21332 20778 21344
rect 21177 21335 21235 21341
rect 21177 21332 21189 21335
rect 20772 21304 21189 21332
rect 20772 21292 20778 21304
rect 21177 21301 21189 21304
rect 21223 21301 21235 21335
rect 21177 21295 21235 21301
rect 22189 21335 22247 21341
rect 22189 21301 22201 21335
rect 22235 21332 22247 21335
rect 22922 21332 22928 21344
rect 22235 21304 22928 21332
rect 22235 21301 22247 21304
rect 22189 21295 22247 21301
rect 22922 21292 22928 21304
rect 22980 21292 22986 21344
rect 23014 21292 23020 21344
rect 23072 21332 23078 21344
rect 23584 21332 23612 21372
rect 23072 21304 23612 21332
rect 23072 21292 23078 21304
rect 23658 21292 23664 21344
rect 23716 21332 23722 21344
rect 24029 21335 24087 21341
rect 24029 21332 24041 21335
rect 23716 21304 24041 21332
rect 23716 21292 23722 21304
rect 24029 21301 24041 21304
rect 24075 21301 24087 21335
rect 24136 21332 24164 21372
rect 26970 21360 26976 21372
rect 27028 21360 27034 21412
rect 28368 21400 28396 21431
rect 29454 21428 29460 21440
rect 29512 21428 29518 21480
rect 29549 21471 29607 21477
rect 29549 21437 29561 21471
rect 29595 21437 29607 21471
rect 29549 21431 29607 21437
rect 29089 21403 29147 21409
rect 27080 21372 27476 21400
rect 28368 21372 29040 21400
rect 27080 21332 27108 21372
rect 24136 21304 27108 21332
rect 27249 21335 27307 21341
rect 24029 21295 24087 21301
rect 27249 21301 27261 21335
rect 27295 21332 27307 21335
rect 27338 21332 27344 21344
rect 27295 21304 27344 21332
rect 27295 21301 27307 21304
rect 27249 21295 27307 21301
rect 27338 21292 27344 21304
rect 27396 21292 27402 21344
rect 27448 21341 27476 21372
rect 27433 21335 27491 21341
rect 27433 21301 27445 21335
rect 27479 21301 27491 21335
rect 28258 21332 28264 21344
rect 28219 21304 28264 21332
rect 27433 21295 27491 21301
rect 28258 21292 28264 21304
rect 28316 21292 28322 21344
rect 28721 21335 28779 21341
rect 28721 21301 28733 21335
rect 28767 21332 28779 21335
rect 28902 21332 28908 21344
rect 28767 21304 28908 21332
rect 28767 21301 28779 21304
rect 28721 21295 28779 21301
rect 28902 21292 28908 21304
rect 28960 21292 28966 21344
rect 29012 21332 29040 21372
rect 29089 21369 29101 21403
rect 29135 21400 29147 21403
rect 29564 21400 29592 21431
rect 30926 21428 30932 21480
rect 30984 21468 30990 21480
rect 31205 21471 31263 21477
rect 31205 21468 31217 21471
rect 30984 21440 31217 21468
rect 30984 21428 30990 21440
rect 31205 21437 31217 21440
rect 31251 21437 31263 21471
rect 32030 21468 32036 21480
rect 31205 21431 31263 21437
rect 31312 21440 32036 21468
rect 31312 21400 31340 21440
rect 32030 21428 32036 21440
rect 32088 21428 32094 21480
rect 32140 21400 32168 21499
rect 32490 21496 32496 21508
rect 32548 21496 32554 21548
rect 32950 21496 32956 21548
rect 33008 21536 33014 21548
rect 33045 21539 33103 21545
rect 33045 21536 33057 21539
rect 33008 21508 33057 21536
rect 33008 21496 33014 21508
rect 33045 21505 33057 21508
rect 33091 21505 33103 21539
rect 33045 21499 33103 21505
rect 36265 21539 36323 21545
rect 36265 21505 36277 21539
rect 36311 21536 36323 21539
rect 36354 21536 36360 21548
rect 36311 21508 36360 21536
rect 36311 21505 36323 21508
rect 36265 21499 36323 21505
rect 36354 21496 36360 21508
rect 36412 21496 36418 21548
rect 37274 21536 37280 21548
rect 37235 21508 37280 21536
rect 37274 21496 37280 21508
rect 37332 21496 37338 21548
rect 32306 21468 32312 21480
rect 32267 21440 32312 21468
rect 32306 21428 32312 21440
rect 32364 21428 32370 21480
rect 33410 21428 33416 21480
rect 33468 21468 33474 21480
rect 33689 21471 33747 21477
rect 33689 21468 33701 21471
rect 33468 21440 33701 21468
rect 33468 21428 33474 21440
rect 33689 21437 33701 21440
rect 33735 21437 33747 21471
rect 33870 21468 33876 21480
rect 33831 21440 33876 21468
rect 33689 21431 33747 21437
rect 33870 21428 33876 21440
rect 33928 21428 33934 21480
rect 35529 21471 35587 21477
rect 35529 21437 35541 21471
rect 35575 21468 35587 21471
rect 45462 21468 45468 21480
rect 35575 21440 45468 21468
rect 35575 21437 35587 21440
rect 35529 21431 35587 21437
rect 45462 21428 45468 21440
rect 45520 21428 45526 21480
rect 48222 21400 48228 21412
rect 29135 21372 31340 21400
rect 31404 21372 48228 21400
rect 29135 21369 29147 21372
rect 29089 21363 29147 21369
rect 29178 21332 29184 21344
rect 29012 21304 29184 21332
rect 29178 21292 29184 21304
rect 29236 21292 29242 21344
rect 29270 21292 29276 21344
rect 29328 21332 29334 21344
rect 29365 21335 29423 21341
rect 29365 21332 29377 21335
rect 29328 21304 29377 21332
rect 29328 21292 29334 21304
rect 29365 21301 29377 21304
rect 29411 21301 29423 21335
rect 29365 21295 29423 21301
rect 29454 21292 29460 21344
rect 29512 21332 29518 21344
rect 30745 21335 30803 21341
rect 30745 21332 30757 21335
rect 29512 21304 30757 21332
rect 29512 21292 29518 21304
rect 30745 21301 30757 21304
rect 30791 21332 30803 21335
rect 30926 21332 30932 21344
rect 30791 21304 30932 21332
rect 30791 21301 30803 21304
rect 30745 21295 30803 21301
rect 30926 21292 30932 21304
rect 30984 21292 30990 21344
rect 31404 21341 31432 21372
rect 48222 21360 48228 21372
rect 48280 21360 48286 21412
rect 31389 21335 31447 21341
rect 31389 21301 31401 21335
rect 31435 21301 31447 21335
rect 31389 21295 31447 21301
rect 31754 21292 31760 21344
rect 31812 21332 31818 21344
rect 32125 21335 32183 21341
rect 32125 21332 32137 21335
rect 31812 21304 32137 21332
rect 31812 21292 31818 21304
rect 32125 21301 32137 21304
rect 32171 21301 32183 21335
rect 32125 21295 32183 21301
rect 32766 21292 32772 21344
rect 32824 21332 32830 21344
rect 39942 21332 39948 21344
rect 32824 21304 39948 21332
rect 32824 21292 32830 21304
rect 39942 21292 39948 21304
rect 40000 21292 40006 21344
rect 48038 21332 48044 21344
rect 47999 21304 48044 21332
rect 48038 21292 48044 21304
rect 48096 21292 48102 21344
rect 1104 21242 48852 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 48852 21242
rect 1104 21168 48852 21190
rect 7466 21088 7472 21140
rect 7524 21128 7530 21140
rect 7561 21131 7619 21137
rect 7561 21128 7573 21131
rect 7524 21100 7573 21128
rect 7524 21088 7530 21100
rect 7561 21097 7573 21100
rect 7607 21097 7619 21131
rect 12158 21128 12164 21140
rect 12119 21100 12164 21128
rect 7561 21091 7619 21097
rect 12158 21088 12164 21100
rect 12216 21088 12222 21140
rect 12250 21088 12256 21140
rect 12308 21128 12314 21140
rect 20622 21128 20628 21140
rect 12308 21100 20628 21128
rect 12308 21088 12314 21100
rect 20622 21088 20628 21100
rect 20680 21088 20686 21140
rect 20806 21088 20812 21140
rect 20864 21128 20870 21140
rect 21266 21128 21272 21140
rect 20864 21100 21272 21128
rect 20864 21088 20870 21100
rect 21266 21088 21272 21100
rect 21324 21088 21330 21140
rect 22370 21088 22376 21140
rect 22428 21128 22434 21140
rect 22465 21131 22523 21137
rect 22465 21128 22477 21131
rect 22428 21100 22477 21128
rect 22428 21088 22434 21100
rect 22465 21097 22477 21100
rect 22511 21097 22523 21131
rect 22465 21091 22523 21097
rect 22554 21088 22560 21140
rect 22612 21128 22618 21140
rect 23658 21128 23664 21140
rect 22612 21100 23664 21128
rect 22612 21088 22618 21100
rect 23658 21088 23664 21100
rect 23716 21088 23722 21140
rect 25774 21088 25780 21140
rect 25832 21128 25838 21140
rect 27430 21128 27436 21140
rect 25832 21100 27436 21128
rect 25832 21088 25838 21100
rect 27430 21088 27436 21100
rect 27488 21088 27494 21140
rect 27522 21088 27528 21140
rect 27580 21128 27586 21140
rect 28353 21131 28411 21137
rect 28353 21128 28365 21131
rect 27580 21100 28365 21128
rect 27580 21088 27586 21100
rect 28353 21097 28365 21100
rect 28399 21128 28411 21131
rect 28442 21128 28448 21140
rect 28399 21100 28448 21128
rect 28399 21097 28411 21100
rect 28353 21091 28411 21097
rect 28442 21088 28448 21100
rect 28500 21088 28506 21140
rect 28810 21128 28816 21140
rect 28771 21100 28816 21128
rect 28810 21088 28816 21100
rect 28868 21088 28874 21140
rect 29825 21131 29883 21137
rect 29825 21097 29837 21131
rect 29871 21097 29883 21131
rect 29825 21091 29883 21097
rect 1394 21020 1400 21072
rect 1452 21060 1458 21072
rect 11606 21060 11612 21072
rect 1452 21032 11612 21060
rect 1452 21020 1458 21032
rect 11606 21020 11612 21032
rect 11664 21020 11670 21072
rect 13446 21060 13452 21072
rect 12406 21032 13452 21060
rect 12406 20992 12434 21032
rect 13446 21020 13452 21032
rect 13504 21020 13510 21072
rect 13538 21020 13544 21072
rect 13596 21060 13602 21072
rect 16666 21060 16672 21072
rect 13596 21032 16672 21060
rect 13596 21020 13602 21032
rect 16666 21020 16672 21032
rect 16724 21020 16730 21072
rect 26694 21060 26700 21072
rect 19306 21032 26700 21060
rect 7484 20964 12434 20992
rect 6822 20884 6828 20936
rect 6880 20924 6886 20936
rect 7484 20933 7512 20964
rect 12802 20952 12808 21004
rect 12860 20992 12866 21004
rect 14461 20995 14519 21001
rect 14461 20992 14473 20995
rect 12860 20964 13308 20992
rect 12860 20952 12866 20964
rect 7469 20927 7527 20933
rect 7469 20924 7481 20927
rect 6880 20896 7481 20924
rect 6880 20884 6886 20896
rect 7469 20893 7481 20896
rect 7515 20893 7527 20927
rect 7469 20887 7527 20893
rect 12069 20927 12127 20933
rect 12069 20893 12081 20927
rect 12115 20893 12127 20927
rect 12069 20887 12127 20893
rect 3970 20816 3976 20868
rect 4028 20856 4034 20868
rect 11606 20856 11612 20868
rect 4028 20828 11612 20856
rect 4028 20816 4034 20828
rect 11606 20816 11612 20828
rect 11664 20816 11670 20868
rect 12084 20856 12112 20887
rect 12342 20884 12348 20936
rect 12400 20924 12406 20936
rect 13280 20933 13308 20964
rect 13464 20964 14473 20992
rect 13153 20927 13211 20933
rect 12400 20921 13032 20924
rect 13153 20921 13165 20927
rect 12400 20896 13165 20921
rect 12400 20884 12406 20896
rect 13004 20893 13165 20896
rect 13199 20924 13211 20927
rect 13262 20927 13320 20933
rect 13199 20893 13216 20924
rect 13262 20893 13274 20927
rect 13308 20893 13320 20927
rect 13153 20887 13211 20893
rect 13262 20887 13320 20893
rect 13378 20927 13436 20933
rect 13378 20893 13390 20927
rect 13424 20924 13436 20927
rect 13464 20924 13492 20964
rect 14461 20961 14473 20964
rect 14507 20961 14519 20995
rect 16850 20992 16856 21004
rect 16811 20964 16856 20992
rect 14461 20955 14519 20961
rect 16850 20952 16856 20964
rect 16908 20952 16914 21004
rect 19306 20992 19334 21032
rect 26694 21020 26700 21032
rect 26752 21020 26758 21072
rect 29840 21060 29868 21091
rect 31018 21088 31024 21140
rect 31076 21128 31082 21140
rect 31205 21131 31263 21137
rect 31205 21128 31217 21131
rect 31076 21100 31217 21128
rect 31076 21088 31082 21100
rect 31205 21097 31217 21100
rect 31251 21097 31263 21131
rect 36170 21128 36176 21140
rect 31205 21091 31263 21097
rect 31352 21100 36176 21128
rect 31352 21060 31380 21100
rect 36170 21088 36176 21100
rect 36228 21088 36234 21140
rect 26804 21032 29776 21060
rect 29840 21032 31380 21060
rect 17880 20964 19334 20992
rect 13538 20933 13544 20936
rect 13424 20896 13492 20924
rect 13424 20893 13436 20896
rect 13378 20887 13436 20893
rect 13535 20887 13544 20933
rect 13538 20884 13544 20887
rect 13596 20884 13602 20936
rect 17402 20924 17408 20936
rect 14016 20896 17408 20924
rect 14016 20856 14044 20896
rect 17402 20884 17408 20896
rect 17460 20884 17466 20936
rect 17586 20884 17592 20936
rect 17644 20924 17650 20936
rect 17880 20924 17908 20964
rect 22370 20952 22376 21004
rect 22428 20992 22434 21004
rect 26804 21001 26832 21032
rect 25593 20995 25651 21001
rect 22428 20964 22876 20992
rect 22428 20952 22434 20964
rect 17644 20896 17908 20924
rect 19705 20927 19763 20933
rect 17644 20884 17650 20896
rect 19705 20893 19717 20927
rect 19751 20924 19763 20927
rect 20162 20924 20168 20936
rect 19751 20896 20168 20924
rect 19751 20893 19763 20896
rect 19705 20887 19763 20893
rect 20162 20884 20168 20896
rect 20220 20884 20226 20936
rect 20990 20924 20996 20936
rect 20951 20896 20996 20924
rect 20990 20884 20996 20896
rect 21048 20884 21054 20936
rect 21266 20924 21272 20936
rect 21227 20896 21272 20924
rect 21266 20884 21272 20896
rect 21324 20884 21330 20936
rect 22848 20933 22876 20964
rect 25593 20961 25605 20995
rect 25639 20992 25651 20995
rect 26789 20995 26847 21001
rect 25639 20964 26096 20992
rect 25639 20961 25651 20964
rect 25593 20955 25651 20961
rect 22741 20927 22799 20933
rect 22741 20893 22753 20927
rect 22787 20893 22799 20927
rect 22741 20887 22799 20893
rect 22833 20927 22891 20933
rect 22833 20893 22845 20927
rect 22879 20893 22891 20927
rect 22833 20887 22891 20893
rect 12084 20828 13216 20856
rect 4062 20748 4068 20800
rect 4120 20788 4126 20800
rect 5534 20788 5540 20800
rect 4120 20760 5540 20788
rect 4120 20748 4126 20760
rect 5534 20748 5540 20760
rect 5592 20748 5598 20800
rect 12894 20788 12900 20800
rect 12855 20760 12900 20788
rect 12894 20748 12900 20760
rect 12952 20748 12958 20800
rect 13188 20788 13216 20828
rect 13372 20828 14044 20856
rect 13372 20788 13400 20828
rect 14090 20816 14096 20868
rect 14148 20856 14154 20868
rect 14277 20859 14335 20865
rect 14148 20828 14193 20856
rect 14148 20816 14154 20828
rect 14277 20825 14289 20859
rect 14323 20856 14335 20859
rect 14366 20856 14372 20868
rect 14323 20828 14372 20856
rect 14323 20825 14335 20828
rect 14277 20819 14335 20825
rect 14366 20816 14372 20828
rect 14424 20816 14430 20868
rect 16758 20856 16764 20868
rect 14476 20828 16764 20856
rect 13188 20760 13400 20788
rect 13446 20748 13452 20800
rect 13504 20788 13510 20800
rect 14476 20788 14504 20828
rect 16758 20816 16764 20828
rect 16816 20816 16822 20868
rect 17120 20859 17178 20865
rect 17120 20825 17132 20859
rect 17166 20856 17178 20859
rect 17494 20856 17500 20868
rect 17166 20828 17500 20856
rect 17166 20825 17178 20828
rect 17120 20819 17178 20825
rect 17494 20816 17500 20828
rect 17552 20816 17558 20868
rect 22554 20856 22560 20868
rect 17604 20828 22560 20856
rect 13504 20760 14504 20788
rect 13504 20748 13510 20760
rect 14550 20748 14556 20800
rect 14608 20788 14614 20800
rect 17604 20788 17632 20828
rect 22554 20816 22560 20828
rect 22612 20816 22618 20868
rect 14608 20760 17632 20788
rect 14608 20748 14614 20760
rect 17770 20748 17776 20800
rect 17828 20788 17834 20800
rect 18233 20791 18291 20797
rect 18233 20788 18245 20791
rect 17828 20760 18245 20788
rect 17828 20748 17834 20760
rect 18233 20757 18245 20760
rect 18279 20757 18291 20791
rect 18233 20751 18291 20757
rect 18322 20748 18328 20800
rect 18380 20788 18386 20800
rect 19797 20791 19855 20797
rect 19797 20788 19809 20791
rect 18380 20760 19809 20788
rect 18380 20748 18386 20760
rect 19797 20757 19809 20760
rect 19843 20757 19855 20791
rect 19797 20751 19855 20757
rect 20990 20748 20996 20800
rect 21048 20788 21054 20800
rect 21358 20788 21364 20800
rect 21048 20760 21364 20788
rect 21048 20748 21054 20760
rect 21358 20748 21364 20760
rect 21416 20748 21422 20800
rect 22756 20788 22784 20887
rect 22922 20884 22928 20936
rect 22980 20924 22986 20936
rect 23109 20927 23167 20933
rect 22980 20896 23025 20924
rect 22980 20884 22986 20896
rect 23109 20893 23121 20927
rect 23155 20924 23167 20927
rect 25038 20924 25044 20936
rect 23155 20896 25044 20924
rect 23155 20893 23167 20896
rect 23109 20887 23167 20893
rect 25038 20884 25044 20896
rect 25096 20884 25102 20936
rect 25501 20927 25559 20933
rect 25501 20893 25513 20927
rect 25547 20893 25559 20927
rect 25501 20887 25559 20893
rect 25685 20927 25743 20933
rect 25685 20893 25697 20927
rect 25731 20924 25743 20927
rect 25774 20924 25780 20936
rect 25731 20896 25780 20924
rect 25731 20893 25743 20896
rect 25685 20887 25743 20893
rect 25516 20856 25544 20887
rect 25774 20884 25780 20896
rect 25832 20884 25838 20936
rect 26068 20924 26096 20964
rect 26789 20961 26801 20995
rect 26835 20961 26847 20995
rect 26789 20955 26847 20961
rect 26878 20952 26884 21004
rect 26936 20992 26942 21004
rect 27614 20992 27620 21004
rect 26936 20964 27476 20992
rect 27575 20964 27620 20992
rect 26936 20952 26942 20964
rect 26142 20924 26148 20936
rect 26055 20896 26148 20924
rect 26142 20884 26148 20896
rect 26200 20924 26206 20936
rect 27448 20933 27476 20964
rect 27614 20952 27620 20964
rect 27672 20952 27678 21004
rect 28445 20995 28503 21001
rect 28445 20961 28457 20995
rect 28491 20992 28503 20995
rect 28718 20992 28724 21004
rect 28491 20964 28724 20992
rect 28491 20961 28503 20964
rect 28445 20955 28503 20961
rect 28718 20952 28724 20964
rect 28776 20952 28782 21004
rect 29086 20952 29092 21004
rect 29144 20992 29150 21004
rect 29641 20995 29699 21001
rect 29641 20992 29653 20995
rect 29144 20964 29653 20992
rect 29144 20952 29150 20964
rect 29641 20961 29653 20964
rect 29687 20961 29699 20995
rect 29748 20992 29776 21032
rect 31570 21020 31576 21072
rect 31628 21060 31634 21072
rect 48038 21060 48044 21072
rect 31628 21032 48044 21060
rect 31628 21020 31634 21032
rect 48038 21020 48044 21032
rect 48096 21020 48102 21072
rect 30650 20992 30656 21004
rect 29748 20964 30656 20992
rect 29641 20955 29699 20961
rect 30650 20952 30656 20964
rect 30708 20952 30714 21004
rect 36078 20992 36084 21004
rect 36039 20964 36084 20992
rect 36078 20952 36084 20964
rect 36136 20952 36142 21004
rect 36262 20992 36268 21004
rect 36223 20964 36268 20992
rect 36262 20952 36268 20964
rect 36320 20952 36326 21004
rect 36354 20952 36360 21004
rect 36412 20992 36418 21004
rect 37826 20992 37832 21004
rect 36412 20964 37832 20992
rect 36412 20952 36418 20964
rect 37826 20952 37832 20964
rect 37884 20992 37890 21004
rect 37884 20964 38424 20992
rect 37884 20952 37890 20964
rect 26421 20927 26479 20933
rect 26421 20924 26433 20927
rect 26200 20896 26433 20924
rect 26200 20884 26206 20896
rect 26421 20893 26433 20896
rect 26467 20893 26479 20927
rect 26421 20887 26479 20893
rect 27433 20927 27491 20933
rect 27433 20893 27445 20927
rect 27479 20893 27491 20927
rect 27433 20887 27491 20893
rect 27709 20927 27767 20933
rect 27709 20893 27721 20927
rect 27755 20924 27767 20927
rect 27798 20924 27804 20936
rect 27755 20896 27804 20924
rect 27755 20893 27767 20896
rect 27709 20887 27767 20893
rect 27798 20884 27804 20896
rect 27856 20884 27862 20936
rect 28166 20884 28172 20936
rect 28224 20924 28230 20936
rect 28353 20927 28411 20933
rect 28353 20924 28365 20927
rect 28224 20896 28365 20924
rect 28224 20884 28230 20896
rect 28353 20893 28365 20896
rect 28399 20893 28411 20927
rect 28353 20887 28411 20893
rect 28534 20884 28540 20936
rect 28592 20924 28598 20936
rect 28629 20927 28687 20933
rect 28629 20924 28641 20927
rect 28592 20896 28641 20924
rect 28592 20884 28598 20896
rect 28629 20893 28641 20896
rect 28675 20893 28687 20927
rect 28629 20887 28687 20893
rect 28810 20884 28816 20936
rect 28868 20924 28874 20936
rect 29825 20927 29883 20933
rect 29825 20924 29837 20927
rect 28868 20896 29837 20924
rect 28868 20884 28874 20896
rect 29825 20893 29837 20896
rect 29871 20893 29883 20927
rect 31386 20924 31392 20936
rect 31347 20896 31392 20924
rect 29825 20887 29883 20893
rect 31386 20884 31392 20896
rect 31444 20884 31450 20936
rect 31481 20927 31539 20933
rect 31481 20893 31493 20927
rect 31527 20918 31539 20927
rect 31662 20924 31668 20936
rect 31588 20918 31668 20924
rect 31527 20896 31668 20918
rect 31527 20893 31616 20896
rect 31481 20890 31616 20893
rect 31481 20887 31539 20890
rect 31662 20884 31668 20896
rect 31720 20884 31726 20936
rect 33226 20884 33232 20936
rect 33284 20924 33290 20936
rect 38396 20933 38424 20964
rect 33413 20927 33471 20933
rect 33413 20924 33425 20927
rect 33284 20896 33425 20924
rect 33284 20884 33290 20896
rect 33413 20893 33425 20896
rect 33459 20893 33471 20927
rect 38381 20927 38439 20933
rect 33413 20887 33471 20893
rect 37476 20896 38056 20924
rect 26234 20856 26240 20868
rect 25516 20828 26240 20856
rect 26234 20816 26240 20828
rect 26292 20816 26298 20868
rect 26329 20859 26387 20865
rect 26329 20825 26341 20859
rect 26375 20856 26387 20859
rect 27246 20856 27252 20868
rect 26375 20828 27252 20856
rect 26375 20825 26387 20828
rect 26329 20819 26387 20825
rect 27246 20816 27252 20828
rect 27304 20816 27310 20868
rect 27724 20828 28028 20856
rect 27724 20788 27752 20828
rect 27890 20788 27896 20800
rect 22756 20760 27752 20788
rect 27851 20760 27896 20788
rect 27890 20748 27896 20760
rect 27948 20748 27954 20800
rect 28000 20788 28028 20828
rect 28902 20816 28908 20868
rect 28960 20856 28966 20868
rect 29549 20859 29607 20865
rect 29549 20856 29561 20859
rect 28960 20828 29561 20856
rect 28960 20816 28966 20828
rect 29549 20825 29561 20828
rect 29595 20825 29607 20859
rect 31202 20856 31208 20868
rect 31115 20828 31208 20856
rect 29549 20819 29607 20825
rect 31202 20816 31208 20828
rect 31260 20856 31266 20868
rect 31754 20856 31760 20868
rect 31260 20828 31760 20856
rect 31260 20816 31266 20828
rect 31754 20816 31760 20828
rect 31812 20816 31818 20868
rect 32030 20816 32036 20868
rect 32088 20856 32094 20868
rect 37476 20856 37504 20896
rect 37918 20856 37924 20868
rect 32088 20828 37504 20856
rect 37879 20828 37924 20856
rect 32088 20816 32094 20828
rect 37918 20816 37924 20828
rect 37976 20816 37982 20868
rect 38028 20856 38056 20896
rect 38381 20893 38393 20927
rect 38427 20893 38439 20927
rect 38381 20887 38439 20893
rect 47670 20856 47676 20868
rect 38028 20828 47676 20856
rect 47670 20816 47676 20828
rect 47728 20816 47734 20868
rect 29914 20788 29920 20800
rect 28000 20760 29920 20788
rect 29914 20748 29920 20760
rect 29972 20748 29978 20800
rect 30006 20748 30012 20800
rect 30064 20788 30070 20800
rect 30064 20760 30109 20788
rect 30064 20748 30070 20760
rect 31110 20748 31116 20800
rect 31168 20788 31174 20800
rect 31665 20791 31723 20797
rect 31665 20788 31677 20791
rect 31168 20760 31677 20788
rect 31168 20748 31174 20760
rect 31665 20757 31677 20760
rect 31711 20757 31723 20791
rect 31665 20751 31723 20757
rect 33505 20791 33563 20797
rect 33505 20757 33517 20791
rect 33551 20788 33563 20791
rect 33686 20788 33692 20800
rect 33551 20760 33692 20788
rect 33551 20757 33563 20760
rect 33505 20751 33563 20757
rect 33686 20748 33692 20760
rect 33744 20748 33750 20800
rect 37458 20748 37464 20800
rect 37516 20788 37522 20800
rect 38473 20791 38531 20797
rect 38473 20788 38485 20791
rect 37516 20760 38485 20788
rect 37516 20748 37522 20760
rect 38473 20757 38485 20760
rect 38519 20757 38531 20791
rect 38473 20751 38531 20757
rect 1104 20698 48852 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 48852 20698
rect 1104 20624 48852 20646
rect 7926 20584 7932 20596
rect 4816 20556 7932 20584
rect 4816 20457 4844 20556
rect 7926 20544 7932 20556
rect 7984 20584 7990 20596
rect 17126 20584 17132 20596
rect 7984 20556 17132 20584
rect 7984 20544 7990 20556
rect 17126 20544 17132 20556
rect 17184 20544 17190 20596
rect 17494 20584 17500 20596
rect 17455 20556 17500 20584
rect 17494 20544 17500 20556
rect 17552 20544 17558 20596
rect 17862 20544 17868 20596
rect 17920 20544 17926 20596
rect 17954 20544 17960 20596
rect 18012 20584 18018 20596
rect 41598 20584 41604 20596
rect 18012 20556 41604 20584
rect 18012 20544 18018 20556
rect 41598 20544 41604 20556
rect 41656 20544 41662 20596
rect 12894 20476 12900 20528
rect 12952 20516 12958 20528
rect 13326 20519 13384 20525
rect 13326 20516 13338 20519
rect 12952 20488 13338 20516
rect 12952 20476 12958 20488
rect 13326 20485 13338 20488
rect 13372 20485 13384 20519
rect 13326 20479 13384 20485
rect 17880 20463 17908 20544
rect 19334 20476 19340 20528
rect 19392 20516 19398 20528
rect 20346 20516 20352 20528
rect 19392 20488 20352 20516
rect 19392 20476 19398 20488
rect 20346 20476 20352 20488
rect 20404 20516 20410 20528
rect 22649 20519 22707 20525
rect 20404 20488 22600 20516
rect 20404 20476 20410 20488
rect 4801 20451 4859 20457
rect 4801 20417 4813 20451
rect 4847 20417 4859 20451
rect 4801 20411 4859 20417
rect 10502 20408 10508 20460
rect 10560 20448 10566 20460
rect 11517 20451 11575 20457
rect 11517 20448 11529 20451
rect 10560 20420 11529 20448
rect 10560 20408 10566 20420
rect 11517 20417 11529 20420
rect 11563 20417 11575 20451
rect 11698 20448 11704 20460
rect 11659 20420 11704 20448
rect 11517 20411 11575 20417
rect 11698 20408 11704 20420
rect 11756 20408 11762 20460
rect 12986 20408 12992 20460
rect 13044 20448 13050 20460
rect 13081 20451 13139 20457
rect 13081 20448 13093 20451
rect 13044 20420 13093 20448
rect 13044 20408 13050 20420
rect 13081 20417 13093 20420
rect 13127 20417 13139 20451
rect 15746 20448 15752 20460
rect 15707 20420 15752 20448
rect 13081 20411 13139 20417
rect 15746 20408 15752 20420
rect 15804 20408 15810 20460
rect 15841 20451 15899 20457
rect 15841 20417 15853 20451
rect 15887 20417 15899 20451
rect 15841 20411 15899 20417
rect 8754 20380 8760 20392
rect 8715 20352 8760 20380
rect 8754 20340 8760 20352
rect 8812 20340 8818 20392
rect 8938 20380 8944 20392
rect 8899 20352 8944 20380
rect 8938 20340 8944 20352
rect 8996 20340 9002 20392
rect 10410 20380 10416 20392
rect 10371 20352 10416 20380
rect 10410 20340 10416 20352
rect 10468 20340 10474 20392
rect 15856 20380 15884 20411
rect 15930 20408 15936 20460
rect 15988 20448 15994 20460
rect 16117 20451 16175 20457
rect 15988 20420 16033 20448
rect 15988 20408 15994 20420
rect 16117 20417 16129 20451
rect 16163 20448 16175 20451
rect 17310 20448 17316 20460
rect 16163 20420 17316 20448
rect 16163 20417 16175 20420
rect 16117 20411 16175 20417
rect 17310 20408 17316 20420
rect 17368 20408 17374 20460
rect 17862 20457 17920 20463
rect 17753 20451 17811 20457
rect 17753 20448 17765 20451
rect 17696 20420 17765 20448
rect 14292 20352 15884 20380
rect 4890 20244 4896 20256
rect 4851 20216 4896 20244
rect 4890 20204 4896 20216
rect 4948 20204 4954 20256
rect 11885 20247 11943 20253
rect 11885 20213 11897 20247
rect 11931 20244 11943 20247
rect 11974 20244 11980 20256
rect 11931 20216 11980 20244
rect 11931 20213 11943 20216
rect 11885 20207 11943 20213
rect 11974 20204 11980 20216
rect 12032 20204 12038 20256
rect 12802 20204 12808 20256
rect 12860 20244 12866 20256
rect 14292 20244 14320 20352
rect 14458 20244 14464 20256
rect 12860 20216 14320 20244
rect 14419 20216 14464 20244
rect 12860 20204 12866 20216
rect 14458 20204 14464 20216
rect 14516 20204 14522 20256
rect 15470 20244 15476 20256
rect 15431 20216 15476 20244
rect 15470 20204 15476 20216
rect 15528 20204 15534 20256
rect 15856 20244 15884 20352
rect 17221 20383 17279 20389
rect 17221 20349 17233 20383
rect 17267 20380 17279 20383
rect 17696 20380 17724 20420
rect 17753 20417 17765 20420
rect 17799 20417 17811 20451
rect 17862 20423 17874 20457
rect 17908 20423 17920 20457
rect 17862 20417 17920 20423
rect 17957 20451 18015 20457
rect 17957 20417 17969 20451
rect 18003 20417 18015 20451
rect 17753 20411 17811 20417
rect 17957 20411 18015 20417
rect 17267 20352 17724 20380
rect 17972 20380 18000 20411
rect 18138 20408 18144 20460
rect 18196 20448 18202 20460
rect 18877 20451 18935 20457
rect 18196 20420 18241 20448
rect 18196 20408 18202 20420
rect 18877 20417 18889 20451
rect 18923 20448 18935 20451
rect 19242 20448 19248 20460
rect 18923 20420 19248 20448
rect 18923 20417 18935 20420
rect 18877 20411 18935 20417
rect 19242 20408 19248 20420
rect 19300 20408 19306 20460
rect 19610 20408 19616 20460
rect 19668 20448 19674 20460
rect 19788 20451 19846 20457
rect 19788 20448 19800 20451
rect 19668 20420 19800 20448
rect 19668 20408 19674 20420
rect 19788 20417 19800 20420
rect 19834 20417 19846 20451
rect 19788 20411 19846 20417
rect 21726 20408 21732 20460
rect 21784 20448 21790 20460
rect 21821 20451 21879 20457
rect 21821 20448 21833 20451
rect 21784 20420 21833 20448
rect 21784 20408 21790 20420
rect 21821 20417 21833 20420
rect 21867 20417 21879 20451
rect 21821 20411 21879 20417
rect 21910 20408 21916 20460
rect 21968 20448 21974 20460
rect 22005 20451 22063 20457
rect 22005 20448 22017 20451
rect 21968 20420 22017 20448
rect 21968 20408 21974 20420
rect 22005 20417 22017 20420
rect 22051 20417 22063 20451
rect 22005 20411 22063 20417
rect 22097 20451 22155 20457
rect 22097 20417 22109 20451
rect 22143 20417 22155 20451
rect 22572 20448 22600 20488
rect 22649 20485 22661 20519
rect 22695 20516 22707 20519
rect 23014 20516 23020 20528
rect 22695 20488 23020 20516
rect 22695 20485 22707 20488
rect 22649 20479 22707 20485
rect 23014 20476 23020 20488
rect 23072 20476 23078 20528
rect 23106 20476 23112 20528
rect 23164 20516 23170 20528
rect 25130 20516 25136 20528
rect 23164 20488 25136 20516
rect 23164 20476 23170 20488
rect 25130 20476 25136 20488
rect 25188 20476 25194 20528
rect 27433 20519 27491 20525
rect 27433 20485 27445 20519
rect 27479 20516 27491 20519
rect 27890 20516 27896 20528
rect 27479 20488 27896 20516
rect 27479 20485 27491 20488
rect 27433 20479 27491 20485
rect 27890 20476 27896 20488
rect 27948 20476 27954 20528
rect 30561 20519 30619 20525
rect 28920 20488 29776 20516
rect 28920 20460 28948 20488
rect 23842 20448 23848 20460
rect 22572 20420 23848 20448
rect 22097 20411 22155 20417
rect 18046 20380 18052 20392
rect 17972 20352 18052 20380
rect 17267 20349 17279 20352
rect 17221 20343 17279 20349
rect 17696 20312 17724 20352
rect 18046 20340 18052 20352
rect 18104 20340 18110 20392
rect 19426 20340 19432 20392
rect 19484 20380 19490 20392
rect 19521 20383 19579 20389
rect 19521 20380 19533 20383
rect 19484 20352 19533 20380
rect 19484 20340 19490 20352
rect 19521 20349 19533 20352
rect 19567 20349 19579 20383
rect 22112 20380 22140 20411
rect 23842 20408 23848 20420
rect 23900 20408 23906 20460
rect 28258 20408 28264 20460
rect 28316 20448 28322 20460
rect 28629 20451 28687 20457
rect 28629 20448 28641 20451
rect 28316 20420 28641 20448
rect 28316 20408 28322 20420
rect 28629 20417 28641 20420
rect 28675 20417 28687 20451
rect 28902 20448 28908 20460
rect 28863 20420 28908 20448
rect 28629 20411 28687 20417
rect 28902 20408 28908 20420
rect 28960 20408 28966 20460
rect 29748 20457 29776 20488
rect 30561 20485 30573 20519
rect 30607 20516 30619 20519
rect 30834 20516 30840 20528
rect 30607 20488 30840 20516
rect 30607 20485 30619 20488
rect 30561 20479 30619 20485
rect 30834 20476 30840 20488
rect 30892 20476 30898 20528
rect 31386 20476 31392 20528
rect 31444 20516 31450 20528
rect 31938 20516 31944 20528
rect 31444 20488 31944 20516
rect 31444 20476 31450 20488
rect 31938 20476 31944 20488
rect 31996 20516 32002 20528
rect 32490 20516 32496 20528
rect 31996 20488 32496 20516
rect 31996 20476 32002 20488
rect 32490 20476 32496 20488
rect 32548 20476 32554 20528
rect 33686 20516 33692 20528
rect 33647 20488 33692 20516
rect 33686 20476 33692 20488
rect 33744 20476 33750 20528
rect 37458 20516 37464 20528
rect 37419 20488 37464 20516
rect 37458 20476 37464 20488
rect 37516 20476 37522 20528
rect 39022 20476 39028 20528
rect 39080 20516 39086 20528
rect 39117 20519 39175 20525
rect 39117 20516 39129 20519
rect 39080 20488 39129 20516
rect 39080 20476 39086 20488
rect 39117 20485 39129 20488
rect 39163 20485 39175 20519
rect 39117 20479 39175 20485
rect 29549 20451 29607 20457
rect 29549 20417 29561 20451
rect 29595 20417 29607 20451
rect 29549 20411 29607 20417
rect 29733 20451 29791 20457
rect 29733 20417 29745 20451
rect 29779 20417 29791 20451
rect 29733 20411 29791 20417
rect 29825 20451 29883 20457
rect 29825 20417 29837 20451
rect 29871 20417 29883 20451
rect 29825 20411 29883 20417
rect 23750 20380 23756 20392
rect 22112 20352 23756 20380
rect 19521 20343 19579 20349
rect 23750 20340 23756 20352
rect 23808 20340 23814 20392
rect 24026 20380 24032 20392
rect 23987 20352 24032 20380
rect 24026 20340 24032 20352
rect 24084 20380 24090 20392
rect 24946 20380 24952 20392
rect 24084 20352 24952 20380
rect 24084 20340 24090 20352
rect 24946 20340 24952 20352
rect 25004 20340 25010 20392
rect 28810 20380 28816 20392
rect 28771 20352 28816 20380
rect 28810 20340 28816 20352
rect 28868 20340 28874 20392
rect 29564 20380 29592 20411
rect 28920 20352 29592 20380
rect 21821 20315 21879 20321
rect 17696 20284 19104 20312
rect 17218 20244 17224 20256
rect 15856 20216 17224 20244
rect 17218 20204 17224 20216
rect 17276 20244 17282 20256
rect 17862 20244 17868 20256
rect 17276 20216 17868 20244
rect 17276 20204 17282 20216
rect 17862 20204 17868 20216
rect 17920 20244 17926 20256
rect 18969 20247 19027 20253
rect 18969 20244 18981 20247
rect 17920 20216 18981 20244
rect 17920 20204 17926 20216
rect 18969 20213 18981 20216
rect 19015 20213 19027 20247
rect 19076 20244 19104 20284
rect 20456 20284 21220 20312
rect 20456 20244 20484 20284
rect 19076 20216 20484 20244
rect 20901 20247 20959 20253
rect 18969 20207 19027 20213
rect 20901 20213 20913 20247
rect 20947 20244 20959 20247
rect 21082 20244 21088 20256
rect 20947 20216 21088 20244
rect 20947 20213 20959 20216
rect 20901 20207 20959 20213
rect 21082 20204 21088 20216
rect 21140 20204 21146 20256
rect 21192 20244 21220 20284
rect 21821 20281 21833 20315
rect 21867 20312 21879 20315
rect 22002 20312 22008 20324
rect 21867 20284 22008 20312
rect 21867 20281 21879 20284
rect 21821 20275 21879 20281
rect 22002 20272 22008 20284
rect 22060 20272 22066 20324
rect 22554 20272 22560 20324
rect 22612 20312 22618 20324
rect 28920 20312 28948 20352
rect 29086 20312 29092 20324
rect 22612 20284 28948 20312
rect 29047 20284 29092 20312
rect 22612 20272 22618 20284
rect 22186 20244 22192 20256
rect 21192 20216 22192 20244
rect 22186 20204 22192 20216
rect 22244 20204 22250 20256
rect 22370 20204 22376 20256
rect 22428 20244 22434 20256
rect 22741 20247 22799 20253
rect 22741 20244 22753 20247
rect 22428 20216 22753 20244
rect 22428 20204 22434 20216
rect 22741 20213 22753 20216
rect 22787 20213 22799 20247
rect 22741 20207 22799 20213
rect 22922 20204 22928 20256
rect 22980 20244 22986 20256
rect 27709 20247 27767 20253
rect 27709 20244 27721 20247
rect 22980 20216 27721 20244
rect 22980 20204 22986 20216
rect 27709 20213 27721 20216
rect 27755 20244 27767 20247
rect 27798 20244 27804 20256
rect 27755 20216 27804 20244
rect 27755 20213 27767 20216
rect 27709 20207 27767 20213
rect 27798 20204 27804 20216
rect 27856 20204 27862 20256
rect 28644 20253 28672 20284
rect 29086 20272 29092 20284
rect 29144 20272 29150 20324
rect 29270 20272 29276 20324
rect 29328 20312 29334 20324
rect 29840 20312 29868 20411
rect 30926 20408 30932 20460
rect 30984 20448 30990 20460
rect 31113 20451 31171 20457
rect 31113 20448 31125 20451
rect 30984 20420 31125 20448
rect 30984 20408 30990 20420
rect 31113 20417 31125 20420
rect 31159 20417 31171 20451
rect 31113 20411 31171 20417
rect 32861 20451 32919 20457
rect 32861 20417 32873 20451
rect 32907 20448 32919 20451
rect 33226 20448 33232 20460
rect 32907 20420 33232 20448
rect 32907 20417 32919 20420
rect 32861 20411 32919 20417
rect 33226 20408 33232 20420
rect 33284 20408 33290 20460
rect 45830 20408 45836 20460
rect 45888 20448 45894 20460
rect 47486 20448 47492 20460
rect 45888 20420 47492 20448
rect 45888 20408 45894 20420
rect 47486 20408 47492 20420
rect 47544 20448 47550 20460
rect 47581 20451 47639 20457
rect 47581 20448 47593 20451
rect 47544 20420 47593 20448
rect 47544 20408 47550 20420
rect 47581 20417 47593 20420
rect 47627 20417 47639 20451
rect 47581 20411 47639 20417
rect 31021 20383 31079 20389
rect 31021 20349 31033 20383
rect 31067 20380 31079 20383
rect 31478 20380 31484 20392
rect 31067 20352 31484 20380
rect 31067 20349 31079 20352
rect 31021 20343 31079 20349
rect 31478 20340 31484 20352
rect 31536 20340 31542 20392
rect 33505 20383 33563 20389
rect 33505 20349 33517 20383
rect 33551 20380 33563 20383
rect 33778 20380 33784 20392
rect 33551 20352 33784 20380
rect 33551 20349 33563 20352
rect 33505 20343 33563 20349
rect 33778 20340 33784 20352
rect 33836 20340 33842 20392
rect 34054 20380 34060 20392
rect 34015 20352 34060 20380
rect 34054 20340 34060 20352
rect 34112 20340 34118 20392
rect 37277 20383 37335 20389
rect 37277 20380 37289 20383
rect 35452 20352 37289 20380
rect 29328 20284 29868 20312
rect 29328 20272 29334 20284
rect 30374 20272 30380 20324
rect 30432 20312 30438 20324
rect 31297 20315 31355 20321
rect 31297 20312 31309 20315
rect 30432 20284 31309 20312
rect 30432 20272 30438 20284
rect 31297 20281 31309 20284
rect 31343 20281 31355 20315
rect 31297 20275 31355 20281
rect 31386 20272 31392 20324
rect 31444 20312 31450 20324
rect 35452 20312 35480 20352
rect 37277 20349 37289 20352
rect 37323 20349 37335 20383
rect 37277 20343 37335 20349
rect 31444 20284 35480 20312
rect 31444 20272 31450 20284
rect 36538 20272 36544 20324
rect 36596 20312 36602 20324
rect 46106 20312 46112 20324
rect 36596 20284 46112 20312
rect 36596 20272 36602 20284
rect 46106 20272 46112 20284
rect 46164 20272 46170 20324
rect 28629 20247 28687 20253
rect 28629 20213 28641 20247
rect 28675 20213 28687 20247
rect 28629 20207 28687 20213
rect 29454 20204 29460 20256
rect 29512 20244 29518 20256
rect 29549 20247 29607 20253
rect 29549 20244 29561 20247
rect 29512 20216 29561 20244
rect 29512 20204 29518 20216
rect 29549 20213 29561 20216
rect 29595 20213 29607 20247
rect 29549 20207 29607 20213
rect 30009 20247 30067 20253
rect 30009 20213 30021 20247
rect 30055 20244 30067 20247
rect 30190 20244 30196 20256
rect 30055 20216 30196 20244
rect 30055 20213 30067 20216
rect 30009 20207 30067 20213
rect 30190 20204 30196 20216
rect 30248 20204 30254 20256
rect 30742 20204 30748 20256
rect 30800 20244 30806 20256
rect 30837 20247 30895 20253
rect 30837 20244 30849 20247
rect 30800 20216 30849 20244
rect 30800 20204 30806 20216
rect 30837 20213 30849 20216
rect 30883 20213 30895 20247
rect 30837 20207 30895 20213
rect 32953 20247 33011 20253
rect 32953 20213 32965 20247
rect 32999 20244 33011 20247
rect 33318 20244 33324 20256
rect 32999 20216 33324 20244
rect 32999 20213 33011 20216
rect 32953 20207 33011 20213
rect 33318 20204 33324 20216
rect 33376 20204 33382 20256
rect 46474 20204 46480 20256
rect 46532 20244 46538 20256
rect 47673 20247 47731 20253
rect 47673 20244 47685 20247
rect 46532 20216 47685 20244
rect 46532 20204 46538 20216
rect 47673 20213 47685 20216
rect 47719 20213 47731 20247
rect 47673 20207 47731 20213
rect 1104 20154 48852 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 48852 20154
rect 1104 20080 48852 20102
rect 8297 20043 8355 20049
rect 8297 20009 8309 20043
rect 8343 20040 8355 20043
rect 8938 20040 8944 20052
rect 8343 20012 8944 20040
rect 8343 20009 8355 20012
rect 8297 20003 8355 20009
rect 8938 20000 8944 20012
rect 8996 20000 9002 20052
rect 11698 20040 11704 20052
rect 9416 20012 11704 20040
rect 9416 19972 9444 20012
rect 11698 20000 11704 20012
rect 11756 20000 11762 20052
rect 14737 20043 14795 20049
rect 14737 20009 14749 20043
rect 14783 20040 14795 20043
rect 15930 20040 15936 20052
rect 14783 20012 15936 20040
rect 14783 20009 14795 20012
rect 14737 20003 14795 20009
rect 15930 20000 15936 20012
rect 15988 20000 15994 20052
rect 16666 20000 16672 20052
rect 16724 20040 16730 20052
rect 16945 20043 17003 20049
rect 16945 20040 16957 20043
rect 16724 20012 16957 20040
rect 16724 20000 16730 20012
rect 16945 20009 16957 20012
rect 16991 20009 17003 20043
rect 16945 20003 17003 20009
rect 17681 20043 17739 20049
rect 17681 20009 17693 20043
rect 17727 20040 17739 20043
rect 18046 20040 18052 20052
rect 17727 20012 18052 20040
rect 17727 20009 17739 20012
rect 17681 20003 17739 20009
rect 18046 20000 18052 20012
rect 18104 20000 18110 20052
rect 19610 20000 19616 20052
rect 19668 20040 19674 20052
rect 19705 20043 19763 20049
rect 19705 20040 19717 20043
rect 19668 20012 19717 20040
rect 19668 20000 19674 20012
rect 19705 20009 19717 20012
rect 19751 20009 19763 20043
rect 24026 20040 24032 20052
rect 19705 20003 19763 20009
rect 19904 20012 24032 20040
rect 15194 19972 15200 19984
rect 4724 19944 9444 19972
rect 12912 19944 15200 19972
rect 4724 19913 4752 19944
rect 4709 19907 4767 19913
rect 4709 19873 4721 19907
rect 4755 19873 4767 19907
rect 4890 19904 4896 19916
rect 4851 19876 4896 19904
rect 4709 19867 4767 19873
rect 4890 19864 4896 19876
rect 4948 19864 4954 19916
rect 5534 19904 5540 19916
rect 5495 19876 5540 19904
rect 5534 19864 5540 19876
rect 5592 19864 5598 19916
rect 8018 19864 8024 19916
rect 8076 19904 8082 19916
rect 10321 19907 10379 19913
rect 10321 19904 10333 19907
rect 8076 19876 10333 19904
rect 8076 19864 8082 19876
rect 10321 19873 10333 19876
rect 10367 19873 10379 19907
rect 12621 19907 12679 19913
rect 12621 19904 12633 19907
rect 10321 19867 10379 19873
rect 11348 19876 12633 19904
rect 1762 19796 1768 19848
rect 1820 19836 1826 19848
rect 2041 19839 2099 19845
rect 2041 19836 2053 19839
rect 1820 19808 2053 19836
rect 1820 19796 1826 19808
rect 2041 19805 2053 19808
rect 2087 19805 2099 19839
rect 2041 19799 2099 19805
rect 8205 19839 8263 19845
rect 8205 19805 8217 19839
rect 8251 19805 8263 19839
rect 8205 19799 8263 19805
rect 8220 19768 8248 19799
rect 9398 19796 9404 19848
rect 9456 19845 9462 19848
rect 9456 19839 9505 19845
rect 9456 19805 9459 19839
rect 9493 19805 9505 19839
rect 9582 19836 9588 19848
rect 9543 19808 9588 19836
rect 9456 19799 9505 19805
rect 9456 19796 9462 19799
rect 9582 19796 9588 19808
rect 9640 19796 9646 19848
rect 9674 19796 9680 19848
rect 9732 19836 9738 19848
rect 9861 19839 9919 19845
rect 9732 19808 9777 19836
rect 9732 19796 9738 19808
rect 9861 19805 9873 19839
rect 9907 19836 9919 19839
rect 10226 19836 10232 19848
rect 9907 19808 10232 19836
rect 9907 19805 9919 19808
rect 9861 19799 9919 19805
rect 10226 19796 10232 19808
rect 10284 19796 10290 19848
rect 10410 19796 10416 19848
rect 10468 19836 10474 19848
rect 11348 19836 11376 19876
rect 12621 19873 12633 19876
rect 12667 19873 12679 19907
rect 12621 19867 12679 19873
rect 10468 19808 11376 19836
rect 12069 19839 12127 19845
rect 10468 19796 10474 19808
rect 12069 19805 12081 19839
rect 12115 19836 12127 19839
rect 12345 19839 12403 19845
rect 12345 19836 12357 19839
rect 12115 19808 12357 19836
rect 12115 19805 12127 19808
rect 12069 19799 12127 19805
rect 12345 19805 12357 19808
rect 12391 19836 12403 19839
rect 12912 19836 12940 19944
rect 15194 19932 15200 19944
rect 15252 19932 15258 19984
rect 17126 19932 17132 19984
rect 17184 19972 17190 19984
rect 19904 19972 19932 20012
rect 24026 20000 24032 20012
rect 24084 20000 24090 20052
rect 28258 20000 28264 20052
rect 28316 20040 28322 20052
rect 28445 20043 28503 20049
rect 28445 20040 28457 20043
rect 28316 20012 28457 20040
rect 28316 20000 28322 20012
rect 28445 20009 28457 20012
rect 28491 20009 28503 20043
rect 28445 20003 28503 20009
rect 28905 20043 28963 20049
rect 28905 20009 28917 20043
rect 28951 20040 28963 20043
rect 29362 20040 29368 20052
rect 28951 20012 29368 20040
rect 28951 20009 28963 20012
rect 28905 20003 28963 20009
rect 29362 20000 29368 20012
rect 29420 20000 29426 20052
rect 30374 20040 30380 20052
rect 30335 20012 30380 20040
rect 30374 20000 30380 20012
rect 30432 20000 30438 20052
rect 30558 20040 30564 20052
rect 30519 20012 30564 20040
rect 30558 20000 30564 20012
rect 30616 20000 30622 20052
rect 30834 20000 30840 20052
rect 30892 20040 30898 20052
rect 33870 20040 33876 20052
rect 30892 20012 31754 20040
rect 33831 20012 33876 20040
rect 30892 20000 30898 20012
rect 20901 19975 20959 19981
rect 20901 19972 20913 19975
rect 17184 19944 19932 19972
rect 19996 19944 20913 19972
rect 17184 19932 17190 19944
rect 16206 19864 16212 19916
rect 16264 19904 16270 19916
rect 19996 19904 20024 19944
rect 20901 19941 20913 19944
rect 20947 19941 20959 19975
rect 20901 19935 20959 19941
rect 21726 19932 21732 19984
rect 21784 19972 21790 19984
rect 22002 19972 22008 19984
rect 21784 19944 22008 19972
rect 21784 19932 21790 19944
rect 22002 19932 22008 19944
rect 22060 19932 22066 19984
rect 31386 19972 31392 19984
rect 22103 19944 31392 19972
rect 21821 19907 21879 19913
rect 21821 19904 21833 19907
rect 16264 19876 20024 19904
rect 20732 19876 21833 19904
rect 16264 19864 16270 19876
rect 12391 19808 12940 19836
rect 12391 19805 12403 19808
rect 12345 19799 12403 19805
rect 12986 19796 12992 19848
rect 13044 19836 13050 19848
rect 15197 19839 15255 19845
rect 15197 19836 15209 19839
rect 13044 19808 15209 19836
rect 13044 19796 13050 19808
rect 15197 19805 15209 19808
rect 15243 19836 15255 19839
rect 15930 19836 15936 19848
rect 15243 19808 15936 19836
rect 15243 19805 15255 19808
rect 15197 19799 15255 19805
rect 15930 19796 15936 19808
rect 15988 19796 15994 19848
rect 18233 19839 18291 19845
rect 18233 19805 18245 19839
rect 18279 19836 18291 19839
rect 19334 19836 19340 19848
rect 18279 19808 19340 19836
rect 18279 19805 18291 19808
rect 18233 19799 18291 19805
rect 19334 19796 19340 19808
rect 19392 19796 19398 19848
rect 19904 19845 19932 19876
rect 20732 19845 20760 19876
rect 19889 19839 19947 19845
rect 19889 19805 19901 19839
rect 19935 19805 19947 19839
rect 19889 19799 19947 19805
rect 20165 19839 20223 19845
rect 20165 19805 20177 19839
rect 20211 19805 20223 19839
rect 20165 19799 20223 19805
rect 20717 19839 20775 19845
rect 20717 19805 20729 19839
rect 20763 19805 20775 19839
rect 20717 19799 20775 19805
rect 10588 19771 10646 19777
rect 8220 19740 9536 19768
rect 9214 19700 9220 19712
rect 9175 19672 9220 19700
rect 9214 19660 9220 19672
rect 9272 19660 9278 19712
rect 9508 19700 9536 19740
rect 10588 19737 10600 19771
rect 10634 19768 10646 19771
rect 11514 19768 11520 19780
rect 10634 19740 11520 19768
rect 10634 19737 10646 19740
rect 10588 19731 10646 19737
rect 11514 19728 11520 19740
rect 11572 19728 11578 19780
rect 14366 19768 14372 19780
rect 14327 19740 14372 19768
rect 14366 19728 14372 19740
rect 14424 19728 14430 19780
rect 14550 19768 14556 19780
rect 14511 19740 14556 19768
rect 14550 19728 14556 19740
rect 14608 19728 14614 19780
rect 15470 19777 15476 19780
rect 15464 19768 15476 19777
rect 15431 19740 15476 19768
rect 15464 19731 15476 19740
rect 15470 19728 15476 19731
rect 15528 19728 15534 19780
rect 16850 19768 16856 19780
rect 16811 19740 16856 19768
rect 16850 19728 16856 19740
rect 16908 19728 16914 19780
rect 16942 19728 16948 19780
rect 17000 19768 17006 19780
rect 17313 19771 17371 19777
rect 17313 19768 17325 19771
rect 17000 19740 17325 19768
rect 17000 19728 17006 19740
rect 17313 19737 17325 19740
rect 17359 19768 17371 19771
rect 17359 19740 17448 19768
rect 17359 19737 17371 19740
rect 17313 19731 17371 19737
rect 10962 19700 10968 19712
rect 9508 19672 10968 19700
rect 10962 19660 10968 19672
rect 11020 19660 11026 19712
rect 15102 19660 15108 19712
rect 15160 19700 15166 19712
rect 16577 19703 16635 19709
rect 16577 19700 16589 19703
rect 15160 19672 16589 19700
rect 15160 19660 15166 19672
rect 16577 19669 16589 19672
rect 16623 19669 16635 19703
rect 17420 19700 17448 19740
rect 17494 19728 17500 19780
rect 17552 19768 17558 19780
rect 17770 19768 17776 19780
rect 17552 19740 17776 19768
rect 17552 19728 17558 19740
rect 17770 19728 17776 19740
rect 17828 19728 17834 19780
rect 18598 19768 18604 19780
rect 18559 19740 18604 19768
rect 18598 19728 18604 19740
rect 18656 19728 18662 19780
rect 20180 19768 20208 19799
rect 21082 19768 21088 19780
rect 20180 19740 21088 19768
rect 21082 19728 21088 19740
rect 21140 19728 21146 19780
rect 21468 19768 21496 19876
rect 21821 19873 21833 19876
rect 21867 19873 21879 19907
rect 21821 19867 21879 19873
rect 21634 19836 21640 19848
rect 21595 19808 21640 19836
rect 21634 19796 21640 19808
rect 21692 19796 21698 19848
rect 21726 19796 21732 19848
rect 21784 19836 21790 19848
rect 22103 19836 22131 19944
rect 31386 19932 31392 19944
rect 31444 19932 31450 19984
rect 31726 19972 31754 20012
rect 33870 20000 33876 20012
rect 33928 20000 33934 20052
rect 36538 19972 36544 19984
rect 31726 19944 36544 19972
rect 36538 19932 36544 19944
rect 36596 19932 36602 19984
rect 27706 19904 27712 19916
rect 27264 19876 27712 19904
rect 21784 19808 22131 19836
rect 22373 19839 22431 19845
rect 21784 19796 21790 19808
rect 22373 19805 22385 19839
rect 22419 19836 22431 19839
rect 26234 19836 26240 19848
rect 22419 19808 26240 19836
rect 22419 19805 22431 19808
rect 22373 19799 22431 19805
rect 26234 19796 26240 19808
rect 26292 19796 26298 19848
rect 27264 19845 27292 19876
rect 27706 19864 27712 19876
rect 27764 19864 27770 19916
rect 28534 19904 28540 19916
rect 28495 19876 28540 19904
rect 28534 19864 28540 19876
rect 28592 19864 28598 19916
rect 30190 19904 30196 19916
rect 30151 19876 30196 19904
rect 30190 19864 30196 19876
rect 30248 19864 30254 19916
rect 30650 19864 30656 19916
rect 30708 19904 30714 19916
rect 32306 19904 32312 19916
rect 30708 19876 32312 19904
rect 30708 19864 30714 19876
rect 32306 19864 32312 19876
rect 32364 19864 32370 19916
rect 46474 19904 46480 19916
rect 46435 19876 46480 19904
rect 46474 19864 46480 19876
rect 46532 19864 46538 19916
rect 27249 19839 27307 19845
rect 27249 19805 27261 19839
rect 27295 19805 27307 19839
rect 27249 19799 27307 19805
rect 27338 19796 27344 19848
rect 27396 19836 27402 19848
rect 28442 19836 28448 19848
rect 27396 19808 27441 19836
rect 28403 19808 28448 19836
rect 27396 19796 27402 19808
rect 28442 19796 28448 19808
rect 28500 19796 28506 19848
rect 28721 19839 28779 19845
rect 28721 19805 28733 19839
rect 28767 19836 28779 19839
rect 28810 19836 28816 19848
rect 28767 19808 28816 19836
rect 28767 19805 28779 19808
rect 28721 19799 28779 19805
rect 28810 19796 28816 19808
rect 28868 19796 28874 19848
rect 28994 19796 29000 19848
rect 29052 19836 29058 19848
rect 30101 19839 30159 19845
rect 30101 19836 30113 19839
rect 29052 19808 30113 19836
rect 29052 19796 29058 19808
rect 30101 19805 30113 19808
rect 30147 19805 30159 19839
rect 30101 19799 30159 19805
rect 30282 19796 30288 19848
rect 30340 19836 30346 19848
rect 30377 19839 30435 19845
rect 30377 19836 30389 19839
rect 30340 19808 30389 19836
rect 30340 19796 30346 19808
rect 30377 19805 30389 19808
rect 30423 19805 30435 19839
rect 30377 19799 30435 19805
rect 33226 19796 33232 19848
rect 33284 19836 33290 19848
rect 33781 19839 33839 19845
rect 33781 19836 33793 19839
rect 33284 19808 33793 19836
rect 33284 19796 33290 19808
rect 33781 19805 33793 19808
rect 33827 19805 33839 19839
rect 33781 19799 33839 19805
rect 46293 19839 46351 19845
rect 46293 19805 46305 19839
rect 46339 19805 46351 19839
rect 46293 19799 46351 19805
rect 21818 19768 21824 19780
rect 21468 19740 21824 19768
rect 21818 19728 21824 19740
rect 21876 19768 21882 19780
rect 21876 19740 23796 19768
rect 21876 19728 21882 19740
rect 19150 19700 19156 19712
rect 17420 19672 19156 19700
rect 16577 19663 16635 19669
rect 19150 19660 19156 19672
rect 19208 19660 19214 19712
rect 20073 19703 20131 19709
rect 20073 19669 20085 19703
rect 20119 19700 20131 19703
rect 20806 19700 20812 19712
rect 20119 19672 20812 19700
rect 20119 19669 20131 19672
rect 20073 19663 20131 19669
rect 20806 19660 20812 19672
rect 20864 19660 20870 19712
rect 20990 19660 20996 19712
rect 21048 19700 21054 19712
rect 22278 19700 22284 19712
rect 21048 19672 22284 19700
rect 21048 19660 21054 19672
rect 22278 19660 22284 19672
rect 22336 19700 22342 19712
rect 22465 19703 22523 19709
rect 22465 19700 22477 19703
rect 22336 19672 22477 19700
rect 22336 19660 22342 19672
rect 22465 19669 22477 19672
rect 22511 19669 22523 19703
rect 23768 19700 23796 19740
rect 23842 19728 23848 19780
rect 23900 19768 23906 19780
rect 31573 19771 31631 19777
rect 31573 19768 31585 19771
rect 23900 19740 31585 19768
rect 23900 19728 23906 19740
rect 31573 19737 31585 19740
rect 31619 19768 31631 19771
rect 32122 19768 32128 19780
rect 31619 19740 32128 19768
rect 31619 19737 31631 19740
rect 31573 19731 31631 19737
rect 32122 19728 32128 19740
rect 32180 19728 32186 19780
rect 46308 19768 46336 19799
rect 47670 19768 47676 19780
rect 46308 19740 47676 19768
rect 47670 19728 47676 19740
rect 47728 19728 47734 19780
rect 48130 19768 48136 19780
rect 48091 19740 48136 19768
rect 48130 19728 48136 19740
rect 48188 19728 48194 19780
rect 23934 19700 23940 19712
rect 23768 19672 23940 19700
rect 22465 19663 22523 19669
rect 23934 19660 23940 19672
rect 23992 19660 23998 19712
rect 26970 19660 26976 19712
rect 27028 19700 27034 19712
rect 27249 19703 27307 19709
rect 27249 19700 27261 19703
rect 27028 19672 27261 19700
rect 27028 19660 27034 19672
rect 27249 19669 27261 19672
rect 27295 19669 27307 19703
rect 27249 19663 27307 19669
rect 27798 19660 27804 19712
rect 27856 19700 27862 19712
rect 31754 19700 31760 19712
rect 27856 19672 31760 19700
rect 27856 19660 27862 19672
rect 31754 19660 31760 19672
rect 31812 19660 31818 19712
rect 32582 19660 32588 19712
rect 32640 19700 32646 19712
rect 32861 19703 32919 19709
rect 32861 19700 32873 19703
rect 32640 19672 32873 19700
rect 32640 19660 32646 19672
rect 32861 19669 32873 19672
rect 32907 19700 32919 19703
rect 35618 19700 35624 19712
rect 32907 19672 35624 19700
rect 32907 19669 32919 19672
rect 32861 19663 32919 19669
rect 35618 19660 35624 19672
rect 35676 19660 35682 19712
rect 1104 19610 48852 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 48852 19610
rect 1104 19536 48852 19558
rect 8754 19456 8760 19508
rect 8812 19496 8818 19508
rect 9401 19499 9459 19505
rect 9401 19496 9413 19499
rect 8812 19468 9413 19496
rect 8812 19456 8818 19468
rect 9401 19465 9413 19468
rect 9447 19465 9459 19499
rect 9401 19459 9459 19465
rect 4062 19388 4068 19440
rect 4120 19428 4126 19440
rect 8288 19431 8346 19437
rect 4120 19400 8156 19428
rect 4120 19388 4126 19400
rect 1762 19360 1768 19372
rect 1723 19332 1768 19360
rect 1762 19320 1768 19332
rect 1820 19320 1826 19372
rect 8018 19360 8024 19372
rect 7979 19332 8024 19360
rect 8018 19320 8024 19332
rect 8076 19320 8082 19372
rect 8128 19360 8156 19400
rect 8288 19397 8300 19431
rect 8334 19428 8346 19431
rect 9214 19428 9220 19440
rect 8334 19400 9220 19428
rect 8334 19397 8346 19400
rect 8288 19391 8346 19397
rect 9214 19388 9220 19400
rect 9272 19388 9278 19440
rect 9416 19428 9444 19459
rect 9674 19456 9680 19508
rect 9732 19496 9738 19508
rect 10229 19499 10287 19505
rect 10229 19496 10241 19499
rect 9732 19468 10241 19496
rect 9732 19456 9738 19468
rect 10229 19465 10241 19468
rect 10275 19465 10287 19499
rect 11514 19496 11520 19508
rect 11475 19468 11520 19496
rect 10229 19459 10287 19465
rect 11514 19456 11520 19468
rect 11572 19456 11578 19508
rect 14090 19456 14096 19508
rect 14148 19496 14154 19508
rect 14366 19496 14372 19508
rect 14148 19468 14372 19496
rect 14148 19456 14154 19468
rect 14366 19456 14372 19468
rect 14424 19496 14430 19508
rect 14424 19468 15516 19496
rect 14424 19456 14430 19468
rect 10045 19431 10103 19437
rect 10045 19428 10057 19431
rect 9416 19400 10057 19428
rect 10045 19397 10057 19400
rect 10091 19397 10103 19431
rect 10045 19391 10103 19397
rect 12713 19431 12771 19437
rect 12713 19397 12725 19431
rect 12759 19428 12771 19431
rect 14182 19428 14188 19440
rect 12759 19400 14188 19428
rect 12759 19397 12771 19400
rect 12713 19391 12771 19397
rect 14182 19388 14188 19400
rect 14240 19388 14246 19440
rect 14550 19388 14556 19440
rect 14608 19428 14614 19440
rect 15488 19428 15516 19468
rect 16850 19456 16856 19508
rect 16908 19496 16914 19508
rect 20990 19496 20996 19508
rect 16908 19468 20996 19496
rect 16908 19456 16914 19468
rect 16942 19428 16948 19440
rect 14608 19400 15424 19428
rect 15488 19400 16948 19428
rect 14608 19388 14614 19400
rect 9766 19360 9772 19372
rect 8128 19332 9772 19360
rect 9766 19320 9772 19332
rect 9824 19320 9830 19372
rect 9861 19363 9919 19369
rect 9861 19329 9873 19363
rect 9907 19360 9919 19363
rect 10502 19360 10508 19372
rect 9907 19332 10508 19360
rect 9907 19329 9919 19332
rect 9861 19323 9919 19329
rect 10502 19320 10508 19332
rect 10560 19320 10566 19372
rect 11790 19360 11796 19372
rect 11751 19332 11796 19360
rect 11790 19320 11796 19332
rect 11848 19320 11854 19372
rect 11885 19363 11943 19369
rect 11885 19329 11897 19363
rect 11931 19329 11943 19363
rect 11885 19323 11943 19329
rect 1946 19292 1952 19304
rect 1907 19264 1952 19292
rect 1946 19252 1952 19264
rect 2004 19252 2010 19304
rect 2222 19292 2228 19304
rect 2183 19264 2228 19292
rect 2222 19252 2228 19264
rect 2280 19252 2286 19304
rect 11900 19292 11928 19323
rect 11974 19320 11980 19372
rect 12032 19360 12038 19372
rect 12032 19332 12077 19360
rect 12032 19320 12038 19332
rect 12158 19320 12164 19372
rect 12216 19360 12222 19372
rect 13538 19360 13544 19372
rect 12216 19332 13544 19360
rect 12216 19320 12222 19332
rect 13538 19320 13544 19332
rect 13596 19320 13602 19372
rect 13633 19363 13691 19369
rect 13633 19329 13645 19363
rect 13679 19360 13691 19363
rect 14277 19363 14335 19369
rect 14277 19360 14289 19363
rect 13679 19332 14289 19360
rect 13679 19329 13691 19332
rect 13633 19323 13691 19329
rect 14277 19329 14289 19332
rect 14323 19360 14335 19363
rect 14366 19360 14372 19372
rect 14323 19332 14372 19360
rect 14323 19329 14335 19332
rect 14277 19323 14335 19329
rect 14366 19320 14372 19332
rect 14424 19320 14430 19372
rect 14461 19363 14519 19369
rect 14461 19329 14473 19363
rect 14507 19360 14519 19363
rect 15102 19360 15108 19372
rect 14507 19332 15108 19360
rect 14507 19329 14519 19332
rect 14461 19323 14519 19329
rect 15102 19320 15108 19332
rect 15160 19320 15166 19372
rect 15396 19304 15424 19400
rect 16942 19388 16948 19400
rect 17000 19388 17006 19440
rect 17236 19437 17264 19468
rect 20990 19456 20996 19468
rect 21048 19456 21054 19508
rect 21269 19499 21327 19505
rect 21269 19465 21281 19499
rect 21315 19496 21327 19499
rect 21910 19496 21916 19508
rect 21315 19468 21916 19496
rect 21315 19465 21327 19468
rect 21269 19459 21327 19465
rect 21910 19456 21916 19468
rect 21968 19456 21974 19508
rect 24762 19496 24768 19508
rect 24723 19468 24768 19496
rect 24762 19456 24768 19468
rect 24820 19456 24826 19508
rect 47762 19496 47768 19508
rect 24872 19468 47768 19496
rect 17221 19431 17279 19437
rect 17221 19397 17233 19431
rect 17267 19397 17279 19431
rect 17221 19391 17279 19397
rect 18785 19431 18843 19437
rect 18785 19397 18797 19431
rect 18831 19428 18843 19431
rect 19334 19428 19340 19440
rect 18831 19400 19340 19428
rect 18831 19397 18843 19400
rect 18785 19391 18843 19397
rect 19334 19388 19340 19400
rect 19392 19388 19398 19440
rect 20441 19431 20499 19437
rect 20441 19397 20453 19431
rect 20487 19428 20499 19431
rect 20806 19428 20812 19440
rect 20487 19400 20812 19428
rect 20487 19397 20499 19400
rect 20441 19391 20499 19397
rect 20806 19388 20812 19400
rect 20864 19388 20870 19440
rect 21726 19428 21732 19440
rect 21192 19400 21732 19428
rect 16482 19320 16488 19372
rect 16540 19360 16546 19372
rect 17494 19360 17500 19372
rect 16540 19332 17500 19360
rect 16540 19320 16546 19332
rect 17494 19320 17500 19332
rect 17552 19320 17558 19372
rect 18138 19320 18144 19372
rect 18196 19360 18202 19372
rect 19705 19363 19763 19369
rect 19705 19360 19717 19363
rect 18196 19332 19717 19360
rect 18196 19320 18202 19332
rect 19705 19329 19717 19332
rect 19751 19329 19763 19363
rect 19705 19323 19763 19329
rect 20341 19363 20399 19369
rect 20341 19329 20353 19363
rect 20387 19329 20399 19363
rect 21082 19360 21088 19372
rect 21043 19332 21088 19360
rect 20341 19323 20399 19329
rect 12250 19292 12256 19304
rect 11900 19264 12256 19292
rect 12250 19252 12256 19264
rect 12308 19292 12314 19304
rect 12897 19295 12955 19301
rect 12897 19292 12909 19295
rect 12308 19264 12909 19292
rect 12308 19252 12314 19264
rect 12897 19261 12909 19264
rect 12943 19261 12955 19295
rect 12897 19255 12955 19261
rect 13814 19252 13820 19304
rect 13872 19292 13878 19304
rect 14645 19295 14703 19301
rect 13872 19264 13917 19292
rect 13872 19252 13878 19264
rect 14645 19261 14657 19295
rect 14691 19292 14703 19295
rect 15286 19292 15292 19304
rect 14691 19264 15292 19292
rect 14691 19261 14703 19264
rect 14645 19255 14703 19261
rect 15286 19252 15292 19264
rect 15344 19252 15350 19304
rect 15378 19252 15384 19304
rect 15436 19292 15442 19304
rect 15436 19264 15481 19292
rect 15436 19252 15442 19264
rect 19334 19252 19340 19304
rect 19392 19292 19398 19304
rect 20364 19292 20392 19323
rect 21082 19320 21088 19332
rect 21140 19320 21146 19372
rect 21192 19360 21220 19400
rect 21726 19388 21732 19400
rect 21784 19388 21790 19440
rect 22186 19388 22192 19440
rect 22244 19428 22250 19440
rect 24872 19428 24900 19468
rect 47762 19456 47768 19468
rect 47820 19456 47826 19508
rect 25869 19431 25927 19437
rect 25869 19428 25881 19431
rect 22244 19400 24900 19428
rect 25148 19400 25881 19428
rect 22244 19388 22250 19400
rect 21269 19363 21327 19369
rect 21269 19360 21281 19363
rect 21192 19332 21281 19360
rect 21192 19292 21220 19332
rect 21269 19329 21281 19332
rect 21315 19329 21327 19363
rect 21818 19360 21824 19372
rect 21779 19332 21824 19360
rect 21269 19323 21327 19329
rect 21818 19320 21824 19332
rect 21876 19320 21882 19372
rect 22002 19320 22008 19372
rect 22060 19360 22066 19372
rect 22060 19332 22416 19360
rect 22060 19320 22066 19332
rect 19392 19264 21220 19292
rect 22388 19292 22416 19332
rect 22462 19320 22468 19372
rect 22520 19360 22526 19372
rect 22833 19363 22891 19369
rect 22833 19360 22845 19363
rect 22520 19332 22845 19360
rect 22520 19320 22526 19332
rect 22833 19329 22845 19332
rect 22879 19329 22891 19363
rect 22833 19323 22891 19329
rect 22922 19320 22928 19372
rect 22980 19360 22986 19372
rect 23089 19363 23147 19369
rect 23089 19360 23101 19363
rect 22980 19332 23101 19360
rect 22980 19320 22986 19332
rect 23089 19329 23101 19332
rect 23135 19329 23147 19363
rect 23089 19323 23147 19329
rect 24673 19363 24731 19369
rect 24673 19329 24685 19363
rect 24719 19360 24731 19363
rect 25038 19360 25044 19372
rect 24719 19332 25044 19360
rect 24719 19329 24731 19332
rect 24673 19323 24731 19329
rect 25038 19320 25044 19332
rect 25096 19320 25102 19372
rect 25148 19292 25176 19400
rect 25869 19397 25881 19400
rect 25915 19397 25927 19431
rect 26970 19428 26976 19440
rect 26931 19400 26976 19428
rect 25869 19391 25927 19397
rect 26970 19388 26976 19400
rect 27028 19388 27034 19440
rect 27154 19428 27160 19440
rect 27115 19400 27160 19428
rect 27154 19388 27160 19400
rect 27212 19388 27218 19440
rect 28442 19388 28448 19440
rect 28500 19428 28506 19440
rect 28902 19428 28908 19440
rect 28500 19400 28908 19428
rect 28500 19388 28506 19400
rect 28902 19388 28908 19400
rect 28960 19388 28966 19440
rect 33134 19428 33140 19440
rect 32324 19400 33140 19428
rect 25685 19363 25743 19369
rect 25685 19329 25697 19363
rect 25731 19360 25743 19363
rect 26988 19360 27016 19388
rect 32122 19360 32128 19372
rect 25731 19332 27016 19360
rect 32083 19332 32128 19360
rect 25731 19329 25743 19332
rect 25685 19323 25743 19329
rect 32122 19320 32128 19332
rect 32180 19320 32186 19372
rect 22388 19264 22876 19292
rect 19392 19252 19398 19264
rect 16114 19184 16120 19236
rect 16172 19224 16178 19236
rect 19061 19227 19119 19233
rect 19061 19224 19073 19227
rect 16172 19196 19073 19224
rect 16172 19184 16178 19196
rect 19061 19193 19073 19196
rect 19107 19224 19119 19227
rect 22186 19224 22192 19236
rect 19107 19196 22192 19224
rect 19107 19193 19119 19196
rect 19061 19187 19119 19193
rect 22186 19184 22192 19196
rect 22244 19184 22250 19236
rect 13538 19116 13544 19168
rect 13596 19156 13602 19168
rect 17310 19156 17316 19168
rect 13596 19128 17316 19156
rect 13596 19116 13602 19128
rect 17310 19116 17316 19128
rect 17368 19156 17374 19168
rect 17494 19156 17500 19168
rect 17368 19128 17500 19156
rect 17368 19116 17374 19128
rect 17494 19116 17500 19128
rect 17552 19116 17558 19168
rect 19426 19116 19432 19168
rect 19484 19156 19490 19168
rect 19794 19156 19800 19168
rect 19484 19128 19800 19156
rect 19484 19116 19490 19128
rect 19794 19116 19800 19128
rect 19852 19116 19858 19168
rect 22002 19156 22008 19168
rect 21963 19128 22008 19156
rect 22002 19116 22008 19128
rect 22060 19116 22066 19168
rect 22848 19156 22876 19264
rect 23860 19264 25176 19292
rect 25501 19295 25559 19301
rect 23106 19156 23112 19168
rect 22848 19128 23112 19156
rect 23106 19116 23112 19128
rect 23164 19116 23170 19168
rect 23566 19116 23572 19168
rect 23624 19156 23630 19168
rect 23860 19156 23888 19264
rect 25501 19261 25513 19295
rect 25547 19292 25559 19295
rect 26234 19292 26240 19304
rect 25547 19264 26240 19292
rect 25547 19261 25559 19264
rect 25501 19255 25559 19261
rect 26234 19252 26240 19264
rect 26292 19292 26298 19304
rect 27062 19292 27068 19304
rect 26292 19264 27068 19292
rect 26292 19252 26298 19264
rect 27062 19252 27068 19264
rect 27120 19252 27126 19304
rect 27341 19227 27399 19233
rect 27341 19193 27353 19227
rect 27387 19224 27399 19227
rect 27614 19224 27620 19236
rect 27387 19196 27620 19224
rect 27387 19193 27399 19196
rect 27341 19187 27399 19193
rect 27614 19184 27620 19196
rect 27672 19184 27678 19236
rect 32324 19233 32352 19400
rect 33134 19388 33140 19400
rect 33192 19388 33198 19440
rect 33318 19428 33324 19440
rect 33279 19400 33324 19428
rect 33318 19388 33324 19400
rect 33376 19388 33382 19440
rect 36449 19363 36507 19369
rect 36449 19329 36461 19363
rect 36495 19360 36507 19363
rect 36630 19360 36636 19372
rect 36495 19332 36636 19360
rect 36495 19329 36507 19332
rect 36449 19323 36507 19329
rect 36630 19320 36636 19332
rect 36688 19360 36694 19372
rect 37277 19363 37335 19369
rect 37277 19360 37289 19363
rect 36688 19332 37289 19360
rect 36688 19320 36694 19332
rect 37277 19329 37289 19332
rect 37323 19329 37335 19363
rect 47854 19360 47860 19372
rect 47815 19332 47860 19360
rect 37277 19323 37335 19329
rect 47854 19320 47860 19332
rect 47912 19320 47918 19372
rect 33137 19295 33195 19301
rect 33137 19261 33149 19295
rect 33183 19292 33195 19295
rect 33594 19292 33600 19304
rect 33183 19264 33600 19292
rect 33183 19261 33195 19264
rect 33137 19255 33195 19261
rect 33594 19252 33600 19264
rect 33652 19252 33658 19304
rect 34146 19292 34152 19304
rect 34107 19264 34152 19292
rect 34146 19252 34152 19264
rect 34204 19252 34210 19304
rect 32309 19227 32367 19233
rect 32309 19193 32321 19227
rect 32355 19193 32367 19227
rect 32309 19187 32367 19193
rect 23624 19128 23888 19156
rect 24213 19159 24271 19165
rect 23624 19116 23630 19128
rect 24213 19125 24225 19159
rect 24259 19156 24271 19159
rect 24578 19156 24584 19168
rect 24259 19128 24584 19156
rect 24259 19125 24271 19128
rect 24213 19119 24271 19125
rect 24578 19116 24584 19128
rect 24636 19116 24642 19168
rect 36538 19156 36544 19168
rect 36499 19128 36544 19156
rect 36538 19116 36544 19128
rect 36596 19116 36602 19168
rect 37369 19159 37427 19165
rect 37369 19125 37381 19159
rect 37415 19156 37427 19159
rect 37458 19156 37464 19168
rect 37415 19128 37464 19156
rect 37415 19125 37427 19128
rect 37369 19119 37427 19125
rect 37458 19116 37464 19128
rect 37516 19116 37522 19168
rect 48038 19156 48044 19168
rect 47999 19128 48044 19156
rect 48038 19116 48044 19128
rect 48096 19116 48102 19168
rect 1104 19066 48852 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 48852 19066
rect 1104 18992 48852 19014
rect 1946 18912 1952 18964
rect 2004 18952 2010 18964
rect 2225 18955 2283 18961
rect 2225 18952 2237 18955
rect 2004 18924 2237 18952
rect 2004 18912 2010 18924
rect 2225 18921 2237 18924
rect 2271 18921 2283 18955
rect 2225 18915 2283 18921
rect 2746 18924 19932 18952
rect 2038 18844 2044 18896
rect 2096 18884 2102 18896
rect 2746 18884 2774 18924
rect 2096 18856 2774 18884
rect 11624 18856 16804 18884
rect 2096 18844 2102 18856
rect 9582 18816 9588 18828
rect 9416 18788 9588 18816
rect 2133 18751 2191 18757
rect 2133 18717 2145 18751
rect 2179 18748 2191 18751
rect 2406 18748 2412 18760
rect 2179 18720 2412 18748
rect 2179 18717 2191 18720
rect 2133 18711 2191 18717
rect 2406 18708 2412 18720
rect 2464 18748 2470 18760
rect 4982 18748 4988 18760
rect 2464 18720 4988 18748
rect 2464 18708 2470 18720
rect 4982 18708 4988 18720
rect 5040 18708 5046 18760
rect 9306 18748 9312 18760
rect 9267 18720 9312 18748
rect 9306 18708 9312 18720
rect 9364 18708 9370 18760
rect 9416 18757 9444 18788
rect 9582 18776 9588 18788
rect 9640 18816 9646 18828
rect 9640 18788 11560 18816
rect 9640 18776 9646 18788
rect 9401 18751 9459 18757
rect 9401 18717 9413 18751
rect 9447 18717 9459 18751
rect 9401 18711 9459 18717
rect 9490 18708 9496 18760
rect 9548 18748 9554 18760
rect 9677 18751 9735 18757
rect 9548 18720 9593 18748
rect 9548 18708 9554 18720
rect 9677 18717 9689 18751
rect 9723 18748 9735 18751
rect 10226 18748 10232 18760
rect 9723 18720 10232 18748
rect 9723 18717 9735 18720
rect 9677 18711 9735 18717
rect 10226 18708 10232 18720
rect 10284 18708 10290 18760
rect 3970 18640 3976 18692
rect 4028 18680 4034 18692
rect 11532 18680 11560 18788
rect 11624 18757 11652 18856
rect 12802 18776 12808 18828
rect 12860 18816 12866 18828
rect 14461 18819 14519 18825
rect 14461 18816 14473 18819
rect 12860 18788 13308 18816
rect 12860 18776 12866 18788
rect 11609 18751 11667 18757
rect 11609 18717 11621 18751
rect 11655 18717 11667 18751
rect 11609 18711 11667 18717
rect 11698 18751 11756 18757
rect 11698 18717 11710 18751
rect 11744 18717 11756 18751
rect 11698 18711 11756 18717
rect 11793 18751 11851 18757
rect 11793 18717 11805 18751
rect 11839 18748 11851 18751
rect 11882 18748 11888 18760
rect 11839 18720 11888 18748
rect 11839 18717 11851 18720
rect 11793 18711 11851 18717
rect 11716 18680 11744 18711
rect 11882 18708 11888 18720
rect 11940 18708 11946 18760
rect 11977 18751 12035 18757
rect 11977 18717 11989 18751
rect 12023 18748 12035 18751
rect 12158 18748 12164 18760
rect 12023 18720 12164 18748
rect 12023 18717 12035 18720
rect 11977 18711 12035 18717
rect 12158 18708 12164 18720
rect 12216 18708 12222 18760
rect 13280 18757 13308 18788
rect 13372 18788 14473 18816
rect 13372 18757 13400 18788
rect 14461 18785 14473 18788
rect 14507 18785 14519 18819
rect 14461 18779 14519 18785
rect 13173 18751 13231 18757
rect 13173 18748 13185 18751
rect 12360 18720 13185 18748
rect 12250 18680 12256 18692
rect 4028 18652 11468 18680
rect 11532 18652 12256 18680
rect 4028 18640 4034 18652
rect 9030 18612 9036 18624
rect 8991 18584 9036 18612
rect 9030 18572 9036 18584
rect 9088 18572 9094 18624
rect 11330 18612 11336 18624
rect 11291 18584 11336 18612
rect 11330 18572 11336 18584
rect 11388 18572 11394 18624
rect 11440 18612 11468 18652
rect 12250 18640 12256 18652
rect 12308 18640 12314 18692
rect 12360 18612 12388 18720
rect 13173 18717 13185 18720
rect 13219 18717 13231 18751
rect 13173 18711 13231 18717
rect 13262 18751 13320 18757
rect 13262 18717 13274 18751
rect 13308 18717 13320 18751
rect 13262 18711 13320 18717
rect 13362 18751 13420 18757
rect 13362 18717 13374 18751
rect 13408 18717 13420 18751
rect 13538 18748 13544 18760
rect 13499 18720 13544 18748
rect 13362 18711 13420 18717
rect 13538 18708 13544 18720
rect 13596 18708 13602 18760
rect 13814 18708 13820 18760
rect 13872 18748 13878 18760
rect 14277 18751 14335 18757
rect 14277 18748 14289 18751
rect 13872 18720 14289 18748
rect 13872 18708 13878 18720
rect 14277 18717 14289 18720
rect 14323 18748 14335 18751
rect 14734 18748 14740 18760
rect 14323 18720 14740 18748
rect 14323 18717 14335 18720
rect 14277 18711 14335 18717
rect 14734 18708 14740 18720
rect 14792 18708 14798 18760
rect 16114 18748 16120 18760
rect 16075 18720 16120 18748
rect 16114 18708 16120 18720
rect 16172 18708 16178 18760
rect 14090 18680 14096 18692
rect 14051 18652 14096 18680
rect 14090 18640 14096 18652
rect 14148 18640 14154 18692
rect 12894 18612 12900 18624
rect 11440 18584 12388 18612
rect 12855 18584 12900 18612
rect 12894 18572 12900 18584
rect 12952 18572 12958 18624
rect 15746 18572 15752 18624
rect 15804 18612 15810 18624
rect 16209 18615 16267 18621
rect 16209 18612 16221 18615
rect 15804 18584 16221 18612
rect 15804 18572 15810 18584
rect 16209 18581 16221 18584
rect 16255 18581 16267 18615
rect 16776 18612 16804 18856
rect 17129 18751 17187 18757
rect 17129 18717 17141 18751
rect 17175 18748 17187 18751
rect 19794 18748 19800 18760
rect 17175 18720 19800 18748
rect 17175 18717 17187 18720
rect 17129 18711 17187 18717
rect 19794 18708 19800 18720
rect 19852 18708 19858 18760
rect 19904 18757 19932 18924
rect 20806 18912 20812 18964
rect 20864 18952 20870 18964
rect 21726 18952 21732 18964
rect 20864 18924 21732 18952
rect 20864 18912 20870 18924
rect 21726 18912 21732 18924
rect 21784 18912 21790 18964
rect 22373 18955 22431 18961
rect 22373 18921 22385 18955
rect 22419 18952 22431 18955
rect 22922 18952 22928 18964
rect 22419 18924 22928 18952
rect 22419 18921 22431 18924
rect 22373 18915 22431 18921
rect 22922 18912 22928 18924
rect 22980 18912 22986 18964
rect 33321 18955 33379 18961
rect 33321 18921 33333 18955
rect 33367 18952 33379 18955
rect 33410 18952 33416 18964
rect 33367 18924 33416 18952
rect 33367 18921 33379 18924
rect 33321 18915 33379 18921
rect 33410 18912 33416 18924
rect 33468 18912 33474 18964
rect 47670 18952 47676 18964
rect 47631 18924 47676 18952
rect 47670 18912 47676 18924
rect 47728 18912 47734 18964
rect 19978 18844 19984 18896
rect 20036 18884 20042 18896
rect 20622 18884 20628 18896
rect 20036 18856 20628 18884
rect 20036 18844 20042 18856
rect 20622 18844 20628 18856
rect 20680 18844 20686 18896
rect 23845 18887 23903 18893
rect 23845 18884 23857 18887
rect 22848 18856 23857 18884
rect 21085 18819 21143 18825
rect 21085 18816 21097 18819
rect 20088 18788 21097 18816
rect 20088 18757 20116 18788
rect 21085 18785 21097 18788
rect 21131 18785 21143 18819
rect 22370 18816 22376 18828
rect 21085 18779 21143 18785
rect 21560 18788 22376 18816
rect 19889 18751 19947 18757
rect 19889 18717 19901 18751
rect 19935 18717 19947 18751
rect 19889 18711 19947 18717
rect 19981 18751 20039 18757
rect 19981 18717 19993 18751
rect 20027 18717 20039 18751
rect 19981 18711 20039 18717
rect 20073 18751 20131 18757
rect 20073 18717 20085 18751
rect 20119 18717 20131 18751
rect 20073 18711 20131 18717
rect 20257 18751 20315 18757
rect 20257 18717 20269 18751
rect 20303 18748 20315 18751
rect 20346 18748 20352 18760
rect 20303 18720 20352 18748
rect 20303 18717 20315 18720
rect 20257 18711 20315 18717
rect 16850 18640 16856 18692
rect 16908 18680 16914 18692
rect 17374 18683 17432 18689
rect 17374 18680 17386 18683
rect 16908 18652 17386 18680
rect 16908 18640 16914 18652
rect 17374 18649 17386 18652
rect 17420 18649 17432 18683
rect 19996 18680 20024 18711
rect 20346 18708 20352 18720
rect 20404 18708 20410 18760
rect 20990 18748 20996 18760
rect 20456 18720 20996 18748
rect 20456 18680 20484 18720
rect 20990 18708 20996 18720
rect 21048 18748 21054 18760
rect 21560 18757 21588 18788
rect 22370 18776 22376 18788
rect 22428 18776 22434 18828
rect 21545 18751 21603 18757
rect 21545 18748 21557 18751
rect 21048 18720 21557 18748
rect 21048 18708 21054 18720
rect 21545 18717 21557 18720
rect 21591 18717 21603 18751
rect 21726 18748 21732 18760
rect 21687 18720 21732 18748
rect 21545 18711 21603 18717
rect 21726 18708 21732 18720
rect 21784 18708 21790 18760
rect 22554 18748 22560 18760
rect 22515 18720 22560 18748
rect 22554 18708 22560 18720
rect 22612 18708 22618 18760
rect 22848 18757 22876 18856
rect 23845 18853 23857 18856
rect 23891 18853 23903 18887
rect 24397 18887 24455 18893
rect 24397 18884 24409 18887
rect 23845 18847 23903 18853
rect 23952 18856 24409 18884
rect 23569 18819 23627 18825
rect 23569 18785 23581 18819
rect 23615 18816 23627 18819
rect 23952 18816 23980 18856
rect 24397 18853 24409 18856
rect 24443 18853 24455 18887
rect 24397 18847 24455 18853
rect 25038 18816 25044 18828
rect 23615 18788 23980 18816
rect 24951 18788 25044 18816
rect 23615 18785 23627 18788
rect 23569 18779 23627 18785
rect 25038 18776 25044 18788
rect 25096 18816 25102 18828
rect 25096 18788 26004 18816
rect 25096 18776 25102 18788
rect 22833 18751 22891 18757
rect 22833 18717 22845 18751
rect 22879 18717 22891 18751
rect 22833 18711 22891 18717
rect 23477 18751 23535 18757
rect 23477 18717 23489 18751
rect 23523 18748 23535 18751
rect 24026 18748 24032 18760
rect 23523 18720 24032 18748
rect 23523 18717 23535 18720
rect 23477 18711 23535 18717
rect 24026 18708 24032 18720
rect 24084 18708 24090 18760
rect 25593 18751 25651 18757
rect 25593 18748 25605 18751
rect 24504 18720 25605 18748
rect 19996 18652 20484 18680
rect 20717 18683 20775 18689
rect 17374 18643 17432 18649
rect 20717 18649 20729 18683
rect 20763 18649 20775 18683
rect 20717 18643 20775 18649
rect 20901 18683 20959 18689
rect 20901 18649 20913 18683
rect 20947 18680 20959 18683
rect 21082 18680 21088 18692
rect 20947 18652 21088 18680
rect 20947 18649 20959 18652
rect 20901 18643 20959 18649
rect 18509 18615 18567 18621
rect 18509 18612 18521 18615
rect 16776 18584 18521 18612
rect 16209 18575 16267 18581
rect 18509 18581 18521 18584
rect 18555 18612 18567 18615
rect 19334 18612 19340 18624
rect 18555 18584 19340 18612
rect 18555 18581 18567 18584
rect 18509 18575 18567 18581
rect 19334 18572 19340 18584
rect 19392 18572 19398 18624
rect 19613 18615 19671 18621
rect 19613 18581 19625 18615
rect 19659 18612 19671 18615
rect 20162 18612 20168 18624
rect 19659 18584 20168 18612
rect 19659 18581 19671 18584
rect 19613 18575 19671 18581
rect 20162 18572 20168 18584
rect 20220 18572 20226 18624
rect 20732 18612 20760 18643
rect 21082 18640 21088 18652
rect 21140 18640 21146 18692
rect 23934 18640 23940 18692
rect 23992 18680 23998 18692
rect 24504 18680 24532 18720
rect 25593 18717 25605 18720
rect 25639 18717 25651 18751
rect 25593 18711 25651 18717
rect 25869 18751 25927 18757
rect 25869 18717 25881 18751
rect 25915 18717 25927 18751
rect 25976 18748 26004 18788
rect 34698 18776 34704 18828
rect 34756 18776 34762 18828
rect 36538 18816 36544 18828
rect 36499 18788 36544 18816
rect 36538 18776 36544 18788
rect 36596 18776 36602 18828
rect 26326 18748 26332 18760
rect 25976 18720 26332 18748
rect 25869 18711 25927 18717
rect 23992 18652 24532 18680
rect 23992 18640 23998 18652
rect 24578 18640 24584 18692
rect 24636 18680 24642 18692
rect 24857 18683 24915 18689
rect 24857 18680 24869 18683
rect 24636 18652 24869 18680
rect 24636 18640 24642 18652
rect 24857 18649 24869 18652
rect 24903 18649 24915 18683
rect 25884 18680 25912 18711
rect 26326 18708 26332 18720
rect 26384 18708 26390 18760
rect 26786 18748 26792 18760
rect 26747 18720 26792 18748
rect 26786 18708 26792 18720
rect 26844 18708 26850 18760
rect 26970 18708 26976 18760
rect 27028 18748 27034 18760
rect 27433 18751 27491 18757
rect 27433 18748 27445 18751
rect 27028 18720 27445 18748
rect 27028 18708 27034 18720
rect 27433 18717 27445 18720
rect 27479 18717 27491 18751
rect 27433 18711 27491 18717
rect 27522 18708 27528 18760
rect 27580 18748 27586 18760
rect 27617 18751 27675 18757
rect 27617 18748 27629 18751
rect 27580 18720 27629 18748
rect 27580 18708 27586 18720
rect 27617 18717 27629 18720
rect 27663 18717 27675 18751
rect 27617 18711 27675 18717
rect 28166 18708 28172 18760
rect 28224 18748 28230 18760
rect 29733 18751 29791 18757
rect 29733 18748 29745 18751
rect 28224 18720 29745 18748
rect 28224 18708 28230 18720
rect 29733 18717 29745 18720
rect 29779 18717 29791 18751
rect 31941 18751 31999 18757
rect 31941 18748 31953 18751
rect 29733 18711 29791 18717
rect 31726 18720 31953 18748
rect 26988 18680 27016 18708
rect 25884 18652 27016 18680
rect 27801 18683 27859 18689
rect 24857 18643 24915 18649
rect 27801 18649 27813 18683
rect 27847 18680 27859 18683
rect 27890 18680 27896 18692
rect 27847 18652 27896 18680
rect 27847 18649 27859 18652
rect 27801 18643 27859 18649
rect 27890 18640 27896 18652
rect 27948 18680 27954 18692
rect 28718 18680 28724 18692
rect 27948 18652 28724 18680
rect 27948 18640 27954 18652
rect 28718 18640 28724 18652
rect 28776 18640 28782 18692
rect 29638 18640 29644 18692
rect 29696 18680 29702 18692
rect 31726 18680 31754 18720
rect 31941 18717 31953 18720
rect 31987 18748 31999 18751
rect 34716 18748 34744 18776
rect 31987 18720 34744 18748
rect 34885 18751 34943 18757
rect 31987 18717 31999 18720
rect 31941 18711 31999 18717
rect 34885 18717 34897 18751
rect 34931 18748 34943 18751
rect 35618 18748 35624 18760
rect 34931 18720 35624 18748
rect 34931 18717 34943 18720
rect 34885 18711 34943 18717
rect 35618 18708 35624 18720
rect 35676 18748 35682 18760
rect 36357 18751 36415 18757
rect 36357 18748 36369 18751
rect 35676 18720 36369 18748
rect 35676 18708 35682 18720
rect 36357 18717 36369 18720
rect 36403 18717 36415 18751
rect 36357 18711 36415 18717
rect 32214 18689 32220 18692
rect 29696 18652 31754 18680
rect 29696 18640 29702 18652
rect 32208 18643 32220 18689
rect 32272 18680 32278 18692
rect 32272 18652 32308 18680
rect 32214 18640 32220 18643
rect 32272 18640 32278 18652
rect 33134 18640 33140 18692
rect 33192 18680 33198 18692
rect 34701 18683 34759 18689
rect 34701 18680 34713 18683
rect 33192 18652 34713 18680
rect 33192 18640 33198 18652
rect 34701 18649 34713 18652
rect 34747 18680 34759 18683
rect 36078 18680 36084 18692
rect 34747 18652 36084 18680
rect 34747 18649 34759 18652
rect 34701 18643 34759 18649
rect 36078 18640 36084 18652
rect 36136 18640 36142 18692
rect 38197 18683 38255 18689
rect 38197 18649 38209 18683
rect 38243 18680 38255 18683
rect 46382 18680 46388 18692
rect 38243 18652 46388 18680
rect 38243 18649 38255 18652
rect 38197 18643 38255 18649
rect 46382 18640 46388 18652
rect 46440 18640 46446 18692
rect 20806 18612 20812 18624
rect 20719 18584 20812 18612
rect 20806 18572 20812 18584
rect 20864 18612 20870 18624
rect 21266 18612 21272 18624
rect 20864 18584 21272 18612
rect 20864 18572 20870 18584
rect 21266 18572 21272 18584
rect 21324 18572 21330 18624
rect 21634 18612 21640 18624
rect 21595 18584 21640 18612
rect 21634 18572 21640 18584
rect 21692 18572 21698 18624
rect 22741 18615 22799 18621
rect 22741 18581 22753 18615
rect 22787 18612 22799 18615
rect 22922 18612 22928 18624
rect 22787 18584 22928 18612
rect 22787 18581 22799 18584
rect 22741 18575 22799 18581
rect 22922 18572 22928 18584
rect 22980 18572 22986 18624
rect 23658 18572 23664 18624
rect 23716 18612 23722 18624
rect 23842 18612 23848 18624
rect 23716 18584 23848 18612
rect 23716 18572 23722 18584
rect 23842 18572 23848 18584
rect 23900 18612 23906 18624
rect 24765 18615 24823 18621
rect 24765 18612 24777 18615
rect 23900 18584 24777 18612
rect 23900 18572 23906 18584
rect 24765 18581 24777 18584
rect 24811 18581 24823 18615
rect 24765 18575 24823 18581
rect 24946 18572 24952 18624
rect 25004 18612 25010 18624
rect 25685 18615 25743 18621
rect 25685 18612 25697 18615
rect 25004 18584 25697 18612
rect 25004 18572 25010 18584
rect 25685 18581 25697 18584
rect 25731 18581 25743 18615
rect 25685 18575 25743 18581
rect 26881 18615 26939 18621
rect 26881 18581 26893 18615
rect 26927 18612 26939 18615
rect 27430 18612 27436 18624
rect 26927 18584 27436 18612
rect 26927 18581 26939 18584
rect 26881 18575 26939 18581
rect 27430 18572 27436 18584
rect 27488 18572 27494 18624
rect 29546 18612 29552 18624
rect 29507 18584 29552 18612
rect 29546 18572 29552 18584
rect 29604 18572 29610 18624
rect 34514 18572 34520 18624
rect 34572 18612 34578 18624
rect 35069 18615 35127 18621
rect 35069 18612 35081 18615
rect 34572 18584 35081 18612
rect 34572 18572 34578 18584
rect 35069 18581 35081 18584
rect 35115 18581 35127 18615
rect 35069 18575 35127 18581
rect 1104 18522 48852 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 48852 18522
rect 1104 18448 48852 18470
rect 9490 18368 9496 18420
rect 9548 18408 9554 18420
rect 10873 18411 10931 18417
rect 10873 18408 10885 18411
rect 9548 18380 10885 18408
rect 9548 18368 9554 18380
rect 10873 18377 10885 18380
rect 10919 18377 10931 18411
rect 11882 18408 11888 18420
rect 11843 18380 11888 18408
rect 10873 18371 10931 18377
rect 11882 18368 11888 18380
rect 11940 18368 11946 18420
rect 14366 18408 14372 18420
rect 14327 18380 14372 18408
rect 14366 18368 14372 18380
rect 14424 18368 14430 18420
rect 15930 18408 15936 18420
rect 15891 18380 15936 18408
rect 15930 18368 15936 18380
rect 15988 18368 15994 18420
rect 16850 18408 16856 18420
rect 16811 18380 16856 18408
rect 16850 18368 16856 18380
rect 16908 18368 16914 18420
rect 17218 18368 17224 18420
rect 17276 18368 17282 18420
rect 22554 18368 22560 18420
rect 22612 18408 22618 18420
rect 24121 18411 24179 18417
rect 24121 18408 24133 18411
rect 22612 18380 24133 18408
rect 22612 18368 22618 18380
rect 24121 18377 24133 18380
rect 24167 18377 24179 18411
rect 26050 18408 26056 18420
rect 26011 18380 26056 18408
rect 24121 18371 24179 18377
rect 26050 18368 26056 18380
rect 26108 18368 26114 18420
rect 26234 18368 26240 18420
rect 26292 18408 26298 18420
rect 27249 18411 27307 18417
rect 27249 18408 27261 18411
rect 26292 18380 27261 18408
rect 26292 18368 26298 18380
rect 27249 18377 27261 18380
rect 27295 18377 27307 18411
rect 28166 18408 28172 18420
rect 28127 18380 28172 18408
rect 27249 18371 27307 18377
rect 28166 18368 28172 18380
rect 28224 18368 28230 18420
rect 32125 18411 32183 18417
rect 28276 18380 32076 18408
rect 8018 18340 8024 18352
rect 7484 18312 8024 18340
rect 7484 18284 7512 18312
rect 8018 18300 8024 18312
rect 8076 18300 8082 18352
rect 10134 18340 10140 18352
rect 9692 18312 10140 18340
rect 2041 18275 2099 18281
rect 2041 18241 2053 18275
rect 2087 18272 2099 18275
rect 2130 18272 2136 18284
rect 2087 18244 2136 18272
rect 2087 18241 2099 18244
rect 2041 18235 2099 18241
rect 2130 18232 2136 18244
rect 2188 18232 2194 18284
rect 6822 18272 6828 18284
rect 6783 18244 6828 18272
rect 6822 18232 6828 18244
rect 6880 18232 6886 18284
rect 7466 18272 7472 18284
rect 7379 18244 7472 18272
rect 7466 18232 7472 18244
rect 7524 18232 7530 18284
rect 7736 18275 7794 18281
rect 7736 18241 7748 18275
rect 7782 18272 7794 18275
rect 9030 18272 9036 18284
rect 7782 18244 9036 18272
rect 7782 18241 7794 18244
rect 7736 18235 7794 18241
rect 9030 18232 9036 18244
rect 9088 18232 9094 18284
rect 9692 18281 9720 18312
rect 10134 18300 10140 18312
rect 10192 18300 10198 18352
rect 11517 18343 11575 18349
rect 11517 18340 11529 18343
rect 10520 18312 11529 18340
rect 10520 18284 10548 18312
rect 11517 18309 11529 18312
rect 11563 18309 11575 18343
rect 11517 18303 11575 18309
rect 12894 18300 12900 18352
rect 12952 18340 12958 18352
rect 13234 18343 13292 18349
rect 13234 18340 13246 18343
rect 12952 18312 13246 18340
rect 12952 18300 12958 18312
rect 13234 18309 13246 18312
rect 13280 18309 13292 18343
rect 17236 18340 17264 18368
rect 21634 18340 21640 18352
rect 13234 18303 13292 18309
rect 17233 18312 17264 18340
rect 17328 18312 21640 18340
rect 17233 18284 17261 18312
rect 17328 18284 17356 18312
rect 21634 18300 21640 18312
rect 21692 18300 21698 18352
rect 22186 18300 22192 18352
rect 22244 18340 22250 18352
rect 28276 18340 28304 18380
rect 22244 18312 28304 18340
rect 22244 18300 22250 18312
rect 29546 18300 29552 18352
rect 29604 18349 29610 18352
rect 29604 18343 29668 18349
rect 29604 18309 29622 18343
rect 29656 18309 29668 18343
rect 32048 18340 32076 18380
rect 32125 18377 32137 18411
rect 32171 18408 32183 18411
rect 32214 18408 32220 18420
rect 32171 18380 32220 18408
rect 32171 18377 32183 18380
rect 32125 18371 32183 18377
rect 32214 18368 32220 18380
rect 32272 18368 32278 18420
rect 35618 18408 35624 18420
rect 32416 18380 35480 18408
rect 35579 18380 35624 18408
rect 32416 18340 32444 18380
rect 33597 18343 33655 18349
rect 33597 18340 33609 18343
rect 32048 18312 32444 18340
rect 32692 18312 33609 18340
rect 29604 18303 29668 18309
rect 29604 18300 29610 18303
rect 9657 18275 9720 18281
rect 9657 18241 9669 18275
rect 9703 18244 9720 18275
rect 9769 18275 9827 18281
rect 9703 18241 9715 18244
rect 9657 18235 9715 18241
rect 9769 18241 9781 18275
rect 9815 18241 9827 18275
rect 9769 18235 9827 18241
rect 8864 18108 9536 18136
rect 1578 18028 1584 18080
rect 1636 18068 1642 18080
rect 2133 18071 2191 18077
rect 2133 18068 2145 18071
rect 1636 18040 2145 18068
rect 1636 18028 1642 18040
rect 2133 18037 2145 18040
rect 2179 18037 2191 18071
rect 2866 18068 2872 18080
rect 2827 18040 2872 18068
rect 2133 18031 2191 18037
rect 2866 18028 2872 18040
rect 2924 18028 2930 18080
rect 4062 18028 4068 18080
rect 4120 18068 4126 18080
rect 6822 18068 6828 18080
rect 4120 18040 6828 18068
rect 4120 18028 4126 18040
rect 6822 18028 6828 18040
rect 6880 18028 6886 18080
rect 6914 18028 6920 18080
rect 6972 18068 6978 18080
rect 6972 18040 7017 18068
rect 6972 18028 6978 18040
rect 8202 18028 8208 18080
rect 8260 18068 8266 18080
rect 8864 18077 8892 18108
rect 8849 18071 8907 18077
rect 8849 18068 8861 18071
rect 8260 18040 8861 18068
rect 8260 18028 8266 18040
rect 8849 18037 8861 18040
rect 8895 18037 8907 18071
rect 9398 18068 9404 18080
rect 9359 18040 9404 18068
rect 8849 18031 8907 18037
rect 9398 18028 9404 18040
rect 9456 18028 9462 18080
rect 9508 18068 9536 18108
rect 9582 18096 9588 18148
rect 9640 18136 9646 18148
rect 9784 18136 9812 18235
rect 9858 18232 9864 18284
rect 9916 18272 9922 18284
rect 10045 18275 10103 18281
rect 9916 18244 9961 18272
rect 9916 18232 9922 18244
rect 10045 18241 10057 18275
rect 10091 18272 10103 18275
rect 10226 18272 10232 18284
rect 10091 18244 10232 18272
rect 10091 18241 10103 18244
rect 10045 18235 10103 18241
rect 10226 18232 10232 18244
rect 10284 18232 10290 18284
rect 10502 18272 10508 18284
rect 10463 18244 10508 18272
rect 10502 18232 10508 18244
rect 10560 18232 10566 18284
rect 10689 18275 10747 18281
rect 10689 18272 10701 18275
rect 10612 18244 10701 18272
rect 9640 18108 9812 18136
rect 9640 18096 9646 18108
rect 10612 18068 10640 18244
rect 10689 18241 10701 18244
rect 10735 18241 10747 18275
rect 11698 18272 11704 18284
rect 11659 18244 11704 18272
rect 10689 18235 10747 18241
rect 11698 18232 11704 18244
rect 11756 18232 11762 18284
rect 12986 18272 12992 18284
rect 12947 18244 12992 18272
rect 12986 18232 12992 18244
rect 13044 18232 13050 18284
rect 15841 18275 15899 18281
rect 15841 18241 15853 18275
rect 15887 18241 15899 18275
rect 15841 18235 15899 18241
rect 15856 18136 15884 18235
rect 17034 18232 17040 18284
rect 17092 18281 17098 18284
rect 17092 18275 17141 18281
rect 17092 18241 17095 18275
rect 17129 18241 17141 18275
rect 17092 18235 17141 18241
rect 17218 18278 17276 18284
rect 17218 18244 17230 18278
rect 17264 18244 17276 18278
rect 17218 18238 17276 18244
rect 17313 18278 17371 18284
rect 17313 18244 17325 18278
rect 17359 18244 17371 18278
rect 17494 18272 17500 18284
rect 17455 18244 17500 18272
rect 17313 18238 17371 18244
rect 17092 18232 17098 18235
rect 17494 18232 17500 18244
rect 17552 18232 17558 18284
rect 19889 18275 19947 18281
rect 19889 18241 19901 18275
rect 19935 18272 19947 18275
rect 19978 18272 19984 18284
rect 19935 18244 19984 18272
rect 19935 18241 19947 18244
rect 19889 18235 19947 18241
rect 19978 18232 19984 18244
rect 20036 18232 20042 18284
rect 20162 18281 20168 18284
rect 20156 18272 20168 18281
rect 20123 18244 20168 18272
rect 20156 18235 20168 18244
rect 20162 18232 20168 18235
rect 20220 18232 20226 18284
rect 23569 18275 23627 18281
rect 23569 18241 23581 18275
rect 23615 18241 23627 18275
rect 23753 18275 23811 18281
rect 23753 18272 23765 18275
rect 23569 18235 23627 18241
rect 23676 18244 23765 18272
rect 18138 18136 18144 18148
rect 15856 18108 18144 18136
rect 18138 18096 18144 18108
rect 18196 18096 18202 18148
rect 9508 18040 10640 18068
rect 20162 18028 20168 18080
rect 20220 18068 20226 18080
rect 20530 18068 20536 18080
rect 20220 18040 20536 18068
rect 20220 18028 20226 18040
rect 20530 18028 20536 18040
rect 20588 18028 20594 18080
rect 21082 18028 21088 18080
rect 21140 18068 21146 18080
rect 21266 18068 21272 18080
rect 21140 18040 21272 18068
rect 21140 18028 21146 18040
rect 21266 18028 21272 18040
rect 21324 18028 21330 18080
rect 23584 18068 23612 18235
rect 23676 18216 23704 18244
rect 23753 18241 23765 18244
rect 23799 18241 23811 18275
rect 23753 18235 23811 18241
rect 23845 18275 23903 18281
rect 23845 18241 23857 18275
rect 23891 18241 23903 18275
rect 23845 18235 23903 18241
rect 23658 18164 23664 18216
rect 23716 18164 23722 18216
rect 23860 18148 23888 18235
rect 23934 18232 23940 18284
rect 23992 18272 23998 18284
rect 23992 18244 24037 18272
rect 23992 18232 23998 18244
rect 24210 18232 24216 18284
rect 24268 18272 24274 18284
rect 24765 18275 24823 18281
rect 24765 18272 24777 18275
rect 24268 18244 24777 18272
rect 24268 18232 24274 18244
rect 24765 18241 24777 18244
rect 24811 18241 24823 18275
rect 25038 18272 25044 18284
rect 24999 18244 25044 18272
rect 24765 18235 24823 18241
rect 25038 18232 25044 18244
rect 25096 18232 25102 18284
rect 25314 18232 25320 18284
rect 25372 18272 25378 18284
rect 25866 18272 25872 18284
rect 25372 18244 25872 18272
rect 25372 18232 25378 18244
rect 25866 18232 25872 18244
rect 25924 18232 25930 18284
rect 26160 18244 27200 18272
rect 26160 18216 26188 18244
rect 24949 18207 25007 18213
rect 24949 18173 24961 18207
rect 24995 18204 25007 18207
rect 26142 18204 26148 18216
rect 24995 18176 25728 18204
rect 26103 18176 26148 18204
rect 24995 18173 25007 18176
rect 24949 18167 25007 18173
rect 23842 18096 23848 18148
rect 23900 18096 23906 18148
rect 24026 18096 24032 18148
rect 24084 18136 24090 18148
rect 25700 18145 25728 18176
rect 26142 18164 26148 18176
rect 26200 18164 26206 18216
rect 26326 18164 26332 18216
rect 26384 18204 26390 18216
rect 26694 18204 26700 18216
rect 26384 18176 26700 18204
rect 26384 18164 26390 18176
rect 26694 18164 26700 18176
rect 26752 18164 26758 18216
rect 27172 18204 27200 18244
rect 27246 18232 27252 18284
rect 27304 18272 27310 18284
rect 27304 18244 27346 18272
rect 27448 18244 28120 18272
rect 27304 18232 27310 18244
rect 27448 18204 27476 18244
rect 27706 18204 27712 18216
rect 27172 18176 27476 18204
rect 27667 18176 27712 18204
rect 27706 18164 27712 18176
rect 27764 18164 27770 18216
rect 28092 18204 28120 18244
rect 28166 18232 28172 18284
rect 28224 18272 28230 18284
rect 28350 18272 28356 18284
rect 28224 18244 28356 18272
rect 28224 18232 28230 18244
rect 28350 18232 28356 18244
rect 28408 18232 28414 18284
rect 28537 18275 28595 18281
rect 28537 18241 28549 18275
rect 28583 18272 28595 18275
rect 28583 18244 30788 18272
rect 28583 18241 28595 18244
rect 28537 18235 28595 18241
rect 28552 18204 28580 18235
rect 28092 18176 28580 18204
rect 28629 18207 28687 18213
rect 28629 18173 28641 18207
rect 28675 18173 28687 18207
rect 28629 18167 28687 18173
rect 25225 18139 25283 18145
rect 25225 18136 25237 18139
rect 24084 18108 25237 18136
rect 24084 18096 24090 18108
rect 25225 18105 25237 18108
rect 25271 18105 25283 18139
rect 25225 18099 25283 18105
rect 25685 18139 25743 18145
rect 25685 18105 25697 18139
rect 25731 18136 25743 18139
rect 25774 18136 25780 18148
rect 25731 18108 25780 18136
rect 25731 18105 25743 18108
rect 25685 18099 25743 18105
rect 25774 18096 25780 18108
rect 25832 18096 25838 18148
rect 27065 18139 27123 18145
rect 27065 18105 27077 18139
rect 27111 18136 27123 18139
rect 28644 18136 28672 18167
rect 28718 18164 28724 18216
rect 28776 18204 28782 18216
rect 29365 18207 29423 18213
rect 28776 18176 28821 18204
rect 28776 18164 28782 18176
rect 29365 18173 29377 18207
rect 29411 18173 29423 18207
rect 29365 18167 29423 18173
rect 27111 18108 28672 18136
rect 27111 18105 27123 18108
rect 27065 18099 27123 18105
rect 24578 18068 24584 18080
rect 23584 18040 24584 18068
rect 24578 18028 24584 18040
rect 24636 18028 24642 18080
rect 25041 18071 25099 18077
rect 25041 18037 25053 18071
rect 25087 18068 25099 18071
rect 25590 18068 25596 18080
rect 25087 18040 25596 18068
rect 25087 18037 25099 18040
rect 25041 18031 25099 18037
rect 25590 18028 25596 18040
rect 25648 18028 25654 18080
rect 27430 18028 27436 18080
rect 27488 18068 27494 18080
rect 27617 18071 27675 18077
rect 27617 18068 27629 18071
rect 27488 18040 27629 18068
rect 27488 18028 27494 18040
rect 27617 18037 27629 18040
rect 27663 18037 27675 18071
rect 27617 18031 27675 18037
rect 27982 18028 27988 18080
rect 28040 18068 28046 18080
rect 28718 18068 28724 18080
rect 28040 18040 28724 18068
rect 28040 18028 28046 18040
rect 28718 18028 28724 18040
rect 28776 18028 28782 18080
rect 29380 18068 29408 18167
rect 30760 18145 30788 18244
rect 30834 18232 30840 18284
rect 30892 18272 30898 18284
rect 32401 18275 32459 18281
rect 32401 18272 32413 18275
rect 30892 18244 32413 18272
rect 30892 18232 30898 18244
rect 32401 18241 32413 18244
rect 32447 18241 32459 18275
rect 32401 18235 32459 18241
rect 32506 18275 32564 18281
rect 32506 18241 32518 18275
rect 32552 18241 32564 18275
rect 32506 18235 32564 18241
rect 32606 18275 32664 18281
rect 32606 18241 32618 18275
rect 32652 18272 32664 18275
rect 32692 18272 32720 18312
rect 33597 18309 33609 18312
rect 33643 18309 33655 18343
rect 35452 18340 35480 18380
rect 35618 18368 35624 18380
rect 35676 18368 35682 18420
rect 36630 18340 36636 18352
rect 35452 18312 36636 18340
rect 33597 18303 33655 18309
rect 36630 18300 36636 18312
rect 36688 18300 36694 18352
rect 37458 18340 37464 18352
rect 37419 18312 37464 18340
rect 37458 18300 37464 18312
rect 37516 18300 37522 18352
rect 39117 18343 39175 18349
rect 39117 18309 39129 18343
rect 39163 18340 39175 18343
rect 40126 18340 40132 18352
rect 39163 18312 40132 18340
rect 39163 18309 39175 18312
rect 39117 18303 39175 18309
rect 40126 18300 40132 18312
rect 40184 18300 40190 18352
rect 32652 18244 32720 18272
rect 32652 18241 32664 18244
rect 32606 18235 32664 18241
rect 32521 18148 32549 18235
rect 32766 18232 32772 18284
rect 32824 18275 32830 18284
rect 32824 18272 32884 18275
rect 32824 18244 32917 18272
rect 32824 18232 32830 18244
rect 32876 18204 32904 18244
rect 33134 18232 33140 18284
rect 33192 18272 33198 18284
rect 33229 18275 33287 18281
rect 33229 18272 33241 18275
rect 33192 18244 33241 18272
rect 33192 18232 33198 18244
rect 33229 18241 33241 18244
rect 33275 18241 33287 18275
rect 33410 18272 33416 18284
rect 33371 18244 33416 18272
rect 33229 18235 33287 18241
rect 33410 18232 33416 18244
rect 33468 18232 33474 18284
rect 34508 18275 34566 18281
rect 34508 18241 34520 18275
rect 34554 18272 34566 18275
rect 34790 18272 34796 18284
rect 34554 18244 34796 18272
rect 34554 18241 34566 18244
rect 34508 18235 34566 18241
rect 34790 18232 34796 18244
rect 34848 18232 34854 18284
rect 36078 18272 36084 18284
rect 36039 18244 36084 18272
rect 36078 18232 36084 18244
rect 36136 18232 36142 18284
rect 36170 18232 36176 18284
rect 36228 18272 36234 18284
rect 36265 18275 36323 18281
rect 36265 18272 36277 18275
rect 36228 18244 36277 18272
rect 36228 18232 36234 18244
rect 36265 18241 36277 18244
rect 36311 18272 36323 18275
rect 37277 18275 37335 18281
rect 37277 18272 37289 18275
rect 36311 18244 37289 18272
rect 36311 18241 36323 18244
rect 36265 18235 36323 18241
rect 37277 18241 37289 18244
rect 37323 18241 37335 18275
rect 37277 18235 37335 18241
rect 33686 18204 33692 18216
rect 32876 18176 33692 18204
rect 33686 18164 33692 18176
rect 33744 18164 33750 18216
rect 34241 18207 34299 18213
rect 34241 18173 34253 18207
rect 34287 18173 34299 18207
rect 34241 18167 34299 18173
rect 30745 18139 30803 18145
rect 30745 18105 30757 18139
rect 30791 18105 30803 18139
rect 30745 18099 30803 18105
rect 32490 18096 32496 18148
rect 32548 18096 32554 18148
rect 29546 18068 29552 18080
rect 29380 18040 29552 18068
rect 29546 18028 29552 18040
rect 29604 18028 29610 18080
rect 34256 18068 34284 18167
rect 34606 18068 34612 18080
rect 34256 18040 34612 18068
rect 34606 18028 34612 18040
rect 34664 18028 34670 18080
rect 35342 18028 35348 18080
rect 35400 18068 35406 18080
rect 36449 18071 36507 18077
rect 36449 18068 36461 18071
rect 35400 18040 36461 18068
rect 35400 18028 35406 18040
rect 36449 18037 36461 18040
rect 36495 18037 36507 18071
rect 36449 18031 36507 18037
rect 1104 17978 48852 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 48852 17978
rect 1104 17904 48852 17926
rect 9950 17824 9956 17876
rect 10008 17864 10014 17876
rect 10008 17836 12434 17864
rect 10008 17824 10014 17836
rect 2866 17796 2872 17808
rect 1412 17768 2872 17796
rect 1412 17737 1440 17768
rect 2866 17756 2872 17768
rect 2924 17756 2930 17808
rect 7466 17796 7472 17808
rect 6748 17768 7472 17796
rect 1397 17731 1455 17737
rect 1397 17697 1409 17731
rect 1443 17697 1455 17731
rect 1578 17728 1584 17740
rect 1539 17700 1584 17728
rect 1397 17691 1455 17697
rect 1578 17688 1584 17700
rect 1636 17688 1642 17740
rect 2774 17688 2780 17740
rect 2832 17728 2838 17740
rect 6748 17737 6776 17768
rect 7466 17756 7472 17768
rect 7524 17756 7530 17808
rect 12406 17796 12434 17836
rect 17862 17824 17868 17876
rect 17920 17864 17926 17876
rect 24765 17867 24823 17873
rect 17920 17836 24164 17864
rect 17920 17824 17926 17836
rect 18138 17796 18144 17808
rect 12406 17768 16068 17796
rect 18099 17768 18144 17796
rect 6733 17731 6791 17737
rect 2832 17700 2877 17728
rect 2832 17688 2838 17700
rect 6733 17697 6745 17731
rect 6779 17697 6791 17731
rect 6733 17691 6791 17697
rect 6822 17688 6828 17740
rect 6880 17728 6886 17740
rect 7009 17731 7067 17737
rect 7009 17728 7021 17731
rect 6880 17700 7021 17728
rect 6880 17688 6886 17700
rect 7009 17697 7021 17700
rect 7055 17697 7067 17731
rect 7484 17728 7512 17756
rect 8941 17731 8999 17737
rect 8941 17728 8953 17731
rect 7484 17700 8953 17728
rect 7009 17691 7067 17697
rect 8941 17697 8953 17700
rect 8987 17697 8999 17731
rect 15746 17728 15752 17740
rect 15707 17700 15752 17728
rect 8941 17691 8999 17697
rect 8956 17660 8984 17691
rect 15746 17688 15752 17700
rect 15804 17688 15810 17740
rect 16040 17737 16068 17768
rect 18138 17756 18144 17768
rect 18196 17756 18202 17808
rect 24136 17796 24164 17836
rect 24765 17833 24777 17867
rect 24811 17864 24823 17867
rect 25222 17864 25228 17876
rect 24811 17836 25228 17864
rect 24811 17833 24823 17836
rect 24765 17827 24823 17833
rect 25222 17824 25228 17836
rect 25280 17824 25286 17876
rect 25590 17864 25596 17876
rect 25551 17836 25596 17864
rect 25590 17824 25596 17836
rect 25648 17824 25654 17876
rect 26234 17864 26240 17876
rect 26195 17836 26240 17864
rect 26234 17824 26240 17836
rect 26292 17824 26298 17876
rect 26418 17824 26424 17876
rect 26476 17864 26482 17876
rect 29914 17864 29920 17876
rect 26476 17836 29920 17864
rect 26476 17824 26482 17836
rect 29914 17824 29920 17836
rect 29972 17824 29978 17876
rect 33137 17867 33195 17873
rect 33137 17833 33149 17867
rect 33183 17864 33195 17867
rect 34790 17864 34796 17876
rect 33183 17836 34796 17864
rect 33183 17833 33195 17836
rect 33137 17827 33195 17833
rect 34790 17824 34796 17836
rect 34848 17824 34854 17876
rect 36170 17864 36176 17876
rect 36131 17836 36176 17864
rect 36170 17824 36176 17836
rect 36228 17824 36234 17876
rect 26326 17796 26332 17808
rect 24136 17768 26332 17796
rect 26326 17756 26332 17768
rect 26384 17756 26390 17808
rect 26605 17799 26663 17805
rect 26605 17796 26617 17799
rect 26436 17768 26617 17796
rect 16025 17731 16083 17737
rect 16025 17697 16037 17731
rect 16071 17697 16083 17731
rect 24578 17728 24584 17740
rect 16025 17691 16083 17697
rect 19260 17700 20484 17728
rect 24539 17700 24584 17728
rect 10781 17663 10839 17669
rect 10781 17660 10793 17663
rect 8956 17632 10793 17660
rect 10781 17629 10793 17632
rect 10827 17660 10839 17663
rect 12434 17660 12440 17672
rect 10827 17632 12440 17660
rect 10827 17629 10839 17632
rect 10781 17623 10839 17629
rect 12434 17620 12440 17632
rect 12492 17660 12498 17672
rect 12986 17660 12992 17672
rect 12492 17632 12992 17660
rect 12492 17620 12498 17632
rect 12986 17620 12992 17632
rect 13044 17620 13050 17672
rect 14921 17663 14979 17669
rect 14921 17629 14933 17663
rect 14967 17660 14979 17663
rect 15562 17660 15568 17672
rect 14967 17632 15568 17660
rect 14967 17629 14979 17632
rect 14921 17623 14979 17629
rect 15562 17620 15568 17632
rect 15620 17620 15626 17672
rect 6825 17595 6883 17601
rect 6825 17561 6837 17595
rect 6871 17592 6883 17595
rect 6914 17592 6920 17604
rect 6871 17564 6920 17592
rect 6871 17561 6883 17564
rect 6825 17555 6883 17561
rect 6914 17552 6920 17564
rect 6972 17552 6978 17604
rect 9208 17595 9266 17601
rect 9208 17561 9220 17595
rect 9254 17592 9266 17595
rect 9398 17592 9404 17604
rect 9254 17564 9404 17592
rect 9254 17561 9266 17564
rect 9208 17555 9266 17561
rect 9398 17552 9404 17564
rect 9456 17552 9462 17604
rect 11048 17595 11106 17601
rect 11048 17561 11060 17595
rect 11094 17592 11106 17595
rect 11330 17592 11336 17604
rect 11094 17564 11336 17592
rect 11094 17561 11106 17564
rect 11048 17555 11106 17561
rect 11330 17552 11336 17564
rect 11388 17552 11394 17604
rect 14737 17595 14795 17601
rect 14737 17561 14749 17595
rect 14783 17592 14795 17595
rect 15194 17592 15200 17604
rect 14783 17564 15200 17592
rect 14783 17561 14795 17564
rect 14737 17555 14795 17561
rect 15194 17552 15200 17564
rect 15252 17552 15258 17604
rect 17954 17592 17960 17604
rect 17915 17564 17960 17592
rect 17954 17552 17960 17564
rect 18012 17552 18018 17604
rect 19260 17592 19288 17700
rect 19334 17620 19340 17672
rect 19392 17660 19398 17672
rect 20349 17663 20407 17669
rect 20349 17660 20361 17663
rect 19392 17632 20361 17660
rect 19392 17620 19398 17632
rect 20349 17629 20361 17632
rect 20395 17629 20407 17663
rect 20456 17660 20484 17700
rect 24578 17688 24584 17700
rect 24636 17688 24642 17740
rect 25777 17731 25835 17737
rect 25777 17697 25789 17731
rect 25823 17697 25835 17731
rect 25777 17691 25835 17697
rect 24765 17663 24823 17669
rect 20456 17632 20852 17660
rect 20349 17623 20407 17629
rect 20824 17604 20852 17632
rect 24765 17629 24777 17663
rect 24811 17660 24823 17663
rect 24854 17660 24860 17672
rect 24811 17632 24860 17660
rect 24811 17629 24823 17632
rect 24765 17623 24823 17629
rect 24854 17620 24860 17632
rect 24912 17620 24918 17672
rect 25038 17620 25044 17672
rect 25096 17660 25102 17672
rect 25498 17660 25504 17672
rect 25096 17632 25504 17660
rect 25096 17620 25102 17632
rect 25498 17620 25504 17632
rect 25556 17620 25562 17672
rect 25792 17660 25820 17691
rect 25866 17688 25872 17740
rect 25924 17728 25930 17740
rect 26436 17728 26464 17768
rect 26605 17765 26617 17768
rect 26651 17765 26663 17799
rect 26605 17759 26663 17765
rect 26694 17756 26700 17808
rect 26752 17796 26758 17808
rect 27338 17796 27344 17808
rect 26752 17768 27344 17796
rect 26752 17756 26758 17768
rect 27338 17756 27344 17768
rect 27396 17796 27402 17808
rect 28721 17799 28779 17805
rect 28721 17796 28733 17799
rect 27396 17768 28733 17796
rect 27396 17756 27402 17768
rect 28721 17765 28733 17768
rect 28767 17765 28779 17799
rect 34422 17796 34428 17808
rect 28721 17759 28779 17765
rect 33520 17768 34428 17796
rect 25924 17700 26464 17728
rect 26513 17731 26571 17737
rect 25924 17688 25930 17700
rect 26513 17697 26525 17731
rect 26559 17728 26571 17731
rect 27249 17731 27307 17737
rect 27249 17728 27261 17731
rect 26559 17700 27261 17728
rect 26559 17697 26571 17700
rect 26513 17691 26571 17697
rect 27249 17697 27261 17700
rect 27295 17728 27307 17731
rect 27706 17728 27712 17740
rect 27295 17700 27712 17728
rect 27295 17697 27307 17700
rect 27249 17691 27307 17697
rect 27706 17688 27712 17700
rect 27764 17688 27770 17740
rect 27798 17688 27804 17740
rect 27856 17728 27862 17740
rect 32125 17731 32183 17737
rect 27856 17700 29684 17728
rect 27856 17688 27862 17700
rect 26234 17660 26240 17672
rect 25792 17632 26240 17660
rect 26234 17620 26240 17632
rect 26292 17620 26298 17672
rect 26418 17660 26424 17672
rect 26379 17632 26424 17660
rect 26418 17620 26424 17632
rect 26476 17620 26482 17672
rect 26697 17663 26755 17669
rect 26697 17629 26709 17663
rect 26743 17660 26755 17663
rect 26786 17660 26792 17672
rect 26743 17632 26792 17660
rect 26743 17629 26755 17632
rect 26697 17623 26755 17629
rect 26786 17620 26792 17632
rect 26844 17620 26850 17672
rect 27062 17620 27068 17672
rect 27120 17660 27126 17672
rect 27525 17663 27583 17669
rect 27525 17660 27537 17663
rect 27120 17632 27537 17660
rect 27120 17620 27126 17632
rect 27525 17629 27537 17632
rect 27571 17629 27583 17663
rect 27525 17623 27583 17629
rect 28537 17663 28595 17669
rect 28537 17629 28549 17663
rect 28583 17660 28595 17663
rect 28626 17660 28632 17672
rect 28583 17632 28632 17660
rect 28583 17629 28595 17632
rect 28537 17623 28595 17629
rect 28626 17620 28632 17632
rect 28684 17620 28690 17672
rect 29546 17660 29552 17672
rect 29507 17632 29552 17660
rect 29546 17620 29552 17632
rect 29604 17620 29610 17672
rect 29656 17660 29684 17700
rect 32125 17697 32137 17731
rect 32171 17728 32183 17731
rect 32490 17728 32496 17740
rect 32171 17700 32496 17728
rect 32171 17697 32183 17700
rect 32125 17691 32183 17697
rect 32490 17688 32496 17700
rect 32548 17728 32554 17740
rect 33520 17728 33548 17768
rect 34422 17756 34428 17768
rect 34480 17756 34486 17808
rect 34514 17728 34520 17740
rect 32548 17700 33548 17728
rect 32548 17688 32554 17700
rect 31662 17660 31668 17672
rect 29656 17632 31668 17660
rect 31662 17620 31668 17632
rect 31720 17620 31726 17672
rect 31754 17620 31760 17672
rect 31812 17660 31818 17672
rect 31849 17663 31907 17669
rect 31849 17660 31861 17663
rect 31812 17632 31861 17660
rect 31812 17620 31818 17632
rect 31849 17629 31861 17632
rect 31895 17629 31907 17663
rect 31849 17623 31907 17629
rect 31938 17620 31944 17672
rect 31996 17660 32002 17672
rect 33520 17669 33548 17700
rect 33612 17700 34520 17728
rect 33612 17669 33640 17700
rect 34514 17688 34520 17700
rect 34572 17688 34578 17740
rect 35894 17688 35900 17740
rect 35952 17728 35958 17740
rect 37277 17731 37335 17737
rect 37277 17728 37289 17731
rect 35952 17700 37289 17728
rect 35952 17688 35958 17700
rect 37277 17697 37289 17700
rect 37323 17697 37335 17731
rect 39114 17728 39120 17740
rect 39075 17700 39120 17728
rect 37277 17691 37335 17697
rect 39114 17688 39120 17700
rect 39172 17688 39178 17740
rect 33413 17663 33471 17669
rect 33413 17660 33425 17663
rect 31996 17632 33425 17660
rect 31996 17620 32002 17632
rect 33413 17629 33425 17632
rect 33459 17629 33471 17663
rect 33413 17623 33471 17629
rect 33505 17663 33563 17669
rect 33505 17629 33517 17663
rect 33551 17629 33563 17663
rect 33505 17623 33563 17629
rect 33597 17663 33655 17669
rect 33597 17629 33609 17663
rect 33643 17629 33655 17663
rect 33597 17623 33655 17629
rect 33686 17620 33692 17672
rect 33744 17660 33750 17672
rect 33781 17663 33839 17669
rect 33781 17660 33793 17663
rect 33744 17632 33793 17660
rect 33744 17620 33750 17632
rect 33781 17629 33793 17632
rect 33827 17629 33839 17663
rect 33781 17623 33839 17629
rect 34606 17620 34612 17672
rect 34664 17660 34670 17672
rect 34793 17663 34851 17669
rect 34793 17660 34805 17663
rect 34664 17632 34805 17660
rect 34664 17620 34670 17632
rect 34793 17629 34805 17632
rect 34839 17629 34851 17663
rect 36630 17660 36636 17672
rect 36591 17632 36636 17660
rect 34793 17623 34851 17629
rect 36630 17620 36636 17632
rect 36688 17620 36694 17672
rect 47118 17620 47124 17672
rect 47176 17660 47182 17672
rect 47673 17663 47731 17669
rect 47673 17660 47685 17663
rect 47176 17632 47685 17660
rect 47176 17620 47182 17632
rect 47673 17629 47685 17632
rect 47719 17629 47731 17663
rect 47673 17623 47731 17629
rect 19521 17595 19579 17601
rect 19521 17592 19533 17595
rect 19260 17564 19533 17592
rect 19521 17561 19533 17564
rect 19567 17561 19579 17595
rect 19521 17555 19579 17561
rect 19705 17595 19763 17601
rect 19705 17561 19717 17595
rect 19751 17561 19763 17595
rect 19705 17555 19763 17561
rect 9582 17484 9588 17536
rect 9640 17524 9646 17536
rect 10321 17527 10379 17533
rect 10321 17524 10333 17527
rect 9640 17496 10333 17524
rect 9640 17484 9646 17496
rect 10321 17493 10333 17496
rect 10367 17493 10379 17527
rect 10321 17487 10379 17493
rect 11514 17484 11520 17536
rect 11572 17524 11578 17536
rect 11698 17524 11704 17536
rect 11572 17496 11704 17524
rect 11572 17484 11578 17496
rect 11698 17484 11704 17496
rect 11756 17524 11762 17536
rect 12161 17527 12219 17533
rect 12161 17524 12173 17527
rect 11756 17496 12173 17524
rect 11756 17484 11762 17496
rect 12161 17493 12173 17496
rect 12207 17493 12219 17527
rect 15102 17524 15108 17536
rect 15063 17496 15108 17524
rect 12161 17487 12219 17493
rect 15102 17484 15108 17496
rect 15160 17484 15166 17536
rect 19426 17484 19432 17536
rect 19484 17524 19490 17536
rect 19720 17524 19748 17555
rect 20070 17552 20076 17604
rect 20128 17592 20134 17604
rect 20594 17595 20652 17601
rect 20594 17592 20606 17595
rect 20128 17564 20606 17592
rect 20128 17552 20134 17564
rect 20594 17561 20606 17564
rect 20640 17561 20652 17595
rect 20594 17555 20652 17561
rect 20806 17552 20812 17604
rect 20864 17552 20870 17604
rect 24486 17592 24492 17604
rect 24447 17564 24492 17592
rect 24486 17552 24492 17564
rect 24544 17552 24550 17604
rect 25777 17595 25835 17601
rect 25777 17561 25789 17595
rect 25823 17592 25835 17595
rect 26878 17592 26884 17604
rect 25823 17564 26884 17592
rect 25823 17561 25835 17564
rect 25777 17555 25835 17561
rect 26878 17552 26884 17564
rect 26936 17552 26942 17604
rect 26970 17552 26976 17604
rect 27028 17592 27034 17604
rect 29454 17592 29460 17604
rect 27028 17564 29460 17592
rect 27028 17552 27034 17564
rect 29454 17552 29460 17564
rect 29512 17552 29518 17604
rect 29822 17601 29828 17604
rect 29794 17595 29828 17601
rect 29794 17561 29806 17595
rect 29794 17555 29828 17561
rect 29822 17552 29828 17555
rect 29880 17552 29886 17604
rect 29914 17552 29920 17604
rect 29972 17592 29978 17604
rect 29972 17564 33640 17592
rect 29972 17552 29978 17564
rect 19484 17496 19748 17524
rect 19889 17527 19947 17533
rect 19484 17484 19490 17496
rect 19889 17493 19901 17527
rect 19935 17524 19947 17527
rect 19978 17524 19984 17536
rect 19935 17496 19984 17524
rect 19935 17493 19947 17496
rect 19889 17487 19947 17493
rect 19978 17484 19984 17496
rect 20036 17484 20042 17536
rect 21726 17524 21732 17536
rect 21687 17496 21732 17524
rect 21726 17484 21732 17496
rect 21784 17484 21790 17536
rect 24118 17484 24124 17536
rect 24176 17524 24182 17536
rect 24578 17524 24584 17536
rect 24176 17496 24584 17524
rect 24176 17484 24182 17496
rect 24578 17484 24584 17496
rect 24636 17484 24642 17536
rect 24854 17484 24860 17536
rect 24912 17524 24918 17536
rect 24949 17527 25007 17533
rect 24949 17524 24961 17527
rect 24912 17496 24961 17524
rect 24912 17484 24918 17496
rect 24949 17493 24961 17496
rect 24995 17493 25007 17527
rect 24949 17487 25007 17493
rect 25222 17484 25228 17536
rect 25280 17524 25286 17536
rect 27982 17524 27988 17536
rect 25280 17496 27988 17524
rect 25280 17484 25286 17496
rect 27982 17484 27988 17496
rect 28040 17484 28046 17536
rect 30926 17524 30932 17536
rect 30887 17496 30932 17524
rect 30926 17484 30932 17496
rect 30984 17484 30990 17536
rect 33612 17524 33640 17564
rect 33962 17552 33968 17604
rect 34020 17592 34026 17604
rect 35038 17595 35096 17601
rect 35038 17592 35050 17595
rect 34020 17564 35050 17592
rect 34020 17552 34026 17564
rect 35038 17561 35050 17564
rect 35084 17561 35096 17595
rect 35038 17555 35096 17561
rect 36725 17595 36783 17601
rect 36725 17561 36737 17595
rect 36771 17592 36783 17595
rect 37461 17595 37519 17601
rect 37461 17592 37473 17595
rect 36771 17564 37473 17592
rect 36771 17561 36783 17564
rect 36725 17555 36783 17561
rect 37461 17561 37473 17564
rect 37507 17561 37519 17595
rect 37461 17555 37519 17561
rect 46842 17524 46848 17536
rect 33612 17496 46848 17524
rect 46842 17484 46848 17496
rect 46900 17484 46906 17536
rect 1104 17434 48852 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 48852 17434
rect 1104 17360 48852 17382
rect 1949 17323 2007 17329
rect 1949 17289 1961 17323
rect 1995 17320 2007 17323
rect 23382 17320 23388 17332
rect 1995 17292 23388 17320
rect 1995 17289 2007 17292
rect 1949 17283 2007 17289
rect 23382 17280 23388 17292
rect 23440 17280 23446 17332
rect 23658 17320 23664 17332
rect 23584 17292 23664 17320
rect 9401 17255 9459 17261
rect 9401 17221 9413 17255
rect 9447 17252 9459 17255
rect 9769 17255 9827 17261
rect 9447 17224 9720 17252
rect 9447 17221 9459 17224
rect 9401 17215 9459 17221
rect 1854 17184 1860 17196
rect 1815 17156 1860 17184
rect 1854 17144 1860 17156
rect 1912 17144 1918 17196
rect 9582 17184 9588 17196
rect 9543 17156 9588 17184
rect 9582 17144 9588 17156
rect 9640 17144 9646 17196
rect 9692 17184 9720 17224
rect 9769 17221 9781 17255
rect 9815 17252 9827 17255
rect 9858 17252 9864 17264
rect 9815 17224 9864 17252
rect 9815 17221 9827 17224
rect 9769 17215 9827 17221
rect 9858 17212 9864 17224
rect 9916 17212 9922 17264
rect 20806 17252 20812 17264
rect 12406 17224 20024 17252
rect 10502 17184 10508 17196
rect 9692 17156 10508 17184
rect 10502 17144 10508 17156
rect 10560 17144 10566 17196
rect 3694 17076 3700 17128
rect 3752 17116 3758 17128
rect 12406 17116 12434 17224
rect 12986 17144 12992 17196
rect 13044 17184 13050 17196
rect 14553 17187 14611 17193
rect 14553 17184 14565 17187
rect 13044 17156 14565 17184
rect 13044 17144 13050 17156
rect 14553 17153 14565 17156
rect 14599 17153 14611 17187
rect 14553 17147 14611 17153
rect 14642 17144 14648 17196
rect 14700 17184 14706 17196
rect 14809 17187 14867 17193
rect 14809 17184 14821 17187
rect 14700 17156 14821 17184
rect 14700 17144 14706 17156
rect 14809 17153 14821 17156
rect 14855 17153 14867 17187
rect 14809 17147 14867 17153
rect 16850 17144 16856 17196
rect 16908 17184 16914 17196
rect 19996 17193 20024 17224
rect 20180 17224 20484 17252
rect 20767 17224 20812 17252
rect 20180 17193 20208 17224
rect 17293 17187 17351 17193
rect 17293 17184 17305 17187
rect 16908 17156 17305 17184
rect 16908 17144 16914 17156
rect 17293 17153 17305 17156
rect 17339 17153 17351 17187
rect 17293 17147 17351 17153
rect 19981 17187 20039 17193
rect 19981 17153 19993 17187
rect 20027 17153 20039 17187
rect 19981 17147 20039 17153
rect 20073 17187 20131 17193
rect 20073 17153 20085 17187
rect 20119 17153 20131 17187
rect 20073 17147 20131 17153
rect 20165 17187 20223 17193
rect 20165 17153 20177 17187
rect 20211 17153 20223 17187
rect 20346 17184 20352 17196
rect 20307 17156 20352 17184
rect 20165 17147 20223 17153
rect 3752 17088 12434 17116
rect 3752 17076 3758 17088
rect 16666 17076 16672 17128
rect 16724 17116 16730 17128
rect 17037 17119 17095 17125
rect 17037 17116 17049 17119
rect 16724 17088 17049 17116
rect 16724 17076 16730 17088
rect 17037 17085 17049 17088
rect 17083 17085 17095 17119
rect 17037 17079 17095 17085
rect 19886 17076 19892 17128
rect 19944 17116 19950 17128
rect 20088 17116 20116 17147
rect 20346 17144 20352 17156
rect 20404 17144 20410 17196
rect 19944 17088 20116 17116
rect 20456 17116 20484 17224
rect 20806 17212 20812 17224
rect 20864 17212 20870 17264
rect 20993 17255 21051 17261
rect 20993 17221 21005 17255
rect 21039 17252 21051 17255
rect 21726 17252 21732 17264
rect 21039 17224 21732 17252
rect 21039 17221 21051 17224
rect 20993 17215 21051 17221
rect 21726 17212 21732 17224
rect 21784 17212 21790 17264
rect 23474 17252 23480 17264
rect 23387 17224 23480 17252
rect 23474 17212 23480 17224
rect 23532 17252 23538 17264
rect 23584 17252 23612 17292
rect 23658 17280 23664 17292
rect 23716 17280 23722 17332
rect 23934 17280 23940 17332
rect 23992 17280 23998 17332
rect 24118 17280 24124 17332
rect 24176 17320 24182 17332
rect 24394 17320 24400 17332
rect 24176 17292 24400 17320
rect 24176 17280 24182 17292
rect 24394 17280 24400 17292
rect 24452 17280 24458 17332
rect 24486 17280 24492 17332
rect 24544 17320 24550 17332
rect 24765 17323 24823 17329
rect 24765 17320 24777 17323
rect 24544 17292 24777 17320
rect 24544 17280 24550 17292
rect 24765 17289 24777 17292
rect 24811 17289 24823 17323
rect 25866 17320 25872 17332
rect 25827 17292 25872 17320
rect 24765 17283 24823 17289
rect 25866 17280 25872 17292
rect 25924 17280 25930 17332
rect 27246 17320 27252 17332
rect 27207 17292 27252 17320
rect 27246 17280 27252 17292
rect 27304 17280 27310 17332
rect 27706 17320 27712 17332
rect 27667 17292 27712 17320
rect 27706 17280 27712 17292
rect 27764 17280 27770 17332
rect 27982 17280 27988 17332
rect 28040 17320 28046 17332
rect 28169 17323 28227 17329
rect 28169 17320 28181 17323
rect 28040 17292 28181 17320
rect 28040 17280 28046 17292
rect 28169 17289 28181 17292
rect 28215 17289 28227 17323
rect 28169 17283 28227 17289
rect 29641 17323 29699 17329
rect 29641 17289 29653 17323
rect 29687 17320 29699 17323
rect 29822 17320 29828 17332
rect 29687 17292 29828 17320
rect 29687 17289 29699 17292
rect 29641 17283 29699 17289
rect 29822 17280 29828 17292
rect 29880 17280 29886 17332
rect 33873 17323 33931 17329
rect 33873 17289 33885 17323
rect 33919 17320 33931 17323
rect 33962 17320 33968 17332
rect 33919 17292 33968 17320
rect 33919 17289 33931 17292
rect 33873 17283 33931 17289
rect 33962 17280 33968 17292
rect 34020 17280 34026 17332
rect 35342 17320 35348 17332
rect 34369 17292 35348 17320
rect 23952 17252 23980 17280
rect 23532 17224 23612 17252
rect 23676 17224 23980 17252
rect 24673 17255 24731 17261
rect 23532 17212 23538 17224
rect 23014 17144 23020 17196
rect 23072 17184 23078 17196
rect 23382 17193 23388 17196
rect 23201 17187 23259 17193
rect 23201 17184 23213 17187
rect 23072 17156 23213 17184
rect 23072 17144 23078 17156
rect 23201 17153 23213 17156
rect 23247 17153 23259 17187
rect 23201 17147 23259 17153
rect 23349 17187 23388 17193
rect 23349 17153 23361 17187
rect 23349 17147 23388 17153
rect 23382 17144 23388 17147
rect 23440 17144 23446 17196
rect 23676 17193 23704 17224
rect 24673 17221 24685 17255
rect 24719 17252 24731 17255
rect 28994 17252 29000 17264
rect 24719 17224 29000 17252
rect 24719 17221 24731 17224
rect 24673 17215 24731 17221
rect 23569 17187 23627 17193
rect 23569 17153 23581 17187
rect 23615 17153 23627 17187
rect 23569 17147 23627 17153
rect 23666 17187 23724 17193
rect 23666 17153 23678 17187
rect 23712 17153 23724 17187
rect 23666 17147 23724 17153
rect 21177 17119 21235 17125
rect 21177 17116 21189 17119
rect 20456 17088 21189 17116
rect 19944 17076 19950 17088
rect 21177 17085 21189 17088
rect 21223 17085 21235 17119
rect 21177 17079 21235 17085
rect 23584 17116 23612 17147
rect 24688 17116 24716 17215
rect 28994 17212 29000 17224
rect 29052 17212 29058 17264
rect 34369 17208 34397 17292
rect 35342 17280 35348 17292
rect 35400 17280 35406 17332
rect 36449 17255 36507 17261
rect 36449 17252 36461 17255
rect 25498 17184 25504 17196
rect 25459 17156 25504 17184
rect 25498 17144 25504 17156
rect 25556 17144 25562 17196
rect 25590 17144 25596 17196
rect 25648 17193 25654 17196
rect 25648 17187 25697 17193
rect 25648 17153 25651 17187
rect 25685 17153 25697 17187
rect 25648 17147 25697 17153
rect 25961 17187 26019 17193
rect 25961 17153 25973 17187
rect 26007 17153 26019 17187
rect 25961 17147 26019 17153
rect 25648 17144 25654 17147
rect 23584 17088 24716 17116
rect 24949 17119 25007 17125
rect 15562 17008 15568 17060
rect 15620 17048 15626 17060
rect 15933 17051 15991 17057
rect 15933 17048 15945 17051
rect 15620 17020 15945 17048
rect 15620 17008 15626 17020
rect 15933 17017 15945 17020
rect 15979 17017 15991 17051
rect 15933 17011 15991 17017
rect 19705 17051 19763 17057
rect 19705 17017 19717 17051
rect 19751 17048 19763 17051
rect 20070 17048 20076 17060
rect 19751 17020 20076 17048
rect 19751 17017 19763 17020
rect 19705 17011 19763 17017
rect 20070 17008 20076 17020
rect 20128 17008 20134 17060
rect 20806 17008 20812 17060
rect 20864 17048 20870 17060
rect 23584 17048 23612 17088
rect 24949 17085 24961 17119
rect 24995 17116 25007 17119
rect 25130 17116 25136 17128
rect 24995 17088 25136 17116
rect 24995 17085 25007 17088
rect 24949 17079 25007 17085
rect 25130 17076 25136 17088
rect 25188 17076 25194 17128
rect 25976 17116 26004 17147
rect 26418 17144 26424 17196
rect 26476 17184 26482 17196
rect 26970 17184 26976 17196
rect 26476 17156 26976 17184
rect 26476 17144 26482 17156
rect 26970 17144 26976 17156
rect 27028 17144 27034 17196
rect 27062 17144 27068 17196
rect 27120 17184 27126 17196
rect 27120 17156 27165 17184
rect 27120 17144 27126 17156
rect 27522 17144 27528 17196
rect 27580 17184 27586 17196
rect 28077 17187 28135 17193
rect 28077 17184 28089 17187
rect 27580 17156 28089 17184
rect 27580 17144 27586 17156
rect 28077 17153 28089 17156
rect 28123 17184 28135 17187
rect 28902 17184 28908 17196
rect 28123 17156 28764 17184
rect 28863 17156 28908 17184
rect 28123 17153 28135 17156
rect 28077 17147 28135 17153
rect 25700 17088 26004 17116
rect 27249 17119 27307 17125
rect 25222 17048 25228 17060
rect 20864 17020 23612 17048
rect 23722 17020 25228 17048
rect 20864 17008 20870 17020
rect 18322 16940 18328 16992
rect 18380 16980 18386 16992
rect 18417 16983 18475 16989
rect 18417 16980 18429 16983
rect 18380 16952 18429 16980
rect 18380 16940 18386 16952
rect 18417 16949 18429 16952
rect 18463 16980 18475 16983
rect 23722 16980 23750 17020
rect 25222 17008 25228 17020
rect 25280 17008 25286 17060
rect 23842 16980 23848 16992
rect 18463 16952 23750 16980
rect 23803 16952 23848 16980
rect 18463 16949 18475 16952
rect 18417 16943 18475 16949
rect 23842 16940 23848 16952
rect 23900 16940 23906 16992
rect 24210 16940 24216 16992
rect 24268 16980 24274 16992
rect 24305 16983 24363 16989
rect 24305 16980 24317 16983
rect 24268 16952 24317 16980
rect 24268 16940 24274 16952
rect 24305 16949 24317 16952
rect 24351 16980 24363 16983
rect 25700 16980 25728 17088
rect 27249 17085 27261 17119
rect 27295 17085 27307 17119
rect 27249 17079 27307 17085
rect 28353 17119 28411 17125
rect 28353 17085 28365 17119
rect 28399 17116 28411 17119
rect 28626 17116 28632 17128
rect 28399 17088 28632 17116
rect 28399 17085 28411 17088
rect 28353 17079 28411 17085
rect 25774 17008 25780 17060
rect 25832 17048 25838 17060
rect 27264 17048 27292 17079
rect 28626 17076 28632 17088
rect 28684 17076 28690 17128
rect 28736 17116 28764 17156
rect 28902 17144 28908 17156
rect 28960 17144 28966 17196
rect 29086 17144 29092 17196
rect 29144 17182 29150 17196
rect 29454 17184 29460 17196
rect 29144 17154 29187 17182
rect 29367 17156 29460 17184
rect 29144 17144 29150 17154
rect 29454 17144 29460 17156
rect 29512 17184 29518 17196
rect 31938 17184 31944 17196
rect 29512 17156 31944 17184
rect 29512 17144 29518 17156
rect 31938 17144 31944 17156
rect 31996 17144 32002 17196
rect 32306 17184 32312 17196
rect 32267 17156 32312 17184
rect 32306 17144 32312 17156
rect 32364 17144 32370 17196
rect 34129 17187 34187 17193
rect 34129 17153 34141 17187
rect 34175 17184 34187 17187
rect 34238 17190 34296 17196
rect 34348 17193 34397 17208
rect 35544 17224 36461 17252
rect 34175 17153 34192 17184
rect 34129 17147 34192 17153
rect 34238 17156 34250 17190
rect 34284 17184 34296 17190
rect 34333 17187 34397 17193
rect 34284 17156 34297 17184
rect 34238 17150 34297 17156
rect 28994 17116 29000 17128
rect 28736 17088 29000 17116
rect 28994 17076 29000 17088
rect 29052 17076 29058 17128
rect 29175 17119 29233 17125
rect 29175 17085 29187 17119
rect 29221 17085 29233 17119
rect 29175 17079 29233 17085
rect 29273 17119 29331 17125
rect 29273 17085 29285 17119
rect 29319 17116 29331 17119
rect 29638 17116 29644 17128
rect 29319 17088 29644 17116
rect 29319 17085 29331 17088
rect 29273 17079 29331 17085
rect 25832 17020 27292 17048
rect 25832 17008 25838 17020
rect 27982 17008 27988 17060
rect 28040 17048 28046 17060
rect 29196 17048 29224 17079
rect 29638 17076 29644 17088
rect 29696 17076 29702 17128
rect 31662 17076 31668 17128
rect 31720 17116 31726 17128
rect 34164 17116 34192 17147
rect 31720 17088 34192 17116
rect 34269 17116 34297 17150
rect 34333 17153 34345 17187
rect 34379 17180 34397 17187
rect 34379 17153 34391 17180
rect 34333 17147 34391 17153
rect 34514 17144 34520 17196
rect 34572 17184 34578 17196
rect 35250 17184 35256 17196
rect 34572 17156 34617 17184
rect 35211 17156 35256 17184
rect 34572 17144 34578 17156
rect 35250 17144 35256 17156
rect 35308 17144 35314 17196
rect 35345 17187 35403 17193
rect 35345 17153 35357 17187
rect 35391 17153 35403 17187
rect 35345 17147 35403 17153
rect 35458 17190 35516 17196
rect 35458 17156 35470 17190
rect 35504 17187 35516 17190
rect 35544 17187 35572 17224
rect 36449 17221 36461 17224
rect 36495 17221 36507 17255
rect 36449 17215 36507 17221
rect 35504 17159 35572 17187
rect 35504 17156 35516 17159
rect 35458 17150 35516 17156
rect 34422 17116 34428 17128
rect 34269 17088 34428 17116
rect 31720 17076 31726 17088
rect 34422 17076 34428 17088
rect 34480 17116 34486 17128
rect 35360 17116 35388 17147
rect 35618 17144 35624 17196
rect 35676 17184 35682 17196
rect 36078 17184 36084 17196
rect 35676 17156 35721 17184
rect 36039 17156 36084 17184
rect 35676 17144 35682 17156
rect 36078 17144 36084 17156
rect 36136 17144 36142 17196
rect 36262 17184 36268 17196
rect 36223 17156 36268 17184
rect 36262 17144 36268 17156
rect 36320 17144 36326 17196
rect 36630 17144 36636 17196
rect 36688 17184 36694 17196
rect 37277 17187 37335 17193
rect 37277 17184 37289 17187
rect 36688 17156 37289 17184
rect 36688 17144 36694 17156
rect 37277 17153 37289 17156
rect 37323 17153 37335 17187
rect 46753 17187 46811 17193
rect 46753 17184 46765 17187
rect 37277 17147 37335 17153
rect 45526 17156 46765 17184
rect 34480 17088 35388 17116
rect 34480 17076 34486 17088
rect 30926 17048 30932 17060
rect 28040 17020 30932 17048
rect 28040 17008 28046 17020
rect 30926 17008 30932 17020
rect 30984 17008 30990 17060
rect 45526 17048 45554 17156
rect 46753 17153 46765 17156
rect 46799 17153 46811 17187
rect 46753 17147 46811 17153
rect 32048 17020 45554 17048
rect 24351 16952 25728 16980
rect 24351 16949 24363 16952
rect 24305 16943 24363 16949
rect 26326 16940 26332 16992
rect 26384 16980 26390 16992
rect 31018 16980 31024 16992
rect 26384 16952 31024 16980
rect 26384 16940 26390 16952
rect 31018 16940 31024 16952
rect 31076 16940 31082 16992
rect 31294 16940 31300 16992
rect 31352 16980 31358 16992
rect 32048 16980 32076 17020
rect 31352 16952 32076 16980
rect 32125 16983 32183 16989
rect 31352 16940 31358 16952
rect 32125 16949 32137 16983
rect 32171 16980 32183 16983
rect 33134 16980 33140 16992
rect 32171 16952 33140 16980
rect 32171 16949 32183 16952
rect 32125 16943 32183 16949
rect 33134 16940 33140 16952
rect 33192 16940 33198 16992
rect 34790 16940 34796 16992
rect 34848 16980 34854 16992
rect 34977 16983 35035 16989
rect 34977 16980 34989 16983
rect 34848 16952 34989 16980
rect 34848 16940 34854 16952
rect 34977 16949 34989 16952
rect 35023 16949 35035 16983
rect 37366 16980 37372 16992
rect 37327 16952 37372 16980
rect 34977 16943 35035 16949
rect 37366 16940 37372 16952
rect 37424 16940 37430 16992
rect 46474 16940 46480 16992
rect 46532 16980 46538 16992
rect 46845 16983 46903 16989
rect 46845 16980 46857 16983
rect 46532 16952 46857 16980
rect 46532 16940 46538 16952
rect 46845 16949 46857 16952
rect 46891 16949 46903 16983
rect 47762 16980 47768 16992
rect 47723 16952 47768 16980
rect 46845 16943 46903 16949
rect 47762 16940 47768 16952
rect 47820 16940 47826 16992
rect 1104 16890 48852 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 48852 16890
rect 1104 16816 48852 16838
rect 14553 16779 14611 16785
rect 14553 16745 14565 16779
rect 14599 16776 14611 16779
rect 14642 16776 14648 16788
rect 14599 16748 14648 16776
rect 14599 16745 14611 16748
rect 14553 16739 14611 16745
rect 14642 16736 14648 16748
rect 14700 16736 14706 16788
rect 16850 16776 16856 16788
rect 14752 16748 16160 16776
rect 16811 16748 16856 16776
rect 12066 16708 12072 16720
rect 2884 16680 12072 16708
rect 2038 16532 2044 16584
rect 2096 16572 2102 16584
rect 2884 16581 2912 16680
rect 12066 16668 12072 16680
rect 12124 16668 12130 16720
rect 14752 16708 14780 16748
rect 13786 16680 14780 16708
rect 9953 16643 10011 16649
rect 9953 16609 9965 16643
rect 9999 16640 10011 16643
rect 13541 16643 13599 16649
rect 9999 16612 12434 16640
rect 9999 16609 10011 16612
rect 9953 16603 10011 16609
rect 2225 16575 2283 16581
rect 2225 16572 2237 16575
rect 2096 16544 2237 16572
rect 2096 16532 2102 16544
rect 2225 16541 2237 16544
rect 2271 16541 2283 16575
rect 2225 16535 2283 16541
rect 2869 16575 2927 16581
rect 2869 16541 2881 16575
rect 2915 16541 2927 16575
rect 2869 16535 2927 16541
rect 11606 16532 11612 16584
rect 11664 16572 11670 16584
rect 11793 16575 11851 16581
rect 11793 16572 11805 16575
rect 11664 16544 11805 16572
rect 11664 16532 11670 16544
rect 11793 16541 11805 16544
rect 11839 16541 11851 16575
rect 12406 16572 12434 16612
rect 13541 16609 13553 16643
rect 13587 16640 13599 16643
rect 13786 16640 13814 16680
rect 14826 16668 14832 16720
rect 14884 16668 14890 16720
rect 13587 16612 13814 16640
rect 13587 16609 13599 16612
rect 13541 16603 13599 16609
rect 14734 16600 14740 16652
rect 14792 16600 14798 16652
rect 14844 16640 14872 16668
rect 14844 16612 14964 16640
rect 13357 16575 13415 16581
rect 13357 16572 13369 16575
rect 12406 16544 13369 16572
rect 11793 16535 11851 16541
rect 13357 16541 13369 16544
rect 13403 16572 13415 16575
rect 13722 16572 13728 16584
rect 13403 16544 13728 16572
rect 13403 16541 13415 16544
rect 13357 16535 13415 16541
rect 13722 16532 13728 16544
rect 13780 16532 13786 16584
rect 14752 16569 14780 16600
rect 14936 16581 14964 16612
rect 14829 16575 14887 16581
rect 14829 16569 14841 16575
rect 14752 16541 14841 16569
rect 14875 16541 14887 16575
rect 14824 16538 14887 16541
rect 14829 16535 14887 16538
rect 14918 16575 14976 16581
rect 14918 16541 14930 16575
rect 14964 16541 14976 16575
rect 14918 16535 14976 16541
rect 15013 16575 15071 16581
rect 15013 16541 15025 16575
rect 15059 16572 15071 16575
rect 15102 16572 15108 16584
rect 15059 16544 15108 16572
rect 15059 16541 15071 16544
rect 15013 16535 15071 16541
rect 15102 16532 15108 16544
rect 15160 16532 15166 16584
rect 15197 16575 15255 16581
rect 15197 16541 15209 16575
rect 15243 16541 15255 16575
rect 15197 16535 15255 16541
rect 10134 16504 10140 16516
rect 10095 16476 10140 16504
rect 10134 16464 10140 16476
rect 10192 16464 10198 16516
rect 13173 16507 13231 16513
rect 13173 16473 13185 16507
rect 13219 16473 13231 16507
rect 15212 16504 15240 16535
rect 15378 16532 15384 16584
rect 15436 16572 15442 16584
rect 16132 16581 16160 16748
rect 16850 16736 16856 16748
rect 16908 16736 16914 16788
rect 17954 16736 17960 16788
rect 18012 16776 18018 16788
rect 18506 16776 18512 16788
rect 18012 16748 18512 16776
rect 18012 16736 18018 16748
rect 18506 16736 18512 16748
rect 18564 16776 18570 16788
rect 18601 16779 18659 16785
rect 18601 16776 18613 16779
rect 18564 16748 18613 16776
rect 18564 16736 18570 16748
rect 18601 16745 18613 16748
rect 18647 16745 18659 16779
rect 18601 16739 18659 16745
rect 19426 16736 19432 16788
rect 19484 16776 19490 16788
rect 20625 16779 20683 16785
rect 20625 16776 20637 16779
rect 19484 16748 20637 16776
rect 19484 16736 19490 16748
rect 20625 16745 20637 16748
rect 20671 16776 20683 16779
rect 20806 16776 20812 16788
rect 20671 16748 20812 16776
rect 20671 16745 20683 16748
rect 20625 16739 20683 16745
rect 20806 16736 20812 16748
rect 20864 16736 20870 16788
rect 23845 16779 23903 16785
rect 23845 16745 23857 16779
rect 23891 16776 23903 16779
rect 24210 16776 24216 16788
rect 23891 16748 24216 16776
rect 23891 16745 23903 16748
rect 23845 16739 23903 16745
rect 24210 16736 24216 16748
rect 24268 16736 24274 16788
rect 24394 16776 24400 16788
rect 24355 16748 24400 16776
rect 24394 16736 24400 16748
rect 24452 16736 24458 16788
rect 26697 16779 26755 16785
rect 26697 16745 26709 16779
rect 26743 16776 26755 16779
rect 28902 16776 28908 16788
rect 26743 16748 28908 16776
rect 26743 16745 26755 16748
rect 26697 16739 26755 16745
rect 28902 16736 28908 16748
rect 28960 16736 28966 16788
rect 35894 16776 35900 16788
rect 31726 16748 35900 16776
rect 16316 16680 17540 16708
rect 16316 16581 16344 16680
rect 16390 16600 16396 16652
rect 16448 16640 16454 16652
rect 16448 16612 17264 16640
rect 16448 16600 16454 16612
rect 17236 16581 17264 16612
rect 15887 16575 15945 16581
rect 15887 16572 15899 16575
rect 15436 16544 15899 16572
rect 15436 16532 15442 16544
rect 15887 16541 15899 16544
rect 15933 16541 15945 16575
rect 15887 16535 15945 16541
rect 16025 16575 16083 16581
rect 16025 16541 16037 16575
rect 16071 16541 16083 16575
rect 16025 16535 16083 16541
rect 16117 16575 16175 16581
rect 16117 16541 16129 16575
rect 16163 16541 16175 16575
rect 16117 16535 16175 16541
rect 16301 16575 16359 16581
rect 16301 16541 16313 16575
rect 16347 16572 16359 16575
rect 17129 16575 17187 16581
rect 16347 16544 16528 16572
rect 16347 16541 16359 16544
rect 16301 16535 16359 16541
rect 16040 16504 16068 16535
rect 16390 16504 16396 16516
rect 15212 16476 15792 16504
rect 16040 16476 16396 16504
rect 13173 16467 13231 16473
rect 2222 16396 2228 16448
rect 2280 16436 2286 16448
rect 2961 16439 3019 16445
rect 2961 16436 2973 16439
rect 2280 16408 2973 16436
rect 2280 16396 2286 16408
rect 2961 16405 2973 16408
rect 3007 16405 3019 16439
rect 13188 16436 13216 16467
rect 15194 16436 15200 16448
rect 13188 16408 15200 16436
rect 2961 16399 3019 16405
rect 15194 16396 15200 16408
rect 15252 16396 15258 16448
rect 15654 16436 15660 16448
rect 15615 16408 15660 16436
rect 15654 16396 15660 16408
rect 15712 16396 15718 16448
rect 15764 16436 15792 16476
rect 16390 16464 16396 16476
rect 16448 16464 16454 16516
rect 16500 16436 16528 16544
rect 17129 16541 17141 16575
rect 17175 16541 17187 16575
rect 17129 16535 17187 16541
rect 17221 16575 17279 16581
rect 17221 16541 17233 16575
rect 17267 16541 17279 16575
rect 17221 16535 17279 16541
rect 17144 16504 17172 16535
rect 17310 16532 17316 16584
rect 17368 16572 17374 16584
rect 17512 16581 17540 16680
rect 25222 16668 25228 16720
rect 25280 16708 25286 16720
rect 31726 16708 31754 16748
rect 35894 16736 35900 16748
rect 35952 16736 35958 16788
rect 36081 16779 36139 16785
rect 36081 16745 36093 16779
rect 36127 16776 36139 16779
rect 36262 16776 36268 16788
rect 36127 16748 36268 16776
rect 36127 16745 36139 16748
rect 36081 16739 36139 16745
rect 36262 16736 36268 16748
rect 36320 16736 36326 16788
rect 25280 16680 31754 16708
rect 25280 16668 25286 16680
rect 19242 16640 19248 16652
rect 19203 16612 19248 16640
rect 19242 16600 19248 16612
rect 19300 16600 19306 16652
rect 22462 16640 22468 16652
rect 22423 16612 22468 16640
rect 22462 16600 22468 16612
rect 22520 16600 22526 16652
rect 27982 16600 27988 16652
rect 28040 16640 28046 16652
rect 31294 16640 31300 16652
rect 28040 16612 31300 16640
rect 28040 16600 28046 16612
rect 31294 16600 31300 16612
rect 31352 16600 31358 16652
rect 32490 16640 32496 16652
rect 32324 16612 32496 16640
rect 17497 16575 17555 16581
rect 17368 16544 17413 16572
rect 17368 16532 17374 16544
rect 17497 16541 17509 16575
rect 17543 16572 17555 16575
rect 17862 16572 17868 16584
rect 17543 16544 17868 16572
rect 17543 16541 17555 16544
rect 17497 16535 17555 16541
rect 17862 16532 17868 16544
rect 17920 16532 17926 16584
rect 22732 16575 22790 16581
rect 18432 16544 22094 16572
rect 18432 16504 18460 16544
rect 17144 16476 18460 16504
rect 18509 16507 18567 16513
rect 18509 16473 18521 16507
rect 18555 16504 18567 16507
rect 19334 16504 19340 16516
rect 18555 16476 19340 16504
rect 18555 16473 18567 16476
rect 18509 16467 18567 16473
rect 19334 16464 19340 16476
rect 19392 16464 19398 16516
rect 19512 16507 19570 16513
rect 19512 16473 19524 16507
rect 19558 16473 19570 16507
rect 19512 16467 19570 16473
rect 15764 16408 16528 16436
rect 19058 16396 19064 16448
rect 19116 16436 19122 16448
rect 19527 16436 19555 16467
rect 19886 16464 19892 16516
rect 19944 16504 19950 16516
rect 20070 16504 20076 16516
rect 19944 16476 20076 16504
rect 19944 16464 19950 16476
rect 20070 16464 20076 16476
rect 20128 16464 20134 16516
rect 22066 16504 22094 16544
rect 22732 16541 22744 16575
rect 22778 16572 22790 16575
rect 23842 16572 23848 16584
rect 22778 16544 23848 16572
rect 22778 16541 22790 16544
rect 22732 16535 22790 16541
rect 23842 16532 23848 16544
rect 23900 16532 23906 16584
rect 24673 16575 24731 16581
rect 24673 16541 24685 16575
rect 24719 16566 24731 16575
rect 24854 16572 24860 16584
rect 24773 16566 24860 16572
rect 24719 16544 24860 16566
rect 24719 16541 24801 16544
rect 24673 16538 24801 16541
rect 24673 16535 24731 16538
rect 24854 16532 24860 16544
rect 24912 16532 24918 16584
rect 26878 16572 26884 16584
rect 26839 16544 26884 16572
rect 26878 16532 26884 16544
rect 26936 16532 26942 16584
rect 27062 16532 27068 16584
rect 27120 16572 27126 16584
rect 27157 16575 27215 16581
rect 27157 16572 27169 16575
rect 27120 16544 27169 16572
rect 27120 16532 27126 16544
rect 27157 16541 27169 16544
rect 27203 16541 27215 16575
rect 27157 16535 27215 16541
rect 27614 16532 27620 16584
rect 27672 16572 27678 16584
rect 27709 16575 27767 16581
rect 27709 16572 27721 16575
rect 27672 16544 27721 16572
rect 27672 16532 27678 16544
rect 27709 16541 27721 16544
rect 27755 16541 27767 16575
rect 27709 16535 27767 16541
rect 28902 16532 28908 16584
rect 28960 16572 28966 16584
rect 32324 16581 32352 16612
rect 32490 16600 32496 16612
rect 32548 16600 32554 16652
rect 34698 16640 34704 16652
rect 34659 16612 34704 16640
rect 34698 16600 34704 16612
rect 34756 16600 34762 16652
rect 36280 16640 36308 16736
rect 47762 16708 47768 16720
rect 46308 16680 47768 16708
rect 36909 16643 36967 16649
rect 36909 16640 36921 16643
rect 36280 16612 36921 16640
rect 36909 16609 36921 16612
rect 36955 16609 36967 16643
rect 38562 16640 38568 16652
rect 38523 16612 38568 16640
rect 36909 16603 36967 16609
rect 38562 16600 38568 16612
rect 38620 16600 38626 16652
rect 46308 16649 46336 16680
rect 47762 16668 47768 16680
rect 47820 16668 47826 16720
rect 46293 16643 46351 16649
rect 46293 16609 46305 16643
rect 46339 16609 46351 16643
rect 46474 16640 46480 16652
rect 46435 16612 46480 16640
rect 46293 16603 46351 16609
rect 46474 16600 46480 16612
rect 46532 16600 46538 16652
rect 48130 16640 48136 16652
rect 48091 16612 48136 16640
rect 48130 16600 48136 16612
rect 48188 16600 48194 16652
rect 32217 16575 32275 16581
rect 32217 16572 32229 16575
rect 28960 16544 32229 16572
rect 28960 16532 28966 16544
rect 32217 16541 32229 16544
rect 32263 16541 32275 16575
rect 32217 16535 32275 16541
rect 32309 16575 32367 16581
rect 32309 16541 32321 16575
rect 32355 16541 32367 16575
rect 32309 16535 32367 16541
rect 32401 16575 32459 16581
rect 32401 16541 32413 16575
rect 32447 16541 32459 16575
rect 32401 16535 32459 16541
rect 32585 16575 32643 16581
rect 32585 16541 32597 16575
rect 32631 16572 32643 16575
rect 32766 16572 32772 16584
rect 32631 16544 32772 16572
rect 32631 16541 32643 16544
rect 32585 16535 32643 16541
rect 23934 16504 23940 16516
rect 22066 16476 23940 16504
rect 23934 16464 23940 16476
rect 23992 16464 23998 16516
rect 24210 16464 24216 16516
rect 24268 16504 24274 16516
rect 24394 16504 24400 16516
rect 24268 16476 24400 16504
rect 24268 16464 24274 16476
rect 24394 16464 24400 16476
rect 24452 16464 24458 16516
rect 24486 16464 24492 16516
rect 24544 16504 24550 16516
rect 24581 16507 24639 16513
rect 24581 16504 24593 16507
rect 24544 16476 24593 16504
rect 24544 16464 24550 16476
rect 24581 16473 24593 16476
rect 24627 16473 24639 16507
rect 24581 16467 24639 16473
rect 19116 16408 19555 16436
rect 19116 16396 19122 16408
rect 23106 16396 23112 16448
rect 23164 16436 23170 16448
rect 23658 16436 23664 16448
rect 23164 16408 23664 16436
rect 23164 16396 23170 16408
rect 23658 16396 23664 16408
rect 23716 16396 23722 16448
rect 25498 16396 25504 16448
rect 25556 16436 25562 16448
rect 26142 16436 26148 16448
rect 25556 16408 26148 16436
rect 25556 16396 25562 16408
rect 26142 16396 26148 16408
rect 26200 16436 26206 16448
rect 27065 16439 27123 16445
rect 27065 16436 27077 16439
rect 26200 16408 27077 16436
rect 26200 16396 26206 16408
rect 27065 16405 27077 16408
rect 27111 16405 27123 16439
rect 27065 16399 27123 16405
rect 27154 16396 27160 16448
rect 27212 16436 27218 16448
rect 27893 16439 27951 16445
rect 27893 16436 27905 16439
rect 27212 16408 27905 16436
rect 27212 16396 27218 16408
rect 27893 16405 27905 16408
rect 27939 16405 27951 16439
rect 31938 16436 31944 16448
rect 31899 16408 31944 16436
rect 27893 16399 27951 16405
rect 31938 16396 31944 16408
rect 31996 16396 32002 16448
rect 32416 16436 32444 16535
rect 32766 16532 32772 16544
rect 32824 16532 32830 16584
rect 32858 16532 32864 16584
rect 32916 16572 32922 16584
rect 33229 16575 33287 16581
rect 33229 16572 33241 16575
rect 32916 16544 33241 16572
rect 32916 16532 32922 16544
rect 33229 16541 33241 16544
rect 33275 16541 33287 16575
rect 33229 16535 33287 16541
rect 34790 16532 34796 16584
rect 34848 16572 34854 16584
rect 34957 16575 35015 16581
rect 34957 16572 34969 16575
rect 34848 16544 34969 16572
rect 34848 16532 34854 16544
rect 34957 16541 34969 16544
rect 35003 16541 35015 16575
rect 34957 16535 35015 16541
rect 33045 16507 33103 16513
rect 33045 16473 33057 16507
rect 33091 16504 33103 16507
rect 33134 16504 33140 16516
rect 33091 16476 33140 16504
rect 33091 16473 33103 16476
rect 33045 16467 33103 16473
rect 33134 16464 33140 16476
rect 33192 16464 33198 16516
rect 37093 16507 37151 16513
rect 37093 16473 37105 16507
rect 37139 16504 37151 16507
rect 37366 16504 37372 16516
rect 37139 16476 37372 16504
rect 37139 16473 37151 16476
rect 37093 16467 37151 16473
rect 37366 16464 37372 16476
rect 37424 16464 37430 16516
rect 33413 16439 33471 16445
rect 33413 16436 33425 16439
rect 32416 16408 33425 16436
rect 33413 16405 33425 16408
rect 33459 16405 33471 16439
rect 33413 16399 33471 16405
rect 1104 16346 48852 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 48852 16346
rect 1104 16272 48852 16294
rect 10134 16232 10140 16244
rect 10095 16204 10140 16232
rect 10134 16192 10140 16204
rect 10192 16192 10198 16244
rect 13722 16232 13728 16244
rect 13683 16204 13728 16232
rect 13722 16192 13728 16204
rect 13780 16192 13786 16244
rect 17221 16235 17279 16241
rect 17221 16201 17233 16235
rect 17267 16232 17279 16235
rect 17310 16232 17316 16244
rect 17267 16204 17316 16232
rect 17267 16201 17279 16204
rect 17221 16195 17279 16201
rect 17310 16192 17316 16204
rect 17368 16192 17374 16244
rect 17862 16232 17868 16244
rect 17823 16204 17868 16232
rect 17862 16192 17868 16204
rect 17920 16192 17926 16244
rect 18969 16235 19027 16241
rect 18969 16201 18981 16235
rect 19015 16232 19027 16235
rect 19058 16232 19064 16244
rect 19015 16204 19064 16232
rect 19015 16201 19027 16204
rect 18969 16195 19027 16201
rect 19058 16192 19064 16204
rect 19116 16192 19122 16244
rect 20070 16232 20076 16244
rect 19352 16204 20076 16232
rect 2222 16164 2228 16176
rect 2183 16136 2228 16164
rect 2222 16124 2228 16136
rect 2280 16124 2286 16176
rect 12434 16164 12440 16176
rect 12360 16136 12440 16164
rect 2038 16096 2044 16108
rect 1999 16068 2044 16096
rect 2038 16056 2044 16068
rect 2096 16056 2102 16108
rect 9674 16056 9680 16108
rect 9732 16096 9738 16108
rect 12360 16105 12388 16136
rect 12434 16124 12440 16136
rect 12492 16124 12498 16176
rect 12612 16167 12670 16173
rect 12612 16133 12624 16167
rect 12658 16164 12670 16167
rect 15654 16164 15660 16176
rect 12658 16136 15660 16164
rect 12658 16133 12670 16136
rect 12612 16127 12670 16133
rect 15654 16124 15660 16136
rect 15712 16124 15718 16176
rect 17037 16167 17095 16173
rect 17037 16133 17049 16167
rect 17083 16164 17095 16167
rect 18322 16164 18328 16176
rect 17083 16136 18328 16164
rect 17083 16133 17095 16136
rect 17037 16127 17095 16133
rect 18322 16124 18328 16136
rect 18380 16124 18386 16176
rect 10045 16099 10103 16105
rect 10045 16096 10057 16099
rect 9732 16068 10057 16096
rect 9732 16056 9738 16068
rect 10045 16065 10057 16068
rect 10091 16065 10103 16099
rect 10045 16059 10103 16065
rect 12345 16099 12403 16105
rect 12345 16065 12357 16099
rect 12391 16065 12403 16099
rect 14458 16096 14464 16108
rect 14371 16068 14464 16096
rect 12345 16059 12403 16065
rect 14458 16056 14464 16068
rect 14516 16096 14522 16108
rect 14826 16096 14832 16108
rect 14516 16068 14832 16096
rect 14516 16056 14522 16068
rect 14826 16056 14832 16068
rect 14884 16096 14890 16108
rect 16390 16096 16396 16108
rect 14884 16068 16396 16096
rect 14884 16056 14890 16068
rect 16390 16056 16396 16068
rect 16448 16056 16454 16108
rect 16853 16099 16911 16105
rect 16853 16065 16865 16099
rect 16899 16096 16911 16099
rect 17310 16096 17316 16108
rect 16899 16068 17316 16096
rect 16899 16065 16911 16068
rect 16853 16059 16911 16065
rect 17310 16056 17316 16068
rect 17368 16056 17374 16108
rect 17681 16099 17739 16105
rect 17681 16065 17693 16099
rect 17727 16096 17739 16099
rect 17862 16096 17868 16108
rect 17727 16068 17868 16096
rect 17727 16065 17739 16068
rect 17681 16059 17739 16065
rect 17862 16056 17868 16068
rect 17920 16056 17926 16108
rect 18414 16056 18420 16108
rect 18472 16096 18478 16108
rect 19352 16105 19380 16204
rect 20070 16192 20076 16204
rect 20128 16192 20134 16244
rect 20898 16232 20904 16244
rect 20859 16204 20904 16232
rect 20898 16192 20904 16204
rect 20956 16232 20962 16244
rect 21266 16232 21272 16244
rect 20956 16204 21272 16232
rect 20956 16192 20962 16204
rect 21266 16192 21272 16204
rect 21324 16192 21330 16244
rect 23750 16192 23756 16244
rect 23808 16232 23814 16244
rect 24765 16235 24823 16241
rect 24765 16232 24777 16235
rect 23808 16204 24777 16232
rect 23808 16192 23814 16204
rect 24765 16201 24777 16204
rect 24811 16201 24823 16235
rect 26694 16232 26700 16244
rect 24765 16195 24823 16201
rect 25056 16204 26700 16232
rect 19978 16164 19984 16176
rect 19444 16136 19984 16164
rect 19444 16105 19472 16136
rect 19978 16124 19984 16136
rect 20036 16124 20042 16176
rect 24305 16167 24363 16173
rect 24305 16133 24317 16167
rect 24351 16164 24363 16167
rect 24946 16164 24952 16176
rect 24351 16136 24952 16164
rect 24351 16133 24363 16136
rect 24305 16127 24363 16133
rect 24946 16124 24952 16136
rect 25004 16124 25010 16176
rect 19245 16099 19303 16105
rect 19245 16096 19257 16099
rect 18472 16068 19257 16096
rect 18472 16056 18478 16068
rect 19245 16065 19257 16068
rect 19291 16065 19303 16099
rect 19245 16059 19303 16065
rect 19337 16099 19395 16105
rect 19337 16065 19349 16099
rect 19383 16065 19395 16099
rect 19337 16059 19395 16065
rect 19429 16099 19487 16105
rect 19429 16065 19441 16099
rect 19475 16065 19487 16099
rect 19429 16059 19487 16065
rect 19518 16056 19524 16108
rect 19576 16096 19582 16108
rect 19613 16099 19671 16105
rect 19613 16096 19625 16099
rect 19576 16068 19625 16096
rect 19576 16056 19582 16068
rect 19613 16065 19625 16068
rect 19659 16096 19671 16099
rect 20346 16096 20352 16108
rect 19659 16068 20352 16096
rect 19659 16065 19671 16068
rect 19613 16059 19671 16065
rect 20346 16056 20352 16068
rect 20404 16056 20410 16108
rect 20714 16096 20720 16108
rect 20675 16068 20720 16096
rect 20714 16056 20720 16068
rect 20772 16096 20778 16108
rect 22278 16096 22284 16108
rect 20772 16068 22284 16096
rect 20772 16056 20778 16068
rect 22278 16056 22284 16068
rect 22336 16056 22342 16108
rect 24581 16099 24639 16105
rect 24581 16065 24593 16099
rect 24627 16096 24639 16099
rect 24762 16096 24768 16108
rect 24627 16068 24768 16096
rect 24627 16065 24639 16068
rect 24581 16059 24639 16065
rect 24762 16056 24768 16068
rect 24820 16056 24826 16108
rect 2774 15988 2780 16040
rect 2832 16028 2838 16040
rect 14182 16028 14188 16040
rect 2832 16000 2877 16028
rect 14095 16000 14188 16028
rect 2832 15988 2838 16000
rect 14182 15988 14188 16000
rect 14240 16028 14246 16040
rect 20070 16028 20076 16040
rect 14240 16000 20076 16028
rect 14240 15988 14246 16000
rect 20070 15988 20076 16000
rect 20128 16028 20134 16040
rect 21450 16028 21456 16040
rect 20128 16000 21456 16028
rect 20128 15988 20134 16000
rect 21450 15988 21456 16000
rect 21508 15988 21514 16040
rect 24486 16028 24492 16040
rect 24447 16000 24492 16028
rect 24486 15988 24492 16000
rect 24544 15988 24550 16040
rect 25056 16028 25084 16204
rect 26694 16192 26700 16204
rect 26752 16232 26758 16244
rect 31018 16232 31024 16244
rect 26752 16204 31024 16232
rect 26752 16192 26758 16204
rect 31018 16192 31024 16204
rect 31076 16192 31082 16244
rect 28537 16167 28595 16173
rect 28537 16133 28549 16167
rect 28583 16164 28595 16167
rect 30285 16167 30343 16173
rect 30285 16164 30297 16167
rect 28583 16136 30297 16164
rect 28583 16133 28595 16136
rect 28537 16127 28595 16133
rect 30285 16133 30297 16136
rect 30331 16164 30343 16167
rect 30374 16164 30380 16176
rect 30331 16136 30380 16164
rect 30331 16133 30343 16136
rect 30285 16127 30343 16133
rect 30374 16124 30380 16136
rect 30432 16124 30438 16176
rect 31938 16124 31944 16176
rect 31996 16164 32002 16176
rect 32370 16167 32428 16173
rect 32370 16164 32382 16167
rect 31996 16136 32382 16164
rect 31996 16124 32002 16136
rect 32370 16133 32382 16136
rect 32416 16133 32428 16167
rect 32370 16127 32428 16133
rect 27246 16096 27252 16108
rect 27207 16068 27252 16096
rect 27246 16056 27252 16068
rect 27304 16056 27310 16108
rect 28350 16096 28356 16108
rect 28311 16068 28356 16096
rect 28350 16056 28356 16068
rect 28408 16056 28414 16108
rect 28994 16096 29000 16108
rect 28955 16068 29000 16096
rect 28994 16056 29000 16068
rect 29052 16056 29058 16108
rect 29086 16056 29092 16108
rect 29144 16096 29150 16108
rect 29181 16099 29239 16105
rect 29181 16096 29193 16099
rect 29144 16068 29193 16096
rect 29144 16056 29150 16068
rect 29181 16065 29193 16068
rect 29227 16065 29239 16099
rect 29546 16096 29552 16108
rect 29459 16068 29552 16096
rect 29181 16059 29239 16065
rect 29546 16056 29552 16068
rect 29604 16096 29610 16108
rect 30834 16096 30840 16108
rect 29604 16068 30840 16096
rect 29604 16056 29610 16068
rect 30834 16056 30840 16068
rect 30892 16056 30898 16108
rect 32125 16099 32183 16105
rect 32125 16065 32137 16099
rect 32171 16096 32183 16099
rect 32950 16096 32956 16108
rect 32171 16068 32956 16096
rect 32171 16065 32183 16068
rect 32125 16059 32183 16065
rect 32950 16056 32956 16068
rect 33008 16056 33014 16108
rect 47578 16096 47584 16108
rect 47539 16068 47584 16096
rect 47578 16056 47584 16068
rect 47636 16056 47642 16108
rect 24596 16000 25084 16028
rect 27525 16031 27583 16037
rect 17862 15920 17868 15972
rect 17920 15960 17926 15972
rect 24596 15960 24624 16000
rect 27525 15997 27537 16031
rect 27571 15997 27583 16031
rect 27525 15991 27583 15997
rect 29273 16031 29331 16037
rect 29273 15997 29285 16031
rect 29319 15997 29331 16031
rect 29273 15991 29331 15997
rect 29365 16031 29423 16037
rect 29365 15997 29377 16031
rect 29411 16028 29423 16031
rect 29638 16028 29644 16040
rect 29411 16000 29644 16028
rect 29411 15997 29423 16000
rect 29365 15991 29423 15997
rect 24854 15960 24860 15972
rect 17920 15932 24624 15960
rect 24688 15932 24860 15960
rect 17920 15920 17926 15932
rect 24581 15895 24639 15901
rect 24581 15861 24593 15895
rect 24627 15892 24639 15895
rect 24688 15892 24716 15932
rect 24854 15920 24860 15932
rect 24912 15920 24918 15972
rect 27540 15960 27568 15991
rect 25056 15932 27568 15960
rect 29288 15960 29316 15991
rect 29638 15988 29644 16000
rect 29696 15988 29702 16040
rect 30466 15960 30472 15972
rect 29288 15932 30472 15960
rect 25056 15904 25084 15932
rect 30466 15920 30472 15932
rect 30524 15920 30530 15972
rect 24627 15864 24716 15892
rect 24627 15861 24639 15864
rect 24581 15855 24639 15861
rect 24762 15852 24768 15904
rect 24820 15892 24826 15904
rect 25038 15892 25044 15904
rect 24820 15864 25044 15892
rect 24820 15852 24826 15864
rect 25038 15852 25044 15864
rect 25096 15852 25102 15904
rect 27338 15892 27344 15904
rect 27299 15864 27344 15892
rect 27338 15852 27344 15864
rect 27396 15852 27402 15904
rect 27433 15895 27491 15901
rect 27433 15861 27445 15895
rect 27479 15892 27491 15895
rect 27890 15892 27896 15904
rect 27479 15864 27896 15892
rect 27479 15861 27491 15864
rect 27433 15855 27491 15861
rect 27890 15852 27896 15864
rect 27948 15852 27954 15904
rect 29730 15892 29736 15904
rect 29691 15864 29736 15892
rect 29730 15852 29736 15864
rect 29788 15852 29794 15904
rect 29822 15852 29828 15904
rect 29880 15892 29886 15904
rect 30377 15895 30435 15901
rect 30377 15892 30389 15895
rect 29880 15864 30389 15892
rect 29880 15852 29886 15864
rect 30377 15861 30389 15864
rect 30423 15861 30435 15895
rect 30377 15855 30435 15861
rect 32858 15852 32864 15904
rect 32916 15892 32922 15904
rect 33505 15895 33563 15901
rect 33505 15892 33517 15895
rect 32916 15864 33517 15892
rect 32916 15852 32922 15864
rect 33505 15861 33517 15864
rect 33551 15861 33563 15895
rect 47026 15892 47032 15904
rect 46987 15864 47032 15892
rect 33505 15855 33563 15861
rect 47026 15852 47032 15864
rect 47084 15852 47090 15904
rect 47670 15892 47676 15904
rect 47631 15864 47676 15892
rect 47670 15852 47676 15864
rect 47728 15852 47734 15904
rect 1104 15802 48852 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 48852 15802
rect 1104 15728 48852 15750
rect 15194 15688 15200 15700
rect 15107 15660 15200 15688
rect 15194 15648 15200 15660
rect 15252 15688 15258 15700
rect 17310 15688 17316 15700
rect 15252 15660 17316 15688
rect 15252 15648 15258 15660
rect 17310 15648 17316 15660
rect 17368 15648 17374 15700
rect 20346 15648 20352 15700
rect 20404 15688 20410 15700
rect 24765 15691 24823 15697
rect 20404 15660 21128 15688
rect 20404 15648 20410 15660
rect 1670 15580 1676 15632
rect 1728 15620 1734 15632
rect 21100 15620 21128 15660
rect 24765 15657 24777 15691
rect 24811 15688 24823 15691
rect 24946 15688 24952 15700
rect 24811 15660 24952 15688
rect 24811 15657 24823 15660
rect 24765 15651 24823 15657
rect 24946 15648 24952 15660
rect 25004 15648 25010 15700
rect 26237 15691 26295 15697
rect 26237 15657 26249 15691
rect 26283 15688 26295 15691
rect 27338 15688 27344 15700
rect 26283 15660 27344 15688
rect 26283 15657 26295 15660
rect 26237 15651 26295 15657
rect 27338 15648 27344 15660
rect 27396 15688 27402 15700
rect 27982 15688 27988 15700
rect 27396 15660 27988 15688
rect 27396 15648 27402 15660
rect 27982 15648 27988 15660
rect 28040 15688 28046 15700
rect 28261 15691 28319 15697
rect 28261 15688 28273 15691
rect 28040 15660 28273 15688
rect 28040 15648 28046 15660
rect 28261 15657 28273 15660
rect 28307 15657 28319 15691
rect 28261 15651 28319 15657
rect 30006 15648 30012 15700
rect 30064 15688 30070 15700
rect 30064 15660 33824 15688
rect 30064 15648 30070 15660
rect 1728 15592 20852 15620
rect 21100 15592 21220 15620
rect 1728 15580 1734 15592
rect 9217 15555 9275 15561
rect 9217 15521 9229 15555
rect 9263 15552 9275 15555
rect 9582 15552 9588 15564
rect 9263 15524 9588 15552
rect 9263 15521 9275 15524
rect 9217 15515 9275 15521
rect 9582 15512 9588 15524
rect 9640 15512 9646 15564
rect 10962 15552 10968 15564
rect 10923 15524 10968 15552
rect 10962 15512 10968 15524
rect 11020 15512 11026 15564
rect 11514 15552 11520 15564
rect 11475 15524 11520 15552
rect 11514 15512 11520 15524
rect 11572 15512 11578 15564
rect 13786 15524 14780 15552
rect 9398 15416 9404 15428
rect 9359 15388 9404 15416
rect 9398 15376 9404 15388
rect 9456 15376 9462 15428
rect 11698 15416 11704 15428
rect 11659 15388 11704 15416
rect 11698 15376 11704 15388
rect 11756 15376 11762 15428
rect 13262 15376 13268 15428
rect 13320 15416 13326 15428
rect 13357 15419 13415 15425
rect 13357 15416 13369 15419
rect 13320 15388 13369 15416
rect 13320 15376 13326 15388
rect 13357 15385 13369 15388
rect 13403 15385 13415 15419
rect 13357 15379 13415 15385
rect 10226 15308 10232 15360
rect 10284 15348 10290 15360
rect 13786 15348 13814 15524
rect 14274 15444 14280 15496
rect 14332 15493 14338 15496
rect 14332 15487 14381 15493
rect 14553 15487 14611 15493
rect 14332 15453 14335 15487
rect 14369 15453 14381 15487
rect 14332 15447 14381 15453
rect 14458 15481 14516 15487
rect 14458 15474 14470 15481
rect 14504 15474 14516 15481
rect 14332 15444 14338 15447
rect 14458 15422 14464 15474
rect 14516 15422 14522 15474
rect 14553 15453 14565 15487
rect 14599 15484 14611 15487
rect 14642 15484 14648 15496
rect 14599 15456 14648 15484
rect 14599 15453 14611 15456
rect 14553 15447 14611 15453
rect 14642 15444 14648 15456
rect 14700 15444 14706 15496
rect 14752 15493 14780 15524
rect 16390 15512 16396 15564
rect 16448 15552 16454 15564
rect 17681 15555 17739 15561
rect 17681 15552 17693 15555
rect 16448 15524 16617 15552
rect 16448 15512 16454 15524
rect 14737 15487 14795 15493
rect 14737 15453 14749 15487
rect 14783 15453 14795 15487
rect 14737 15447 14795 15453
rect 14752 15416 14780 15447
rect 15286 15444 15292 15496
rect 15344 15484 15350 15496
rect 15381 15487 15439 15493
rect 15381 15484 15393 15487
rect 15344 15456 15393 15484
rect 15344 15444 15350 15456
rect 15381 15453 15393 15456
rect 15427 15453 15439 15487
rect 16482 15484 16488 15496
rect 16443 15456 16488 15484
rect 15381 15447 15439 15453
rect 16482 15444 16488 15456
rect 16540 15444 16546 15496
rect 16589 15493 16617 15524
rect 16776 15524 17693 15552
rect 16574 15487 16632 15493
rect 16574 15453 16586 15487
rect 16620 15453 16632 15487
rect 16574 15447 16632 15453
rect 16690 15487 16748 15493
rect 16690 15453 16702 15487
rect 16736 15484 16748 15487
rect 16776 15484 16804 15524
rect 17681 15521 17693 15524
rect 17727 15521 17739 15555
rect 17681 15515 17739 15521
rect 19245 15555 19303 15561
rect 19245 15521 19257 15555
rect 19291 15552 19303 15555
rect 20714 15552 20720 15564
rect 19291 15524 20720 15552
rect 19291 15521 19303 15524
rect 19245 15515 19303 15521
rect 20714 15512 20720 15524
rect 20772 15512 20778 15564
rect 16736 15456 16804 15484
rect 16853 15487 16911 15493
rect 16736 15453 16748 15456
rect 16690 15447 16748 15453
rect 16853 15453 16865 15487
rect 16899 15484 16911 15487
rect 18417 15487 18475 15493
rect 18417 15484 18429 15487
rect 16899 15456 18429 15484
rect 16899 15453 16911 15456
rect 16853 15447 16911 15453
rect 18417 15453 18429 15456
rect 18463 15453 18475 15487
rect 19518 15484 19524 15496
rect 19479 15456 19524 15484
rect 18417 15447 18475 15453
rect 16868 15416 16896 15447
rect 19518 15444 19524 15456
rect 19576 15444 19582 15496
rect 20824 15493 20852 15592
rect 21192 15493 21220 15592
rect 26142 15580 26148 15632
rect 26200 15620 26206 15632
rect 27111 15623 27169 15629
rect 27111 15620 27123 15623
rect 26200 15592 27123 15620
rect 26200 15580 26206 15592
rect 27111 15589 27123 15592
rect 27157 15589 27169 15623
rect 27111 15583 27169 15589
rect 28626 15580 28632 15632
rect 28684 15620 28690 15632
rect 28684 15592 28856 15620
rect 28684 15580 28690 15592
rect 24118 15512 24124 15564
rect 24176 15552 24182 15564
rect 26421 15555 26479 15561
rect 24176 15524 25176 15552
rect 24176 15512 24182 15524
rect 20809 15487 20867 15493
rect 20993 15487 21051 15493
rect 20809 15453 20821 15487
rect 20855 15453 20867 15487
rect 20809 15447 20867 15453
rect 20898 15481 20956 15487
rect 20898 15474 20910 15481
rect 20944 15474 20956 15481
rect 17310 15416 17316 15428
rect 14752 15388 16896 15416
rect 17271 15388 17316 15416
rect 17310 15376 17316 15388
rect 17368 15376 17374 15428
rect 17494 15416 17500 15428
rect 17455 15388 17500 15416
rect 17494 15376 17500 15388
rect 17552 15376 17558 15428
rect 17862 15376 17868 15428
rect 17920 15416 17926 15428
rect 18233 15419 18291 15425
rect 20898 15422 20904 15474
rect 20956 15422 20962 15474
rect 20993 15453 21005 15487
rect 21039 15453 21051 15487
rect 20993 15447 21051 15453
rect 21177 15487 21235 15493
rect 21177 15453 21189 15487
rect 21223 15453 21235 15487
rect 21177 15447 21235 15453
rect 21637 15487 21695 15493
rect 21637 15453 21649 15487
rect 21683 15484 21695 15487
rect 21910 15484 21916 15496
rect 21683 15456 21916 15484
rect 21683 15453 21695 15456
rect 21637 15447 21695 15453
rect 18233 15416 18245 15419
rect 17920 15388 18245 15416
rect 17920 15376 17926 15388
rect 18233 15385 18245 15388
rect 18279 15385 18291 15419
rect 21008 15416 21036 15447
rect 21910 15444 21916 15456
rect 21968 15444 21974 15496
rect 23658 15444 23664 15496
rect 23716 15484 23722 15496
rect 24673 15487 24731 15493
rect 24673 15484 24685 15487
rect 23716 15456 24685 15484
rect 23716 15444 23722 15456
rect 24673 15453 24685 15456
rect 24719 15484 24731 15487
rect 24762 15484 24768 15496
rect 24719 15456 24768 15484
rect 24719 15453 24731 15456
rect 24673 15447 24731 15453
rect 24762 15444 24768 15456
rect 24820 15444 24826 15496
rect 24857 15487 24915 15493
rect 24857 15453 24869 15487
rect 24903 15453 24915 15487
rect 24857 15447 24915 15453
rect 21542 15416 21548 15428
rect 21008 15388 21548 15416
rect 18233 15379 18291 15385
rect 21542 15376 21548 15388
rect 21600 15376 21606 15428
rect 21818 15416 21824 15428
rect 21779 15388 21824 15416
rect 21818 15376 21824 15388
rect 21876 15376 21882 15428
rect 24486 15376 24492 15428
rect 24544 15416 24550 15428
rect 24872 15416 24900 15447
rect 24946 15444 24952 15496
rect 25004 15484 25010 15496
rect 25148 15493 25176 15524
rect 26421 15521 26433 15555
rect 26467 15552 26479 15555
rect 27522 15552 27528 15564
rect 26467 15524 27528 15552
rect 26467 15521 26479 15524
rect 26421 15515 26479 15521
rect 27522 15512 27528 15524
rect 27580 15512 27586 15564
rect 28828 15561 28856 15592
rect 28813 15555 28871 15561
rect 28813 15521 28825 15555
rect 28859 15552 28871 15555
rect 29454 15552 29460 15564
rect 28859 15524 29460 15552
rect 28859 15521 28871 15524
rect 28813 15515 28871 15521
rect 29454 15512 29460 15524
rect 29512 15512 29518 15564
rect 29730 15512 29736 15564
rect 29788 15552 29794 15564
rect 29788 15524 29960 15552
rect 29788 15512 29794 15524
rect 25133 15487 25191 15493
rect 25004 15456 25049 15484
rect 25004 15444 25010 15456
rect 25133 15453 25145 15487
rect 25179 15453 25191 15487
rect 25133 15447 25191 15453
rect 26145 15487 26203 15493
rect 26145 15453 26157 15487
rect 26191 15484 26203 15487
rect 26510 15484 26516 15496
rect 26191 15456 26516 15484
rect 26191 15453 26203 15456
rect 26145 15447 26203 15453
rect 26510 15444 26516 15456
rect 26568 15444 26574 15496
rect 26878 15484 26884 15496
rect 26839 15456 26884 15484
rect 26878 15444 26884 15456
rect 26936 15444 26942 15496
rect 27062 15444 27068 15496
rect 27120 15484 27126 15496
rect 29822 15484 29828 15496
rect 27120 15456 28672 15484
rect 29783 15456 29828 15484
rect 27120 15444 27126 15456
rect 27798 15416 27804 15428
rect 24544 15388 27804 15416
rect 24544 15376 24550 15388
rect 27798 15376 27804 15388
rect 27856 15376 27862 15428
rect 28644 15425 28672 15456
rect 29822 15444 29828 15456
rect 29880 15444 29886 15496
rect 29932 15484 29960 15524
rect 30081 15487 30139 15493
rect 30081 15484 30093 15487
rect 29932 15456 30093 15484
rect 30081 15453 30093 15456
rect 30127 15453 30139 15487
rect 30081 15447 30139 15453
rect 30374 15444 30380 15496
rect 30432 15484 30438 15496
rect 32493 15487 32551 15493
rect 32493 15484 32505 15487
rect 30432 15456 32505 15484
rect 30432 15444 30438 15456
rect 32493 15453 32505 15456
rect 32539 15453 32551 15487
rect 33796 15484 33824 15660
rect 47118 15620 47124 15632
rect 46308 15592 47124 15620
rect 46308 15561 46336 15592
rect 47118 15580 47124 15592
rect 47176 15580 47182 15632
rect 46293 15555 46351 15561
rect 46293 15521 46305 15555
rect 46339 15521 46351 15555
rect 46293 15515 46351 15521
rect 46477 15555 46535 15561
rect 46477 15521 46489 15555
rect 46523 15552 46535 15555
rect 47670 15552 47676 15564
rect 46523 15524 47676 15552
rect 46523 15521 46535 15524
rect 46477 15515 46535 15521
rect 47670 15512 47676 15524
rect 47728 15512 47734 15564
rect 48130 15552 48136 15564
rect 48091 15524 48136 15552
rect 48130 15512 48136 15524
rect 48188 15512 48194 15564
rect 34514 15484 34520 15496
rect 33796 15456 34520 15484
rect 32493 15447 32551 15453
rect 34514 15444 34520 15456
rect 34572 15484 34578 15496
rect 34977 15487 35035 15493
rect 34977 15484 34989 15487
rect 34572 15456 34989 15484
rect 34572 15444 34578 15456
rect 34977 15453 34989 15456
rect 35023 15453 35035 15487
rect 34977 15447 35035 15453
rect 28629 15419 28687 15425
rect 28629 15385 28641 15419
rect 28675 15416 28687 15419
rect 29546 15416 29552 15428
rect 28675 15388 29552 15416
rect 28675 15385 28687 15388
rect 28629 15379 28687 15385
rect 29546 15376 29552 15388
rect 29604 15376 29610 15428
rect 31018 15376 31024 15428
rect 31076 15416 31082 15428
rect 31757 15419 31815 15425
rect 31757 15416 31769 15419
rect 31076 15388 31769 15416
rect 31076 15376 31082 15388
rect 31757 15385 31769 15388
rect 31803 15385 31815 15419
rect 31757 15379 31815 15385
rect 32677 15419 32735 15425
rect 32677 15385 32689 15419
rect 32723 15416 32735 15419
rect 32950 15416 32956 15428
rect 32723 15388 32956 15416
rect 32723 15385 32735 15388
rect 32677 15379 32735 15385
rect 32950 15376 32956 15388
rect 33008 15376 33014 15428
rect 35161 15419 35219 15425
rect 35161 15385 35173 15419
rect 35207 15416 35219 15419
rect 36538 15416 36544 15428
rect 35207 15388 36544 15416
rect 35207 15385 35219 15388
rect 35161 15379 35219 15385
rect 36538 15376 36544 15388
rect 36596 15376 36602 15428
rect 14090 15348 14096 15360
rect 10284 15320 13814 15348
rect 14051 15320 14096 15348
rect 10284 15308 10290 15320
rect 14090 15308 14096 15320
rect 14148 15308 14154 15360
rect 16209 15351 16267 15357
rect 16209 15317 16221 15351
rect 16255 15348 16267 15351
rect 16942 15348 16948 15360
rect 16255 15320 16948 15348
rect 16255 15317 16267 15320
rect 16209 15311 16267 15317
rect 16942 15308 16948 15320
rect 17000 15308 17006 15360
rect 17218 15308 17224 15360
rect 17276 15348 17282 15360
rect 17880 15348 17908 15376
rect 17276 15320 17908 15348
rect 20533 15351 20591 15357
rect 17276 15308 17282 15320
rect 20533 15317 20545 15351
rect 20579 15348 20591 15351
rect 20898 15348 20904 15360
rect 20579 15320 20904 15348
rect 20579 15317 20591 15320
rect 20533 15311 20591 15317
rect 20898 15308 20904 15320
rect 20956 15308 20962 15360
rect 22002 15348 22008 15360
rect 21963 15320 22008 15348
rect 22002 15308 22008 15320
rect 22060 15308 22066 15360
rect 24394 15348 24400 15360
rect 24355 15320 24400 15348
rect 24394 15308 24400 15320
rect 24452 15308 24458 15360
rect 26418 15348 26424 15360
rect 26379 15320 26424 15348
rect 26418 15308 26424 15320
rect 26476 15308 26482 15360
rect 26510 15308 26516 15360
rect 26568 15348 26574 15360
rect 27246 15348 27252 15360
rect 26568 15320 27252 15348
rect 26568 15308 26574 15320
rect 27246 15308 27252 15320
rect 27304 15308 27310 15360
rect 28721 15351 28779 15357
rect 28721 15317 28733 15351
rect 28767 15348 28779 15351
rect 30466 15348 30472 15360
rect 28767 15320 30472 15348
rect 28767 15317 28779 15320
rect 28721 15311 28779 15317
rect 30466 15308 30472 15320
rect 30524 15348 30530 15360
rect 31205 15351 31263 15357
rect 31205 15348 31217 15351
rect 30524 15320 31217 15348
rect 30524 15308 30530 15320
rect 31205 15317 31217 15320
rect 31251 15317 31263 15351
rect 31205 15311 31263 15317
rect 31849 15351 31907 15357
rect 31849 15317 31861 15351
rect 31895 15348 31907 15351
rect 32766 15348 32772 15360
rect 31895 15320 32772 15348
rect 31895 15317 31907 15320
rect 31849 15311 31907 15317
rect 32766 15308 32772 15320
rect 32824 15348 32830 15360
rect 33134 15348 33140 15360
rect 32824 15320 33140 15348
rect 32824 15308 32830 15320
rect 33134 15308 33140 15320
rect 33192 15308 33198 15360
rect 35345 15351 35403 15357
rect 35345 15317 35357 15351
rect 35391 15348 35403 15351
rect 35618 15348 35624 15360
rect 35391 15320 35624 15348
rect 35391 15317 35403 15320
rect 35345 15311 35403 15317
rect 35618 15308 35624 15320
rect 35676 15308 35682 15360
rect 1104 15258 48852 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 48852 15258
rect 1104 15184 48852 15206
rect 9398 15104 9404 15156
rect 9456 15144 9462 15156
rect 9585 15147 9643 15153
rect 9585 15144 9597 15147
rect 9456 15116 9597 15144
rect 9456 15104 9462 15116
rect 9585 15113 9597 15116
rect 9631 15113 9643 15147
rect 9585 15107 9643 15113
rect 10597 15147 10655 15153
rect 10597 15113 10609 15147
rect 10643 15144 10655 15147
rect 11698 15144 11704 15156
rect 10643 15116 11704 15144
rect 10643 15113 10655 15116
rect 10597 15107 10655 15113
rect 11698 15104 11704 15116
rect 11756 15104 11762 15156
rect 13722 15104 13728 15156
rect 13780 15144 13786 15156
rect 14553 15147 14611 15153
rect 13780 15116 14412 15144
rect 13780 15104 13786 15116
rect 7926 15036 7932 15088
rect 7984 15076 7990 15088
rect 14274 15076 14280 15088
rect 7984 15048 10548 15076
rect 7984 15036 7990 15048
rect 9493 15011 9551 15017
rect 9493 14977 9505 15011
rect 9539 15008 9551 15011
rect 9674 15008 9680 15020
rect 9539 14980 9680 15008
rect 9539 14977 9551 14980
rect 9493 14971 9551 14977
rect 9674 14968 9680 14980
rect 9732 14968 9738 15020
rect 10520 15017 10548 15048
rect 12360 15048 14280 15076
rect 12360 15017 12388 15048
rect 14274 15036 14280 15048
rect 14332 15036 14338 15088
rect 14384 15085 14412 15116
rect 14553 15113 14565 15147
rect 14599 15144 14611 15147
rect 14642 15144 14648 15156
rect 14599 15116 14648 15144
rect 14599 15113 14611 15116
rect 14553 15107 14611 15113
rect 14642 15104 14648 15116
rect 14700 15104 14706 15156
rect 17494 15104 17500 15156
rect 17552 15144 17558 15156
rect 18049 15147 18107 15153
rect 18049 15144 18061 15147
rect 17552 15116 18061 15144
rect 17552 15104 17558 15116
rect 18049 15113 18061 15116
rect 18095 15113 18107 15147
rect 18049 15107 18107 15113
rect 21542 15104 21548 15156
rect 21600 15144 21606 15156
rect 22189 15147 22247 15153
rect 22189 15144 22201 15147
rect 21600 15116 22201 15144
rect 21600 15104 21606 15116
rect 22189 15113 22201 15116
rect 22235 15113 22247 15147
rect 22189 15107 22247 15113
rect 25498 15104 25504 15156
rect 25556 15144 25562 15156
rect 25869 15147 25927 15153
rect 25869 15144 25881 15147
rect 25556 15116 25881 15144
rect 25556 15104 25562 15116
rect 25869 15113 25881 15116
rect 25915 15113 25927 15147
rect 25869 15107 25927 15113
rect 26234 15104 26240 15156
rect 26292 15144 26298 15156
rect 27154 15144 27160 15156
rect 26292 15116 27160 15144
rect 26292 15104 26298 15116
rect 27154 15104 27160 15116
rect 27212 15144 27218 15156
rect 27522 15144 27528 15156
rect 27212 15116 27384 15144
rect 27483 15116 27528 15144
rect 27212 15104 27218 15116
rect 16942 15085 16948 15088
rect 14369 15079 14427 15085
rect 14369 15045 14381 15079
rect 14415 15045 14427 15079
rect 16936 15076 16948 15085
rect 16903 15048 16948 15076
rect 14369 15039 14427 15045
rect 16936 15039 16948 15048
rect 16942 15036 16948 15039
rect 17000 15036 17006 15088
rect 27062 15076 27068 15088
rect 22020 15048 27068 15076
rect 10505 15011 10563 15017
rect 10505 14977 10517 15011
rect 10551 14977 10563 15011
rect 10505 14971 10563 14977
rect 12345 15011 12403 15017
rect 12345 14977 12357 15011
rect 12391 14977 12403 15011
rect 12345 14971 12403 14977
rect 12612 15011 12670 15017
rect 12612 14977 12624 15011
rect 12658 15008 12670 15011
rect 14090 15008 14096 15020
rect 12658 14980 14096 15008
rect 12658 14977 12670 14980
rect 12612 14971 12670 14977
rect 14090 14968 14096 14980
rect 14148 14968 14154 15020
rect 14185 15011 14243 15017
rect 14185 14977 14197 15011
rect 14231 14977 14243 15011
rect 14292 15006 14320 15036
rect 16666 15008 16672 15020
rect 14384 15006 16672 15008
rect 14292 14980 16672 15006
rect 14292 14978 14412 14980
rect 14185 14971 14243 14977
rect 14200 14940 14228 14971
rect 16666 14968 16672 14980
rect 16724 14968 16730 15020
rect 17954 14968 17960 15020
rect 18012 15008 18018 15020
rect 18509 15011 18567 15017
rect 18509 15008 18521 15011
rect 18012 14980 18521 15008
rect 18012 14968 18018 14980
rect 18509 14977 18521 14980
rect 18555 15008 18567 15011
rect 18598 15008 18604 15020
rect 18555 14980 18604 15008
rect 18555 14977 18567 14980
rect 18509 14971 18567 14977
rect 18598 14968 18604 14980
rect 18656 14968 18662 15020
rect 19426 14968 19432 15020
rect 19484 15008 19490 15020
rect 19886 15008 19892 15020
rect 19484 14980 19892 15008
rect 19484 14968 19490 14980
rect 19886 14968 19892 14980
rect 19944 14968 19950 15020
rect 19978 14968 19984 15020
rect 20036 15008 20042 15020
rect 20145 15011 20203 15017
rect 20145 15008 20157 15011
rect 20036 14980 20157 15008
rect 20036 14968 20042 14980
rect 20145 14977 20157 14980
rect 20191 14977 20203 15011
rect 20145 14971 20203 14977
rect 21821 15011 21879 15017
rect 21821 14977 21833 15011
rect 21867 15008 21879 15011
rect 21910 15008 21916 15020
rect 21867 14980 21916 15008
rect 21867 14977 21879 14980
rect 21821 14971 21879 14977
rect 21910 14968 21916 14980
rect 21968 14968 21974 15020
rect 22020 15017 22048 15048
rect 27062 15036 27068 15048
rect 27120 15036 27126 15088
rect 27356 15076 27384 15116
rect 27522 15104 27528 15116
rect 27580 15104 27586 15156
rect 27798 15104 27804 15156
rect 27856 15144 27862 15156
rect 27893 15147 27951 15153
rect 27893 15144 27905 15147
rect 27856 15116 27905 15144
rect 27856 15104 27862 15116
rect 27893 15113 27905 15116
rect 27939 15144 27951 15147
rect 28902 15144 28908 15156
rect 27939 15116 28908 15144
rect 27939 15113 27951 15116
rect 27893 15107 27951 15113
rect 28902 15104 28908 15116
rect 28960 15104 28966 15156
rect 30834 15144 30840 15156
rect 29288 15116 30840 15144
rect 28718 15076 28724 15088
rect 27356 15048 28724 15076
rect 28718 15036 28724 15048
rect 28776 15036 28782 15088
rect 22005 15011 22063 15017
rect 22005 14977 22017 15011
rect 22051 15008 22063 15011
rect 22186 15008 22192 15020
rect 22051 14980 22192 15008
rect 22051 14977 22063 14980
rect 22005 14971 22063 14977
rect 22186 14968 22192 14980
rect 22244 14968 22250 15020
rect 22278 14968 22284 15020
rect 22336 15008 22342 15020
rect 22649 15011 22707 15017
rect 22649 15008 22661 15011
rect 22336 14980 22661 15008
rect 22336 14968 22342 14980
rect 22649 14977 22661 14980
rect 22695 14977 22707 15011
rect 26050 15008 26056 15020
rect 26011 14980 26056 15008
rect 22649 14971 22707 14977
rect 26050 14968 26056 14980
rect 26108 14968 26114 15020
rect 26145 15011 26203 15017
rect 26145 14977 26157 15011
rect 26191 15008 26203 15011
rect 26418 15008 26424 15020
rect 26191 14980 26424 15008
rect 26191 14977 26203 14980
rect 26145 14971 26203 14977
rect 26418 14968 26424 14980
rect 26476 14968 26482 15020
rect 26602 14968 26608 15020
rect 26660 15008 26666 15020
rect 27798 15008 27804 15020
rect 26660 14980 27804 15008
rect 26660 14968 26666 14980
rect 27798 14968 27804 14980
rect 27856 14968 27862 15020
rect 27985 15011 28043 15017
rect 27985 14977 27997 15011
rect 28031 15008 28043 15011
rect 29178 15008 29184 15020
rect 28031 14980 29184 15008
rect 28031 14977 28043 14980
rect 27985 14971 28043 14977
rect 15194 14940 15200 14952
rect 14200 14912 15200 14940
rect 15194 14900 15200 14912
rect 15252 14900 15258 14952
rect 20990 14900 20996 14952
rect 21048 14940 21054 14952
rect 26234 14940 26240 14952
rect 21048 14912 26004 14940
rect 26195 14912 26240 14940
rect 21048 14900 21054 14912
rect 21269 14875 21327 14881
rect 21269 14841 21281 14875
rect 21315 14872 21327 14875
rect 21818 14872 21824 14884
rect 21315 14844 21824 14872
rect 21315 14841 21327 14844
rect 21269 14835 21327 14841
rect 21818 14832 21824 14844
rect 21876 14872 21882 14884
rect 21876 14844 22094 14872
rect 21876 14832 21882 14844
rect 13722 14804 13728 14816
rect 13683 14776 13728 14804
rect 13722 14764 13728 14776
rect 13780 14764 13786 14816
rect 18598 14804 18604 14816
rect 18559 14776 18604 14804
rect 18598 14764 18604 14776
rect 18656 14764 18662 14816
rect 22066 14804 22094 14844
rect 22462 14832 22468 14884
rect 22520 14872 22526 14884
rect 22833 14875 22891 14881
rect 22833 14872 22845 14875
rect 22520 14844 22845 14872
rect 22520 14832 22526 14844
rect 22833 14841 22845 14844
rect 22879 14872 22891 14875
rect 25976 14872 26004 14912
rect 26234 14900 26240 14912
rect 26292 14900 26298 14952
rect 26326 14900 26332 14952
rect 26384 14940 26390 14952
rect 26384 14912 26429 14940
rect 26384 14900 26390 14912
rect 26510 14900 26516 14952
rect 26568 14940 26574 14952
rect 28000 14940 28028 14971
rect 29178 14968 29184 14980
rect 29236 14968 29242 15020
rect 29288 15017 29316 15116
rect 30834 15104 30840 15116
rect 30892 15104 30898 15156
rect 30926 15104 30932 15156
rect 30984 15144 30990 15156
rect 30984 15116 31029 15144
rect 30984 15104 30990 15116
rect 31110 15104 31116 15156
rect 31168 15144 31174 15156
rect 31168 15116 41414 15144
rect 31168 15104 31174 15116
rect 30466 15076 30472 15088
rect 30427 15048 30472 15076
rect 30466 15036 30472 15048
rect 30524 15036 30530 15088
rect 41386 15076 41414 15116
rect 47946 15104 47952 15156
rect 48004 15144 48010 15156
rect 48041 15147 48099 15153
rect 48041 15144 48053 15147
rect 48004 15116 48053 15144
rect 48004 15104 48010 15116
rect 48041 15113 48053 15116
rect 48087 15113 48099 15147
rect 48041 15107 48099 15113
rect 47854 15076 47860 15088
rect 30576 15048 32536 15076
rect 41386 15048 47860 15076
rect 29273 15011 29331 15017
rect 29273 14977 29285 15011
rect 29319 14977 29331 15011
rect 29457 15011 29515 15017
rect 29457 15008 29469 15011
rect 29273 14971 29331 14977
rect 29380 14980 29469 15008
rect 26568 14912 28028 14940
rect 28169 14943 28227 14949
rect 26568 14900 26574 14912
rect 28169 14909 28181 14943
rect 28215 14940 28227 14943
rect 28626 14940 28632 14952
rect 28215 14912 28632 14940
rect 28215 14909 28227 14912
rect 28169 14903 28227 14909
rect 28626 14900 28632 14912
rect 28684 14900 28690 14952
rect 29086 14900 29092 14952
rect 29144 14940 29150 14952
rect 29380 14940 29408 14980
rect 29457 14977 29469 14980
rect 29503 14977 29515 15011
rect 29457 14971 29515 14977
rect 29825 15011 29883 15017
rect 29825 14977 29837 15011
rect 29871 15008 29883 15011
rect 30576 15008 30604 15048
rect 32508 15020 32536 15048
rect 47854 15036 47860 15048
rect 47912 15036 47918 15088
rect 29871 14980 30604 15008
rect 29871 14977 29883 14980
rect 29825 14971 29883 14977
rect 29546 14940 29552 14952
rect 29144 14912 29408 14940
rect 29507 14912 29552 14940
rect 29144 14900 29150 14912
rect 29546 14900 29552 14912
rect 29604 14900 29610 14952
rect 29638 14900 29644 14952
rect 29696 14940 29702 14952
rect 29696 14912 29741 14940
rect 29696 14900 29702 14912
rect 29730 14872 29736 14884
rect 22879 14844 25912 14872
rect 25976 14844 29736 14872
rect 22879 14841 22891 14844
rect 22833 14835 22891 14841
rect 25130 14804 25136 14816
rect 22066 14776 25136 14804
rect 25130 14764 25136 14776
rect 25188 14764 25194 14816
rect 25884 14804 25912 14844
rect 29730 14832 29736 14844
rect 29788 14832 29794 14884
rect 26786 14804 26792 14816
rect 25884 14776 26792 14804
rect 26786 14764 26792 14776
rect 26844 14764 26850 14816
rect 26970 14764 26976 14816
rect 27028 14804 27034 14816
rect 27614 14804 27620 14816
rect 27028 14776 27620 14804
rect 27028 14764 27034 14776
rect 27614 14764 27620 14776
rect 27672 14764 27678 14816
rect 29270 14764 29276 14816
rect 29328 14804 29334 14816
rect 29840 14804 29868 14971
rect 30650 14968 30656 15020
rect 30708 15008 30714 15020
rect 30745 15011 30803 15017
rect 30745 15008 30757 15011
rect 30708 14980 30757 15008
rect 30708 14968 30714 14980
rect 30745 14977 30757 14980
rect 30791 14977 30803 15011
rect 30745 14971 30803 14977
rect 32490 14968 32496 15020
rect 32548 15008 32554 15020
rect 32677 15011 32735 15017
rect 32677 15008 32689 15011
rect 32548 14980 32689 15008
rect 32548 14968 32554 14980
rect 32677 14977 32689 14980
rect 32723 14977 32735 15011
rect 32677 14971 32735 14977
rect 32782 15011 32840 15017
rect 32782 14977 32794 15011
rect 32828 14977 32840 15011
rect 32782 14971 32840 14977
rect 32882 15011 32940 15017
rect 32882 14977 32894 15011
rect 32928 15008 32940 15011
rect 33045 15011 33103 15017
rect 32928 14980 32996 15008
rect 32928 14977 32940 14980
rect 32882 14971 32940 14977
rect 30282 14900 30288 14952
rect 30340 14940 30346 14952
rect 30561 14943 30619 14949
rect 30561 14940 30573 14943
rect 30340 14912 30573 14940
rect 30340 14900 30346 14912
rect 30561 14909 30573 14912
rect 30607 14909 30619 14943
rect 30561 14903 30619 14909
rect 31662 14900 31668 14952
rect 31720 14940 31726 14952
rect 32214 14940 32220 14952
rect 31720 14912 32220 14940
rect 31720 14900 31726 14912
rect 32214 14900 32220 14912
rect 32272 14900 32278 14952
rect 32582 14900 32588 14952
rect 32640 14940 32646 14952
rect 32784 14940 32812 14971
rect 32640 14912 32812 14940
rect 32640 14900 32646 14912
rect 32306 14832 32312 14884
rect 32364 14872 32370 14884
rect 32364 14844 32628 14872
rect 32364 14832 32370 14844
rect 29328 14776 29868 14804
rect 30009 14807 30067 14813
rect 29328 14764 29334 14776
rect 30009 14773 30021 14807
rect 30055 14804 30067 14807
rect 30098 14804 30104 14816
rect 30055 14776 30104 14804
rect 30055 14773 30067 14776
rect 30009 14767 30067 14773
rect 30098 14764 30104 14776
rect 30156 14764 30162 14816
rect 30374 14764 30380 14816
rect 30432 14804 30438 14816
rect 30469 14807 30527 14813
rect 30469 14804 30481 14807
rect 30432 14776 30481 14804
rect 30432 14764 30438 14776
rect 30469 14773 30481 14776
rect 30515 14773 30527 14807
rect 30469 14767 30527 14773
rect 32401 14807 32459 14813
rect 32401 14773 32413 14807
rect 32447 14804 32459 14807
rect 32490 14804 32496 14816
rect 32447 14776 32496 14804
rect 32447 14773 32459 14776
rect 32401 14767 32459 14773
rect 32490 14764 32496 14776
rect 32548 14764 32554 14816
rect 32600 14804 32628 14844
rect 32968 14804 32996 14980
rect 33045 14977 33057 15011
rect 33091 15008 33103 15011
rect 33134 15008 33140 15020
rect 33091 14980 33140 15008
rect 33091 14977 33103 14980
rect 33045 14971 33103 14977
rect 33134 14968 33140 14980
rect 33192 14968 33198 15020
rect 35434 15017 35440 15020
rect 35428 14971 35440 15017
rect 35492 15008 35498 15020
rect 35492 14980 35528 15008
rect 35434 14968 35440 14971
rect 35492 14968 35498 14980
rect 43530 14968 43536 15020
rect 43588 15008 43594 15020
rect 46845 15011 46903 15017
rect 46845 15008 46857 15011
rect 43588 14980 46857 15008
rect 43588 14968 43594 14980
rect 46845 14977 46857 14980
rect 46891 15008 46903 15011
rect 47578 15008 47584 15020
rect 46891 14980 47584 15008
rect 46891 14977 46903 14980
rect 46845 14971 46903 14977
rect 47578 14968 47584 14980
rect 47636 14968 47642 15020
rect 47946 15008 47952 15020
rect 47907 14980 47952 15008
rect 47946 14968 47952 14980
rect 48004 14968 48010 15020
rect 34606 14900 34612 14952
rect 34664 14940 34670 14952
rect 35161 14943 35219 14949
rect 35161 14940 35173 14943
rect 34664 14912 35173 14940
rect 34664 14900 34670 14912
rect 35161 14909 35173 14912
rect 35207 14909 35219 14943
rect 35161 14903 35219 14909
rect 36538 14804 36544 14816
rect 32600 14776 32996 14804
rect 36499 14776 36544 14804
rect 36538 14764 36544 14776
rect 36596 14764 36602 14816
rect 46474 14764 46480 14816
rect 46532 14804 46538 14816
rect 46937 14807 46995 14813
rect 46937 14804 46949 14807
rect 46532 14776 46949 14804
rect 46532 14764 46538 14776
rect 46937 14773 46949 14776
rect 46983 14773 46995 14807
rect 46937 14767 46995 14773
rect 1104 14714 48852 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 48852 14714
rect 1104 14640 48852 14662
rect 19334 14560 19340 14612
rect 19392 14600 19398 14612
rect 19392 14572 22876 14600
rect 19392 14560 19398 14572
rect 3142 14492 3148 14544
rect 3200 14532 3206 14544
rect 19705 14535 19763 14541
rect 3200 14504 18644 14532
rect 3200 14492 3206 14504
rect 9674 14424 9680 14476
rect 9732 14464 9738 14476
rect 12526 14464 12532 14476
rect 9732 14436 12532 14464
rect 9732 14424 9738 14436
rect 12452 14405 12480 14436
rect 12526 14424 12532 14436
rect 12584 14464 12590 14476
rect 17954 14464 17960 14476
rect 12584 14436 17960 14464
rect 12584 14424 12590 14436
rect 17954 14424 17960 14436
rect 18012 14424 18018 14476
rect 12437 14399 12495 14405
rect 12437 14365 12449 14399
rect 12483 14396 12495 14399
rect 14737 14399 14795 14405
rect 12483 14368 12517 14396
rect 12483 14365 12495 14368
rect 12437 14359 12495 14365
rect 14737 14365 14749 14399
rect 14783 14365 14795 14399
rect 14918 14396 14924 14408
rect 14879 14368 14924 14396
rect 14737 14359 14795 14365
rect 14752 14328 14780 14359
rect 14918 14356 14924 14368
rect 14976 14356 14982 14408
rect 18506 14396 18512 14408
rect 18467 14368 18512 14396
rect 18506 14356 18512 14368
rect 18564 14356 18570 14408
rect 18616 14396 18644 14504
rect 19705 14501 19717 14535
rect 19751 14532 19763 14535
rect 19978 14532 19984 14544
rect 19751 14504 19984 14532
rect 19751 14501 19763 14504
rect 19705 14495 19763 14501
rect 19978 14492 19984 14504
rect 20036 14492 20042 14544
rect 22186 14532 22192 14544
rect 22147 14504 22192 14532
rect 22186 14492 22192 14504
rect 22244 14492 22250 14544
rect 19886 14424 19892 14476
rect 19944 14464 19950 14476
rect 20809 14467 20867 14473
rect 20809 14464 20821 14467
rect 19944 14436 20821 14464
rect 19944 14424 19950 14436
rect 20809 14433 20821 14436
rect 20855 14433 20867 14467
rect 20809 14427 20867 14433
rect 19981 14399 20039 14405
rect 19981 14396 19993 14399
rect 18616 14368 19993 14396
rect 19981 14365 19993 14368
rect 20027 14365 20039 14399
rect 19981 14359 20039 14365
rect 20073 14399 20131 14405
rect 20073 14365 20085 14399
rect 20119 14365 20131 14399
rect 20073 14359 20131 14365
rect 20165 14399 20223 14405
rect 20165 14365 20177 14399
rect 20211 14365 20223 14399
rect 20346 14396 20352 14408
rect 20307 14368 20352 14396
rect 20165 14359 20223 14365
rect 15194 14328 15200 14340
rect 14752 14300 15200 14328
rect 15194 14288 15200 14300
rect 15252 14288 15258 14340
rect 18690 14328 18696 14340
rect 18651 14300 18696 14328
rect 18690 14288 18696 14300
rect 18748 14288 18754 14340
rect 12529 14263 12587 14269
rect 12529 14229 12541 14263
rect 12575 14260 12587 14263
rect 12618 14260 12624 14272
rect 12575 14232 12624 14260
rect 12575 14229 12587 14232
rect 12529 14223 12587 14229
rect 12618 14220 12624 14232
rect 12676 14220 12682 14272
rect 14090 14220 14096 14272
rect 14148 14260 14154 14272
rect 14829 14263 14887 14269
rect 14829 14260 14841 14263
rect 14148 14232 14841 14260
rect 14148 14220 14154 14232
rect 14829 14229 14841 14232
rect 14875 14229 14887 14263
rect 20088 14260 20116 14359
rect 20180 14328 20208 14359
rect 20346 14356 20352 14368
rect 20404 14356 20410 14408
rect 20898 14356 20904 14408
rect 20956 14396 20962 14408
rect 21065 14399 21123 14405
rect 21065 14396 21077 14399
rect 20956 14368 21077 14396
rect 20956 14356 20962 14368
rect 21065 14365 21077 14368
rect 21111 14365 21123 14399
rect 22738 14396 22744 14408
rect 22699 14368 22744 14396
rect 21065 14359 21123 14365
rect 22738 14356 22744 14368
rect 22796 14356 22802 14408
rect 22002 14328 22008 14340
rect 20180 14300 22008 14328
rect 22002 14288 22008 14300
rect 22060 14288 22066 14340
rect 22848 14272 22876 14572
rect 23014 14560 23020 14612
rect 23072 14600 23078 14612
rect 27709 14603 27767 14609
rect 23072 14572 27108 14600
rect 23072 14560 23078 14572
rect 23474 14492 23480 14544
rect 23532 14532 23538 14544
rect 24762 14532 24768 14544
rect 23532 14504 24768 14532
rect 23532 14492 23538 14504
rect 24762 14492 24768 14504
rect 24820 14492 24826 14544
rect 26329 14535 26387 14541
rect 26329 14501 26341 14535
rect 26375 14532 26387 14535
rect 26510 14532 26516 14544
rect 26375 14504 26516 14532
rect 26375 14501 26387 14504
rect 26329 14495 26387 14501
rect 26510 14492 26516 14504
rect 26568 14492 26574 14544
rect 27080 14532 27108 14572
rect 27709 14569 27721 14603
rect 27755 14600 27767 14603
rect 28994 14600 29000 14612
rect 27755 14572 29000 14600
rect 27755 14569 27767 14572
rect 27709 14563 27767 14569
rect 28994 14560 29000 14572
rect 29052 14560 29058 14612
rect 29546 14560 29552 14612
rect 29604 14600 29610 14612
rect 30650 14600 30656 14612
rect 29604 14572 30656 14600
rect 29604 14560 29610 14572
rect 30650 14560 30656 14572
rect 30708 14600 30714 14612
rect 31389 14603 31447 14609
rect 31389 14600 31401 14603
rect 30708 14572 31401 14600
rect 30708 14560 30714 14572
rect 31389 14569 31401 14572
rect 31435 14569 31447 14603
rect 31389 14563 31447 14569
rect 35161 14603 35219 14609
rect 35161 14569 35173 14603
rect 35207 14600 35219 14603
rect 35434 14600 35440 14612
rect 35207 14572 35440 14600
rect 35207 14569 35219 14572
rect 35161 14563 35219 14569
rect 35434 14560 35440 14572
rect 35492 14560 35498 14612
rect 35526 14560 35532 14612
rect 35584 14600 35590 14612
rect 35584 14572 36676 14600
rect 35584 14560 35590 14572
rect 30006 14532 30012 14544
rect 27080 14504 30012 14532
rect 30006 14492 30012 14504
rect 30064 14492 30070 14544
rect 31938 14492 31944 14544
rect 31996 14532 32002 14544
rect 32674 14532 32680 14544
rect 31996 14504 32680 14532
rect 31996 14492 32002 14504
rect 32674 14492 32680 14504
rect 32732 14492 32738 14544
rect 34698 14532 34704 14544
rect 32784 14504 34704 14532
rect 29822 14464 29828 14476
rect 27172 14436 29828 14464
rect 23382 14356 23388 14408
rect 23440 14396 23446 14408
rect 24949 14399 25007 14405
rect 24949 14396 24961 14399
rect 23440 14368 24961 14396
rect 23440 14356 23446 14368
rect 24949 14365 24961 14368
rect 24995 14396 25007 14399
rect 27172 14396 27200 14436
rect 29822 14424 29828 14436
rect 29880 14424 29886 14476
rect 24995 14368 27200 14396
rect 27249 14399 27307 14405
rect 24995 14365 25007 14368
rect 24949 14359 25007 14365
rect 27249 14365 27261 14399
rect 27295 14396 27307 14399
rect 27614 14396 27620 14408
rect 27295 14368 27620 14396
rect 27295 14365 27307 14368
rect 27249 14359 27307 14365
rect 27614 14356 27620 14368
rect 27672 14356 27678 14408
rect 27890 14396 27896 14408
rect 27851 14368 27896 14396
rect 27890 14356 27896 14368
rect 27948 14356 27954 14408
rect 27982 14356 27988 14408
rect 28040 14396 28046 14408
rect 28169 14399 28227 14405
rect 28169 14396 28181 14399
rect 28040 14368 28181 14396
rect 28040 14356 28046 14368
rect 28169 14365 28181 14368
rect 28215 14365 28227 14399
rect 28902 14396 28908 14408
rect 28169 14359 28227 14365
rect 28644 14368 28908 14396
rect 25216 14331 25274 14337
rect 25216 14297 25228 14331
rect 25262 14328 25274 14331
rect 26142 14328 26148 14340
rect 25262 14300 26148 14328
rect 25262 14297 25274 14300
rect 25216 14291 25274 14297
rect 26142 14288 26148 14300
rect 26200 14288 26206 14340
rect 26970 14328 26976 14340
rect 26931 14300 26976 14328
rect 26970 14288 26976 14300
rect 27028 14288 27034 14340
rect 27632 14328 27660 14356
rect 28644 14337 28672 14368
rect 28902 14356 28908 14368
rect 28960 14356 28966 14408
rect 30006 14396 30012 14408
rect 29967 14368 30012 14396
rect 30006 14356 30012 14368
rect 30064 14356 30070 14408
rect 30098 14356 30104 14408
rect 30156 14396 30162 14408
rect 30265 14399 30323 14405
rect 30265 14396 30277 14399
rect 30156 14368 30277 14396
rect 30156 14356 30162 14368
rect 30265 14365 30277 14368
rect 30311 14365 30323 14399
rect 30265 14359 30323 14365
rect 30558 14356 30564 14408
rect 30616 14396 30622 14408
rect 32784 14405 32812 14504
rect 34698 14492 34704 14504
rect 34756 14492 34762 14544
rect 33965 14467 34023 14473
rect 33965 14464 33977 14467
rect 32968 14436 33977 14464
rect 32968 14405 32996 14436
rect 33965 14433 33977 14436
rect 34011 14433 34023 14467
rect 33965 14427 34023 14433
rect 34790 14424 34796 14476
rect 34848 14464 34854 14476
rect 34848 14436 35848 14464
rect 34848 14424 34854 14436
rect 32769 14399 32827 14405
rect 32769 14396 32781 14399
rect 30616 14368 32781 14396
rect 30616 14356 30622 14368
rect 32769 14365 32781 14368
rect 32815 14365 32827 14399
rect 32769 14359 32827 14365
rect 32861 14399 32919 14405
rect 32861 14365 32873 14399
rect 32907 14365 32919 14399
rect 32861 14359 32919 14365
rect 32953 14399 33011 14405
rect 32953 14365 32965 14399
rect 32999 14365 33011 14399
rect 33134 14396 33140 14408
rect 33095 14368 33140 14396
rect 32953 14359 33011 14365
rect 28629 14331 28687 14337
rect 28629 14328 28641 14331
rect 27632 14300 28641 14328
rect 28629 14297 28641 14300
rect 28675 14297 28687 14331
rect 28629 14291 28687 14297
rect 28718 14288 28724 14340
rect 28776 14328 28782 14340
rect 28813 14331 28871 14337
rect 28813 14328 28825 14331
rect 28776 14300 28825 14328
rect 28776 14288 28782 14300
rect 28813 14297 28825 14300
rect 28859 14297 28871 14331
rect 28813 14291 28871 14297
rect 32582 14288 32588 14340
rect 32640 14328 32646 14340
rect 32876 14328 32904 14359
rect 33134 14356 33140 14368
rect 33192 14356 33198 14408
rect 33778 14396 33784 14408
rect 33739 14368 33784 14396
rect 33778 14356 33784 14368
rect 33836 14356 33842 14408
rect 35342 14356 35348 14408
rect 35400 14405 35406 14408
rect 35400 14399 35449 14405
rect 35400 14365 35403 14399
rect 35437 14365 35449 14399
rect 35526 14396 35532 14408
rect 35487 14368 35532 14396
rect 35400 14359 35449 14365
rect 35400 14356 35406 14359
rect 35526 14356 35532 14368
rect 35584 14356 35590 14408
rect 35618 14356 35624 14408
rect 35676 14396 35682 14408
rect 35820 14405 35848 14436
rect 36648 14405 36676 14572
rect 47026 14532 47032 14544
rect 46308 14504 47032 14532
rect 46308 14473 46336 14504
rect 47026 14492 47032 14504
rect 47084 14492 47090 14544
rect 46293 14467 46351 14473
rect 46293 14433 46305 14467
rect 46339 14433 46351 14467
rect 46474 14464 46480 14476
rect 46435 14436 46480 14464
rect 46293 14427 46351 14433
rect 46474 14424 46480 14436
rect 46532 14424 46538 14476
rect 35805 14399 35863 14405
rect 35676 14368 35721 14396
rect 35676 14356 35682 14368
rect 35805 14365 35817 14399
rect 35851 14365 35863 14399
rect 36541 14399 36599 14405
rect 36541 14396 36553 14399
rect 35805 14359 35863 14365
rect 36464 14368 36553 14396
rect 32640 14300 32904 14328
rect 33597 14331 33655 14337
rect 32640 14288 32646 14300
rect 33597 14297 33609 14331
rect 33643 14297 33655 14331
rect 33597 14291 33655 14297
rect 20990 14260 20996 14272
rect 20088 14232 20996 14260
rect 14829 14223 14887 14229
rect 20990 14220 20996 14232
rect 21048 14220 21054 14272
rect 22830 14260 22836 14272
rect 22791 14232 22836 14260
rect 22830 14220 22836 14232
rect 22888 14220 22894 14272
rect 25130 14220 25136 14272
rect 25188 14260 25194 14272
rect 26602 14260 26608 14272
rect 25188 14232 26608 14260
rect 25188 14220 25194 14232
rect 26602 14220 26608 14232
rect 26660 14220 26666 14272
rect 27062 14260 27068 14272
rect 27120 14269 27126 14272
rect 27029 14232 27068 14260
rect 27062 14220 27068 14232
rect 27120 14223 27129 14269
rect 27157 14263 27215 14269
rect 27157 14229 27169 14263
rect 27203 14260 27215 14263
rect 27798 14260 27804 14272
rect 27203 14232 27804 14260
rect 27203 14229 27215 14232
rect 27157 14223 27215 14229
rect 27120 14220 27126 14223
rect 27798 14220 27804 14232
rect 27856 14220 27862 14272
rect 27890 14220 27896 14272
rect 27948 14260 27954 14272
rect 28077 14263 28135 14269
rect 28077 14260 28089 14263
rect 27948 14232 28089 14260
rect 27948 14220 27954 14232
rect 28077 14229 28089 14232
rect 28123 14260 28135 14263
rect 28997 14263 29055 14269
rect 28997 14260 29009 14263
rect 28123 14232 29009 14260
rect 28123 14229 28135 14232
rect 28077 14223 28135 14229
rect 28997 14229 29009 14232
rect 29043 14260 29055 14263
rect 30926 14260 30932 14272
rect 29043 14232 30932 14260
rect 29043 14229 29055 14232
rect 28997 14223 29055 14229
rect 30926 14220 30932 14232
rect 30984 14220 30990 14272
rect 32493 14263 32551 14269
rect 32493 14229 32505 14263
rect 32539 14260 32551 14263
rect 32674 14260 32680 14272
rect 32539 14232 32680 14260
rect 32539 14229 32551 14232
rect 32493 14223 32551 14229
rect 32674 14220 32680 14232
rect 32732 14220 32738 14272
rect 32766 14220 32772 14272
rect 32824 14260 32830 14272
rect 33612 14260 33640 14291
rect 35710 14288 35716 14340
rect 35768 14328 35774 14340
rect 35820 14328 35848 14359
rect 36464 14328 36492 14368
rect 36541 14365 36553 14368
rect 36587 14365 36599 14399
rect 36541 14359 36599 14365
rect 36630 14399 36688 14405
rect 36630 14365 36642 14399
rect 36676 14365 36688 14399
rect 36630 14359 36688 14365
rect 36722 14356 36728 14408
rect 36780 14396 36786 14408
rect 36780 14368 36825 14396
rect 36780 14356 36786 14368
rect 36906 14356 36912 14408
rect 36964 14396 36970 14408
rect 36964 14368 37009 14396
rect 36964 14356 36970 14368
rect 47210 14328 47216 14340
rect 35768 14300 36400 14328
rect 36464 14300 47216 14328
rect 35768 14288 35774 14300
rect 36262 14260 36268 14272
rect 32824 14232 33640 14260
rect 36223 14232 36268 14260
rect 32824 14220 32830 14232
rect 36262 14220 36268 14232
rect 36320 14220 36326 14272
rect 36372 14260 36400 14300
rect 47210 14288 47216 14300
rect 47268 14288 47274 14340
rect 48130 14328 48136 14340
rect 48091 14300 48136 14328
rect 48130 14288 48136 14300
rect 48188 14288 48194 14340
rect 36906 14260 36912 14272
rect 36372 14232 36912 14260
rect 36906 14220 36912 14232
rect 36964 14220 36970 14272
rect 36998 14220 37004 14272
rect 37056 14260 37062 14272
rect 43990 14260 43996 14272
rect 37056 14232 43996 14260
rect 37056 14220 37062 14232
rect 43990 14220 43996 14232
rect 44048 14220 44054 14272
rect 1104 14170 48852 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 48852 14170
rect 1104 14096 48852 14118
rect 13722 14056 13728 14068
rect 12452 14028 13728 14056
rect 14 13948 20 14000
rect 72 13988 78 14000
rect 72 13960 10088 13988
rect 72 13948 78 13960
rect 1670 13880 1676 13932
rect 1728 13920 1734 13932
rect 2041 13923 2099 13929
rect 2041 13920 2053 13923
rect 1728 13892 2053 13920
rect 1728 13880 1734 13892
rect 2041 13889 2053 13892
rect 2087 13920 2099 13923
rect 2130 13920 2136 13932
rect 2087 13892 2136 13920
rect 2087 13889 2099 13892
rect 2041 13883 2099 13889
rect 2130 13880 2136 13892
rect 2188 13880 2194 13932
rect 8110 13920 8116 13932
rect 8071 13892 8116 13920
rect 8110 13880 8116 13892
rect 8168 13880 8174 13932
rect 8294 13852 8300 13864
rect 8255 13824 8300 13852
rect 8294 13812 8300 13824
rect 8352 13812 8358 13864
rect 8573 13855 8631 13861
rect 8573 13821 8585 13855
rect 8619 13821 8631 13855
rect 10060 13852 10088 13960
rect 12452 13929 12480 14028
rect 13722 14016 13728 14028
rect 13780 14016 13786 14068
rect 16666 14016 16672 14068
rect 16724 14056 16730 14068
rect 16853 14059 16911 14065
rect 16853 14056 16865 14059
rect 16724 14028 16865 14056
rect 16724 14016 16730 14028
rect 16853 14025 16865 14028
rect 16899 14025 16911 14059
rect 16853 14019 16911 14025
rect 20533 14059 20591 14065
rect 20533 14025 20545 14059
rect 20579 14056 20591 14059
rect 20990 14056 20996 14068
rect 20579 14028 20996 14056
rect 20579 14025 20591 14028
rect 20533 14019 20591 14025
rect 20990 14016 20996 14028
rect 21048 14016 21054 14068
rect 21910 14016 21916 14068
rect 21968 14056 21974 14068
rect 22373 14059 22431 14065
rect 22373 14056 22385 14059
rect 21968 14028 22385 14056
rect 21968 14016 21974 14028
rect 22373 14025 22385 14028
rect 22419 14056 22431 14059
rect 23014 14056 23020 14068
rect 22419 14028 23020 14056
rect 22419 14025 22431 14028
rect 22373 14019 22431 14025
rect 23014 14016 23020 14028
rect 23072 14016 23078 14068
rect 25498 14056 25504 14068
rect 25459 14028 25504 14056
rect 25498 14016 25504 14028
rect 25556 14016 25562 14068
rect 26142 14056 26148 14068
rect 26103 14028 26148 14056
rect 26142 14016 26148 14028
rect 26200 14016 26206 14068
rect 27062 14016 27068 14068
rect 27120 14056 27126 14068
rect 27890 14056 27896 14068
rect 27120 14028 27896 14056
rect 27120 14016 27126 14028
rect 27890 14016 27896 14028
rect 27948 14016 27954 14068
rect 28350 14016 28356 14068
rect 28408 14056 28414 14068
rect 28902 14056 28908 14068
rect 28408 14028 28908 14056
rect 28408 14016 28414 14028
rect 28902 14016 28908 14028
rect 28960 14056 28966 14068
rect 30285 14059 30343 14065
rect 30285 14056 30297 14059
rect 28960 14028 30297 14056
rect 28960 14016 28966 14028
rect 30285 14025 30297 14028
rect 30331 14025 30343 14059
rect 30285 14019 30343 14025
rect 31573 14059 31631 14065
rect 31573 14025 31585 14059
rect 31619 14056 31631 14059
rect 32306 14056 32312 14068
rect 31619 14028 32312 14056
rect 31619 14025 31631 14028
rect 31573 14019 31631 14025
rect 32306 14016 32312 14028
rect 32364 14016 32370 14068
rect 32766 14056 32772 14068
rect 32508 14028 32772 14056
rect 12618 13988 12624 14000
rect 12579 13960 12624 13988
rect 12618 13948 12624 13960
rect 12676 13948 12682 14000
rect 13170 13948 13176 14000
rect 13228 13988 13234 14000
rect 15657 13991 15715 13997
rect 15657 13988 15669 13991
rect 13228 13960 14872 13988
rect 13228 13948 13234 13960
rect 14844 13929 14872 13960
rect 14936 13960 15669 13988
rect 14936 13932 14964 13960
rect 15657 13957 15669 13960
rect 15703 13957 15715 13991
rect 15657 13951 15715 13957
rect 16761 13991 16819 13997
rect 16761 13957 16773 13991
rect 16807 13988 16819 13991
rect 18690 13988 18696 14000
rect 16807 13960 18696 13988
rect 16807 13957 16819 13960
rect 16761 13951 16819 13957
rect 18690 13948 18696 13960
rect 18748 13948 18754 14000
rect 21358 13948 21364 14000
rect 21416 13988 21422 14000
rect 22281 13991 22339 13997
rect 22281 13988 22293 13991
rect 21416 13960 22293 13988
rect 21416 13948 21422 13960
rect 22281 13957 22293 13960
rect 22327 13957 22339 13991
rect 22281 13951 22339 13957
rect 22830 13948 22836 14000
rect 22888 13988 22894 14000
rect 30193 13991 30251 13997
rect 30193 13988 30205 13991
rect 22888 13960 30205 13988
rect 22888 13948 22894 13960
rect 30193 13957 30205 13960
rect 30239 13957 30251 13991
rect 30193 13951 30251 13957
rect 31205 13991 31263 13997
rect 31205 13957 31217 13991
rect 31251 13988 31263 13991
rect 32508 13988 32536 14028
rect 32766 14016 32772 14028
rect 32824 14016 32830 14068
rect 33778 14016 33784 14068
rect 33836 14056 33842 14068
rect 33965 14059 34023 14065
rect 33965 14056 33977 14059
rect 33836 14028 33977 14056
rect 33836 14016 33842 14028
rect 33965 14025 33977 14028
rect 34011 14025 34023 14059
rect 33965 14019 34023 14025
rect 47854 14016 47860 14068
rect 47912 14056 47918 14068
rect 48041 14059 48099 14065
rect 48041 14056 48053 14059
rect 47912 14028 48053 14056
rect 47912 14016 47918 14028
rect 48041 14025 48053 14028
rect 48087 14025 48099 14059
rect 48041 14019 48099 14025
rect 32950 13988 32956 14000
rect 31251 13960 32536 13988
rect 32600 13960 32956 13988
rect 31251 13957 31263 13960
rect 31205 13951 31263 13957
rect 12437 13923 12495 13929
rect 12437 13889 12449 13923
rect 12483 13889 12495 13923
rect 12437 13883 12495 13889
rect 14829 13923 14887 13929
rect 14829 13889 14841 13923
rect 14875 13889 14887 13923
rect 14829 13883 14887 13889
rect 14918 13880 14924 13932
rect 14976 13920 14982 13932
rect 14976 13892 15021 13920
rect 14976 13880 14982 13892
rect 15470 13880 15476 13932
rect 15528 13920 15534 13932
rect 15565 13923 15623 13929
rect 15565 13920 15577 13923
rect 15528 13892 15577 13920
rect 15528 13880 15534 13892
rect 15565 13889 15577 13892
rect 15611 13889 15623 13923
rect 15565 13883 15623 13889
rect 17494 13880 17500 13932
rect 17552 13920 17558 13932
rect 17773 13923 17831 13929
rect 17773 13920 17785 13923
rect 17552 13892 17785 13920
rect 17552 13880 17558 13892
rect 17773 13889 17785 13892
rect 17819 13889 17831 13923
rect 17773 13883 17831 13889
rect 20349 13923 20407 13929
rect 20349 13889 20361 13923
rect 20395 13920 20407 13923
rect 20622 13920 20628 13932
rect 20395 13892 20628 13920
rect 20395 13889 20407 13892
rect 20349 13883 20407 13889
rect 20622 13880 20628 13892
rect 20680 13880 20686 13932
rect 23382 13920 23388 13932
rect 23343 13892 23388 13920
rect 23382 13880 23388 13892
rect 23440 13880 23446 13932
rect 23652 13923 23710 13929
rect 23652 13889 23664 13923
rect 23698 13920 23710 13923
rect 24394 13920 24400 13932
rect 23698 13892 24400 13920
rect 23698 13889 23710 13892
rect 23652 13883 23710 13889
rect 24394 13880 24400 13892
rect 24452 13880 24458 13932
rect 25869 13923 25927 13929
rect 25869 13889 25881 13923
rect 25915 13920 25927 13923
rect 26510 13920 26516 13932
rect 25915 13892 26516 13920
rect 25915 13889 25927 13892
rect 25869 13883 25927 13889
rect 26510 13880 26516 13892
rect 26568 13880 26574 13932
rect 27522 13920 27528 13932
rect 27483 13892 27528 13920
rect 27522 13880 27528 13892
rect 27580 13880 27586 13932
rect 27798 13920 27804 13932
rect 27711 13892 27804 13920
rect 27798 13880 27804 13892
rect 27856 13920 27862 13932
rect 28718 13920 28724 13932
rect 27856 13892 28724 13920
rect 27856 13880 27862 13892
rect 28718 13880 28724 13892
rect 28776 13880 28782 13932
rect 29270 13920 29276 13932
rect 29231 13892 29276 13920
rect 29270 13880 29276 13892
rect 29328 13880 29334 13932
rect 29365 13923 29423 13929
rect 29365 13889 29377 13923
rect 29411 13920 29423 13923
rect 29546 13920 29552 13932
rect 29411 13892 29552 13920
rect 29411 13889 29423 13892
rect 29365 13883 29423 13889
rect 29546 13880 29552 13892
rect 29604 13880 29610 13932
rect 32600 13929 32628 13960
rect 32950 13948 32956 13960
rect 33008 13988 33014 14000
rect 34606 13988 34612 14000
rect 33008 13960 34612 13988
rect 33008 13948 33014 13960
rect 34606 13948 34612 13960
rect 34664 13988 34670 14000
rect 34790 13988 34796 14000
rect 34664 13960 34796 13988
rect 34664 13948 34670 13960
rect 34790 13948 34796 13960
rect 34848 13988 34854 14000
rect 35336 13991 35394 13997
rect 34848 13960 35112 13988
rect 34848 13948 34854 13960
rect 31389 13923 31447 13929
rect 31389 13889 31401 13923
rect 31435 13920 31447 13923
rect 32585 13923 32643 13929
rect 32585 13920 32597 13923
rect 31435 13892 32076 13920
rect 31435 13889 31447 13892
rect 31389 13883 31447 13889
rect 12897 13855 12955 13861
rect 12897 13852 12909 13855
rect 10060 13824 12434 13852
rect 8573 13815 8631 13821
rect 4062 13744 4068 13796
rect 4120 13784 4126 13796
rect 8588 13784 8616 13815
rect 4120 13756 8616 13784
rect 12406 13784 12434 13824
rect 12544 13824 12909 13852
rect 12544 13784 12572 13824
rect 12897 13821 12909 13824
rect 12943 13821 12955 13855
rect 12897 13815 12955 13821
rect 15105 13855 15163 13861
rect 15105 13821 15117 13855
rect 15151 13852 15163 13855
rect 15194 13852 15200 13864
rect 15151 13824 15200 13852
rect 15151 13821 15163 13824
rect 15105 13815 15163 13821
rect 15194 13812 15200 13824
rect 15252 13812 15258 13864
rect 17957 13855 18015 13861
rect 17957 13821 17969 13855
rect 18003 13852 18015 13855
rect 18598 13852 18604 13864
rect 18003 13824 18604 13852
rect 18003 13821 18015 13824
rect 17957 13815 18015 13821
rect 18598 13812 18604 13824
rect 18656 13812 18662 13864
rect 19426 13852 19432 13864
rect 19387 13824 19432 13852
rect 19426 13812 19432 13824
rect 19484 13812 19490 13864
rect 24762 13812 24768 13864
rect 24820 13852 24826 13864
rect 25961 13855 26019 13861
rect 25961 13852 25973 13855
rect 24820 13824 25973 13852
rect 24820 13812 24826 13824
rect 25961 13821 25973 13824
rect 26007 13821 26019 13855
rect 25961 13815 26019 13821
rect 26878 13812 26884 13864
rect 26936 13852 26942 13864
rect 27709 13855 27767 13861
rect 26936 13824 27660 13852
rect 26936 13812 26942 13824
rect 12406 13756 12572 13784
rect 27632 13784 27660 13824
rect 27709 13821 27721 13855
rect 27755 13852 27767 13855
rect 27982 13852 27988 13864
rect 27755 13824 27988 13852
rect 27755 13821 27767 13824
rect 27709 13815 27767 13821
rect 27982 13812 27988 13824
rect 28040 13812 28046 13864
rect 29454 13852 29460 13864
rect 29415 13824 29460 13852
rect 29454 13812 29460 13824
rect 29512 13812 29518 13864
rect 28905 13787 28963 13793
rect 27632 13756 28028 13784
rect 4120 13744 4126 13756
rect 1578 13676 1584 13728
rect 1636 13716 1642 13728
rect 2133 13719 2191 13725
rect 2133 13716 2145 13719
rect 1636 13688 2145 13716
rect 1636 13676 1642 13688
rect 2133 13685 2145 13688
rect 2179 13685 2191 13719
rect 2866 13716 2872 13728
rect 2827 13688 2872 13716
rect 2133 13679 2191 13685
rect 2866 13676 2872 13688
rect 2924 13676 2930 13728
rect 15010 13676 15016 13728
rect 15068 13716 15074 13728
rect 15068 13688 15113 13716
rect 15068 13676 15074 13688
rect 19702 13676 19708 13728
rect 19760 13716 19766 13728
rect 20070 13716 20076 13728
rect 19760 13688 20076 13716
rect 19760 13676 19766 13688
rect 20070 13676 20076 13688
rect 20128 13676 20134 13728
rect 24765 13719 24823 13725
rect 24765 13685 24777 13719
rect 24811 13716 24823 13719
rect 25222 13716 25228 13728
rect 24811 13688 25228 13716
rect 24811 13685 24823 13688
rect 24765 13679 24823 13685
rect 25222 13676 25228 13688
rect 25280 13676 25286 13728
rect 27522 13716 27528 13728
rect 27483 13688 27528 13716
rect 27522 13676 27528 13688
rect 27580 13676 27586 13728
rect 28000 13725 28028 13756
rect 28905 13753 28917 13787
rect 28951 13784 28963 13787
rect 28994 13784 29000 13796
rect 28951 13756 29000 13784
rect 28951 13753 28963 13756
rect 28905 13747 28963 13753
rect 28994 13744 29000 13756
rect 29052 13744 29058 13796
rect 31202 13744 31208 13796
rect 31260 13784 31266 13796
rect 31570 13784 31576 13796
rect 31260 13756 31576 13784
rect 31260 13744 31266 13756
rect 31570 13744 31576 13756
rect 31628 13744 31634 13796
rect 27985 13719 28043 13725
rect 27985 13685 27997 13719
rect 28031 13685 28043 13719
rect 32048 13716 32076 13892
rect 32505 13892 32597 13920
rect 32398 13812 32404 13864
rect 32456 13852 32462 13864
rect 32505 13852 32533 13892
rect 32585 13889 32597 13892
rect 32631 13889 32643 13923
rect 32585 13883 32643 13889
rect 32674 13880 32680 13932
rect 32732 13920 32738 13932
rect 35084 13929 35112 13960
rect 35336 13957 35348 13991
rect 35382 13988 35394 13991
rect 36262 13988 36268 14000
rect 35382 13960 36268 13988
rect 35382 13957 35394 13960
rect 35336 13951 35394 13957
rect 36262 13948 36268 13960
rect 36320 13948 36326 14000
rect 32841 13923 32899 13929
rect 32841 13920 32853 13923
rect 32732 13892 32853 13920
rect 32732 13880 32738 13892
rect 32841 13889 32853 13892
rect 32887 13889 32899 13923
rect 32841 13883 32899 13889
rect 35069 13923 35127 13929
rect 35069 13889 35081 13923
rect 35115 13889 35127 13923
rect 47854 13920 47860 13932
rect 47815 13892 47860 13920
rect 35069 13883 35127 13889
rect 47854 13880 47860 13892
rect 47912 13880 47918 13932
rect 32456 13824 32533 13852
rect 32456 13812 32462 13824
rect 32122 13744 32128 13796
rect 32180 13784 32186 13796
rect 32306 13784 32312 13796
rect 32180 13756 32312 13784
rect 32180 13744 32186 13756
rect 32306 13744 32312 13756
rect 32364 13744 32370 13796
rect 33594 13716 33600 13728
rect 32048 13688 33600 13716
rect 27985 13679 28043 13685
rect 33594 13676 33600 13688
rect 33652 13676 33658 13728
rect 34698 13676 34704 13728
rect 34756 13716 34762 13728
rect 36354 13716 36360 13728
rect 34756 13688 36360 13716
rect 34756 13676 34762 13688
rect 36354 13676 36360 13688
rect 36412 13716 36418 13728
rect 36449 13719 36507 13725
rect 36449 13716 36461 13719
rect 36412 13688 36461 13716
rect 36412 13676 36418 13688
rect 36449 13685 36461 13688
rect 36495 13685 36507 13719
rect 36449 13679 36507 13685
rect 1104 13626 48852 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 48852 13626
rect 1104 13552 48852 13574
rect 8294 13512 8300 13524
rect 8255 13484 8300 13512
rect 8294 13472 8300 13484
rect 8352 13472 8358 13524
rect 15562 13472 15568 13524
rect 15620 13512 15626 13524
rect 16025 13515 16083 13521
rect 16025 13512 16037 13515
rect 15620 13484 16037 13512
rect 15620 13472 15626 13484
rect 16025 13481 16037 13484
rect 16071 13481 16083 13515
rect 23566 13512 23572 13524
rect 16025 13475 16083 13481
rect 18156 13484 23572 13512
rect 2866 13444 2872 13456
rect 1412 13416 2872 13444
rect 1412 13385 1440 13416
rect 2866 13404 2872 13416
rect 2924 13404 2930 13456
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13345 1455 13379
rect 1578 13376 1584 13388
rect 1539 13348 1584 13376
rect 1397 13339 1455 13345
rect 1578 13336 1584 13348
rect 1636 13336 1642 13388
rect 2774 13336 2780 13388
rect 2832 13376 2838 13388
rect 2832 13348 2877 13376
rect 2832 13336 2838 13348
rect 14274 13336 14280 13388
rect 14332 13376 14338 13388
rect 14645 13379 14703 13385
rect 14645 13376 14657 13379
rect 14332 13348 14657 13376
rect 14332 13336 14338 13348
rect 14645 13345 14657 13348
rect 14691 13345 14703 13379
rect 14645 13339 14703 13345
rect 7926 13268 7932 13320
rect 7984 13308 7990 13320
rect 8110 13308 8116 13320
rect 7984 13280 8116 13308
rect 7984 13268 7990 13280
rect 8110 13268 8116 13280
rect 8168 13308 8174 13320
rect 8205 13311 8263 13317
rect 8205 13308 8217 13311
rect 8168 13280 8217 13308
rect 8168 13268 8174 13280
rect 8205 13277 8217 13280
rect 8251 13277 8263 13311
rect 8205 13271 8263 13277
rect 15194 13268 15200 13320
rect 15252 13308 15258 13320
rect 18156 13317 18184 13484
rect 23566 13472 23572 13484
rect 23624 13472 23630 13524
rect 26326 13472 26332 13524
rect 26384 13512 26390 13524
rect 26881 13515 26939 13521
rect 26881 13512 26893 13515
rect 26384 13484 26893 13512
rect 26384 13472 26390 13484
rect 26881 13481 26893 13484
rect 26927 13481 26939 13515
rect 26881 13475 26939 13481
rect 27154 13472 27160 13524
rect 27212 13512 27218 13524
rect 27614 13512 27620 13524
rect 27212 13484 27620 13512
rect 27212 13472 27218 13484
rect 27614 13472 27620 13484
rect 27672 13472 27678 13524
rect 28813 13515 28871 13521
rect 28813 13481 28825 13515
rect 28859 13512 28871 13515
rect 29454 13512 29460 13524
rect 28859 13484 29460 13512
rect 28859 13481 28871 13484
rect 28813 13475 28871 13481
rect 29454 13472 29460 13484
rect 29512 13472 29518 13524
rect 29914 13472 29920 13524
rect 29972 13512 29978 13524
rect 29972 13484 30768 13512
rect 29972 13472 29978 13484
rect 27890 13404 27896 13456
rect 27948 13444 27954 13456
rect 27948 13416 30696 13444
rect 27948 13404 27954 13416
rect 18598 13376 18604 13388
rect 18248 13348 18604 13376
rect 18248 13317 18276 13348
rect 18598 13336 18604 13348
rect 18656 13376 18662 13388
rect 19889 13379 19947 13385
rect 19889 13376 19901 13379
rect 18656 13348 19901 13376
rect 18656 13336 18662 13348
rect 19889 13345 19901 13348
rect 19935 13345 19947 13379
rect 19889 13339 19947 13345
rect 23934 13336 23940 13388
rect 23992 13376 23998 13388
rect 26145 13379 26203 13385
rect 26145 13376 26157 13379
rect 23992 13348 26157 13376
rect 23992 13336 23998 13348
rect 26145 13345 26157 13348
rect 26191 13345 26203 13379
rect 26145 13339 26203 13345
rect 26973 13379 27031 13385
rect 26973 13345 26985 13379
rect 27019 13376 27031 13379
rect 27706 13376 27712 13388
rect 27019 13348 27712 13376
rect 27019 13345 27031 13348
rect 26973 13339 27031 13345
rect 27706 13336 27712 13348
rect 27764 13336 27770 13388
rect 29825 13379 29883 13385
rect 29825 13345 29837 13379
rect 29871 13376 29883 13379
rect 30374 13376 30380 13388
rect 29871 13348 30380 13376
rect 29871 13345 29883 13348
rect 29825 13339 29883 13345
rect 30374 13336 30380 13348
rect 30432 13336 30438 13388
rect 18141 13311 18199 13317
rect 15252 13280 17448 13308
rect 15252 13268 15258 13280
rect 14912 13243 14970 13249
rect 14912 13209 14924 13243
rect 14958 13240 14970 13243
rect 15010 13240 15016 13252
rect 14958 13212 15016 13240
rect 14958 13209 14970 13212
rect 14912 13203 14970 13209
rect 15010 13200 15016 13212
rect 15068 13200 15074 13252
rect 17218 13240 17224 13252
rect 17179 13212 17224 13240
rect 17218 13200 17224 13212
rect 17276 13200 17282 13252
rect 17420 13249 17448 13280
rect 18141 13277 18153 13311
rect 18187 13277 18199 13311
rect 18141 13271 18199 13277
rect 18233 13311 18291 13317
rect 18233 13277 18245 13311
rect 18279 13277 18291 13311
rect 18233 13271 18291 13277
rect 18322 13268 18328 13320
rect 18380 13308 18386 13320
rect 18380 13280 18425 13308
rect 18380 13268 18386 13280
rect 18506 13268 18512 13320
rect 18564 13308 18570 13320
rect 19702 13308 19708 13320
rect 18564 13280 18609 13308
rect 19663 13280 19708 13308
rect 18564 13268 18570 13280
rect 19702 13268 19708 13280
rect 19760 13268 19766 13320
rect 20349 13311 20407 13317
rect 20349 13277 20361 13311
rect 20395 13308 20407 13311
rect 20714 13308 20720 13320
rect 20395 13280 20720 13308
rect 20395 13277 20407 13280
rect 20349 13271 20407 13277
rect 20714 13268 20720 13280
rect 20772 13268 20778 13320
rect 22465 13311 22523 13317
rect 22465 13277 22477 13311
rect 22511 13308 22523 13311
rect 23014 13308 23020 13320
rect 22511 13280 23020 13308
rect 22511 13277 22523 13280
rect 22465 13271 22523 13277
rect 23014 13268 23020 13280
rect 23072 13268 23078 13320
rect 25222 13308 25228 13320
rect 25183 13280 25228 13308
rect 25222 13268 25228 13280
rect 25280 13308 25286 13320
rect 25961 13311 26019 13317
rect 25961 13308 25973 13311
rect 25280 13280 25973 13308
rect 25280 13268 25286 13280
rect 25961 13277 25973 13280
rect 26007 13277 26019 13311
rect 25961 13271 26019 13277
rect 26602 13268 26608 13320
rect 26660 13308 26666 13320
rect 26697 13311 26755 13317
rect 26697 13308 26709 13311
rect 26660 13280 26709 13308
rect 26660 13268 26666 13280
rect 26697 13277 26709 13280
rect 26743 13277 26755 13311
rect 26697 13271 26755 13277
rect 26789 13311 26847 13317
rect 26789 13277 26801 13311
rect 26835 13308 26847 13311
rect 26878 13308 26884 13320
rect 26835 13280 26884 13308
rect 26835 13277 26847 13280
rect 26789 13271 26847 13277
rect 26878 13268 26884 13280
rect 26936 13308 26942 13320
rect 27985 13311 28043 13317
rect 27985 13308 27997 13311
rect 26936 13280 27997 13308
rect 26936 13268 26942 13280
rect 27985 13277 27997 13280
rect 28031 13277 28043 13311
rect 27985 13271 28043 13277
rect 28994 13268 29000 13320
rect 29052 13308 29058 13320
rect 29549 13311 29607 13317
rect 29549 13308 29561 13311
rect 29052 13280 29561 13308
rect 29052 13268 29058 13280
rect 29549 13277 29561 13280
rect 29595 13277 29607 13311
rect 29730 13308 29736 13320
rect 29691 13280 29736 13308
rect 29549 13271 29607 13277
rect 29730 13268 29736 13280
rect 29788 13268 29794 13320
rect 29917 13311 29975 13317
rect 29917 13277 29929 13311
rect 29963 13308 29975 13311
rect 30006 13308 30012 13320
rect 29963 13280 30012 13308
rect 29963 13277 29975 13280
rect 29917 13271 29975 13277
rect 17405 13243 17463 13249
rect 17405 13209 17417 13243
rect 17451 13240 17463 13243
rect 18524 13240 18552 13268
rect 17451 13212 18552 13240
rect 22732 13243 22790 13249
rect 17451 13209 17463 13212
rect 17405 13203 17463 13209
rect 22732 13209 22744 13243
rect 22778 13240 22790 13243
rect 25130 13240 25136 13252
rect 22778 13212 25136 13240
rect 22778 13209 22790 13212
rect 22732 13203 22790 13209
rect 25130 13200 25136 13212
rect 25188 13200 25194 13252
rect 28721 13243 28779 13249
rect 28721 13240 28733 13243
rect 25332 13212 28733 13240
rect 17862 13172 17868 13184
rect 17823 13144 17868 13172
rect 17862 13132 17868 13144
rect 17920 13132 17926 13184
rect 20254 13132 20260 13184
rect 20312 13172 20318 13184
rect 20441 13175 20499 13181
rect 20441 13172 20453 13175
rect 20312 13144 20453 13172
rect 20312 13132 20318 13144
rect 20441 13141 20453 13144
rect 20487 13141 20499 13175
rect 20441 13135 20499 13141
rect 23750 13132 23756 13184
rect 23808 13172 23814 13184
rect 23845 13175 23903 13181
rect 23845 13172 23857 13175
rect 23808 13144 23857 13172
rect 23808 13132 23814 13144
rect 23845 13141 23857 13144
rect 23891 13141 23903 13175
rect 23845 13135 23903 13141
rect 25038 13132 25044 13184
rect 25096 13172 25102 13184
rect 25332 13181 25360 13212
rect 28721 13209 28733 13212
rect 28767 13240 28779 13243
rect 29454 13240 29460 13252
rect 28767 13212 29460 13240
rect 28767 13209 28779 13212
rect 28721 13203 28779 13209
rect 29454 13200 29460 13212
rect 29512 13200 29518 13252
rect 25317 13175 25375 13181
rect 25317 13172 25329 13175
rect 25096 13144 25329 13172
rect 25096 13132 25102 13144
rect 25317 13141 25329 13144
rect 25363 13141 25375 13175
rect 25317 13135 25375 13141
rect 28077 13175 28135 13181
rect 28077 13141 28089 13175
rect 28123 13172 28135 13175
rect 29638 13172 29644 13184
rect 28123 13144 29644 13172
rect 28123 13141 28135 13144
rect 28077 13135 28135 13141
rect 29638 13132 29644 13144
rect 29696 13172 29702 13184
rect 29932 13172 29960 13271
rect 30006 13268 30012 13280
rect 30064 13268 30070 13320
rect 30101 13311 30159 13317
rect 30101 13277 30113 13311
rect 30147 13308 30159 13311
rect 30558 13308 30564 13320
rect 30147 13280 30564 13308
rect 30147 13277 30159 13280
rect 30101 13271 30159 13277
rect 30116 13240 30144 13271
rect 30558 13268 30564 13280
rect 30616 13268 30622 13320
rect 30668 13308 30696 13416
rect 30740 13376 30768 13484
rect 33594 13472 33600 13524
rect 33652 13512 33658 13524
rect 33781 13515 33839 13521
rect 33781 13512 33793 13515
rect 33652 13484 33793 13512
rect 33652 13472 33658 13484
rect 33781 13481 33793 13484
rect 33827 13481 33839 13515
rect 33781 13475 33839 13481
rect 36541 13515 36599 13521
rect 36541 13481 36553 13515
rect 36587 13512 36599 13515
rect 36722 13512 36728 13524
rect 36587 13484 36728 13512
rect 36587 13481 36599 13484
rect 36541 13475 36599 13481
rect 36722 13472 36728 13484
rect 36780 13472 36786 13524
rect 30834 13404 30840 13456
rect 30892 13444 30898 13456
rect 30892 13416 30937 13444
rect 30892 13404 30898 13416
rect 35526 13404 35532 13456
rect 35584 13404 35590 13456
rect 32398 13376 32404 13388
rect 30740 13348 32404 13376
rect 32398 13336 32404 13348
rect 32456 13336 32462 13388
rect 35544 13376 35572 13404
rect 35452 13348 35572 13376
rect 30745 13311 30803 13317
rect 30745 13308 30757 13311
rect 30668 13280 30757 13308
rect 30745 13277 30757 13280
rect 30791 13277 30803 13311
rect 30926 13308 30932 13320
rect 30887 13280 30932 13308
rect 30745 13271 30803 13277
rect 30926 13268 30932 13280
rect 30984 13268 30990 13320
rect 31754 13268 31760 13320
rect 31812 13308 31818 13320
rect 31812 13280 31857 13308
rect 31812 13268 31818 13280
rect 32490 13268 32496 13320
rect 32548 13308 32554 13320
rect 32657 13311 32715 13317
rect 32657 13308 32669 13311
rect 32548 13280 32669 13308
rect 32548 13268 32554 13280
rect 32657 13277 32669 13280
rect 32703 13277 32715 13311
rect 35342 13308 35348 13320
rect 35303 13280 35348 13308
rect 32657 13271 32715 13277
rect 35342 13268 35348 13280
rect 35400 13268 35406 13320
rect 35452 13317 35480 13348
rect 35434 13311 35492 13317
rect 35434 13277 35446 13311
rect 35480 13277 35492 13311
rect 35434 13271 35492 13277
rect 35526 13268 35532 13320
rect 35584 13308 35590 13320
rect 35710 13308 35716 13320
rect 35584 13280 35629 13308
rect 35671 13280 35716 13308
rect 35584 13268 35590 13280
rect 35710 13268 35716 13280
rect 35768 13268 35774 13320
rect 36354 13308 36360 13320
rect 36315 13280 36360 13308
rect 36354 13268 36360 13280
rect 36412 13268 36418 13320
rect 30024 13212 30144 13240
rect 30024 13184 30052 13212
rect 34514 13200 34520 13252
rect 34572 13240 34578 13252
rect 36173 13243 36231 13249
rect 36173 13240 36185 13243
rect 34572 13212 36185 13240
rect 34572 13200 34578 13212
rect 36173 13209 36185 13212
rect 36219 13209 36231 13243
rect 36173 13203 36231 13209
rect 29696 13144 29960 13172
rect 29696 13132 29702 13144
rect 30006 13132 30012 13184
rect 30064 13132 30070 13184
rect 30190 13132 30196 13184
rect 30248 13172 30254 13184
rect 30285 13175 30343 13181
rect 30285 13172 30297 13175
rect 30248 13144 30297 13172
rect 30248 13132 30254 13144
rect 30285 13141 30297 13144
rect 30331 13141 30343 13175
rect 30285 13135 30343 13141
rect 31849 13175 31907 13181
rect 31849 13141 31861 13175
rect 31895 13172 31907 13175
rect 32490 13172 32496 13184
rect 31895 13144 32496 13172
rect 31895 13141 31907 13144
rect 31849 13135 31907 13141
rect 32490 13132 32496 13144
rect 32548 13132 32554 13184
rect 35066 13172 35072 13184
rect 35027 13144 35072 13172
rect 35066 13132 35072 13144
rect 35124 13132 35130 13184
rect 1104 13082 48852 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 48852 13082
rect 1104 13008 48852 13030
rect 19334 12928 19340 12980
rect 19392 12968 19398 12980
rect 19978 12968 19984 12980
rect 19392 12940 19984 12968
rect 19392 12928 19398 12940
rect 19978 12928 19984 12940
rect 20036 12928 20042 12980
rect 23566 12928 23572 12980
rect 23624 12968 23630 12980
rect 23661 12971 23719 12977
rect 23661 12968 23673 12971
rect 23624 12940 23673 12968
rect 23624 12928 23630 12940
rect 23661 12937 23673 12940
rect 23707 12968 23719 12971
rect 23707 12940 24992 12968
rect 23707 12937 23719 12940
rect 23661 12931 23719 12937
rect 15286 12860 15292 12912
rect 15344 12900 15350 12912
rect 16936 12903 16994 12909
rect 15344 12872 16896 12900
rect 15344 12860 15350 12872
rect 1673 12835 1731 12841
rect 1673 12801 1685 12835
rect 1719 12832 1731 12835
rect 3970 12832 3976 12844
rect 1719 12804 3976 12832
rect 1719 12801 1731 12804
rect 1673 12795 1731 12801
rect 3970 12792 3976 12804
rect 4028 12792 4034 12844
rect 14090 12832 14096 12844
rect 14051 12804 14096 12832
rect 14090 12792 14096 12804
rect 14148 12792 14154 12844
rect 16666 12832 16672 12844
rect 16627 12804 16672 12832
rect 16666 12792 16672 12804
rect 16724 12792 16730 12844
rect 16868 12832 16896 12872
rect 16936 12869 16948 12903
rect 16982 12900 16994 12903
rect 17862 12900 17868 12912
rect 16982 12872 17868 12900
rect 16982 12869 16994 12872
rect 16936 12863 16994 12869
rect 17862 12860 17868 12872
rect 17920 12860 17926 12912
rect 18690 12860 18696 12912
rect 18748 12900 18754 12912
rect 19889 12903 19947 12909
rect 19889 12900 19901 12903
rect 18748 12872 19901 12900
rect 18748 12860 18754 12872
rect 19889 12869 19901 12872
rect 19935 12869 19947 12903
rect 19889 12863 19947 12869
rect 20717 12903 20775 12909
rect 20717 12869 20729 12903
rect 20763 12900 20775 12903
rect 20990 12900 20996 12912
rect 20763 12872 20996 12900
rect 20763 12869 20775 12872
rect 20717 12863 20775 12869
rect 20990 12860 20996 12872
rect 21048 12900 21054 12912
rect 21358 12900 21364 12912
rect 21048 12872 21364 12900
rect 21048 12860 21054 12872
rect 21358 12860 21364 12872
rect 21416 12860 21422 12912
rect 23750 12860 23756 12912
rect 23808 12900 23814 12912
rect 23808 12872 24808 12900
rect 23808 12860 23814 12872
rect 18509 12835 18567 12841
rect 18509 12832 18521 12835
rect 16868 12804 18521 12832
rect 18509 12801 18521 12804
rect 18555 12832 18567 12835
rect 23566 12832 23572 12844
rect 18555 12804 23572 12832
rect 18555 12801 18567 12804
rect 18509 12795 18567 12801
rect 23566 12792 23572 12804
rect 23624 12792 23630 12844
rect 24486 12832 24492 12844
rect 24447 12804 24492 12832
rect 24486 12792 24492 12804
rect 24544 12792 24550 12844
rect 24780 12841 24808 12872
rect 24673 12835 24731 12841
rect 24673 12801 24685 12835
rect 24719 12801 24731 12835
rect 24673 12795 24731 12801
rect 24765 12835 24823 12841
rect 24765 12801 24777 12835
rect 24811 12801 24823 12835
rect 24964 12832 24992 12940
rect 27246 12928 27252 12980
rect 27304 12968 27310 12980
rect 29086 12968 29092 12980
rect 27304 12940 29092 12968
rect 27304 12928 27310 12940
rect 29086 12928 29092 12940
rect 29144 12928 29150 12980
rect 29273 12971 29331 12977
rect 29273 12937 29285 12971
rect 29319 12968 29331 12971
rect 30006 12968 30012 12980
rect 29319 12940 30012 12968
rect 29319 12937 29331 12940
rect 29273 12931 29331 12937
rect 30006 12928 30012 12940
rect 30064 12928 30070 12980
rect 26786 12860 26792 12912
rect 26844 12900 26850 12912
rect 29730 12900 29736 12912
rect 26844 12872 29736 12900
rect 26844 12860 26850 12872
rect 29288 12844 29316 12872
rect 29730 12860 29736 12872
rect 29788 12860 29794 12912
rect 35066 12860 35072 12912
rect 35124 12900 35130 12912
rect 35222 12903 35280 12909
rect 35222 12900 35234 12903
rect 35124 12872 35234 12900
rect 35124 12860 35130 12872
rect 35222 12869 35234 12872
rect 35268 12869 35280 12903
rect 35222 12863 35280 12869
rect 25041 12835 25099 12841
rect 25041 12832 25053 12835
rect 24964 12804 25053 12832
rect 24765 12795 24823 12801
rect 25041 12801 25053 12804
rect 25087 12801 25099 12835
rect 25041 12795 25099 12801
rect 1394 12764 1400 12776
rect 1355 12736 1400 12764
rect 1394 12724 1400 12736
rect 1452 12724 1458 12776
rect 14274 12764 14280 12776
rect 14235 12736 14280 12764
rect 14274 12724 14280 12736
rect 14332 12724 14338 12776
rect 14553 12767 14611 12773
rect 14553 12733 14565 12767
rect 14599 12733 14611 12767
rect 14553 12727 14611 12733
rect 18785 12767 18843 12773
rect 18785 12733 18797 12767
rect 18831 12764 18843 12767
rect 19150 12764 19156 12776
rect 18831 12736 19156 12764
rect 18831 12733 18843 12736
rect 18785 12727 18843 12733
rect 12434 12656 12440 12708
rect 12492 12696 12498 12708
rect 14568 12696 14596 12727
rect 19150 12724 19156 12736
rect 19208 12724 19214 12776
rect 23750 12764 23756 12776
rect 23711 12736 23756 12764
rect 23750 12724 23756 12736
rect 23808 12724 23814 12776
rect 23934 12764 23940 12776
rect 23895 12736 23940 12764
rect 23934 12724 23940 12736
rect 23992 12724 23998 12776
rect 12492 12668 14596 12696
rect 12492 12656 12498 12668
rect 18046 12628 18052 12640
rect 18007 12600 18052 12628
rect 18046 12588 18052 12600
rect 18104 12588 18110 12640
rect 19242 12588 19248 12640
rect 19300 12628 19306 12640
rect 20070 12628 20076 12640
rect 19300 12600 20076 12628
rect 19300 12588 19306 12600
rect 20070 12588 20076 12600
rect 20128 12628 20134 12640
rect 20809 12631 20867 12637
rect 20809 12628 20821 12631
rect 20128 12600 20821 12628
rect 20128 12588 20134 12600
rect 20809 12597 20821 12600
rect 20855 12597 20867 12631
rect 20809 12591 20867 12597
rect 23293 12631 23351 12637
rect 23293 12597 23305 12631
rect 23339 12628 23351 12631
rect 23474 12628 23480 12640
rect 23339 12600 23480 12628
rect 23339 12597 23351 12600
rect 23293 12591 23351 12597
rect 23474 12588 23480 12600
rect 23532 12588 23538 12640
rect 24688 12628 24716 12795
rect 25130 12792 25136 12844
rect 25188 12832 25194 12844
rect 25225 12835 25283 12841
rect 25225 12832 25237 12835
rect 25188 12804 25237 12832
rect 25188 12792 25194 12804
rect 25225 12801 25237 12804
rect 25271 12801 25283 12835
rect 25225 12795 25283 12801
rect 27706 12792 27712 12844
rect 27764 12832 27770 12844
rect 27801 12835 27859 12841
rect 27801 12832 27813 12835
rect 27764 12804 27813 12832
rect 27764 12792 27770 12804
rect 27801 12801 27813 12804
rect 27847 12801 27859 12835
rect 27801 12795 27859 12801
rect 29270 12792 29276 12844
rect 29328 12792 29334 12844
rect 29365 12835 29423 12841
rect 29365 12801 29377 12835
rect 29411 12832 29423 12835
rect 30374 12832 30380 12844
rect 29411 12804 30380 12832
rect 29411 12801 29423 12804
rect 29365 12795 29423 12801
rect 30374 12792 30380 12804
rect 30432 12832 30438 12844
rect 31294 12832 31300 12844
rect 30432 12804 31300 12832
rect 30432 12792 30438 12804
rect 31294 12792 31300 12804
rect 31352 12792 31358 12844
rect 32398 12832 32404 12844
rect 32311 12804 32404 12832
rect 32398 12792 32404 12804
rect 32456 12832 32462 12844
rect 32766 12832 32772 12844
rect 32456 12804 32772 12832
rect 32456 12792 32462 12804
rect 32766 12792 32772 12804
rect 32824 12792 32830 12844
rect 34790 12792 34796 12844
rect 34848 12832 34854 12844
rect 34977 12835 35035 12841
rect 34977 12832 34989 12835
rect 34848 12804 34989 12832
rect 34848 12792 34854 12804
rect 34977 12801 34989 12804
rect 35023 12801 35035 12835
rect 34977 12795 35035 12801
rect 24857 12767 24915 12773
rect 24857 12733 24869 12767
rect 24903 12764 24915 12767
rect 26326 12764 26332 12776
rect 24903 12736 26332 12764
rect 24903 12733 24915 12736
rect 24857 12727 24915 12733
rect 26326 12724 26332 12736
rect 26384 12764 26390 12776
rect 28350 12764 28356 12776
rect 26384 12736 28356 12764
rect 26384 12724 26390 12736
rect 28350 12724 28356 12736
rect 28408 12724 28414 12776
rect 29454 12764 29460 12776
rect 29415 12736 29460 12764
rect 29454 12724 29460 12736
rect 29512 12724 29518 12776
rect 31754 12764 31760 12776
rect 29564 12736 31760 12764
rect 25130 12656 25136 12708
rect 25188 12696 25194 12708
rect 29564 12696 29592 12736
rect 31754 12724 31760 12736
rect 31812 12764 31818 12776
rect 32125 12767 32183 12773
rect 32125 12764 32137 12767
rect 31812 12736 32137 12764
rect 31812 12724 31818 12736
rect 32125 12733 32137 12736
rect 32171 12733 32183 12767
rect 32125 12727 32183 12733
rect 25188 12668 29592 12696
rect 25188 12656 25194 12668
rect 26786 12628 26792 12640
rect 24688 12600 26792 12628
rect 26786 12588 26792 12600
rect 26844 12588 26850 12640
rect 27246 12588 27252 12640
rect 27304 12628 27310 12640
rect 27893 12631 27951 12637
rect 27893 12628 27905 12631
rect 27304 12600 27905 12628
rect 27304 12588 27310 12600
rect 27893 12597 27905 12600
rect 27939 12597 27951 12631
rect 27893 12591 27951 12597
rect 27982 12588 27988 12640
rect 28040 12628 28046 12640
rect 28905 12631 28963 12637
rect 28905 12628 28917 12631
rect 28040 12600 28917 12628
rect 28040 12588 28046 12600
rect 28905 12597 28917 12600
rect 28951 12597 28963 12631
rect 36354 12628 36360 12640
rect 36315 12600 36360 12628
rect 28905 12591 28963 12597
rect 36354 12588 36360 12600
rect 36412 12588 36418 12640
rect 1104 12538 48852 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 48852 12538
rect 1104 12464 48852 12486
rect 14274 12424 14280 12436
rect 14235 12396 14280 12424
rect 14274 12384 14280 12396
rect 14332 12384 14338 12436
rect 18322 12384 18328 12436
rect 18380 12424 18386 12436
rect 18693 12427 18751 12433
rect 18693 12424 18705 12427
rect 18380 12396 18705 12424
rect 18380 12384 18386 12396
rect 18693 12393 18705 12396
rect 18739 12393 18751 12427
rect 18693 12387 18751 12393
rect 18874 12384 18880 12436
rect 18932 12424 18938 12436
rect 20714 12424 20720 12436
rect 18932 12396 20720 12424
rect 18932 12384 18938 12396
rect 20714 12384 20720 12396
rect 20772 12384 20778 12436
rect 23569 12427 23627 12433
rect 23569 12393 23581 12427
rect 23615 12424 23627 12427
rect 24486 12424 24492 12436
rect 23615 12396 24492 12424
rect 23615 12393 23627 12396
rect 23569 12387 23627 12393
rect 24486 12384 24492 12396
rect 24544 12384 24550 12436
rect 26694 12384 26700 12436
rect 26752 12424 26758 12436
rect 26881 12427 26939 12433
rect 26881 12424 26893 12427
rect 26752 12396 26893 12424
rect 26752 12384 26758 12396
rect 26881 12393 26893 12396
rect 26927 12393 26939 12427
rect 31294 12424 31300 12436
rect 31255 12396 31300 12424
rect 26881 12387 26939 12393
rect 31294 12384 31300 12396
rect 31352 12384 31358 12436
rect 35345 12427 35403 12433
rect 35345 12393 35357 12427
rect 35391 12424 35403 12427
rect 35526 12424 35532 12436
rect 35391 12396 35532 12424
rect 35391 12393 35403 12396
rect 35345 12387 35403 12393
rect 35526 12384 35532 12396
rect 35584 12384 35590 12436
rect 40770 12384 40776 12436
rect 40828 12424 40834 12436
rect 46842 12424 46848 12436
rect 40828 12396 46848 12424
rect 40828 12384 40834 12396
rect 46842 12384 46848 12396
rect 46900 12384 46906 12436
rect 16025 12291 16083 12297
rect 16025 12257 16037 12291
rect 16071 12288 16083 12291
rect 18046 12288 18052 12300
rect 16071 12260 18052 12288
rect 16071 12257 16083 12260
rect 16025 12251 16083 12257
rect 18046 12248 18052 12260
rect 18104 12288 18110 12300
rect 20254 12288 20260 12300
rect 18104 12260 18552 12288
rect 20215 12260 20260 12288
rect 18104 12248 18110 12260
rect 18524 12229 18552 12260
rect 20254 12248 20260 12260
rect 20312 12248 20318 12300
rect 26878 12288 26884 12300
rect 26712 12260 26884 12288
rect 26712 12232 26740 12260
rect 26878 12248 26884 12260
rect 26936 12288 26942 12300
rect 27709 12291 27767 12297
rect 27709 12288 27721 12291
rect 26936 12260 27721 12288
rect 26936 12248 26942 12260
rect 27709 12257 27721 12260
rect 27755 12257 27767 12291
rect 29914 12288 29920 12300
rect 29875 12260 29920 12288
rect 27709 12251 27767 12257
rect 29914 12248 29920 12260
rect 29972 12248 29978 12300
rect 33410 12248 33416 12300
rect 33468 12288 33474 12300
rect 33468 12260 35204 12288
rect 33468 12248 33474 12260
rect 14185 12223 14243 12229
rect 14185 12189 14197 12223
rect 14231 12220 14243 12223
rect 15381 12223 15439 12229
rect 15381 12220 15393 12223
rect 14231 12192 15393 12220
rect 14231 12189 14243 12192
rect 14185 12183 14243 12189
rect 15381 12189 15393 12192
rect 15427 12189 15439 12223
rect 15381 12183 15439 12189
rect 18509 12223 18567 12229
rect 18509 12189 18521 12223
rect 18555 12189 18567 12223
rect 18509 12183 18567 12189
rect 19429 12223 19487 12229
rect 19429 12189 19441 12223
rect 19475 12220 19487 12223
rect 20070 12220 20076 12232
rect 19475 12192 20076 12220
rect 19475 12189 19487 12192
rect 19429 12183 19487 12189
rect 15396 12084 15424 12183
rect 20070 12180 20076 12192
rect 20128 12180 20134 12232
rect 23474 12220 23480 12232
rect 23435 12192 23480 12220
rect 23474 12180 23480 12192
rect 23532 12180 23538 12232
rect 23658 12220 23664 12232
rect 23619 12192 23664 12220
rect 23658 12180 23664 12192
rect 23716 12180 23722 12232
rect 26694 12220 26700 12232
rect 26655 12192 26700 12220
rect 26694 12180 26700 12192
rect 26752 12180 26758 12232
rect 27433 12223 27491 12229
rect 27433 12189 27445 12223
rect 27479 12220 27491 12223
rect 27522 12220 27528 12232
rect 27479 12192 27528 12220
rect 27479 12189 27491 12192
rect 27433 12183 27491 12189
rect 27522 12180 27528 12192
rect 27580 12180 27586 12232
rect 28997 12223 29055 12229
rect 27632 12192 28948 12220
rect 15473 12155 15531 12161
rect 15473 12121 15485 12155
rect 15519 12152 15531 12155
rect 16209 12155 16267 12161
rect 16209 12152 16221 12155
rect 15519 12124 16221 12152
rect 15519 12121 15531 12124
rect 15473 12115 15531 12121
rect 16209 12121 16221 12124
rect 16255 12121 16267 12155
rect 17862 12152 17868 12164
rect 17823 12124 17868 12152
rect 16209 12115 16267 12121
rect 17862 12112 17868 12124
rect 17920 12112 17926 12164
rect 18325 12155 18383 12161
rect 18325 12121 18337 12155
rect 18371 12152 18383 12155
rect 19150 12152 19156 12164
rect 18371 12124 19156 12152
rect 18371 12121 18383 12124
rect 18325 12115 18383 12121
rect 19150 12112 19156 12124
rect 19208 12152 19214 12164
rect 19245 12155 19303 12161
rect 19245 12152 19257 12155
rect 19208 12124 19257 12152
rect 19208 12112 19214 12124
rect 19245 12121 19257 12124
rect 19291 12121 19303 12155
rect 19245 12115 19303 12121
rect 19518 12112 19524 12164
rect 19576 12152 19582 12164
rect 20254 12152 20260 12164
rect 19576 12124 20260 12152
rect 19576 12112 19582 12124
rect 20254 12112 20260 12124
rect 20312 12112 20318 12164
rect 21910 12152 21916 12164
rect 21871 12124 21916 12152
rect 21910 12112 21916 12124
rect 21968 12112 21974 12164
rect 26878 12112 26884 12164
rect 26936 12152 26942 12164
rect 27632 12152 27660 12192
rect 26936 12124 27660 12152
rect 26936 12112 26942 12124
rect 27706 12112 27712 12164
rect 27764 12152 27770 12164
rect 28813 12155 28871 12161
rect 28813 12152 28825 12155
rect 27764 12124 28825 12152
rect 27764 12112 27770 12124
rect 28813 12121 28825 12124
rect 28859 12121 28871 12155
rect 28920 12152 28948 12192
rect 28997 12189 29009 12223
rect 29043 12220 29055 12223
rect 29362 12220 29368 12232
rect 29043 12192 29368 12220
rect 29043 12189 29055 12192
rect 28997 12183 29055 12189
rect 29362 12180 29368 12192
rect 29420 12220 29426 12232
rect 30006 12220 30012 12232
rect 29420 12192 30012 12220
rect 29420 12180 29426 12192
rect 30006 12180 30012 12192
rect 30064 12180 30070 12232
rect 30190 12229 30196 12232
rect 30184 12183 30196 12229
rect 30248 12220 30254 12232
rect 30248 12192 30284 12220
rect 30190 12180 30196 12183
rect 30248 12180 30254 12192
rect 34514 12180 34520 12232
rect 34572 12220 34578 12232
rect 35176 12229 35204 12260
rect 34977 12223 35035 12229
rect 34977 12220 34989 12223
rect 34572 12192 34989 12220
rect 34572 12180 34578 12192
rect 34977 12189 34989 12192
rect 35023 12189 35035 12223
rect 34977 12183 35035 12189
rect 35161 12223 35219 12229
rect 35161 12189 35173 12223
rect 35207 12220 35219 12223
rect 36354 12220 36360 12232
rect 35207 12192 36360 12220
rect 35207 12189 35219 12192
rect 35161 12183 35219 12189
rect 36354 12180 36360 12192
rect 36412 12180 36418 12232
rect 28920 12124 31754 12152
rect 28813 12115 28871 12121
rect 18230 12084 18236 12096
rect 15396 12056 18236 12084
rect 18230 12044 18236 12056
rect 18288 12044 18294 12096
rect 19613 12087 19671 12093
rect 19613 12053 19625 12087
rect 19659 12084 19671 12087
rect 19978 12084 19984 12096
rect 19659 12056 19984 12084
rect 19659 12053 19671 12056
rect 19613 12047 19671 12053
rect 19978 12044 19984 12056
rect 20036 12044 20042 12096
rect 28258 12044 28264 12096
rect 28316 12084 28322 12096
rect 28534 12084 28540 12096
rect 28316 12056 28540 12084
rect 28316 12044 28322 12056
rect 28534 12044 28540 12056
rect 28592 12044 28598 12096
rect 28828 12084 28856 12115
rect 29638 12084 29644 12096
rect 28828 12056 29644 12084
rect 29638 12044 29644 12056
rect 29696 12044 29702 12096
rect 31726 12084 31754 12124
rect 32582 12084 32588 12096
rect 31726 12056 32588 12084
rect 32582 12044 32588 12056
rect 32640 12044 32646 12096
rect 1104 11994 48852 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 48852 11994
rect 1104 11920 48852 11942
rect 19889 11883 19947 11889
rect 19889 11849 19901 11883
rect 19935 11880 19947 11883
rect 20070 11880 20076 11892
rect 19935 11852 20076 11880
rect 19935 11849 19947 11852
rect 19889 11843 19947 11849
rect 20070 11840 20076 11852
rect 20128 11840 20134 11892
rect 20530 11880 20536 11892
rect 20180 11852 20536 11880
rect 17218 11704 17224 11756
rect 17276 11744 17282 11756
rect 17773 11747 17831 11753
rect 17773 11744 17785 11747
rect 17276 11716 17785 11744
rect 17276 11704 17282 11716
rect 17773 11713 17785 11716
rect 17819 11713 17831 11747
rect 17773 11707 17831 11713
rect 18776 11747 18834 11753
rect 18776 11713 18788 11747
rect 18822 11744 18834 11747
rect 19242 11744 19248 11756
rect 18822 11716 19248 11744
rect 18822 11713 18834 11716
rect 18776 11707 18834 11713
rect 19242 11704 19248 11716
rect 19300 11704 19306 11756
rect 19886 11704 19892 11756
rect 19944 11744 19950 11756
rect 20180 11744 20208 11852
rect 20530 11840 20536 11852
rect 20588 11840 20594 11892
rect 21910 11840 21916 11892
rect 21968 11880 21974 11892
rect 46750 11880 46756 11892
rect 21968 11852 46756 11880
rect 21968 11840 21974 11852
rect 46750 11840 46756 11852
rect 46808 11840 46814 11892
rect 23474 11772 23480 11824
rect 23532 11812 23538 11824
rect 24762 11812 24768 11824
rect 23532 11784 24768 11812
rect 23532 11772 23538 11784
rect 24762 11772 24768 11784
rect 24820 11812 24826 11824
rect 27065 11815 27123 11821
rect 24820 11784 26096 11812
rect 24820 11772 24826 11784
rect 20530 11744 20536 11756
rect 19944 11716 20208 11744
rect 20491 11716 20536 11744
rect 19944 11704 19950 11716
rect 20530 11704 20536 11716
rect 20588 11704 20594 11756
rect 20990 11704 20996 11756
rect 21048 11744 21054 11756
rect 21821 11747 21879 11753
rect 21821 11744 21833 11747
rect 21048 11716 21833 11744
rect 21048 11704 21054 11716
rect 21821 11713 21833 11716
rect 21867 11713 21879 11747
rect 21821 11707 21879 11713
rect 25777 11747 25835 11753
rect 25777 11713 25789 11747
rect 25823 11713 25835 11747
rect 25958 11744 25964 11756
rect 25919 11716 25964 11744
rect 25777 11707 25835 11713
rect 16666 11636 16672 11688
rect 16724 11676 16730 11688
rect 17034 11676 17040 11688
rect 16724 11648 17040 11676
rect 16724 11636 16730 11648
rect 17034 11636 17040 11648
rect 17092 11676 17098 11688
rect 18509 11679 18567 11685
rect 18509 11676 18521 11679
rect 17092 11648 18521 11676
rect 17092 11636 17098 11648
rect 18509 11645 18521 11648
rect 18555 11645 18567 11679
rect 18509 11639 18567 11645
rect 20349 11679 20407 11685
rect 20349 11645 20361 11679
rect 20395 11676 20407 11679
rect 20622 11676 20628 11688
rect 20395 11648 20628 11676
rect 20395 11645 20407 11648
rect 20349 11639 20407 11645
rect 20622 11636 20628 11648
rect 20680 11636 20686 11688
rect 20714 11636 20720 11688
rect 20772 11636 20778 11688
rect 22097 11679 22155 11685
rect 22097 11645 22109 11679
rect 22143 11676 22155 11679
rect 22186 11676 22192 11688
rect 22143 11648 22192 11676
rect 22143 11645 22155 11648
rect 22097 11639 22155 11645
rect 22186 11636 22192 11648
rect 22244 11636 22250 11688
rect 25792 11676 25820 11707
rect 25958 11704 25964 11716
rect 26016 11704 26022 11756
rect 26068 11753 26096 11784
rect 27065 11781 27077 11815
rect 27111 11812 27123 11815
rect 28902 11812 28908 11824
rect 27111 11784 28908 11812
rect 27111 11781 27123 11784
rect 27065 11775 27123 11781
rect 28902 11772 28908 11784
rect 28960 11772 28966 11824
rect 26053 11747 26111 11753
rect 26053 11713 26065 11747
rect 26099 11713 26111 11747
rect 26053 11707 26111 11713
rect 27522 11704 27528 11756
rect 27580 11744 27586 11756
rect 27709 11747 27767 11753
rect 27709 11744 27721 11747
rect 27580 11716 27721 11744
rect 27580 11704 27586 11716
rect 27709 11713 27721 11716
rect 27755 11713 27767 11747
rect 28442 11744 28448 11756
rect 28403 11716 28448 11744
rect 27709 11707 27767 11713
rect 28442 11704 28448 11716
rect 28500 11704 28506 11756
rect 28626 11744 28632 11756
rect 28587 11716 28632 11744
rect 28626 11704 28632 11716
rect 28684 11704 28690 11756
rect 29457 11747 29515 11753
rect 29457 11713 29469 11747
rect 29503 11744 29515 11747
rect 29822 11744 29828 11756
rect 29503 11716 29828 11744
rect 29503 11713 29515 11716
rect 29457 11707 29515 11713
rect 29822 11704 29828 11716
rect 29880 11704 29886 11756
rect 26418 11676 26424 11688
rect 25792 11648 26424 11676
rect 26418 11636 26424 11648
rect 26476 11636 26482 11688
rect 28258 11636 28264 11688
rect 28316 11676 28322 11688
rect 29549 11679 29607 11685
rect 29549 11676 29561 11679
rect 28316 11648 29561 11676
rect 28316 11636 28322 11648
rect 29549 11645 29561 11648
rect 29595 11645 29607 11679
rect 29549 11639 29607 11645
rect 29638 11636 29644 11688
rect 29696 11676 29702 11688
rect 29696 11648 29741 11676
rect 29696 11636 29702 11648
rect 20732 11608 20760 11636
rect 26878 11608 26884 11620
rect 20732 11580 26884 11608
rect 26878 11568 26884 11580
rect 26936 11568 26942 11620
rect 28537 11611 28595 11617
rect 28537 11577 28549 11611
rect 28583 11608 28595 11611
rect 28994 11608 29000 11620
rect 28583 11580 29000 11608
rect 28583 11577 28595 11580
rect 28537 11571 28595 11577
rect 28994 11568 29000 11580
rect 29052 11568 29058 11620
rect 17957 11543 18015 11549
rect 17957 11509 17969 11543
rect 18003 11540 18015 11543
rect 18414 11540 18420 11552
rect 18003 11512 18420 11540
rect 18003 11509 18015 11512
rect 17957 11503 18015 11509
rect 18414 11500 18420 11512
rect 18472 11500 18478 11552
rect 20717 11543 20775 11549
rect 20717 11509 20729 11543
rect 20763 11540 20775 11543
rect 20898 11540 20904 11552
rect 20763 11512 20904 11540
rect 20763 11509 20775 11512
rect 20717 11503 20775 11509
rect 20898 11500 20904 11512
rect 20956 11500 20962 11552
rect 25498 11500 25504 11552
rect 25556 11540 25562 11552
rect 25593 11543 25651 11549
rect 25593 11540 25605 11543
rect 25556 11512 25605 11540
rect 25556 11500 25562 11512
rect 25593 11509 25605 11512
rect 25639 11509 25651 11543
rect 27154 11540 27160 11552
rect 27115 11512 27160 11540
rect 25593 11503 25651 11509
rect 27154 11500 27160 11512
rect 27212 11500 27218 11552
rect 27614 11500 27620 11552
rect 27672 11540 27678 11552
rect 27890 11540 27896 11552
rect 27672 11512 27896 11540
rect 27672 11500 27678 11512
rect 27890 11500 27896 11512
rect 27948 11500 27954 11552
rect 29089 11543 29147 11549
rect 29089 11509 29101 11543
rect 29135 11540 29147 11543
rect 30006 11540 30012 11552
rect 29135 11512 30012 11540
rect 29135 11509 29147 11512
rect 29089 11503 29147 11509
rect 30006 11500 30012 11512
rect 30064 11500 30070 11552
rect 1104 11450 48852 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 48852 11450
rect 1104 11376 48852 11398
rect 17954 11296 17960 11348
rect 18012 11336 18018 11348
rect 18417 11339 18475 11345
rect 18417 11336 18429 11339
rect 18012 11308 18429 11336
rect 18012 11296 18018 11308
rect 18417 11305 18429 11308
rect 18463 11336 18475 11339
rect 18874 11336 18880 11348
rect 18463 11308 18880 11336
rect 18463 11305 18475 11308
rect 18417 11299 18475 11305
rect 18874 11296 18880 11308
rect 18932 11296 18938 11348
rect 19242 11336 19248 11348
rect 19203 11308 19248 11336
rect 19242 11296 19248 11308
rect 19300 11296 19306 11348
rect 19352 11308 19653 11336
rect 18598 11228 18604 11280
rect 18656 11268 18662 11280
rect 19352 11268 19380 11308
rect 18656 11240 19380 11268
rect 18656 11228 18662 11240
rect 2041 11203 2099 11209
rect 2041 11169 2053 11203
rect 2087 11200 2099 11203
rect 2087 11172 6914 11200
rect 2087 11169 2099 11172
rect 2041 11163 2099 11169
rect 1762 11092 1768 11144
rect 1820 11132 1826 11144
rect 2501 11135 2559 11141
rect 2501 11132 2513 11135
rect 1820 11104 2513 11132
rect 1820 11092 1826 11104
rect 2501 11101 2513 11104
rect 2547 11101 2559 11135
rect 6886 11132 6914 11172
rect 17126 11132 17132 11144
rect 6886 11104 17132 11132
rect 2501 11095 2559 11101
rect 17126 11092 17132 11104
rect 17184 11092 17190 11144
rect 18230 11092 18236 11144
rect 18288 11132 18294 11144
rect 19625 11141 19653 11308
rect 25130 11296 25136 11348
rect 25188 11336 25194 11348
rect 25958 11336 25964 11348
rect 25188 11308 25964 11336
rect 25188 11296 25194 11308
rect 25958 11296 25964 11308
rect 26016 11336 26022 11348
rect 26605 11339 26663 11345
rect 26605 11336 26617 11339
rect 26016 11308 26617 11336
rect 26016 11296 26022 11308
rect 26605 11305 26617 11308
rect 26651 11305 26663 11339
rect 26605 11299 26663 11305
rect 27525 11339 27583 11345
rect 27525 11305 27537 11339
rect 27571 11336 27583 11339
rect 28442 11336 28448 11348
rect 27571 11308 28448 11336
rect 27571 11305 27583 11308
rect 27525 11299 27583 11305
rect 28442 11296 28448 11308
rect 28500 11296 28506 11348
rect 29914 11296 29920 11348
rect 29972 11336 29978 11348
rect 31849 11339 31907 11345
rect 31849 11336 31861 11339
rect 29972 11308 31861 11336
rect 29972 11296 29978 11308
rect 31849 11305 31861 11308
rect 31895 11305 31907 11339
rect 31849 11299 31907 11305
rect 23842 11268 23848 11280
rect 21008 11240 23848 11268
rect 19978 11200 19984 11212
rect 19720 11172 19984 11200
rect 19720 11141 19748 11172
rect 19978 11160 19984 11172
rect 20036 11160 20042 11212
rect 20070 11160 20076 11212
rect 20128 11200 20134 11212
rect 20438 11200 20444 11212
rect 20128 11172 20444 11200
rect 20128 11160 20134 11172
rect 20438 11160 20444 11172
rect 20496 11160 20502 11212
rect 18325 11135 18383 11141
rect 18325 11132 18337 11135
rect 18288 11104 18337 11132
rect 18288 11092 18294 11104
rect 18325 11101 18337 11104
rect 18371 11101 18383 11135
rect 19521 11135 19579 11141
rect 19521 11110 19533 11135
rect 18325 11095 18383 11101
rect 19516 11101 19533 11110
rect 19567 11101 19579 11135
rect 19516 11098 19579 11101
rect 19444 11095 19579 11098
rect 19610 11135 19668 11141
rect 19610 11101 19622 11135
rect 19656 11101 19668 11135
rect 19610 11095 19668 11101
rect 19705 11135 19763 11141
rect 19705 11101 19717 11135
rect 19751 11101 19763 11135
rect 19705 11095 19763 11101
rect 19889 11135 19947 11141
rect 19889 11101 19901 11135
rect 19935 11101 19947 11135
rect 19889 11095 19947 11101
rect 19444 11082 19564 11095
rect 19444 11076 19544 11082
rect 1854 11064 1860 11076
rect 1815 11036 1860 11064
rect 1854 11024 1860 11036
rect 1912 11024 1918 11076
rect 1946 11024 1952 11076
rect 2004 11064 2010 11076
rect 2593 11067 2651 11073
rect 2593 11064 2605 11067
rect 2004 11036 2605 11064
rect 2004 11024 2010 11036
rect 2593 11033 2605 11036
rect 2639 11033 2651 11067
rect 2593 11027 2651 11033
rect 19426 11024 19432 11076
rect 19484 11070 19544 11076
rect 19484 11024 19490 11070
rect 18506 10956 18512 11008
rect 18564 10996 18570 11008
rect 18874 10996 18880 11008
rect 18564 10968 18880 10996
rect 18564 10956 18570 10968
rect 18874 10956 18880 10968
rect 18932 10996 18938 11008
rect 19904 10996 19932 11095
rect 20162 11092 20168 11144
rect 20220 11132 20226 11144
rect 20625 11135 20683 11141
rect 20625 11132 20637 11135
rect 20220 11104 20637 11132
rect 20220 11092 20226 11104
rect 20625 11101 20637 11104
rect 20671 11101 20683 11135
rect 20625 11095 20683 11101
rect 20717 11135 20775 11141
rect 20717 11101 20729 11135
rect 20763 11101 20775 11135
rect 20898 11132 20904 11144
rect 20859 11104 20904 11132
rect 20717 11095 20775 11101
rect 20732 11064 20760 11095
rect 20898 11092 20904 11104
rect 20956 11092 20962 11144
rect 21008 11141 21036 11240
rect 23842 11228 23848 11240
rect 23900 11228 23906 11280
rect 24210 11228 24216 11280
rect 24268 11268 24274 11280
rect 28258 11268 28264 11280
rect 24268 11240 24624 11268
rect 28219 11240 28264 11268
rect 24268 11228 24274 11240
rect 24489 11203 24547 11209
rect 24489 11200 24501 11203
rect 23216 11172 24501 11200
rect 20993 11135 21051 11141
rect 20993 11101 21005 11135
rect 21039 11101 21051 11135
rect 20993 11095 21051 11101
rect 21821 11135 21879 11141
rect 21821 11101 21833 11135
rect 21867 11132 21879 11135
rect 22186 11132 22192 11144
rect 21867 11104 22192 11132
rect 21867 11101 21879 11104
rect 21821 11095 21879 11101
rect 22186 11092 22192 11104
rect 22244 11092 22250 11144
rect 23216 11141 23244 11172
rect 24489 11169 24501 11172
rect 24535 11169 24547 11203
rect 24489 11163 24547 11169
rect 23201 11135 23259 11141
rect 23201 11101 23213 11135
rect 23247 11101 23259 11135
rect 23201 11095 23259 11101
rect 23349 11135 23407 11141
rect 23349 11101 23361 11135
rect 23395 11132 23407 11135
rect 23395 11101 23428 11132
rect 23349 11095 23428 11101
rect 21450 11064 21456 11076
rect 20732 11036 21456 11064
rect 21450 11024 21456 11036
rect 21508 11024 21514 11076
rect 22005 11067 22063 11073
rect 22005 11033 22017 11067
rect 22051 11064 22063 11067
rect 22370 11064 22376 11076
rect 22051 11036 22376 11064
rect 22051 11033 22063 11036
rect 22005 11027 22063 11033
rect 22370 11024 22376 11036
rect 22428 11024 22434 11076
rect 23400 11064 23428 11095
rect 23474 11092 23480 11144
rect 23532 11132 23538 11144
rect 23707 11135 23765 11141
rect 23532 11104 23577 11132
rect 23532 11092 23538 11104
rect 23707 11101 23719 11135
rect 23753 11132 23765 11135
rect 23842 11132 23848 11144
rect 23753 11104 23848 11132
rect 23753 11101 23765 11104
rect 23707 11095 23765 11101
rect 23842 11092 23848 11104
rect 23900 11092 23906 11144
rect 24394 11132 24400 11144
rect 24355 11104 24400 11132
rect 24394 11092 24400 11104
rect 24452 11092 24458 11144
rect 24596 11141 24624 11240
rect 28258 11228 28264 11240
rect 28316 11228 28322 11280
rect 29825 11271 29883 11277
rect 29825 11237 29837 11271
rect 29871 11237 29883 11271
rect 29825 11231 29883 11237
rect 27522 11160 27528 11212
rect 27580 11200 27586 11212
rect 28813 11203 28871 11209
rect 28813 11200 28825 11203
rect 27580 11172 28825 11200
rect 27580 11160 27586 11172
rect 28813 11169 28825 11172
rect 28859 11169 28871 11203
rect 29840 11200 29868 11231
rect 32582 11228 32588 11280
rect 32640 11268 32646 11280
rect 33134 11268 33140 11280
rect 32640 11240 33140 11268
rect 32640 11228 32646 11240
rect 33134 11228 33140 11240
rect 33192 11228 33198 11280
rect 29840 11172 30604 11200
rect 28813 11163 28871 11169
rect 24581 11135 24639 11141
rect 24581 11101 24593 11135
rect 24627 11101 24639 11135
rect 25222 11132 25228 11144
rect 25183 11104 25228 11132
rect 24581 11095 24639 11101
rect 25222 11092 25228 11104
rect 25280 11092 25286 11144
rect 25498 11141 25504 11144
rect 25492 11132 25504 11141
rect 25459 11104 25504 11132
rect 25492 11095 25504 11104
rect 25498 11092 25504 11095
rect 25556 11092 25562 11144
rect 27801 11135 27859 11141
rect 27801 11101 27813 11135
rect 27847 11132 27859 11135
rect 27982 11132 27988 11144
rect 27847 11104 27988 11132
rect 27847 11101 27859 11104
rect 27801 11095 27859 11101
rect 27982 11092 27988 11104
rect 28040 11092 28046 11144
rect 28258 11092 28264 11144
rect 28316 11132 28322 11144
rect 28718 11132 28724 11144
rect 28316 11104 28724 11132
rect 28316 11092 28322 11104
rect 28718 11092 28724 11104
rect 28776 11092 28782 11144
rect 30006 11132 30012 11144
rect 29967 11104 30012 11132
rect 30006 11092 30012 11104
rect 30064 11092 30070 11144
rect 30469 11135 30527 11141
rect 30469 11101 30481 11135
rect 30515 11101 30527 11135
rect 30576 11132 30604 11172
rect 33042 11160 33048 11212
rect 33100 11200 33106 11212
rect 33100 11172 41414 11200
rect 33100 11160 33106 11172
rect 30725 11135 30783 11141
rect 30725 11132 30737 11135
rect 30576 11104 30737 11132
rect 30469 11095 30527 11101
rect 30725 11101 30737 11104
rect 30771 11101 30783 11135
rect 30725 11095 30783 11101
rect 23569 11067 23627 11073
rect 23400 11036 23520 11064
rect 20438 10996 20444 11008
rect 18932 10968 19932 10996
rect 20399 10968 20444 10996
rect 18932 10956 18938 10968
rect 20438 10956 20444 10968
rect 20496 10956 20502 11008
rect 22189 10999 22247 11005
rect 22189 10965 22201 10999
rect 22235 10996 22247 10999
rect 22278 10996 22284 11008
rect 22235 10968 22284 10996
rect 22235 10965 22247 10968
rect 22189 10959 22247 10965
rect 22278 10956 22284 10968
rect 22336 10956 22342 11008
rect 23492 10996 23520 11036
rect 23569 11033 23581 11067
rect 23615 11064 23627 11067
rect 24026 11064 24032 11076
rect 23615 11036 24032 11064
rect 23615 11033 23627 11036
rect 23569 11027 23627 11033
rect 24026 11024 24032 11036
rect 24084 11024 24090 11076
rect 26970 11024 26976 11076
rect 27028 11064 27034 11076
rect 27522 11064 27528 11076
rect 27028 11036 27528 11064
rect 27028 11024 27034 11036
rect 27522 11024 27528 11036
rect 27580 11024 27586 11076
rect 27890 11024 27896 11076
rect 27948 11064 27954 11076
rect 28534 11064 28540 11076
rect 27948 11036 28540 11064
rect 27948 11024 27954 11036
rect 28534 11024 28540 11036
rect 28592 11024 28598 11076
rect 28629 11067 28687 11073
rect 28629 11033 28641 11067
rect 28675 11064 28687 11067
rect 29914 11064 29920 11076
rect 28675 11036 29920 11064
rect 28675 11033 28687 11036
rect 28629 11027 28687 11033
rect 29914 11024 29920 11036
rect 29972 11024 29978 11076
rect 23658 10996 23664 11008
rect 23492 10968 23664 10996
rect 23658 10956 23664 10968
rect 23716 10956 23722 11008
rect 23842 10996 23848 11008
rect 23803 10968 23848 10996
rect 23842 10956 23848 10968
rect 23900 10956 23906 11008
rect 26326 10956 26332 11008
rect 26384 10996 26390 11008
rect 27246 10996 27252 11008
rect 26384 10968 27252 10996
rect 26384 10956 26390 10968
rect 27246 10956 27252 10968
rect 27304 10956 27310 11008
rect 27706 10996 27712 11008
rect 27667 10968 27712 10996
rect 27706 10956 27712 10968
rect 27764 10956 27770 11008
rect 28718 10956 28724 11008
rect 28776 10996 28782 11008
rect 28776 10968 28821 10996
rect 28776 10956 28782 10968
rect 30006 10956 30012 11008
rect 30064 10996 30070 11008
rect 30484 10996 30512 11095
rect 32398 11092 32404 11144
rect 32456 11132 32462 11144
rect 32677 11135 32735 11141
rect 32677 11132 32689 11135
rect 32456 11104 32689 11132
rect 32456 11092 32462 11104
rect 32677 11101 32689 11104
rect 32723 11132 32735 11135
rect 32950 11132 32956 11144
rect 32723 11104 32956 11132
rect 32723 11101 32735 11104
rect 32677 11095 32735 11101
rect 32950 11092 32956 11104
rect 33008 11092 33014 11144
rect 33134 11092 33140 11144
rect 33192 11132 33198 11144
rect 33505 11135 33563 11141
rect 33505 11132 33517 11135
rect 33192 11104 33517 11132
rect 33192 11092 33198 11104
rect 33505 11101 33517 11104
rect 33551 11101 33563 11135
rect 41386 11132 41414 11172
rect 47210 11132 47216 11144
rect 41386 11104 47216 11132
rect 33505 11095 33563 11101
rect 47210 11092 47216 11104
rect 47268 11092 47274 11144
rect 48038 11132 48044 11144
rect 47999 11104 48044 11132
rect 48038 11092 48044 11104
rect 48096 11092 48102 11144
rect 32861 11067 32919 11073
rect 32861 11033 32873 11067
rect 32907 11064 32919 11067
rect 33410 11064 33416 11076
rect 32907 11036 33416 11064
rect 32907 11033 32919 11036
rect 32861 11027 32919 11033
rect 33410 11024 33416 11036
rect 33468 11024 33474 11076
rect 30064 10968 30512 10996
rect 30064 10956 30070 10968
rect 32582 10956 32588 11008
rect 32640 10996 32646 11008
rect 33045 10999 33103 11005
rect 33045 10996 33057 10999
rect 32640 10968 33057 10996
rect 32640 10956 32646 10968
rect 33045 10965 33057 10968
rect 33091 10965 33103 10999
rect 33045 10959 33103 10965
rect 33597 10999 33655 11005
rect 33597 10965 33609 10999
rect 33643 10996 33655 10999
rect 33778 10996 33784 11008
rect 33643 10968 33784 10996
rect 33643 10965 33655 10968
rect 33597 10959 33655 10965
rect 33778 10956 33784 10968
rect 33836 10956 33842 11008
rect 47302 10996 47308 11008
rect 47263 10968 47308 10996
rect 47302 10956 47308 10968
rect 47360 10956 47366 11008
rect 1104 10906 48852 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 48852 10906
rect 1104 10832 48852 10854
rect 20622 10792 20628 10804
rect 18708 10764 20628 10792
rect 18708 10724 18736 10764
rect 20622 10752 20628 10764
rect 20680 10752 20686 10804
rect 26234 10792 26240 10804
rect 22112 10764 25636 10792
rect 18616 10696 18736 10724
rect 19880 10727 19938 10733
rect 2130 10656 2136 10668
rect 2091 10628 2136 10656
rect 2130 10616 2136 10628
rect 2188 10616 2194 10668
rect 18616 10665 18644 10696
rect 19880 10693 19892 10727
rect 19926 10724 19938 10727
rect 20438 10724 20444 10736
rect 19926 10696 20444 10724
rect 19926 10693 19938 10696
rect 19880 10687 19938 10693
rect 20438 10684 20444 10696
rect 20496 10684 20502 10736
rect 18601 10659 18659 10665
rect 18601 10625 18613 10659
rect 18647 10625 18659 10659
rect 18601 10619 18659 10625
rect 18693 10659 18751 10665
rect 18693 10625 18705 10659
rect 18739 10625 18751 10659
rect 18693 10619 18751 10625
rect 18708 10588 18736 10619
rect 18782 10616 18788 10668
rect 18840 10656 18846 10668
rect 18969 10659 19027 10665
rect 18840 10628 18885 10656
rect 18840 10616 18846 10628
rect 18969 10625 18981 10659
rect 19015 10656 19027 10659
rect 19058 10656 19064 10668
rect 19015 10628 19064 10656
rect 19015 10625 19027 10628
rect 18969 10619 19027 10625
rect 19058 10616 19064 10628
rect 19116 10616 19122 10668
rect 19334 10616 19340 10668
rect 19392 10656 19398 10668
rect 22112 10665 22140 10764
rect 23474 10724 23480 10736
rect 23032 10696 23480 10724
rect 23032 10668 23060 10696
rect 23474 10684 23480 10696
rect 23532 10724 23538 10736
rect 25222 10724 25228 10736
rect 23532 10696 25228 10724
rect 23532 10684 23538 10696
rect 25222 10684 25228 10696
rect 25280 10684 25286 10736
rect 19613 10659 19671 10665
rect 19613 10656 19625 10659
rect 19392 10628 19625 10656
rect 19392 10616 19398 10628
rect 19613 10625 19625 10628
rect 19659 10625 19671 10659
rect 19613 10619 19671 10625
rect 22097 10659 22155 10665
rect 22097 10625 22109 10659
rect 22143 10625 22155 10659
rect 22097 10619 22155 10625
rect 22189 10659 22247 10665
rect 22189 10625 22201 10659
rect 22235 10625 22247 10659
rect 22189 10619 22247 10625
rect 18616 10560 18736 10588
rect 18616 10532 18644 10560
rect 18598 10480 18604 10532
rect 18656 10480 18662 10532
rect 20622 10480 20628 10532
rect 20680 10520 20686 10532
rect 20993 10523 21051 10529
rect 20993 10520 21005 10523
rect 20680 10492 21005 10520
rect 20680 10480 20686 10492
rect 20993 10489 21005 10492
rect 21039 10520 21051 10523
rect 22002 10520 22008 10532
rect 21039 10492 22008 10520
rect 21039 10489 21051 10492
rect 20993 10483 21051 10489
rect 22002 10480 22008 10492
rect 22060 10480 22066 10532
rect 22204 10520 22232 10619
rect 22278 10616 22284 10668
rect 22336 10656 22342 10668
rect 22336 10628 22381 10656
rect 22336 10616 22342 10628
rect 22462 10616 22468 10668
rect 22520 10656 22526 10668
rect 23014 10656 23020 10668
rect 22520 10628 22784 10656
rect 22975 10628 23020 10656
rect 22520 10616 22526 10628
rect 22278 10520 22284 10532
rect 22204 10492 22284 10520
rect 22278 10480 22284 10492
rect 22336 10480 22342 10532
rect 1394 10412 1400 10464
rect 1452 10452 1458 10464
rect 1673 10455 1731 10461
rect 1673 10452 1685 10455
rect 1452 10424 1685 10452
rect 1452 10412 1458 10424
rect 1673 10421 1685 10424
rect 1719 10421 1731 10455
rect 2222 10452 2228 10464
rect 2183 10424 2228 10452
rect 1673 10415 1731 10421
rect 2222 10412 2228 10424
rect 2280 10412 2286 10464
rect 2958 10452 2964 10464
rect 2919 10424 2964 10452
rect 2958 10412 2964 10424
rect 3016 10412 3022 10464
rect 18322 10452 18328 10464
rect 18283 10424 18328 10452
rect 18322 10412 18328 10424
rect 18380 10412 18386 10464
rect 18414 10412 18420 10464
rect 18472 10452 18478 10464
rect 19058 10452 19064 10464
rect 18472 10424 19064 10452
rect 18472 10412 18478 10424
rect 19058 10412 19064 10424
rect 19116 10412 19122 10464
rect 21818 10452 21824 10464
rect 21779 10424 21824 10452
rect 21818 10412 21824 10424
rect 21876 10412 21882 10464
rect 22756 10452 22784 10628
rect 23014 10616 23020 10628
rect 23072 10616 23078 10668
rect 23284 10659 23342 10665
rect 23284 10625 23296 10659
rect 23330 10656 23342 10659
rect 23842 10656 23848 10668
rect 23330 10628 23848 10656
rect 23330 10625 23342 10628
rect 23284 10619 23342 10625
rect 23842 10616 23848 10628
rect 23900 10616 23906 10668
rect 24854 10656 24860 10668
rect 24815 10628 24860 10656
rect 24854 10616 24860 10628
rect 24912 10616 24918 10668
rect 25041 10659 25099 10665
rect 25041 10625 25053 10659
rect 25087 10656 25099 10659
rect 25498 10656 25504 10668
rect 25087 10628 25504 10656
rect 25087 10625 25099 10628
rect 25041 10619 25099 10625
rect 25498 10616 25504 10628
rect 25556 10616 25562 10668
rect 24946 10548 24952 10600
rect 25004 10588 25010 10600
rect 25225 10591 25283 10597
rect 25225 10588 25237 10591
rect 25004 10560 25237 10588
rect 25004 10548 25010 10560
rect 25225 10557 25237 10560
rect 25271 10557 25283 10591
rect 25225 10551 25283 10557
rect 23382 10452 23388 10464
rect 22756 10424 23388 10452
rect 23382 10412 23388 10424
rect 23440 10412 23446 10464
rect 23658 10412 23664 10464
rect 23716 10452 23722 10464
rect 24397 10455 24455 10461
rect 24397 10452 24409 10455
rect 23716 10424 24409 10452
rect 23716 10412 23722 10424
rect 24397 10421 24409 10424
rect 24443 10452 24455 10455
rect 24486 10452 24492 10464
rect 24443 10424 24492 10452
rect 24443 10421 24455 10424
rect 24397 10415 24455 10421
rect 24486 10412 24492 10424
rect 24544 10412 24550 10464
rect 25608 10452 25636 10764
rect 25884 10764 26240 10792
rect 25884 10724 25912 10764
rect 26234 10752 26240 10764
rect 26292 10752 26298 10804
rect 26418 10792 26424 10804
rect 26379 10764 26424 10792
rect 26418 10752 26424 10764
rect 26476 10752 26482 10804
rect 27154 10752 27160 10804
rect 27212 10752 27218 10804
rect 27985 10795 28043 10801
rect 27985 10761 27997 10795
rect 28031 10792 28043 10795
rect 28626 10792 28632 10804
rect 28031 10764 28632 10792
rect 28031 10761 28043 10764
rect 27985 10755 28043 10761
rect 28626 10752 28632 10764
rect 28684 10752 28690 10804
rect 32398 10752 32404 10804
rect 32456 10752 32462 10804
rect 32490 10752 32496 10804
rect 32548 10752 32554 10804
rect 32582 10752 32588 10804
rect 32640 10752 32646 10804
rect 26694 10724 26700 10736
rect 25700 10696 25912 10724
rect 26068 10696 26700 10724
rect 25700 10665 25728 10696
rect 25685 10659 25743 10665
rect 25685 10625 25697 10659
rect 25731 10625 25743 10659
rect 25685 10619 25743 10625
rect 25866 10616 25872 10668
rect 25924 10656 25930 10668
rect 26068 10665 26096 10696
rect 26694 10684 26700 10696
rect 26752 10724 26758 10736
rect 27172 10724 27200 10752
rect 28997 10727 29055 10733
rect 28997 10724 29009 10727
rect 26752 10696 27108 10724
rect 27172 10696 29009 10724
rect 26752 10684 26758 10696
rect 26053 10659 26111 10665
rect 25924 10628 25969 10656
rect 25924 10616 25930 10628
rect 26053 10625 26065 10659
rect 26099 10625 26111 10659
rect 26234 10656 26240 10668
rect 26195 10628 26240 10656
rect 26053 10619 26111 10625
rect 26234 10616 26240 10628
rect 26292 10616 26298 10668
rect 26970 10656 26976 10668
rect 26931 10628 26976 10656
rect 26970 10616 26976 10628
rect 27028 10616 27034 10668
rect 27080 10656 27108 10696
rect 28997 10693 29009 10696
rect 29043 10693 29055 10727
rect 28997 10687 29055 10693
rect 27157 10659 27215 10665
rect 27157 10656 27169 10659
rect 27080 10628 27169 10656
rect 27157 10625 27169 10628
rect 27203 10625 27215 10659
rect 27157 10619 27215 10625
rect 27617 10659 27675 10665
rect 27617 10625 27629 10659
rect 27663 10656 27675 10659
rect 27982 10656 27988 10668
rect 27663 10628 27988 10656
rect 27663 10625 27675 10628
rect 27617 10619 27675 10625
rect 27982 10616 27988 10628
rect 28040 10616 28046 10668
rect 32416 10665 32444 10752
rect 32508 10665 32536 10752
rect 32600 10671 32628 10752
rect 47946 10724 47952 10736
rect 33152 10696 47952 10724
rect 32585 10665 32643 10671
rect 32381 10659 32444 10665
rect 32381 10625 32393 10659
rect 32427 10628 32444 10659
rect 32490 10659 32548 10665
rect 32427 10625 32439 10628
rect 32381 10619 32439 10625
rect 32490 10625 32502 10659
rect 32536 10625 32548 10659
rect 32585 10631 32597 10665
rect 32631 10631 32643 10665
rect 32766 10656 32772 10668
rect 32585 10625 32643 10631
rect 32727 10628 32772 10656
rect 32490 10619 32548 10625
rect 32766 10616 32772 10628
rect 32824 10616 32830 10668
rect 25961 10591 26019 10597
rect 25961 10557 25973 10591
rect 26007 10557 26019 10591
rect 25961 10551 26019 10557
rect 25976 10520 26004 10551
rect 26786 10548 26792 10600
rect 26844 10588 26850 10600
rect 27709 10591 27767 10597
rect 27709 10588 27721 10591
rect 26844 10560 27721 10588
rect 26844 10548 26850 10560
rect 27709 10557 27721 10560
rect 27755 10557 27767 10591
rect 33152 10588 33180 10696
rect 47946 10684 47952 10696
rect 48004 10684 48010 10736
rect 33410 10616 33416 10668
rect 33468 10656 33474 10668
rect 33597 10659 33655 10665
rect 33597 10656 33609 10659
rect 33468 10628 33609 10656
rect 33468 10616 33474 10628
rect 33597 10625 33609 10628
rect 33643 10625 33655 10659
rect 33597 10619 33655 10625
rect 35437 10659 35495 10665
rect 35437 10625 35449 10659
rect 35483 10656 35495 10659
rect 40678 10656 40684 10668
rect 35483 10628 40684 10656
rect 35483 10625 35495 10628
rect 35437 10619 35495 10625
rect 40678 10616 40684 10628
rect 40736 10616 40742 10668
rect 47762 10656 47768 10668
rect 47723 10628 47768 10656
rect 47762 10616 47768 10628
rect 47820 10616 47826 10668
rect 33778 10588 33784 10600
rect 27709 10551 27767 10557
rect 27816 10560 33180 10588
rect 33739 10560 33784 10588
rect 27065 10523 27123 10529
rect 27065 10520 27077 10523
rect 25976 10492 27077 10520
rect 27065 10489 27077 10492
rect 27111 10489 27123 10523
rect 27816 10520 27844 10560
rect 33778 10548 33784 10560
rect 33836 10548 33842 10600
rect 27065 10483 27123 10489
rect 27632 10492 27844 10520
rect 29181 10523 29239 10529
rect 27632 10452 27660 10492
rect 29181 10489 29193 10523
rect 29227 10520 29239 10523
rect 30006 10520 30012 10532
rect 29227 10492 30012 10520
rect 29227 10489 29239 10492
rect 29181 10483 29239 10489
rect 30006 10480 30012 10492
rect 30064 10480 30070 10532
rect 47949 10523 48007 10529
rect 47949 10520 47961 10523
rect 31726 10492 47961 10520
rect 27798 10452 27804 10464
rect 25608 10424 27660 10452
rect 27759 10424 27804 10452
rect 27798 10412 27804 10424
rect 27856 10412 27862 10464
rect 27890 10412 27896 10464
rect 27948 10452 27954 10464
rect 31726 10452 31754 10492
rect 47949 10489 47961 10492
rect 47995 10489 48007 10523
rect 47949 10483 48007 10489
rect 27948 10424 31754 10452
rect 32125 10455 32183 10461
rect 27948 10412 27954 10424
rect 32125 10421 32137 10455
rect 32171 10452 32183 10455
rect 32490 10452 32496 10464
rect 32171 10424 32496 10452
rect 32171 10421 32183 10424
rect 32125 10415 32183 10421
rect 32490 10412 32496 10424
rect 32548 10412 32554 10464
rect 1104 10362 48852 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 48852 10362
rect 1104 10288 48852 10310
rect 18782 10208 18788 10260
rect 18840 10248 18846 10260
rect 19613 10251 19671 10257
rect 19613 10248 19625 10251
rect 18840 10220 19625 10248
rect 18840 10208 18846 10220
rect 19613 10217 19625 10220
rect 19659 10217 19671 10251
rect 22370 10248 22376 10260
rect 22331 10220 22376 10248
rect 19613 10211 19671 10217
rect 22370 10208 22376 10220
rect 22428 10208 22434 10260
rect 25222 10208 25228 10260
rect 25280 10248 25286 10260
rect 26053 10251 26111 10257
rect 26053 10248 26065 10251
rect 25280 10220 26065 10248
rect 25280 10208 25286 10220
rect 26053 10217 26065 10220
rect 26099 10217 26111 10251
rect 26053 10211 26111 10217
rect 27706 10208 27712 10260
rect 27764 10248 27770 10260
rect 27801 10251 27859 10257
rect 27801 10248 27813 10251
rect 27764 10220 27813 10248
rect 27764 10208 27770 10220
rect 27801 10217 27813 10220
rect 27847 10248 27859 10251
rect 27847 10220 28304 10248
rect 27847 10217 27859 10220
rect 27801 10211 27859 10217
rect 22388 10180 22416 10208
rect 25406 10180 25412 10192
rect 22388 10152 25412 10180
rect 25406 10140 25412 10152
rect 25464 10140 25470 10192
rect 25590 10140 25596 10192
rect 25648 10180 25654 10192
rect 27430 10180 27436 10192
rect 25648 10152 27436 10180
rect 25648 10140 25654 10152
rect 27430 10140 27436 10152
rect 27488 10140 27494 10192
rect 1394 10112 1400 10124
rect 1355 10084 1400 10112
rect 1394 10072 1400 10084
rect 1452 10072 1458 10124
rect 1581 10115 1639 10121
rect 1581 10081 1593 10115
rect 1627 10112 1639 10115
rect 2222 10112 2228 10124
rect 1627 10084 2228 10112
rect 1627 10081 1639 10084
rect 1581 10075 1639 10081
rect 2222 10072 2228 10084
rect 2280 10072 2286 10124
rect 2774 10112 2780 10124
rect 2735 10084 2780 10112
rect 2774 10072 2780 10084
rect 2832 10072 2838 10124
rect 17034 10112 17040 10124
rect 16995 10084 17040 10112
rect 17034 10072 17040 10084
rect 17092 10072 17098 10124
rect 19334 10072 19340 10124
rect 19392 10112 19398 10124
rect 20993 10115 21051 10121
rect 20993 10112 21005 10115
rect 19392 10084 21005 10112
rect 19392 10072 19398 10084
rect 20993 10081 21005 10084
rect 21039 10081 21051 10115
rect 20993 10075 21051 10081
rect 23569 10115 23627 10121
rect 23569 10081 23581 10115
rect 23615 10112 23627 10115
rect 23658 10112 23664 10124
rect 23615 10084 23664 10112
rect 23615 10081 23627 10084
rect 23569 10075 23627 10081
rect 23658 10072 23664 10084
rect 23716 10072 23722 10124
rect 23753 10115 23811 10121
rect 23753 10081 23765 10115
rect 23799 10112 23811 10115
rect 24118 10112 24124 10124
rect 23799 10084 24124 10112
rect 23799 10081 23811 10084
rect 23753 10075 23811 10081
rect 24118 10072 24124 10084
rect 24176 10072 24182 10124
rect 24946 10072 24952 10124
rect 25004 10112 25010 10124
rect 25225 10115 25283 10121
rect 25225 10112 25237 10115
rect 25004 10084 25237 10112
rect 25004 10072 25010 10084
rect 25225 10081 25237 10084
rect 25271 10081 25283 10115
rect 26234 10112 26240 10124
rect 25225 10075 25283 10081
rect 25884 10084 26240 10112
rect 17304 10047 17362 10053
rect 17304 10013 17316 10047
rect 17350 10044 17362 10047
rect 18322 10044 18328 10056
rect 17350 10016 18328 10044
rect 17350 10013 17362 10016
rect 17304 10007 17362 10013
rect 18322 10004 18328 10016
rect 18380 10004 18386 10056
rect 20349 10047 20407 10053
rect 20349 10013 20361 10047
rect 20395 10044 20407 10047
rect 20438 10044 20444 10056
rect 20395 10016 20444 10044
rect 20395 10013 20407 10016
rect 20349 10007 20407 10013
rect 20438 10004 20444 10016
rect 20496 10004 20502 10056
rect 21260 10047 21318 10053
rect 21260 10013 21272 10047
rect 21306 10044 21318 10047
rect 21818 10044 21824 10056
rect 21306 10016 21824 10044
rect 21306 10013 21318 10016
rect 21260 10007 21318 10013
rect 21818 10004 21824 10016
rect 21876 10004 21882 10056
rect 22002 10004 22008 10056
rect 22060 10044 22066 10056
rect 25041 10047 25099 10053
rect 25041 10044 25053 10047
rect 22060 10016 25053 10044
rect 22060 10004 22066 10016
rect 25041 10013 25053 10016
rect 25087 10044 25099 10047
rect 25884 10044 25912 10084
rect 26234 10072 26240 10084
rect 26292 10072 26298 10124
rect 28276 10121 28304 10220
rect 28718 10208 28724 10260
rect 28776 10248 28782 10260
rect 28905 10251 28963 10257
rect 28905 10248 28917 10251
rect 28776 10220 28917 10248
rect 28776 10208 28782 10220
rect 28905 10217 28917 10220
rect 28951 10217 28963 10251
rect 28905 10211 28963 10217
rect 33410 10208 33416 10260
rect 33468 10248 33474 10260
rect 33781 10251 33839 10257
rect 33781 10248 33793 10251
rect 33468 10220 33793 10248
rect 33468 10208 33474 10220
rect 33781 10217 33793 10220
rect 33827 10217 33839 10251
rect 33781 10211 33839 10217
rect 48038 10180 48044 10192
rect 46308 10152 48044 10180
rect 28261 10115 28319 10121
rect 28261 10081 28273 10115
rect 28307 10081 28319 10115
rect 28261 10075 28319 10081
rect 28629 10115 28687 10121
rect 28629 10081 28641 10115
rect 28675 10112 28687 10115
rect 28902 10112 28908 10124
rect 28675 10084 28908 10112
rect 28675 10081 28687 10084
rect 28629 10075 28687 10081
rect 28902 10072 28908 10084
rect 28960 10072 28966 10124
rect 29454 10072 29460 10124
rect 29512 10112 29518 10124
rect 46308 10121 46336 10152
rect 48038 10140 48044 10152
rect 48096 10140 48102 10192
rect 30101 10115 30159 10121
rect 30101 10112 30113 10115
rect 29512 10084 30113 10112
rect 29512 10072 29518 10084
rect 30101 10081 30113 10084
rect 30147 10081 30159 10115
rect 30101 10075 30159 10081
rect 46293 10115 46351 10121
rect 46293 10081 46305 10115
rect 46339 10081 46351 10115
rect 46293 10075 46351 10081
rect 46477 10115 46535 10121
rect 46477 10081 46489 10115
rect 46523 10112 46535 10115
rect 47302 10112 47308 10124
rect 46523 10084 47308 10112
rect 46523 10081 46535 10084
rect 46477 10075 46535 10081
rect 47302 10072 47308 10084
rect 47360 10072 47366 10124
rect 48130 10112 48136 10124
rect 48091 10084 48136 10112
rect 48130 10072 48136 10084
rect 48188 10072 48194 10124
rect 25087 10016 25912 10044
rect 25961 10047 26019 10053
rect 25087 10013 25099 10016
rect 25041 10007 25099 10013
rect 25961 10013 25973 10047
rect 26007 10044 26019 10047
rect 27154 10044 27160 10056
rect 26007 10016 27160 10044
rect 26007 10013 26019 10016
rect 25961 10007 26019 10013
rect 27154 10004 27160 10016
rect 27212 10004 27218 10056
rect 27433 10047 27491 10053
rect 27433 10013 27445 10047
rect 27479 10044 27491 10047
rect 27798 10044 27804 10056
rect 27479 10016 27804 10044
rect 27479 10013 27491 10016
rect 27433 10007 27491 10013
rect 27798 10004 27804 10016
rect 27856 10044 27862 10056
rect 28074 10044 28080 10056
rect 27856 10016 28080 10044
rect 27856 10004 27862 10016
rect 28074 10004 28080 10016
rect 28132 10004 28138 10056
rect 28721 10047 28779 10053
rect 28721 10013 28733 10047
rect 28767 10013 28779 10047
rect 29914 10044 29920 10056
rect 29875 10016 29920 10044
rect 28721 10007 28779 10013
rect 19242 9976 19248 9988
rect 19203 9948 19248 9976
rect 19242 9936 19248 9948
rect 19300 9936 19306 9988
rect 19429 9979 19487 9985
rect 19429 9945 19441 9979
rect 19475 9945 19487 9979
rect 19429 9939 19487 9945
rect 20533 9979 20591 9985
rect 20533 9945 20545 9979
rect 20579 9976 20591 9979
rect 22278 9976 22284 9988
rect 20579 9948 22284 9976
rect 20579 9945 20591 9948
rect 20533 9939 20591 9945
rect 18414 9908 18420 9920
rect 18327 9880 18420 9908
rect 18414 9868 18420 9880
rect 18472 9908 18478 9920
rect 19444 9908 19472 9939
rect 22278 9936 22284 9948
rect 22336 9936 22342 9988
rect 23477 9979 23535 9985
rect 23477 9945 23489 9979
rect 23523 9976 23535 9979
rect 23842 9976 23848 9988
rect 23523 9948 23848 9976
rect 23523 9945 23535 9948
rect 23477 9939 23535 9945
rect 23842 9936 23848 9948
rect 23900 9976 23906 9988
rect 24026 9976 24032 9988
rect 23900 9948 24032 9976
rect 23900 9936 23906 9948
rect 24026 9936 24032 9948
rect 24084 9936 24090 9988
rect 24578 9936 24584 9988
rect 24636 9976 24642 9988
rect 26786 9976 26792 9988
rect 24636 9948 25268 9976
rect 26747 9948 26792 9976
rect 24636 9936 24642 9948
rect 18472 9880 19472 9908
rect 23109 9911 23167 9917
rect 18472 9868 18478 9880
rect 23109 9877 23121 9911
rect 23155 9908 23167 9911
rect 23290 9908 23296 9920
rect 23155 9880 23296 9908
rect 23155 9877 23167 9880
rect 23109 9871 23167 9877
rect 23290 9868 23296 9880
rect 23348 9868 23354 9920
rect 24673 9911 24731 9917
rect 24673 9877 24685 9911
rect 24719 9908 24731 9911
rect 24762 9908 24768 9920
rect 24719 9880 24768 9908
rect 24719 9877 24731 9880
rect 24673 9871 24731 9877
rect 24762 9868 24768 9880
rect 24820 9868 24826 9920
rect 25130 9908 25136 9920
rect 25091 9880 25136 9908
rect 25130 9868 25136 9880
rect 25188 9868 25194 9920
rect 25240 9908 25268 9948
rect 26786 9936 26792 9948
rect 26844 9936 26850 9988
rect 26970 9936 26976 9988
rect 27028 9976 27034 9988
rect 27614 9976 27620 9988
rect 27028 9948 27620 9976
rect 27028 9936 27034 9948
rect 27614 9936 27620 9948
rect 27672 9936 27678 9988
rect 27706 9936 27712 9988
rect 27764 9976 27770 9988
rect 28736 9976 28764 10007
rect 29914 10004 29920 10016
rect 29972 10004 29978 10056
rect 30006 10004 30012 10056
rect 30064 10044 30070 10056
rect 32401 10047 32459 10053
rect 32401 10044 32413 10047
rect 30064 10016 32413 10044
rect 30064 10004 30070 10016
rect 32401 10013 32413 10016
rect 32447 10013 32459 10047
rect 32401 10007 32459 10013
rect 32490 10004 32496 10056
rect 32548 10044 32554 10056
rect 32657 10047 32715 10053
rect 32657 10044 32669 10047
rect 32548 10016 32669 10044
rect 32548 10004 32554 10016
rect 32657 10013 32669 10016
rect 32703 10013 32715 10047
rect 32657 10007 32715 10013
rect 27764 9948 29592 9976
rect 27764 9936 27770 9948
rect 27890 9908 27896 9920
rect 25240 9880 27896 9908
rect 27890 9868 27896 9880
rect 27948 9868 27954 9920
rect 29564 9917 29592 9948
rect 29549 9911 29607 9917
rect 29549 9877 29561 9911
rect 29595 9877 29607 9911
rect 29549 9871 29607 9877
rect 29822 9868 29828 9920
rect 29880 9908 29886 9920
rect 30009 9911 30067 9917
rect 30009 9908 30021 9911
rect 29880 9880 30021 9908
rect 29880 9868 29886 9880
rect 30009 9877 30021 9880
rect 30055 9877 30067 9911
rect 30009 9871 30067 9877
rect 1104 9818 48852 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 48852 9818
rect 1104 9744 48852 9766
rect 24854 9704 24860 9716
rect 24815 9676 24860 9704
rect 24854 9664 24860 9676
rect 24912 9664 24918 9716
rect 29914 9664 29920 9716
rect 29972 9664 29978 9716
rect 32122 9704 32128 9716
rect 31404 9676 32128 9704
rect 2958 9636 2964 9648
rect 1780 9608 2964 9636
rect 1780 9577 1808 9608
rect 2958 9596 2964 9608
rect 3016 9596 3022 9648
rect 3418 9596 3424 9648
rect 3476 9636 3482 9648
rect 12434 9636 12440 9648
rect 3476 9608 12440 9636
rect 3476 9596 3482 9608
rect 12434 9596 12440 9608
rect 12492 9596 12498 9648
rect 18414 9636 18420 9648
rect 17604 9608 18420 9636
rect 17604 9577 17632 9608
rect 18414 9596 18420 9608
rect 18472 9596 18478 9648
rect 23750 9596 23756 9648
rect 23808 9636 23814 9648
rect 24213 9639 24271 9645
rect 24213 9636 24225 9639
rect 23808 9608 24225 9636
rect 23808 9596 23814 9608
rect 24213 9605 24225 9608
rect 24259 9605 24271 9639
rect 24394 9636 24400 9648
rect 24213 9599 24271 9605
rect 24320 9608 24400 9636
rect 1765 9571 1823 9577
rect 1765 9537 1777 9571
rect 1811 9537 1823 9571
rect 1765 9531 1823 9537
rect 17589 9571 17647 9577
rect 17589 9537 17601 9571
rect 17635 9537 17647 9571
rect 23198 9568 23204 9580
rect 23159 9540 23204 9568
rect 17589 9531 17647 9537
rect 23198 9528 23204 9540
rect 23256 9528 23262 9580
rect 1946 9500 1952 9512
rect 1907 9472 1952 9500
rect 1946 9460 1952 9472
rect 2004 9460 2010 9512
rect 2774 9500 2780 9512
rect 2735 9472 2780 9500
rect 2774 9460 2780 9472
rect 2832 9460 2838 9512
rect 17770 9500 17776 9512
rect 17731 9472 17776 9500
rect 17770 9460 17776 9472
rect 17828 9460 17834 9512
rect 17926 9472 18184 9500
rect 17926 9432 17954 9472
rect 6886 9404 17954 9432
rect 18156 9432 18184 9472
rect 18230 9460 18236 9512
rect 18288 9500 18294 9512
rect 23290 9500 23296 9512
rect 18288 9472 18333 9500
rect 23251 9472 23296 9500
rect 18288 9460 18294 9472
rect 23290 9460 23296 9472
rect 23348 9460 23354 9512
rect 23569 9503 23627 9509
rect 23569 9469 23581 9503
rect 23615 9500 23627 9503
rect 24320 9500 24348 9608
rect 24394 9596 24400 9608
rect 24452 9596 24458 9648
rect 24762 9596 24768 9648
rect 24820 9636 24826 9648
rect 25317 9639 25375 9645
rect 25317 9636 25329 9639
rect 24820 9608 25329 9636
rect 24820 9596 24826 9608
rect 25317 9605 25329 9608
rect 25363 9605 25375 9639
rect 25317 9599 25375 9605
rect 25406 9596 25412 9648
rect 25464 9636 25470 9648
rect 29932 9636 29960 9664
rect 31404 9636 31432 9676
rect 32122 9664 32128 9676
rect 32180 9704 32186 9716
rect 32180 9676 32904 9704
rect 32180 9664 32186 9676
rect 25464 9608 28994 9636
rect 29932 9608 31432 9636
rect 31481 9639 31539 9645
rect 25464 9596 25470 9608
rect 24486 9568 24492 9580
rect 24447 9540 24492 9568
rect 24486 9528 24492 9540
rect 24544 9528 24550 9580
rect 24578 9528 24584 9580
rect 24636 9568 24642 9580
rect 24673 9571 24731 9577
rect 24673 9568 24685 9571
rect 24636 9540 24685 9568
rect 24636 9528 24642 9540
rect 24673 9537 24685 9540
rect 24719 9537 24731 9571
rect 24673 9531 24731 9537
rect 24854 9528 24860 9580
rect 24912 9568 24918 9580
rect 25593 9571 25651 9577
rect 25593 9568 25605 9571
rect 24912 9540 25605 9568
rect 24912 9528 24918 9540
rect 25593 9537 25605 9540
rect 25639 9537 25651 9571
rect 25593 9531 25651 9537
rect 27154 9528 27160 9580
rect 27212 9568 27218 9580
rect 27801 9571 27859 9577
rect 27801 9568 27813 9571
rect 27212 9540 27813 9568
rect 27212 9528 27218 9540
rect 27801 9537 27813 9540
rect 27847 9537 27859 9571
rect 27982 9568 27988 9580
rect 27943 9540 27988 9568
rect 27801 9531 27859 9537
rect 27982 9528 27988 9540
rect 28040 9528 28046 9580
rect 28077 9571 28135 9577
rect 28077 9537 28089 9571
rect 28123 9568 28135 9571
rect 28534 9568 28540 9580
rect 28123 9540 28540 9568
rect 28123 9537 28135 9540
rect 28077 9531 28135 9537
rect 28534 9528 28540 9540
rect 28592 9528 28598 9580
rect 28966 9568 28994 9608
rect 31481 9605 31493 9639
rect 31527 9636 31539 9639
rect 32769 9639 32827 9645
rect 32769 9636 32781 9639
rect 31527 9608 32781 9636
rect 31527 9605 31539 9608
rect 31481 9599 31539 9605
rect 32769 9605 32781 9608
rect 32815 9605 32827 9639
rect 32876 9636 32904 9676
rect 36538 9636 36544 9648
rect 32876 9608 36544 9636
rect 32769 9599 32827 9605
rect 36538 9596 36544 9608
rect 36596 9596 36602 9648
rect 29089 9571 29147 9577
rect 29089 9568 29101 9571
rect 28966 9540 29101 9568
rect 29089 9537 29101 9540
rect 29135 9537 29147 9571
rect 29089 9531 29147 9537
rect 29181 9571 29239 9577
rect 29181 9537 29193 9571
rect 29227 9568 29239 9571
rect 29227 9540 29868 9568
rect 29227 9537 29239 9540
rect 29181 9531 29239 9537
rect 23615 9472 24348 9500
rect 23615 9469 23627 9472
rect 23569 9463 23627 9469
rect 24394 9460 24400 9512
rect 24452 9500 24458 9512
rect 25130 9500 25136 9512
rect 24452 9472 25136 9500
rect 24452 9460 24458 9472
rect 25130 9460 25136 9472
rect 25188 9460 25194 9512
rect 25406 9500 25412 9512
rect 25367 9472 25412 9500
rect 25406 9460 25412 9472
rect 25464 9460 25470 9512
rect 29104 9500 29132 9531
rect 29365 9503 29423 9509
rect 29104 9472 29224 9500
rect 28994 9432 29000 9444
rect 18156 9404 29000 9432
rect 658 9324 664 9376
rect 716 9364 722 9376
rect 6886 9364 6914 9404
rect 28994 9392 29000 9404
rect 29052 9392 29058 9444
rect 29196 9432 29224 9472
rect 29365 9469 29377 9503
rect 29411 9500 29423 9503
rect 29454 9500 29460 9512
rect 29411 9472 29460 9500
rect 29411 9469 29423 9472
rect 29365 9463 29423 9469
rect 29454 9460 29460 9472
rect 29512 9460 29518 9512
rect 29840 9500 29868 9540
rect 29914 9528 29920 9580
rect 29972 9568 29978 9580
rect 29972 9540 30017 9568
rect 29972 9528 29978 9540
rect 30098 9528 30104 9580
rect 30156 9568 30162 9580
rect 30282 9568 30288 9580
rect 30156 9540 30201 9568
rect 30243 9540 30288 9568
rect 30156 9528 30162 9540
rect 30282 9528 30288 9540
rect 30340 9528 30346 9580
rect 30469 9571 30527 9577
rect 30469 9537 30481 9571
rect 30515 9537 30527 9571
rect 31386 9568 31392 9580
rect 31347 9540 31392 9568
rect 30469 9531 30527 9537
rect 30190 9500 30196 9512
rect 29840 9472 30196 9500
rect 30190 9460 30196 9472
rect 30248 9460 30254 9512
rect 30484 9500 30512 9531
rect 31386 9528 31392 9540
rect 31444 9528 31450 9580
rect 32398 9500 32404 9512
rect 30291 9472 32404 9500
rect 30291 9432 30319 9472
rect 32398 9460 32404 9472
rect 32456 9460 32462 9512
rect 32585 9503 32643 9509
rect 32585 9469 32597 9503
rect 32631 9500 32643 9503
rect 32858 9500 32864 9512
rect 32631 9472 32864 9500
rect 32631 9469 32643 9472
rect 32585 9463 32643 9469
rect 32858 9460 32864 9472
rect 32916 9460 32922 9512
rect 33134 9500 33140 9512
rect 33095 9472 33140 9500
rect 33134 9460 33140 9472
rect 33192 9460 33198 9512
rect 29196 9404 30319 9432
rect 30834 9392 30840 9444
rect 30892 9432 30898 9444
rect 32674 9432 32680 9444
rect 30892 9404 32680 9432
rect 30892 9392 30898 9404
rect 32674 9392 32680 9404
rect 32732 9392 32738 9444
rect 716 9336 6914 9364
rect 716 9324 722 9336
rect 16574 9324 16580 9376
rect 16632 9364 16638 9376
rect 18230 9364 18236 9376
rect 16632 9336 18236 9364
rect 16632 9324 16638 9336
rect 18230 9324 18236 9336
rect 18288 9324 18294 9376
rect 24394 9364 24400 9376
rect 24355 9336 24400 9364
rect 24394 9324 24400 9336
rect 24452 9324 24458 9376
rect 24486 9324 24492 9376
rect 24544 9364 24550 9376
rect 25317 9367 25375 9373
rect 25317 9364 25329 9367
rect 24544 9336 25329 9364
rect 24544 9324 24550 9336
rect 25317 9333 25329 9336
rect 25363 9333 25375 9367
rect 25317 9327 25375 9333
rect 25777 9367 25835 9373
rect 25777 9333 25789 9367
rect 25823 9364 25835 9367
rect 26786 9364 26792 9376
rect 25823 9336 26792 9364
rect 25823 9333 25835 9336
rect 25777 9327 25835 9333
rect 26786 9324 26792 9336
rect 26844 9324 26850 9376
rect 26970 9324 26976 9376
rect 27028 9364 27034 9376
rect 27801 9367 27859 9373
rect 27801 9364 27813 9367
rect 27028 9336 27813 9364
rect 27028 9324 27034 9336
rect 27801 9333 27813 9336
rect 27847 9333 27859 9367
rect 27801 9327 27859 9333
rect 28534 9324 28540 9376
rect 28592 9364 28598 9376
rect 28721 9367 28779 9373
rect 28721 9364 28733 9367
rect 28592 9336 28733 9364
rect 28592 9324 28598 9336
rect 28721 9333 28733 9336
rect 28767 9333 28779 9367
rect 30650 9364 30656 9376
rect 30611 9336 30656 9364
rect 28721 9327 28779 9333
rect 30650 9324 30656 9336
rect 30708 9324 30714 9376
rect 31386 9324 31392 9376
rect 31444 9364 31450 9376
rect 33226 9364 33232 9376
rect 31444 9336 33232 9364
rect 31444 9324 31450 9336
rect 33226 9324 33232 9336
rect 33284 9324 33290 9376
rect 1104 9274 48852 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 48852 9274
rect 1104 9200 48852 9222
rect 17770 9120 17776 9172
rect 17828 9160 17834 9172
rect 18049 9163 18107 9169
rect 18049 9160 18061 9163
rect 17828 9132 18061 9160
rect 17828 9120 17834 9132
rect 18049 9129 18061 9132
rect 18095 9129 18107 9163
rect 18049 9123 18107 9129
rect 23198 9120 23204 9172
rect 23256 9160 23262 9172
rect 23845 9163 23903 9169
rect 23845 9160 23857 9163
rect 23256 9132 23857 9160
rect 23256 9120 23262 9132
rect 23845 9129 23857 9132
rect 23891 9160 23903 9163
rect 24394 9160 24400 9172
rect 23891 9132 24400 9160
rect 23891 9129 23903 9132
rect 23845 9123 23903 9129
rect 24394 9120 24400 9132
rect 24452 9160 24458 9172
rect 27890 9160 27896 9172
rect 24452 9132 24900 9160
rect 27851 9132 27896 9160
rect 24452 9120 24458 9132
rect 24762 9052 24768 9104
rect 24820 9052 24826 9104
rect 23566 8984 23572 9036
rect 23624 9024 23630 9036
rect 24486 9024 24492 9036
rect 23624 8996 24492 9024
rect 23624 8984 23630 8996
rect 24486 8984 24492 8996
rect 24544 8984 24550 9036
rect 24780 9024 24808 9052
rect 24872 9033 24900 9132
rect 27890 9120 27896 9132
rect 27948 9120 27954 9172
rect 28074 9160 28080 9172
rect 28035 9132 28080 9160
rect 28074 9120 28080 9132
rect 28132 9120 28138 9172
rect 30190 9120 30196 9172
rect 30248 9160 30254 9172
rect 31389 9163 31447 9169
rect 31389 9160 31401 9163
rect 30248 9132 31401 9160
rect 30248 9120 30254 9132
rect 31389 9129 31401 9132
rect 31435 9129 31447 9163
rect 31389 9123 31447 9129
rect 32214 9120 32220 9172
rect 32272 9160 32278 9172
rect 32674 9160 32680 9172
rect 32272 9132 32680 9160
rect 32272 9120 32278 9132
rect 32674 9120 32680 9132
rect 32732 9120 32738 9172
rect 39298 9120 39304 9172
rect 39356 9160 39362 9172
rect 46842 9160 46848 9172
rect 39356 9132 46848 9160
rect 39356 9120 39362 9132
rect 46842 9120 46848 9132
rect 46900 9120 46906 9172
rect 27065 9095 27123 9101
rect 27065 9061 27077 9095
rect 27111 9092 27123 9095
rect 29914 9092 29920 9104
rect 27111 9064 29920 9092
rect 27111 9061 27123 9064
rect 27065 9055 27123 9061
rect 29914 9052 29920 9064
rect 29972 9052 29978 9104
rect 31478 9052 31484 9104
rect 31536 9092 31542 9104
rect 48133 9095 48191 9101
rect 48133 9092 48145 9095
rect 31536 9064 48145 9092
rect 31536 9052 31542 9064
rect 48133 9061 48145 9064
rect 48179 9061 48191 9095
rect 48133 9055 48191 9061
rect 24596 8996 24808 9024
rect 24857 9027 24915 9033
rect 17954 8956 17960 8968
rect 17915 8928 17960 8956
rect 17954 8916 17960 8928
rect 18012 8916 18018 8968
rect 23290 8916 23296 8968
rect 23348 8956 23354 8968
rect 24596 8965 24624 8996
rect 24857 8993 24869 9027
rect 24903 8993 24915 9027
rect 24857 8987 24915 8993
rect 27801 9027 27859 9033
rect 27801 8993 27813 9027
rect 27847 9024 27859 9027
rect 33134 9024 33140 9036
rect 27847 8996 28580 9024
rect 27847 8993 27859 8996
rect 27801 8987 27859 8993
rect 28552 8968 28580 8996
rect 32692 8996 33140 9024
rect 24581 8959 24639 8965
rect 23348 8928 24532 8956
rect 23348 8916 23354 8928
rect 23477 8891 23535 8897
rect 23477 8857 23489 8891
rect 23523 8888 23535 8891
rect 23566 8888 23572 8900
rect 23523 8860 23572 8888
rect 23523 8857 23535 8860
rect 23477 8851 23535 8857
rect 23566 8848 23572 8860
rect 23624 8848 23630 8900
rect 23661 8891 23719 8897
rect 23661 8857 23673 8891
rect 23707 8888 23719 8891
rect 23750 8888 23756 8900
rect 23707 8860 23756 8888
rect 23707 8857 23719 8860
rect 23661 8851 23719 8857
rect 23750 8848 23756 8860
rect 23808 8848 23814 8900
rect 24504 8888 24532 8928
rect 24581 8925 24593 8959
rect 24627 8925 24639 8959
rect 24581 8919 24639 8925
rect 24765 8959 24823 8965
rect 24765 8925 24777 8959
rect 24811 8956 24823 8959
rect 25406 8956 25412 8968
rect 24811 8928 25412 8956
rect 24811 8925 24823 8928
rect 24765 8919 24823 8925
rect 24780 8888 24808 8919
rect 25406 8916 25412 8928
rect 25464 8916 25470 8968
rect 26970 8956 26976 8968
rect 26931 8928 26976 8956
rect 26970 8916 26976 8928
rect 27028 8916 27034 8968
rect 27157 8959 27215 8965
rect 27157 8925 27169 8959
rect 27203 8925 27215 8959
rect 27157 8919 27215 8925
rect 27617 8959 27675 8965
rect 27617 8925 27629 8959
rect 27663 8956 27675 8959
rect 27706 8956 27712 8968
rect 27663 8928 27712 8956
rect 27663 8925 27675 8928
rect 27617 8919 27675 8925
rect 24504 8860 24808 8888
rect 24397 8823 24455 8829
rect 24397 8789 24409 8823
rect 24443 8820 24455 8823
rect 25866 8820 25872 8832
rect 24443 8792 25872 8820
rect 24443 8789 24455 8792
rect 24397 8783 24455 8789
rect 25866 8780 25872 8792
rect 25924 8780 25930 8832
rect 27172 8820 27200 8919
rect 27706 8916 27712 8928
rect 27764 8916 27770 8968
rect 27893 8959 27951 8965
rect 27893 8956 27905 8959
rect 27816 8928 27905 8956
rect 27816 8900 27844 8928
rect 27893 8925 27905 8928
rect 27939 8925 27951 8959
rect 28534 8956 28540 8968
rect 28495 8928 28540 8956
rect 27893 8919 27951 8925
rect 28534 8916 28540 8928
rect 28592 8916 28598 8968
rect 29546 8916 29552 8968
rect 29604 8956 29610 8968
rect 30006 8956 30012 8968
rect 29604 8928 30012 8956
rect 29604 8916 29610 8928
rect 30006 8916 30012 8928
rect 30064 8916 30070 8968
rect 30276 8959 30334 8965
rect 30276 8925 30288 8959
rect 30322 8956 30334 8959
rect 30650 8956 30656 8968
rect 30322 8928 30656 8956
rect 30322 8925 30334 8928
rect 30276 8919 30334 8925
rect 30650 8916 30656 8928
rect 30708 8916 30714 8968
rect 32122 8916 32128 8968
rect 32180 8956 32186 8968
rect 32447 8959 32505 8965
rect 32447 8956 32459 8959
rect 32180 8928 32459 8956
rect 32180 8916 32186 8928
rect 32447 8925 32459 8928
rect 32493 8925 32505 8959
rect 32582 8956 32588 8968
rect 32543 8928 32588 8956
rect 32447 8919 32505 8925
rect 32582 8916 32588 8928
rect 32640 8916 32646 8968
rect 32692 8965 32720 8996
rect 33134 8984 33140 8996
rect 33192 8984 33198 9036
rect 33226 8984 33232 9036
rect 33284 8984 33290 9036
rect 32682 8959 32740 8965
rect 32682 8925 32694 8959
rect 32728 8925 32740 8959
rect 32861 8959 32919 8965
rect 32861 8956 32873 8959
rect 32682 8919 32740 8925
rect 32784 8928 32873 8956
rect 32784 8900 32812 8928
rect 32861 8925 32873 8928
rect 32907 8925 32919 8959
rect 33244 8956 33272 8984
rect 33321 8959 33379 8965
rect 33321 8956 33333 8959
rect 33244 8928 33333 8956
rect 32861 8919 32919 8925
rect 33321 8925 33333 8928
rect 33367 8925 33379 8959
rect 33321 8919 33379 8925
rect 33410 8916 33416 8968
rect 33468 8956 33474 8968
rect 46753 8959 46811 8965
rect 46753 8956 46765 8959
rect 33468 8928 33513 8956
rect 41386 8928 46765 8956
rect 33468 8916 33474 8928
rect 27798 8848 27804 8900
rect 27856 8848 27862 8900
rect 27982 8848 27988 8900
rect 28040 8888 28046 8900
rect 28626 8888 28632 8900
rect 28040 8860 28632 8888
rect 28040 8848 28046 8860
rect 28626 8848 28632 8860
rect 28684 8888 28690 8900
rect 28721 8891 28779 8897
rect 28721 8888 28733 8891
rect 28684 8860 28733 8888
rect 28684 8848 28690 8860
rect 28721 8857 28733 8860
rect 28767 8857 28779 8891
rect 28721 8851 28779 8857
rect 29454 8848 29460 8900
rect 29512 8888 29518 8900
rect 30098 8888 30104 8900
rect 29512 8860 30104 8888
rect 29512 8848 29518 8860
rect 30098 8848 30104 8860
rect 30156 8848 30162 8900
rect 31938 8848 31944 8900
rect 31996 8888 32002 8900
rect 31996 8860 32352 8888
rect 31996 8848 32002 8860
rect 28902 8820 28908 8832
rect 27172 8792 28908 8820
rect 28902 8780 28908 8792
rect 28960 8780 28966 8832
rect 32214 8820 32220 8832
rect 32175 8792 32220 8820
rect 32214 8780 32220 8792
rect 32272 8780 32278 8832
rect 32324 8820 32352 8860
rect 32766 8848 32772 8900
rect 32824 8848 32830 8900
rect 41386 8888 41414 8928
rect 46753 8925 46765 8928
rect 46799 8925 46811 8959
rect 46753 8919 46811 8925
rect 47946 8888 47952 8900
rect 33336 8860 41414 8888
rect 47907 8860 47952 8888
rect 33336 8820 33364 8860
rect 47946 8848 47952 8860
rect 48004 8848 48010 8900
rect 32324 8792 33364 8820
rect 46474 8780 46480 8832
rect 46532 8820 46538 8832
rect 46845 8823 46903 8829
rect 46845 8820 46857 8823
rect 46532 8792 46857 8820
rect 46532 8780 46538 8792
rect 46845 8789 46857 8792
rect 46891 8789 46903 8823
rect 46845 8783 46903 8789
rect 1104 8730 48852 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 48852 8730
rect 1104 8656 48852 8678
rect 23569 8619 23627 8625
rect 18248 8588 19625 8616
rect 18248 8557 18276 8588
rect 18233 8551 18291 8557
rect 18233 8517 18245 8551
rect 18279 8517 18291 8551
rect 18233 8511 18291 8517
rect 18414 8508 18420 8560
rect 18472 8548 18478 8560
rect 19597 8557 19625 8588
rect 23569 8585 23581 8619
rect 23615 8616 23627 8619
rect 23750 8616 23756 8628
rect 23615 8588 23756 8616
rect 23615 8585 23627 8588
rect 23569 8579 23627 8585
rect 23750 8576 23756 8588
rect 23808 8616 23814 8628
rect 24762 8616 24768 8628
rect 23808 8588 24768 8616
rect 23808 8576 23814 8588
rect 24762 8576 24768 8588
rect 24820 8576 24826 8628
rect 27430 8576 27436 8628
rect 27488 8616 27494 8628
rect 28537 8619 28595 8625
rect 27488 8588 28396 8616
rect 27488 8576 27494 8588
rect 19582 8551 19640 8557
rect 18472 8520 18644 8548
rect 18472 8508 18478 8520
rect 18616 8492 18644 8520
rect 19582 8517 19594 8551
rect 19628 8517 19640 8551
rect 19582 8511 19640 8517
rect 23385 8551 23443 8557
rect 23385 8517 23397 8551
rect 23431 8548 23443 8551
rect 24210 8548 24216 8560
rect 23431 8520 24216 8548
rect 23431 8517 23443 8520
rect 23385 8511 23443 8517
rect 24210 8508 24216 8520
rect 24268 8548 24274 8560
rect 27154 8548 27160 8560
rect 24268 8520 27160 8548
rect 24268 8508 24274 8520
rect 27154 8508 27160 8520
rect 27212 8508 27218 8560
rect 28258 8508 28264 8560
rect 28316 8508 28322 8560
rect 28368 8548 28396 8588
rect 28537 8585 28549 8619
rect 28583 8616 28595 8619
rect 28626 8616 28632 8628
rect 28583 8588 28632 8616
rect 28583 8585 28595 8588
rect 28537 8579 28595 8585
rect 28626 8576 28632 8588
rect 28684 8576 28690 8628
rect 29549 8619 29607 8625
rect 29549 8616 29561 8619
rect 28736 8588 29561 8616
rect 28736 8548 28764 8588
rect 29549 8585 29561 8588
rect 29595 8585 29607 8619
rect 29549 8579 29607 8585
rect 28368 8520 28764 8548
rect 29089 8551 29147 8557
rect 29089 8517 29101 8551
rect 29135 8548 29147 8551
rect 30190 8548 30196 8560
rect 29135 8520 30196 8548
rect 29135 8517 29147 8520
rect 29089 8511 29147 8517
rect 30190 8508 30196 8520
rect 30248 8508 30254 8560
rect 32214 8508 32220 8560
rect 32272 8548 32278 8560
rect 32646 8551 32704 8557
rect 32646 8548 32658 8551
rect 32272 8520 32658 8548
rect 32272 8508 32278 8520
rect 32646 8517 32658 8520
rect 32692 8517 32704 8551
rect 32646 8511 32704 8517
rect 1854 8480 1860 8492
rect 1815 8452 1860 8480
rect 1854 8440 1860 8452
rect 1912 8440 1918 8492
rect 18509 8483 18567 8489
rect 18509 8449 18521 8483
rect 18555 8449 18567 8483
rect 18509 8443 18567 8449
rect 18598 8486 18656 8492
rect 18598 8452 18610 8486
rect 18644 8452 18656 8486
rect 18598 8446 18656 8452
rect 18693 8483 18751 8489
rect 18782 8483 18788 8492
rect 18693 8449 18705 8483
rect 18739 8455 18788 8483
rect 18739 8449 18751 8455
rect 18693 8443 18751 8449
rect 18322 8372 18328 8424
rect 18380 8412 18386 8424
rect 18524 8412 18552 8443
rect 18782 8440 18788 8455
rect 18840 8440 18846 8492
rect 18874 8440 18880 8492
rect 18932 8480 18938 8492
rect 19334 8480 19340 8492
rect 18932 8452 18977 8480
rect 19295 8452 19340 8480
rect 18932 8440 18938 8452
rect 19334 8440 19340 8452
rect 19392 8440 19398 8492
rect 23658 8440 23664 8492
rect 23716 8480 23722 8492
rect 24121 8483 24179 8489
rect 23716 8452 23761 8480
rect 23716 8440 23722 8452
rect 24121 8449 24133 8483
rect 24167 8449 24179 8483
rect 24121 8443 24179 8449
rect 24305 8483 24363 8489
rect 24305 8449 24317 8483
rect 24351 8480 24363 8483
rect 24394 8480 24400 8492
rect 24351 8452 24400 8480
rect 24351 8449 24363 8452
rect 24305 8443 24363 8449
rect 18380 8384 18552 8412
rect 18380 8372 18386 8384
rect 2133 8347 2191 8353
rect 2133 8313 2145 8347
rect 2179 8344 2191 8347
rect 17678 8344 17684 8356
rect 2179 8316 17684 8344
rect 2179 8313 2191 8316
rect 2133 8307 2191 8313
rect 17678 8304 17684 8316
rect 17736 8304 17742 8356
rect 18782 8304 18788 8356
rect 18840 8344 18846 8356
rect 20714 8344 20720 8356
rect 18840 8316 19380 8344
rect 20675 8316 20720 8344
rect 18840 8304 18846 8316
rect 19352 8276 19380 8316
rect 20714 8304 20720 8316
rect 20772 8304 20778 8356
rect 23385 8347 23443 8353
rect 23385 8313 23397 8347
rect 23431 8344 23443 8347
rect 24136 8344 24164 8443
rect 24394 8440 24400 8452
rect 24452 8440 24458 8492
rect 27433 8483 27491 8489
rect 27433 8449 27445 8483
rect 27479 8480 27491 8483
rect 27890 8480 27896 8492
rect 27479 8452 27896 8480
rect 27479 8449 27491 8452
rect 27433 8443 27491 8449
rect 27890 8440 27896 8452
rect 27948 8480 27954 8492
rect 28169 8483 28227 8489
rect 28169 8480 28181 8483
rect 27948 8452 28181 8480
rect 27948 8440 27954 8452
rect 28169 8449 28181 8452
rect 28215 8480 28227 8483
rect 28276 8480 28304 8508
rect 28215 8452 28304 8480
rect 29365 8483 29423 8489
rect 28215 8449 28227 8452
rect 28169 8443 28227 8449
rect 29365 8449 29377 8483
rect 29411 8449 29423 8483
rect 29365 8443 29423 8449
rect 26050 8372 26056 8424
rect 26108 8412 26114 8424
rect 27614 8412 27620 8424
rect 26108 8384 27620 8412
rect 26108 8372 26114 8384
rect 27614 8372 27620 8384
rect 27672 8412 27678 8424
rect 27709 8415 27767 8421
rect 27709 8412 27721 8415
rect 27672 8384 27721 8412
rect 27672 8372 27678 8384
rect 27709 8381 27721 8384
rect 27755 8412 27767 8415
rect 28261 8415 28319 8421
rect 28261 8412 28273 8415
rect 27755 8384 28273 8412
rect 27755 8381 27767 8384
rect 27709 8375 27767 8381
rect 28261 8381 28273 8384
rect 28307 8381 28319 8415
rect 28261 8375 28319 8381
rect 29273 8415 29331 8421
rect 29273 8381 29285 8415
rect 29319 8381 29331 8415
rect 29380 8412 29408 8443
rect 29546 8440 29552 8492
rect 29604 8480 29610 8492
rect 32401 8483 32459 8489
rect 32401 8480 32413 8483
rect 29604 8452 32413 8480
rect 29604 8440 29610 8452
rect 32401 8449 32413 8452
rect 32447 8449 32459 8483
rect 47854 8480 47860 8492
rect 47815 8452 47860 8480
rect 32401 8443 32459 8449
rect 47854 8440 47860 8452
rect 47912 8440 47918 8492
rect 29638 8412 29644 8424
rect 29380 8384 29644 8412
rect 29273 8375 29331 8381
rect 23431 8316 24164 8344
rect 27249 8347 27307 8353
rect 23431 8313 23443 8316
rect 23385 8307 23443 8313
rect 27249 8313 27261 8347
rect 27295 8344 27307 8347
rect 28074 8344 28080 8356
rect 27295 8316 28080 8344
rect 27295 8313 27307 8316
rect 27249 8307 27307 8313
rect 28074 8304 28080 8316
rect 28132 8304 28138 8356
rect 29288 8344 29316 8375
rect 29638 8372 29644 8384
rect 29696 8372 29702 8424
rect 29822 8344 29828 8356
rect 29288 8316 29828 8344
rect 29822 8304 29828 8316
rect 29880 8304 29886 8356
rect 35802 8304 35808 8356
rect 35860 8344 35866 8356
rect 48041 8347 48099 8353
rect 48041 8344 48053 8347
rect 35860 8316 48053 8344
rect 35860 8304 35866 8316
rect 48041 8313 48053 8316
rect 48087 8313 48099 8347
rect 48041 8307 48099 8313
rect 19610 8276 19616 8288
rect 19352 8248 19616 8276
rect 19610 8236 19616 8248
rect 19668 8236 19674 8288
rect 24213 8279 24271 8285
rect 24213 8245 24225 8279
rect 24259 8276 24271 8279
rect 24394 8276 24400 8288
rect 24259 8248 24400 8276
rect 24259 8245 24271 8248
rect 24213 8239 24271 8245
rect 24394 8236 24400 8248
rect 24452 8236 24458 8288
rect 27614 8276 27620 8288
rect 27575 8248 27620 8276
rect 27614 8236 27620 8248
rect 27672 8276 27678 8288
rect 27798 8276 27804 8288
rect 27672 8248 27804 8276
rect 27672 8236 27678 8248
rect 27798 8236 27804 8248
rect 27856 8276 27862 8288
rect 28169 8279 28227 8285
rect 28169 8276 28181 8279
rect 27856 8248 28181 8276
rect 27856 8236 27862 8248
rect 28169 8245 28181 8248
rect 28215 8245 28227 8279
rect 28169 8239 28227 8245
rect 28902 8236 28908 8288
rect 28960 8276 28966 8288
rect 29089 8279 29147 8285
rect 29089 8276 29101 8279
rect 28960 8248 29101 8276
rect 28960 8236 28966 8248
rect 29089 8245 29101 8248
rect 29135 8245 29147 8279
rect 33778 8276 33784 8288
rect 33739 8248 33784 8276
rect 29089 8239 29147 8245
rect 33778 8236 33784 8248
rect 33836 8236 33842 8288
rect 47026 8276 47032 8288
rect 46987 8248 47032 8276
rect 47026 8236 47032 8248
rect 47084 8236 47090 8288
rect 1104 8186 48852 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 48852 8186
rect 1104 8112 48852 8134
rect 18966 8072 18972 8084
rect 6886 8044 18972 8072
rect 2133 7939 2191 7945
rect 2133 7905 2145 7939
rect 2179 7936 2191 7939
rect 6886 7936 6914 8044
rect 18966 8032 18972 8044
rect 19024 8032 19030 8084
rect 19610 8072 19616 8084
rect 19571 8044 19616 8072
rect 19610 8032 19616 8044
rect 19668 8032 19674 8084
rect 20714 8032 20720 8084
rect 20772 8072 20778 8084
rect 20772 8044 25360 8072
rect 20772 8032 20778 8044
rect 24578 8004 24584 8016
rect 2179 7908 6914 7936
rect 17236 7976 18828 8004
rect 2179 7905 2191 7908
rect 2133 7899 2191 7905
rect 17236 7877 17264 7976
rect 17589 7939 17647 7945
rect 17589 7905 17601 7939
rect 17635 7936 17647 7939
rect 17635 7908 18657 7936
rect 17635 7905 17647 7908
rect 17589 7899 17647 7905
rect 17221 7871 17279 7877
rect 17221 7837 17233 7871
rect 17267 7837 17279 7871
rect 18046 7868 18052 7880
rect 17221 7831 17279 7837
rect 17420 7840 18052 7868
rect 1854 7800 1860 7812
rect 1815 7772 1860 7800
rect 1854 7760 1860 7772
rect 1912 7760 1918 7812
rect 17420 7809 17448 7840
rect 18046 7828 18052 7840
rect 18104 7828 18110 7880
rect 18325 7871 18383 7877
rect 18325 7837 18337 7871
rect 18371 7837 18383 7871
rect 18430 7865 18488 7871
rect 18430 7858 18442 7865
rect 18325 7831 18383 7837
rect 17405 7803 17463 7809
rect 17405 7769 17417 7803
rect 17451 7769 17463 7803
rect 17405 7763 17463 7769
rect 17678 7692 17684 7744
rect 17736 7732 17742 7744
rect 18049 7735 18107 7741
rect 18049 7732 18061 7735
rect 17736 7704 18061 7732
rect 17736 7692 17742 7704
rect 18049 7701 18061 7704
rect 18095 7701 18107 7735
rect 18340 7732 18368 7831
rect 18414 7806 18420 7858
rect 18476 7831 18488 7865
rect 18472 7825 18488 7831
rect 18530 7868 18588 7874
rect 18530 7834 18542 7868
rect 18576 7865 18588 7868
rect 18629 7865 18657 7908
rect 18576 7837 18657 7865
rect 18693 7871 18751 7877
rect 18693 7837 18705 7871
rect 18739 7837 18751 7871
rect 18800 7868 18828 7976
rect 23584 7976 24584 8004
rect 20346 7896 20352 7948
rect 20404 7936 20410 7948
rect 23584 7945 23612 7976
rect 24578 7964 24584 7976
rect 24636 8004 24642 8016
rect 24636 7976 24716 8004
rect 24636 7964 24642 7976
rect 20809 7939 20867 7945
rect 20809 7936 20821 7939
rect 20404 7908 20821 7936
rect 20404 7896 20410 7908
rect 20809 7905 20821 7908
rect 20855 7905 20867 7939
rect 20809 7899 20867 7905
rect 23569 7939 23627 7945
rect 23569 7905 23581 7939
rect 23615 7905 23627 7939
rect 23569 7899 23627 7905
rect 23753 7939 23811 7945
rect 23753 7905 23765 7939
rect 23799 7936 23811 7939
rect 24118 7936 24124 7948
rect 23799 7908 24124 7936
rect 23799 7905 23811 7908
rect 23753 7899 23811 7905
rect 24118 7896 24124 7908
rect 24176 7896 24182 7948
rect 24688 7945 24716 7976
rect 24673 7939 24731 7945
rect 24673 7905 24685 7939
rect 24719 7905 24731 7939
rect 25332 7936 25360 8044
rect 27522 8032 27528 8084
rect 27580 8072 27586 8084
rect 28077 8075 28135 8081
rect 28077 8072 28089 8075
rect 27580 8044 28089 8072
rect 27580 8032 27586 8044
rect 28077 8041 28089 8044
rect 28123 8041 28135 8075
rect 28077 8035 28135 8041
rect 33134 8032 33140 8084
rect 33192 8072 33198 8084
rect 33413 8075 33471 8081
rect 33413 8072 33425 8075
rect 33192 8044 33425 8072
rect 33192 8032 33198 8044
rect 33413 8041 33425 8044
rect 33459 8041 33471 8075
rect 33413 8035 33471 8041
rect 25685 7939 25743 7945
rect 25685 7936 25697 7939
rect 24673 7899 24731 7905
rect 24872 7908 25268 7936
rect 25332 7908 25697 7936
rect 19242 7868 19248 7880
rect 18800 7840 19248 7868
rect 18576 7834 18588 7837
rect 18530 7828 18588 7834
rect 18693 7831 18751 7837
rect 18472 7806 18478 7825
rect 18708 7800 18736 7831
rect 19242 7828 19248 7840
rect 19300 7828 19306 7880
rect 19429 7871 19487 7877
rect 19429 7837 19441 7871
rect 19475 7868 19487 7871
rect 20714 7868 20720 7880
rect 19475 7840 20720 7868
rect 19475 7837 19487 7840
rect 19429 7831 19487 7837
rect 20714 7828 20720 7840
rect 20772 7828 20778 7880
rect 24394 7868 24400 7880
rect 24355 7840 24400 7868
rect 24394 7828 24400 7840
rect 24452 7828 24458 7880
rect 24486 7828 24492 7880
rect 24544 7868 24550 7880
rect 24581 7871 24639 7877
rect 24581 7868 24593 7871
rect 24544 7840 24593 7868
rect 24544 7828 24550 7840
rect 24581 7837 24593 7840
rect 24627 7837 24639 7871
rect 24581 7831 24639 7837
rect 24765 7871 24823 7877
rect 24765 7837 24777 7871
rect 24811 7868 24823 7871
rect 24872 7868 24900 7908
rect 24811 7840 24900 7868
rect 24949 7871 25007 7877
rect 24811 7837 24823 7840
rect 24765 7831 24823 7837
rect 24949 7837 24961 7871
rect 24995 7837 25007 7871
rect 24949 7831 25007 7837
rect 18782 7800 18788 7812
rect 18708 7772 18788 7800
rect 18782 7760 18788 7772
rect 18840 7800 18846 7812
rect 19058 7800 19064 7812
rect 18840 7772 19064 7800
rect 18840 7760 18846 7772
rect 19058 7760 19064 7772
rect 19116 7760 19122 7812
rect 20990 7800 20996 7812
rect 20951 7772 20996 7800
rect 20990 7760 20996 7772
rect 21048 7760 21054 7812
rect 22649 7803 22707 7809
rect 22649 7769 22661 7803
rect 22695 7800 22707 7803
rect 22830 7800 22836 7812
rect 22695 7772 22836 7800
rect 22695 7769 22707 7772
rect 22649 7763 22707 7769
rect 22830 7760 22836 7772
rect 22888 7760 22894 7812
rect 23477 7803 23535 7809
rect 23477 7800 23489 7803
rect 23032 7772 23489 7800
rect 20254 7732 20260 7744
rect 18340 7704 20260 7732
rect 18049 7695 18107 7701
rect 20254 7692 20260 7704
rect 20312 7692 20318 7744
rect 21082 7692 21088 7744
rect 21140 7732 21146 7744
rect 21634 7732 21640 7744
rect 21140 7704 21640 7732
rect 21140 7692 21146 7704
rect 21634 7692 21640 7704
rect 21692 7732 21698 7744
rect 23032 7732 23060 7772
rect 23477 7769 23489 7772
rect 23523 7800 23535 7803
rect 24964 7800 24992 7831
rect 23523 7772 24992 7800
rect 23523 7769 23535 7772
rect 23477 7763 23535 7769
rect 21692 7704 23060 7732
rect 23109 7735 23167 7741
rect 21692 7692 21698 7704
rect 23109 7701 23121 7735
rect 23155 7732 23167 7735
rect 23658 7732 23664 7744
rect 23155 7704 23664 7732
rect 23155 7701 23167 7704
rect 23109 7695 23167 7701
rect 23658 7692 23664 7704
rect 23716 7692 23722 7744
rect 25130 7732 25136 7744
rect 25091 7704 25136 7732
rect 25130 7692 25136 7704
rect 25188 7692 25194 7744
rect 25240 7732 25268 7908
rect 25685 7905 25697 7908
rect 25731 7905 25743 7939
rect 25685 7899 25743 7905
rect 28074 7896 28080 7948
rect 28132 7936 28138 7948
rect 28261 7939 28319 7945
rect 28261 7936 28273 7939
rect 28132 7908 28273 7936
rect 28132 7896 28138 7908
rect 28261 7905 28273 7908
rect 28307 7905 28319 7939
rect 28261 7899 28319 7905
rect 29546 7896 29552 7948
rect 29604 7936 29610 7948
rect 31205 7939 31263 7945
rect 31205 7936 31217 7939
rect 29604 7908 31217 7936
rect 29604 7896 29610 7908
rect 31205 7905 31217 7908
rect 31251 7905 31263 7939
rect 31205 7899 31263 7905
rect 46293 7939 46351 7945
rect 46293 7905 46305 7939
rect 46339 7936 46351 7939
rect 47026 7936 47032 7948
rect 46339 7908 47032 7936
rect 46339 7905 46351 7908
rect 46293 7899 46351 7905
rect 47026 7896 47032 7908
rect 47084 7896 47090 7948
rect 27982 7868 27988 7880
rect 27943 7840 27988 7868
rect 27982 7828 27988 7840
rect 28040 7828 28046 7880
rect 33226 7868 33232 7880
rect 33139 7840 33232 7868
rect 33226 7828 33232 7840
rect 33284 7868 33290 7880
rect 33778 7868 33784 7880
rect 33284 7840 33784 7868
rect 33284 7828 33290 7840
rect 33778 7828 33784 7840
rect 33836 7828 33842 7880
rect 25314 7760 25320 7812
rect 25372 7800 25378 7812
rect 25869 7803 25927 7809
rect 25869 7800 25881 7803
rect 25372 7772 25881 7800
rect 25372 7760 25378 7772
rect 25869 7769 25881 7772
rect 25915 7769 25927 7803
rect 27522 7800 27528 7812
rect 27483 7772 27528 7800
rect 25869 7763 25927 7769
rect 27522 7760 27528 7772
rect 27580 7760 27586 7812
rect 30926 7760 30932 7812
rect 30984 7800 30990 7812
rect 31450 7803 31508 7809
rect 31450 7800 31462 7803
rect 30984 7772 31462 7800
rect 30984 7760 30990 7772
rect 31450 7769 31462 7772
rect 31496 7769 31508 7803
rect 31450 7763 31508 7769
rect 32214 7760 32220 7812
rect 32272 7800 32278 7812
rect 32950 7800 32956 7812
rect 32272 7772 32956 7800
rect 32272 7760 32278 7772
rect 32950 7760 32956 7772
rect 33008 7800 33014 7812
rect 33045 7803 33103 7809
rect 33045 7800 33057 7803
rect 33008 7772 33057 7800
rect 33008 7760 33014 7772
rect 33045 7769 33057 7772
rect 33091 7769 33103 7803
rect 46474 7800 46480 7812
rect 46435 7772 46480 7800
rect 33045 7763 33103 7769
rect 46474 7760 46480 7772
rect 46532 7760 46538 7812
rect 48130 7800 48136 7812
rect 48091 7772 48136 7800
rect 48130 7760 48136 7772
rect 48188 7760 48194 7812
rect 26142 7732 26148 7744
rect 25240 7704 26148 7732
rect 26142 7692 26148 7704
rect 26200 7732 26206 7744
rect 27798 7732 27804 7744
rect 26200 7704 27804 7732
rect 26200 7692 26206 7704
rect 27798 7692 27804 7704
rect 27856 7692 27862 7744
rect 28537 7735 28595 7741
rect 28537 7701 28549 7735
rect 28583 7732 28595 7735
rect 29362 7732 29368 7744
rect 28583 7704 29368 7732
rect 28583 7701 28595 7704
rect 28537 7695 28595 7701
rect 29362 7692 29368 7704
rect 29420 7692 29426 7744
rect 32582 7732 32588 7744
rect 32543 7704 32588 7732
rect 32582 7692 32588 7704
rect 32640 7692 32646 7744
rect 1104 7642 48852 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 48852 7642
rect 1104 7568 48852 7590
rect 18046 7488 18052 7540
rect 18104 7528 18110 7540
rect 18230 7528 18236 7540
rect 18104 7500 18236 7528
rect 18104 7488 18110 7500
rect 18230 7488 18236 7500
rect 18288 7528 18294 7540
rect 18509 7531 18567 7537
rect 18509 7528 18521 7531
rect 18288 7500 18521 7528
rect 18288 7488 18294 7500
rect 18509 7497 18521 7500
rect 18555 7497 18567 7531
rect 18509 7491 18567 7497
rect 19426 7488 19432 7540
rect 19484 7528 19490 7540
rect 20990 7528 20996 7540
rect 19484 7500 20392 7528
rect 20951 7500 20996 7528
rect 19484 7488 19490 7500
rect 19334 7460 19340 7472
rect 17144 7432 19340 7460
rect 17144 7401 17172 7432
rect 19334 7420 19340 7432
rect 19392 7420 19398 7472
rect 20254 7460 20260 7472
rect 20215 7432 20260 7460
rect 20254 7420 20260 7432
rect 20312 7420 20318 7472
rect 20364 7460 20392 7500
rect 20990 7488 20996 7500
rect 21048 7488 21054 7540
rect 24578 7488 24584 7540
rect 24636 7528 24642 7540
rect 24857 7531 24915 7537
rect 24857 7528 24869 7531
rect 24636 7500 24869 7528
rect 24636 7488 24642 7500
rect 24857 7497 24869 7500
rect 24903 7497 24915 7531
rect 28169 7531 28227 7537
rect 24857 7491 24915 7497
rect 25240 7500 26234 7528
rect 23744 7463 23802 7469
rect 20364 7432 20944 7460
rect 20916 7404 20944 7432
rect 23744 7429 23756 7463
rect 23790 7460 23802 7463
rect 25130 7460 25136 7472
rect 23790 7432 25136 7460
rect 23790 7429 23802 7432
rect 23744 7423 23802 7429
rect 25130 7420 25136 7432
rect 25188 7420 25194 7472
rect 17129 7395 17187 7401
rect 17129 7361 17141 7395
rect 17175 7361 17187 7395
rect 17129 7355 17187 7361
rect 17396 7395 17454 7401
rect 17396 7361 17408 7395
rect 17442 7392 17454 7395
rect 17678 7392 17684 7404
rect 17442 7364 17684 7392
rect 17442 7361 17454 7364
rect 17396 7355 17454 7361
rect 17678 7352 17684 7364
rect 17736 7352 17742 7404
rect 20073 7395 20131 7401
rect 20073 7361 20085 7395
rect 20119 7361 20131 7395
rect 20898 7392 20904 7404
rect 20859 7364 20904 7392
rect 20073 7355 20131 7361
rect 20088 7324 20116 7355
rect 20898 7352 20904 7364
rect 20956 7352 20962 7404
rect 23474 7392 23480 7404
rect 23435 7364 23480 7392
rect 23474 7352 23480 7364
rect 23532 7352 23538 7404
rect 25240 7392 25268 7500
rect 26206 7460 26234 7500
rect 28169 7497 28181 7531
rect 28215 7528 28227 7531
rect 28258 7528 28264 7540
rect 28215 7500 28264 7528
rect 28215 7497 28227 7500
rect 28169 7491 28227 7497
rect 28258 7488 28264 7500
rect 28316 7488 28322 7540
rect 30926 7528 30932 7540
rect 30887 7500 30932 7528
rect 30926 7488 30932 7500
rect 30984 7488 30990 7540
rect 31570 7528 31576 7540
rect 31220 7500 31576 7528
rect 31220 7460 31248 7500
rect 31570 7488 31576 7500
rect 31628 7528 31634 7540
rect 32766 7528 32772 7540
rect 31628 7500 32772 7528
rect 31628 7488 31634 7500
rect 32766 7488 32772 7500
rect 32824 7488 32830 7540
rect 32950 7528 32956 7540
rect 32876 7500 32956 7528
rect 32490 7460 32496 7472
rect 26206 7432 31248 7460
rect 31312 7432 32496 7460
rect 26050 7392 26056 7404
rect 23584 7364 25268 7392
rect 26011 7364 26056 7392
rect 22186 7324 22192 7336
rect 20088 7296 22192 7324
rect 22186 7284 22192 7296
rect 22244 7284 22250 7336
rect 23584 7324 23612 7364
rect 26050 7352 26056 7364
rect 26108 7352 26114 7404
rect 26234 7352 26240 7404
rect 26292 7392 26298 7404
rect 27341 7395 27399 7401
rect 27341 7392 27353 7395
rect 26292 7364 27353 7392
rect 26292 7352 26298 7364
rect 27341 7361 27353 7364
rect 27387 7361 27399 7395
rect 28534 7392 28540 7404
rect 28495 7364 28540 7392
rect 27341 7355 27399 7361
rect 28534 7352 28540 7364
rect 28592 7352 28598 7404
rect 28629 7395 28687 7401
rect 28629 7361 28641 7395
rect 28675 7392 28687 7395
rect 29362 7392 29368 7404
rect 28675 7364 29224 7392
rect 29323 7364 29368 7392
rect 28675 7361 28687 7364
rect 28629 7355 28687 7361
rect 26142 7324 26148 7336
rect 23492 7296 23612 7324
rect 26103 7296 26148 7324
rect 18782 7216 18788 7268
rect 18840 7256 18846 7268
rect 23492 7256 23520 7296
rect 26142 7284 26148 7296
rect 26200 7284 26206 7336
rect 27430 7324 27436 7336
rect 26252 7296 27292 7324
rect 27391 7296 27436 7324
rect 26252 7256 26280 7296
rect 18840 7228 23520 7256
rect 26068 7228 26280 7256
rect 26421 7259 26479 7265
rect 18840 7216 18846 7228
rect 2038 7188 2044 7200
rect 1999 7160 2044 7188
rect 2038 7148 2044 7160
rect 2096 7148 2102 7200
rect 20441 7191 20499 7197
rect 20441 7157 20453 7191
rect 20487 7188 20499 7191
rect 21082 7188 21088 7200
rect 20487 7160 21088 7188
rect 20487 7157 20499 7160
rect 20441 7151 20499 7157
rect 21082 7148 21088 7160
rect 21140 7148 21146 7200
rect 24118 7148 24124 7200
rect 24176 7188 24182 7200
rect 26068 7188 26096 7228
rect 26421 7225 26433 7259
rect 26467 7256 26479 7259
rect 27062 7256 27068 7268
rect 26467 7228 27068 7256
rect 26467 7225 26479 7228
rect 26421 7219 26479 7225
rect 27062 7216 27068 7228
rect 27120 7216 27126 7268
rect 27264 7256 27292 7296
rect 27430 7284 27436 7296
rect 27488 7284 27494 7336
rect 27525 7327 27583 7333
rect 27525 7293 27537 7327
rect 27571 7324 27583 7327
rect 28721 7327 28779 7333
rect 28721 7324 28733 7327
rect 27571 7296 28733 7324
rect 27571 7293 27583 7296
rect 27525 7287 27583 7293
rect 28721 7293 28733 7296
rect 28767 7293 28779 7327
rect 29196 7324 29224 7364
rect 29362 7352 29368 7364
rect 29420 7352 29426 7404
rect 29454 7352 29460 7404
rect 29512 7392 29518 7404
rect 31312 7401 31340 7432
rect 32490 7420 32496 7432
rect 32548 7420 32554 7472
rect 29549 7395 29607 7401
rect 29549 7392 29561 7395
rect 29512 7364 29561 7392
rect 29512 7352 29518 7364
rect 29549 7361 29561 7364
rect 29595 7361 29607 7395
rect 29549 7355 29607 7361
rect 29733 7395 29791 7401
rect 29733 7361 29745 7395
rect 29779 7361 29791 7395
rect 29917 7395 29975 7401
rect 29917 7392 29929 7395
rect 29733 7355 29791 7361
rect 29840 7364 29929 7392
rect 29638 7324 29644 7336
rect 29196 7296 29644 7324
rect 28721 7287 28779 7293
rect 27540 7256 27568 7287
rect 29638 7284 29644 7296
rect 29696 7284 29702 7336
rect 27264 7228 27568 7256
rect 27798 7216 27804 7268
rect 27856 7256 27862 7268
rect 29748 7256 29776 7355
rect 27856 7228 29776 7256
rect 27856 7216 27862 7228
rect 24176 7160 26096 7188
rect 24176 7148 24182 7160
rect 26142 7148 26148 7200
rect 26200 7188 26206 7200
rect 26973 7191 27031 7197
rect 26973 7188 26985 7191
rect 26200 7160 26985 7188
rect 26200 7148 26206 7160
rect 26973 7157 26985 7160
rect 27019 7188 27031 7191
rect 27614 7188 27620 7200
rect 27019 7160 27620 7188
rect 27019 7157 27031 7160
rect 26973 7151 27031 7157
rect 27614 7148 27620 7160
rect 27672 7148 27678 7200
rect 28534 7148 28540 7200
rect 28592 7188 28598 7200
rect 29840 7188 29868 7364
rect 29917 7361 29929 7364
rect 29963 7392 29975 7395
rect 31185 7395 31243 7401
rect 31185 7392 31197 7395
rect 29963 7364 31197 7392
rect 29963 7361 29975 7364
rect 29917 7355 29975 7361
rect 31185 7361 31197 7364
rect 31231 7361 31243 7395
rect 31185 7355 31243 7361
rect 31297 7395 31355 7401
rect 31297 7361 31309 7395
rect 31343 7361 31355 7395
rect 31297 7355 31355 7361
rect 31389 7395 31447 7401
rect 31389 7361 31401 7395
rect 31435 7361 31447 7395
rect 31389 7355 31447 7361
rect 31404 7324 31432 7355
rect 31570 7352 31576 7404
rect 31628 7392 31634 7404
rect 32125 7395 32183 7401
rect 31628 7364 31673 7392
rect 31628 7352 31634 7364
rect 32125 7361 32137 7395
rect 32171 7392 32183 7395
rect 32876 7392 32904 7500
rect 32950 7488 32956 7500
rect 33008 7488 33014 7540
rect 33045 7463 33103 7469
rect 33045 7429 33057 7463
rect 33091 7460 33103 7463
rect 33410 7460 33416 7472
rect 33091 7432 33416 7460
rect 33091 7429 33103 7432
rect 33045 7423 33103 7429
rect 33410 7420 33416 7432
rect 33468 7420 33474 7472
rect 32171 7364 32904 7392
rect 32171 7361 32183 7364
rect 32125 7355 32183 7361
rect 32490 7324 32496 7336
rect 31404 7296 32496 7324
rect 32490 7284 32496 7296
rect 32548 7284 32554 7336
rect 32861 7327 32919 7333
rect 32861 7293 32873 7327
rect 32907 7324 32919 7327
rect 33226 7324 33232 7336
rect 32907 7296 33232 7324
rect 32907 7293 32919 7296
rect 32861 7287 32919 7293
rect 33226 7284 33232 7296
rect 33284 7284 33290 7336
rect 33321 7327 33379 7333
rect 33321 7293 33333 7327
rect 33367 7293 33379 7327
rect 33321 7287 33379 7293
rect 29914 7216 29920 7268
rect 29972 7256 29978 7268
rect 33336 7256 33364 7287
rect 29972 7228 33364 7256
rect 29972 7216 29978 7228
rect 30098 7188 30104 7200
rect 28592 7160 29868 7188
rect 30059 7160 30104 7188
rect 28592 7148 28598 7160
rect 30098 7148 30104 7160
rect 30156 7148 30162 7200
rect 31846 7148 31852 7200
rect 31904 7188 31910 7200
rect 32217 7191 32275 7197
rect 32217 7188 32229 7191
rect 31904 7160 32229 7188
rect 31904 7148 31910 7160
rect 32217 7157 32229 7160
rect 32263 7157 32275 7191
rect 32217 7151 32275 7157
rect 1104 7098 48852 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 48852 7098
rect 1104 7024 48852 7046
rect 20898 6944 20904 6996
rect 20956 6984 20962 6996
rect 29270 6984 29276 6996
rect 20956 6956 29276 6984
rect 20956 6944 20962 6956
rect 29270 6944 29276 6956
rect 29328 6944 29334 6996
rect 24486 6876 24492 6928
rect 24544 6916 24550 6928
rect 29362 6916 29368 6928
rect 24544 6888 29368 6916
rect 24544 6876 24550 6888
rect 29362 6876 29368 6888
rect 29420 6876 29426 6928
rect 1397 6851 1455 6857
rect 1397 6817 1409 6851
rect 1443 6848 1455 6851
rect 2038 6848 2044 6860
rect 1443 6820 2044 6848
rect 1443 6817 1455 6820
rect 1397 6811 1455 6817
rect 2038 6808 2044 6820
rect 2096 6808 2102 6860
rect 2222 6808 2228 6860
rect 2280 6848 2286 6860
rect 2406 6848 2412 6860
rect 2280 6820 2412 6848
rect 2280 6808 2286 6820
rect 2406 6808 2412 6820
rect 2464 6808 2470 6860
rect 2774 6848 2780 6860
rect 2735 6820 2780 6848
rect 2774 6808 2780 6820
rect 2832 6808 2838 6860
rect 19334 6808 19340 6860
rect 19392 6848 19398 6860
rect 20254 6848 20260 6860
rect 19392 6820 20260 6848
rect 19392 6808 19398 6820
rect 20254 6808 20260 6820
rect 20312 6808 20318 6860
rect 26326 6808 26332 6860
rect 26384 6848 26390 6860
rect 27249 6851 27307 6857
rect 27249 6848 27261 6851
rect 26384 6820 27261 6848
rect 26384 6808 26390 6820
rect 27249 6817 27261 6820
rect 27295 6817 27307 6851
rect 28718 6848 28724 6860
rect 27249 6811 27307 6817
rect 27356 6820 28724 6848
rect 17954 6740 17960 6792
rect 18012 6780 18018 6792
rect 18325 6783 18383 6789
rect 18325 6780 18337 6783
rect 18012 6752 18337 6780
rect 18012 6740 18018 6752
rect 18325 6749 18337 6752
rect 18371 6749 18383 6783
rect 26234 6780 26240 6792
rect 18325 6743 18383 6749
rect 21652 6752 26240 6780
rect 1581 6715 1639 6721
rect 1581 6681 1593 6715
rect 1627 6712 1639 6715
rect 2222 6712 2228 6724
rect 1627 6684 2228 6712
rect 1627 6681 1639 6684
rect 1581 6675 1639 6681
rect 2222 6672 2228 6684
rect 2280 6672 2286 6724
rect 20524 6715 20582 6721
rect 20524 6681 20536 6715
rect 20570 6712 20582 6715
rect 20622 6712 20628 6724
rect 20570 6684 20628 6712
rect 20570 6681 20582 6684
rect 20524 6675 20582 6681
rect 20622 6672 20628 6684
rect 20680 6672 20686 6724
rect 18322 6604 18328 6656
rect 18380 6644 18386 6656
rect 18417 6647 18475 6653
rect 18417 6644 18429 6647
rect 18380 6616 18429 6644
rect 18380 6604 18386 6616
rect 18417 6613 18429 6616
rect 18463 6613 18475 6647
rect 18417 6607 18475 6613
rect 20346 6604 20352 6656
rect 20404 6644 20410 6656
rect 21652 6653 21680 6752
rect 26234 6740 26240 6752
rect 26292 6740 26298 6792
rect 26421 6783 26479 6789
rect 26421 6749 26433 6783
rect 26467 6780 26479 6783
rect 26881 6783 26939 6789
rect 26881 6780 26893 6783
rect 26467 6752 26893 6780
rect 26467 6749 26479 6752
rect 26421 6743 26479 6749
rect 26881 6749 26893 6752
rect 26927 6749 26939 6783
rect 27062 6780 27068 6792
rect 27023 6752 27068 6780
rect 26881 6743 26939 6749
rect 27062 6740 27068 6752
rect 27120 6740 27126 6792
rect 27154 6740 27160 6792
rect 27212 6780 27218 6792
rect 27212 6752 27257 6780
rect 27212 6740 27218 6752
rect 22186 6672 22192 6724
rect 22244 6712 22250 6724
rect 22649 6715 22707 6721
rect 22649 6712 22661 6715
rect 22244 6684 22661 6712
rect 22244 6672 22250 6684
rect 22649 6681 22661 6684
rect 22695 6681 22707 6715
rect 22649 6675 22707 6681
rect 22833 6715 22891 6721
rect 22833 6681 22845 6715
rect 22879 6712 22891 6715
rect 24762 6712 24768 6724
rect 22879 6684 24768 6712
rect 22879 6681 22891 6684
rect 22833 6675 22891 6681
rect 24762 6672 24768 6684
rect 24820 6672 24826 6724
rect 26053 6715 26111 6721
rect 26053 6681 26065 6715
rect 26099 6712 26111 6715
rect 27356 6712 27384 6820
rect 28718 6808 28724 6820
rect 28776 6808 28782 6860
rect 31846 6848 31852 6860
rect 31807 6820 31852 6848
rect 31846 6808 31852 6820
rect 31904 6808 31910 6860
rect 32122 6848 32128 6860
rect 32083 6820 32128 6848
rect 32122 6808 32128 6820
rect 32180 6808 32186 6860
rect 27430 6740 27436 6792
rect 27488 6780 27494 6792
rect 28902 6780 28908 6792
rect 27488 6752 28908 6780
rect 27488 6740 27494 6752
rect 28902 6740 28908 6752
rect 28960 6740 28966 6792
rect 29546 6780 29552 6792
rect 29507 6752 29552 6780
rect 29546 6740 29552 6752
rect 29604 6740 29610 6792
rect 29816 6783 29874 6789
rect 29816 6749 29828 6783
rect 29862 6780 29874 6783
rect 30098 6780 30104 6792
rect 29862 6752 30104 6780
rect 29862 6749 29874 6752
rect 29816 6743 29874 6749
rect 30098 6740 30104 6752
rect 30156 6740 30162 6792
rect 31665 6783 31723 6789
rect 31665 6749 31677 6783
rect 31711 6749 31723 6783
rect 31665 6743 31723 6749
rect 28534 6712 28540 6724
rect 26099 6684 27384 6712
rect 27540 6684 28540 6712
rect 26099 6681 26111 6684
rect 26053 6675 26111 6681
rect 21637 6647 21695 6653
rect 21637 6644 21649 6647
rect 20404 6616 21649 6644
rect 20404 6604 20410 6616
rect 21637 6613 21649 6616
rect 21683 6613 21695 6647
rect 21637 6607 21695 6613
rect 23017 6647 23075 6653
rect 23017 6613 23029 6647
rect 23063 6644 23075 6647
rect 23198 6644 23204 6656
rect 23063 6616 23204 6644
rect 23063 6613 23075 6616
rect 23017 6607 23075 6613
rect 23198 6604 23204 6616
rect 23256 6604 23262 6656
rect 24780 6644 24808 6672
rect 27540 6644 27568 6684
rect 28534 6672 28540 6684
rect 28592 6672 28598 6724
rect 31680 6712 31708 6743
rect 32582 6712 32588 6724
rect 31680 6684 32588 6712
rect 32582 6672 32588 6684
rect 32640 6672 32646 6724
rect 24780 6616 27568 6644
rect 27617 6647 27675 6653
rect 27617 6613 27629 6647
rect 27663 6644 27675 6647
rect 27706 6644 27712 6656
rect 27663 6616 27712 6644
rect 27663 6613 27675 6616
rect 27617 6607 27675 6613
rect 27706 6604 27712 6616
rect 27764 6604 27770 6656
rect 29638 6604 29644 6656
rect 29696 6644 29702 6656
rect 30929 6647 30987 6653
rect 30929 6644 30941 6647
rect 29696 6616 30941 6644
rect 29696 6604 29702 6616
rect 30929 6613 30941 6616
rect 30975 6613 30987 6647
rect 30929 6607 30987 6613
rect 1104 6554 48852 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 48852 6554
rect 1104 6480 48852 6502
rect 2222 6440 2228 6452
rect 2183 6412 2228 6440
rect 2222 6400 2228 6412
rect 2280 6400 2286 6452
rect 28813 6443 28871 6449
rect 20824 6412 22324 6440
rect 18322 6372 18328 6384
rect 18283 6344 18328 6372
rect 18322 6332 18328 6344
rect 18380 6332 18386 6384
rect 2130 6304 2136 6316
rect 2091 6276 2136 6304
rect 2130 6264 2136 6276
rect 2188 6264 2194 6316
rect 18138 6304 18144 6316
rect 18099 6276 18144 6304
rect 18138 6264 18144 6276
rect 18196 6264 18202 6316
rect 20824 6313 20852 6412
rect 22296 6384 22324 6412
rect 28813 6409 28825 6443
rect 28859 6440 28871 6443
rect 28902 6440 28908 6452
rect 28859 6412 28908 6440
rect 28859 6409 28871 6412
rect 28813 6403 28871 6409
rect 28902 6400 28908 6412
rect 28960 6400 28966 6452
rect 46842 6440 46848 6452
rect 31726 6412 46848 6440
rect 22189 6375 22247 6381
rect 22189 6372 22201 6375
rect 20916 6344 22201 6372
rect 20916 6313 20944 6344
rect 22189 6341 22201 6344
rect 22235 6341 22247 6375
rect 22189 6335 22247 6341
rect 22278 6332 22284 6384
rect 22336 6372 22342 6384
rect 22462 6372 22468 6384
rect 22336 6344 22468 6372
rect 22336 6332 22342 6344
rect 22462 6332 22468 6344
rect 22520 6372 22526 6384
rect 29546 6372 29552 6384
rect 22520 6344 23152 6372
rect 22520 6332 22526 6344
rect 20717 6307 20775 6313
rect 20717 6304 20729 6307
rect 19628 6276 20729 6304
rect 19521 6239 19579 6245
rect 19521 6236 19533 6239
rect 19444 6208 19533 6236
rect 19444 6180 19472 6208
rect 19521 6205 19533 6208
rect 19567 6205 19579 6239
rect 19521 6199 19579 6205
rect 19426 6128 19432 6180
rect 19484 6128 19490 6180
rect 15194 6060 15200 6112
rect 15252 6100 15258 6112
rect 19628 6100 19656 6276
rect 20717 6273 20729 6276
rect 20763 6273 20775 6307
rect 20717 6267 20775 6273
rect 20809 6307 20867 6313
rect 20809 6273 20821 6307
rect 20855 6273 20867 6307
rect 20809 6267 20867 6273
rect 20901 6307 20959 6313
rect 20901 6273 20913 6307
rect 20947 6273 20959 6307
rect 20901 6267 20959 6273
rect 21085 6307 21143 6313
rect 21085 6273 21097 6307
rect 21131 6304 21143 6307
rect 21266 6304 21272 6316
rect 21131 6276 21272 6304
rect 21131 6273 21143 6276
rect 21085 6267 21143 6273
rect 21266 6264 21272 6276
rect 21324 6264 21330 6316
rect 21818 6304 21824 6316
rect 21779 6276 21824 6304
rect 21818 6264 21824 6276
rect 21876 6264 21882 6316
rect 21910 6264 21916 6316
rect 21968 6304 21974 6316
rect 23124 6313 23152 6344
rect 27448 6344 29552 6372
rect 22005 6307 22063 6313
rect 22005 6304 22017 6307
rect 21968 6276 22017 6304
rect 21968 6264 21974 6276
rect 22005 6273 22017 6276
rect 22051 6273 22063 6307
rect 22005 6267 22063 6273
rect 23017 6307 23075 6313
rect 23017 6273 23029 6307
rect 23063 6273 23075 6307
rect 23017 6267 23075 6273
rect 23109 6307 23167 6313
rect 23109 6273 23121 6307
rect 23155 6273 23167 6307
rect 23109 6267 23167 6273
rect 21836 6236 21864 6264
rect 22186 6236 22192 6248
rect 21836 6208 22192 6236
rect 22186 6196 22192 6208
rect 22244 6196 22250 6248
rect 23032 6236 23060 6267
rect 23198 6264 23204 6316
rect 23256 6304 23262 6316
rect 23256 6276 23301 6304
rect 23256 6264 23262 6276
rect 23382 6264 23388 6316
rect 23440 6304 23446 6316
rect 27448 6313 27476 6344
rect 29546 6332 29552 6344
rect 29604 6332 29610 6384
rect 27706 6313 27712 6316
rect 27433 6307 27491 6313
rect 23440 6276 23485 6304
rect 23440 6264 23446 6276
rect 27433 6273 27445 6307
rect 27479 6273 27491 6307
rect 27700 6304 27712 6313
rect 27667 6276 27712 6304
rect 27433 6267 27491 6273
rect 27700 6267 27712 6276
rect 27706 6264 27712 6267
rect 27764 6264 27770 6316
rect 26142 6236 26148 6248
rect 23032 6208 26148 6236
rect 26142 6196 26148 6208
rect 26200 6196 26206 6248
rect 22830 6128 22836 6180
rect 22888 6168 22894 6180
rect 22888 6140 27476 6168
rect 22888 6128 22894 6140
rect 15252 6072 19656 6100
rect 20441 6103 20499 6109
rect 15252 6060 15258 6072
rect 20441 6069 20453 6103
rect 20487 6100 20499 6103
rect 20530 6100 20536 6112
rect 20487 6072 20536 6100
rect 20487 6069 20499 6072
rect 20441 6063 20499 6069
rect 20530 6060 20536 6072
rect 20588 6060 20594 6112
rect 22741 6103 22799 6109
rect 22741 6069 22753 6103
rect 22787 6100 22799 6103
rect 23658 6100 23664 6112
rect 22787 6072 23664 6100
rect 22787 6069 22799 6072
rect 22741 6063 22799 6069
rect 23658 6060 23664 6072
rect 23716 6060 23722 6112
rect 27448 6100 27476 6140
rect 31726 6100 31754 6412
rect 46842 6400 46848 6412
rect 46900 6400 46906 6452
rect 32125 6375 32183 6381
rect 32125 6341 32137 6375
rect 32171 6372 32183 6375
rect 32214 6372 32220 6384
rect 32171 6344 32220 6372
rect 32171 6341 32183 6344
rect 32125 6335 32183 6341
rect 32214 6332 32220 6344
rect 32272 6332 32278 6384
rect 32490 6372 32496 6384
rect 32451 6344 32496 6372
rect 32490 6332 32496 6344
rect 32548 6332 32554 6384
rect 32309 6307 32367 6313
rect 32309 6273 32321 6307
rect 32355 6304 32367 6307
rect 32582 6304 32588 6316
rect 32355 6276 32588 6304
rect 32355 6273 32367 6276
rect 32309 6267 32367 6273
rect 32582 6264 32588 6276
rect 32640 6264 32646 6316
rect 27448 6072 31754 6100
rect 1104 6010 48852 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 48852 6010
rect 1104 5936 48852 5958
rect 3418 5856 3424 5908
rect 3476 5896 3482 5908
rect 32122 5896 32128 5908
rect 3476 5868 32128 5896
rect 3476 5856 3482 5868
rect 32122 5856 32128 5868
rect 32180 5856 32186 5908
rect 21634 5828 21640 5840
rect 21595 5800 21640 5828
rect 21634 5788 21640 5800
rect 21692 5788 21698 5840
rect 20254 5760 20260 5772
rect 20215 5732 20260 5760
rect 20254 5720 20260 5732
rect 20312 5720 20318 5772
rect 2133 5695 2191 5701
rect 2133 5661 2145 5695
rect 2179 5692 2191 5695
rect 2314 5692 2320 5704
rect 2179 5664 2320 5692
rect 2179 5661 2191 5664
rect 2133 5655 2191 5661
rect 2314 5652 2320 5664
rect 2372 5652 2378 5704
rect 2958 5692 2964 5704
rect 2919 5664 2964 5692
rect 2958 5652 2964 5664
rect 3016 5652 3022 5704
rect 3789 5695 3847 5701
rect 3789 5661 3801 5695
rect 3835 5661 3847 5695
rect 3789 5655 3847 5661
rect 19245 5695 19303 5701
rect 19245 5661 19257 5695
rect 19291 5692 19303 5695
rect 20070 5692 20076 5704
rect 19291 5664 20076 5692
rect 19291 5661 19303 5664
rect 19245 5655 19303 5661
rect 3804 5624 3832 5655
rect 20070 5652 20076 5664
rect 20128 5652 20134 5704
rect 20530 5701 20536 5704
rect 20524 5692 20536 5701
rect 20491 5664 20536 5692
rect 20524 5655 20536 5664
rect 20530 5652 20536 5655
rect 20588 5652 20594 5704
rect 22465 5695 22523 5701
rect 22465 5661 22477 5695
rect 22511 5692 22523 5695
rect 23474 5692 23480 5704
rect 22511 5664 23480 5692
rect 22511 5661 22523 5664
rect 22465 5655 22523 5661
rect 23474 5652 23480 5664
rect 23532 5652 23538 5704
rect 47854 5692 47860 5704
rect 47815 5664 47860 5692
rect 47854 5652 47860 5664
rect 47912 5652 47918 5704
rect 4798 5624 4804 5636
rect 3804 5596 4804 5624
rect 4798 5584 4804 5596
rect 4856 5624 4862 5636
rect 4856 5596 22094 5624
rect 4856 5584 4862 5596
rect 1578 5516 1584 5568
rect 1636 5556 1642 5568
rect 2225 5559 2283 5565
rect 2225 5556 2237 5559
rect 1636 5528 2237 5556
rect 1636 5516 1642 5528
rect 2225 5525 2237 5528
rect 2271 5525 2283 5559
rect 3878 5556 3884 5568
rect 3839 5528 3884 5556
rect 2225 5519 2283 5525
rect 3878 5516 3884 5528
rect 3936 5516 3942 5568
rect 19334 5556 19340 5568
rect 19295 5528 19340 5556
rect 19334 5516 19340 5528
rect 19392 5516 19398 5568
rect 22066 5556 22094 5596
rect 22186 5584 22192 5636
rect 22244 5624 22250 5636
rect 22710 5627 22768 5633
rect 22710 5624 22722 5627
rect 22244 5596 22722 5624
rect 22244 5584 22250 5596
rect 22710 5593 22722 5596
rect 22756 5593 22768 5627
rect 32030 5624 32036 5636
rect 22710 5587 22768 5593
rect 22848 5596 32036 5624
rect 22848 5556 22876 5596
rect 32030 5584 32036 5596
rect 32088 5624 32094 5636
rect 33042 5624 33048 5636
rect 32088 5596 33048 5624
rect 32088 5584 32094 5596
rect 33042 5584 33048 5596
rect 33100 5584 33106 5636
rect 23842 5556 23848 5568
rect 22066 5528 22876 5556
rect 23803 5528 23848 5556
rect 23842 5516 23848 5528
rect 23900 5516 23906 5568
rect 28626 5516 28632 5568
rect 28684 5556 28690 5568
rect 48041 5559 48099 5565
rect 48041 5556 48053 5559
rect 28684 5528 48053 5556
rect 28684 5516 28690 5528
rect 48041 5525 48053 5528
rect 48087 5525 48099 5559
rect 48041 5519 48099 5525
rect 1104 5466 48852 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 48852 5466
rect 1104 5392 48852 5414
rect 2958 5352 2964 5364
rect 2148 5324 2964 5352
rect 2148 5225 2176 5324
rect 2958 5312 2964 5324
rect 3016 5312 3022 5364
rect 3418 5312 3424 5364
rect 3476 5352 3482 5364
rect 10962 5352 10968 5364
rect 3476 5324 10968 5352
rect 3476 5312 3482 5324
rect 10962 5312 10968 5324
rect 11020 5312 11026 5364
rect 20622 5352 20628 5364
rect 20583 5324 20628 5352
rect 20622 5312 20628 5324
rect 20680 5312 20686 5364
rect 22097 5355 22155 5361
rect 22097 5321 22109 5355
rect 22143 5352 22155 5355
rect 22186 5352 22192 5364
rect 22143 5324 22192 5352
rect 22143 5321 22155 5324
rect 22097 5315 22155 5321
rect 22186 5312 22192 5324
rect 22244 5312 22250 5364
rect 24762 5352 24768 5364
rect 24723 5324 24768 5352
rect 24762 5312 24768 5324
rect 24820 5312 24826 5364
rect 38562 5312 38568 5364
rect 38620 5352 38626 5364
rect 46842 5352 46848 5364
rect 38620 5324 46848 5352
rect 38620 5312 38626 5324
rect 46842 5312 46848 5324
rect 46900 5312 46906 5364
rect 2317 5287 2375 5293
rect 2317 5253 2329 5287
rect 2363 5284 2375 5287
rect 3878 5284 3884 5296
rect 2363 5256 3884 5284
rect 2363 5253 2375 5256
rect 2317 5247 2375 5253
rect 3878 5244 3884 5256
rect 3936 5244 3942 5296
rect 18509 5287 18567 5293
rect 18509 5253 18521 5287
rect 18555 5284 18567 5287
rect 19334 5284 19340 5296
rect 18555 5256 19340 5284
rect 18555 5253 18567 5256
rect 18509 5247 18567 5253
rect 19334 5244 19340 5256
rect 19392 5244 19398 5296
rect 20165 5287 20223 5293
rect 20165 5253 20177 5287
rect 20211 5284 20223 5287
rect 46750 5284 46756 5296
rect 20211 5256 46756 5284
rect 20211 5253 20223 5256
rect 20165 5247 20223 5253
rect 46750 5244 46756 5256
rect 46808 5244 46814 5296
rect 2133 5219 2191 5225
rect 2133 5185 2145 5219
rect 2179 5185 2191 5219
rect 2133 5179 2191 5185
rect 20901 5219 20959 5225
rect 20901 5185 20913 5219
rect 20947 5185 20959 5219
rect 20901 5179 20959 5185
rect 20993 5219 21051 5225
rect 20993 5185 21005 5219
rect 21039 5185 21051 5219
rect 20993 5179 21051 5185
rect 2774 5148 2780 5160
rect 2735 5120 2780 5148
rect 2774 5108 2780 5120
rect 2832 5108 2838 5160
rect 18325 5151 18383 5157
rect 18325 5117 18337 5151
rect 18371 5148 18383 5151
rect 18690 5148 18696 5160
rect 18371 5120 18696 5148
rect 18371 5117 18383 5120
rect 18325 5111 18383 5117
rect 18690 5108 18696 5120
rect 18748 5108 18754 5160
rect 18782 5108 18788 5160
rect 18840 5148 18846 5160
rect 20916 5148 20944 5179
rect 18840 5120 20944 5148
rect 18840 5108 18846 5120
rect 21008 5080 21036 5179
rect 21082 5176 21088 5228
rect 21140 5216 21146 5228
rect 21140 5188 21185 5216
rect 21140 5176 21146 5188
rect 21266 5176 21272 5228
rect 21324 5216 21330 5228
rect 21324 5188 21369 5216
rect 21324 5176 21330 5188
rect 22278 5176 22284 5228
rect 22336 5225 22342 5228
rect 22336 5219 22385 5225
rect 22336 5185 22339 5219
rect 22373 5185 22385 5219
rect 22462 5216 22468 5228
rect 22423 5188 22468 5216
rect 22336 5179 22385 5185
rect 22336 5176 22342 5179
rect 22462 5176 22468 5188
rect 22520 5176 22526 5228
rect 22554 5176 22560 5228
rect 22612 5216 22618 5228
rect 22741 5219 22799 5225
rect 22612 5188 22657 5216
rect 22612 5176 22618 5188
rect 22741 5185 22753 5219
rect 22787 5185 22799 5219
rect 22741 5179 22799 5185
rect 23385 5219 23443 5225
rect 23385 5185 23397 5219
rect 23431 5216 23443 5219
rect 23474 5216 23480 5228
rect 23431 5188 23480 5216
rect 23431 5185 23443 5188
rect 23385 5179 23443 5185
rect 22462 5080 22468 5092
rect 21008 5052 22468 5080
rect 22462 5040 22468 5052
rect 22520 5040 22526 5092
rect 1394 4972 1400 5024
rect 1452 5012 1458 5024
rect 1673 5015 1731 5021
rect 1673 5012 1685 5015
rect 1452 4984 1685 5012
rect 1452 4972 1458 4984
rect 1673 4981 1685 4984
rect 1719 4981 1731 5015
rect 1673 4975 1731 4981
rect 21266 4972 21272 5024
rect 21324 5012 21330 5024
rect 22756 5012 22784 5179
rect 23474 5176 23480 5188
rect 23532 5176 23538 5228
rect 23658 5225 23664 5228
rect 23652 5216 23664 5225
rect 23619 5188 23664 5216
rect 23652 5179 23664 5188
rect 23658 5176 23664 5179
rect 23716 5176 23722 5228
rect 45646 5176 45652 5228
rect 45704 5216 45710 5228
rect 47581 5219 47639 5225
rect 47581 5216 47593 5219
rect 45704 5188 47593 5216
rect 45704 5176 45710 5188
rect 47581 5185 47593 5188
rect 47627 5185 47639 5219
rect 47581 5179 47639 5185
rect 21324 4984 22784 5012
rect 21324 4972 21330 4984
rect 46290 4972 46296 5024
rect 46348 5012 46354 5024
rect 47029 5015 47087 5021
rect 47029 5012 47041 5015
rect 46348 4984 47041 5012
rect 46348 4972 46354 4984
rect 47029 4981 47041 4984
rect 47075 4981 47087 5015
rect 47670 5012 47676 5024
rect 47631 4984 47676 5012
rect 47029 4975 47087 4981
rect 47670 4972 47676 4984
rect 47728 4972 47734 5024
rect 1104 4922 48852 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 48852 4922
rect 1104 4848 48852 4870
rect 22281 4811 22339 4817
rect 22281 4777 22293 4811
rect 22327 4808 22339 4811
rect 22554 4808 22560 4820
rect 22327 4780 22560 4808
rect 22327 4777 22339 4780
rect 22281 4771 22339 4777
rect 22554 4768 22560 4780
rect 22612 4768 22618 4820
rect 2498 4700 2504 4752
rect 2556 4740 2562 4752
rect 2556 4712 12388 4740
rect 2556 4700 2562 4712
rect 1394 4672 1400 4684
rect 1355 4644 1400 4672
rect 1394 4632 1400 4644
rect 1452 4632 1458 4684
rect 1578 4672 1584 4684
rect 1539 4644 1584 4672
rect 1578 4632 1584 4644
rect 1636 4632 1642 4684
rect 2774 4672 2780 4684
rect 2735 4644 2780 4672
rect 2774 4632 2780 4644
rect 2832 4632 2838 4684
rect 4614 4604 4620 4616
rect 4575 4576 4620 4604
rect 4614 4564 4620 4576
rect 4672 4564 4678 4616
rect 12360 4613 12388 4712
rect 20162 4700 20168 4752
rect 20220 4740 20226 4752
rect 32214 4740 32220 4752
rect 20220 4712 32220 4740
rect 20220 4700 20226 4712
rect 32214 4700 32220 4712
rect 32272 4700 32278 4752
rect 27890 4632 27896 4684
rect 27948 4672 27954 4684
rect 46290 4672 46296 4684
rect 27948 4644 31754 4672
rect 46251 4644 46296 4672
rect 27948 4632 27954 4644
rect 11701 4607 11759 4613
rect 11701 4573 11713 4607
rect 11747 4573 11759 4607
rect 11701 4567 11759 4573
rect 12345 4607 12403 4613
rect 12345 4573 12357 4607
rect 12391 4573 12403 4607
rect 12345 4567 12403 4573
rect 18509 4607 18567 4613
rect 18509 4573 18521 4607
rect 18555 4604 18567 4607
rect 20070 4604 20076 4616
rect 18555 4576 20076 4604
rect 18555 4573 18567 4576
rect 18509 4567 18567 4573
rect 11716 4536 11744 4567
rect 20070 4564 20076 4576
rect 20128 4564 20134 4616
rect 21818 4564 21824 4616
rect 21876 4604 21882 4616
rect 21913 4607 21971 4613
rect 21913 4604 21925 4607
rect 21876 4576 21925 4604
rect 21876 4564 21882 4576
rect 21913 4573 21925 4576
rect 21959 4573 21971 4607
rect 21913 4567 21971 4573
rect 22097 4607 22155 4613
rect 22097 4573 22109 4607
rect 22143 4604 22155 4607
rect 23842 4604 23848 4616
rect 22143 4576 23848 4604
rect 22143 4573 22155 4576
rect 22097 4567 22155 4573
rect 23842 4564 23848 4576
rect 23900 4564 23906 4616
rect 31202 4564 31208 4616
rect 31260 4604 31266 4616
rect 31481 4607 31539 4613
rect 31481 4604 31493 4607
rect 31260 4576 31493 4604
rect 31260 4564 31266 4576
rect 31481 4573 31493 4576
rect 31527 4573 31539 4607
rect 31726 4604 31754 4644
rect 46290 4632 46296 4644
rect 46348 4632 46354 4684
rect 46477 4675 46535 4681
rect 46477 4641 46489 4675
rect 46523 4672 46535 4675
rect 47670 4672 47676 4684
rect 46523 4644 47676 4672
rect 46523 4641 46535 4644
rect 46477 4635 46535 4641
rect 47670 4632 47676 4644
rect 47728 4632 47734 4684
rect 48130 4672 48136 4684
rect 48091 4644 48136 4672
rect 48130 4632 48136 4644
rect 48188 4632 48194 4684
rect 39853 4607 39911 4613
rect 39853 4604 39865 4607
rect 31726 4576 39865 4604
rect 31481 4567 31539 4573
rect 39853 4573 39865 4576
rect 39899 4573 39911 4607
rect 39853 4567 39911 4573
rect 14090 4536 14096 4548
rect 11716 4508 14096 4536
rect 14090 4496 14096 4508
rect 14148 4496 14154 4548
rect 11698 4428 11704 4480
rect 11756 4468 11762 4480
rect 11793 4471 11851 4477
rect 11793 4468 11805 4471
rect 11756 4440 11805 4468
rect 11756 4428 11762 4440
rect 11793 4437 11805 4440
rect 11839 4437 11851 4471
rect 11793 4431 11851 4437
rect 12434 4428 12440 4480
rect 12492 4468 12498 4480
rect 12492 4440 12537 4468
rect 12492 4428 12498 4440
rect 18138 4428 18144 4480
rect 18196 4468 18202 4480
rect 18601 4471 18659 4477
rect 18601 4468 18613 4471
rect 18196 4440 18613 4468
rect 18196 4428 18202 4440
rect 18601 4437 18613 4440
rect 18647 4437 18659 4471
rect 18601 4431 18659 4437
rect 39945 4471 40003 4477
rect 39945 4437 39957 4471
rect 39991 4468 40003 4471
rect 40218 4468 40224 4480
rect 39991 4440 40224 4468
rect 39991 4437 40003 4440
rect 39945 4431 40003 4437
rect 40218 4428 40224 4440
rect 40276 4428 40282 4480
rect 40494 4468 40500 4480
rect 40455 4440 40500 4468
rect 40494 4428 40500 4440
rect 40552 4428 40558 4480
rect 1104 4378 48852 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 48852 4378
rect 1104 4304 48852 4326
rect 19334 4224 19340 4276
rect 19392 4264 19398 4276
rect 37274 4264 37280 4276
rect 19392 4236 21036 4264
rect 19392 4224 19398 4236
rect 11698 4196 11704 4208
rect 11659 4168 11704 4196
rect 11698 4156 11704 4168
rect 11756 4156 11762 4208
rect 18616 4168 20116 4196
rect 4157 4131 4215 4137
rect 4157 4097 4169 4131
rect 4203 4097 4215 4131
rect 4798 4128 4804 4140
rect 4759 4100 4804 4128
rect 4157 4091 4215 4097
rect 4172 4060 4200 4091
rect 4798 4088 4804 4100
rect 4856 4088 4862 4140
rect 11517 4131 11575 4137
rect 11517 4128 11529 4131
rect 10520 4100 11529 4128
rect 8110 4060 8116 4072
rect 4172 4032 8116 4060
rect 8110 4020 8116 4032
rect 8168 4020 8174 4072
rect 9125 4063 9183 4069
rect 9125 4029 9137 4063
rect 9171 4029 9183 4063
rect 9306 4060 9312 4072
rect 9267 4032 9312 4060
rect 9125 4023 9183 4029
rect 2590 3952 2596 4004
rect 2648 3992 2654 4004
rect 8018 3992 8024 4004
rect 2648 3964 8024 3992
rect 2648 3952 2654 3964
rect 8018 3952 8024 3964
rect 8076 3952 8082 4004
rect 9140 3992 9168 4023
rect 9306 4020 9312 4032
rect 9364 4020 9370 4072
rect 9398 4020 9404 4072
rect 9456 4060 9462 4072
rect 9585 4063 9643 4069
rect 9585 4060 9597 4063
rect 9456 4032 9597 4060
rect 9456 4020 9462 4032
rect 9585 4029 9597 4032
rect 9631 4029 9643 4063
rect 9585 4023 9643 4029
rect 10134 4020 10140 4072
rect 10192 4060 10198 4072
rect 10520 4060 10548 4100
rect 11517 4097 11529 4100
rect 11563 4097 11575 4131
rect 11517 4091 11575 4097
rect 13817 4131 13875 4137
rect 13817 4097 13829 4131
rect 13863 4097 13875 4131
rect 13817 4091 13875 4097
rect 15197 4131 15255 4137
rect 15197 4097 15209 4131
rect 15243 4128 15255 4131
rect 18616 4128 18644 4168
rect 15243 4100 18644 4128
rect 15243 4097 15255 4100
rect 15197 4091 15255 4097
rect 12526 4060 12532 4072
rect 10192 4032 10548 4060
rect 12487 4032 12532 4060
rect 10192 4020 10198 4032
rect 12526 4020 12532 4032
rect 12584 4020 12590 4072
rect 13832 4060 13860 4091
rect 18690 4088 18696 4140
rect 18748 4128 18754 4140
rect 19426 4128 19432 4140
rect 18748 4100 19432 4128
rect 18748 4088 18754 4100
rect 19426 4088 19432 4100
rect 19484 4088 19490 4140
rect 19981 4131 20039 4137
rect 19981 4097 19993 4131
rect 20027 4097 20039 4131
rect 20088 4128 20116 4168
rect 20898 4128 20904 4140
rect 20088 4100 20904 4128
rect 19981 4091 20039 4097
rect 19334 4060 19340 4072
rect 13832 4032 19340 4060
rect 19334 4020 19340 4032
rect 19392 4020 19398 4072
rect 19996 4060 20024 4091
rect 20898 4088 20904 4100
rect 20956 4088 20962 4140
rect 20806 4060 20812 4072
rect 19996 4032 20812 4060
rect 20806 4020 20812 4032
rect 20864 4020 20870 4072
rect 21008 4060 21036 4236
rect 29104 4236 37280 4264
rect 23293 4131 23351 4137
rect 23293 4097 23305 4131
rect 23339 4128 23351 4131
rect 23934 4128 23940 4140
rect 23339 4100 23940 4128
rect 23339 4097 23351 4100
rect 23293 4091 23351 4097
rect 23934 4088 23940 4100
rect 23992 4088 23998 4140
rect 26053 4131 26111 4137
rect 26053 4097 26065 4131
rect 26099 4128 26111 4131
rect 28902 4128 28908 4140
rect 26099 4100 28908 4128
rect 26099 4097 26111 4100
rect 26053 4091 26111 4097
rect 28902 4088 28908 4100
rect 28960 4088 28966 4140
rect 29104 4060 29132 4236
rect 37274 4224 37280 4236
rect 37332 4264 37338 4276
rect 37734 4264 37740 4276
rect 37332 4236 37740 4264
rect 37332 4224 37338 4236
rect 37734 4224 37740 4236
rect 37792 4224 37798 4276
rect 29454 4156 29460 4208
rect 29512 4196 29518 4208
rect 29512 4168 32168 4196
rect 29512 4156 29518 4168
rect 29178 4088 29184 4140
rect 29236 4128 29242 4140
rect 29822 4128 29828 4140
rect 29236 4100 29828 4128
rect 29236 4088 29242 4100
rect 29822 4088 29828 4100
rect 29880 4088 29886 4140
rect 30926 4128 30932 4140
rect 30839 4100 30932 4128
rect 30926 4088 30932 4100
rect 30984 4128 30990 4140
rect 31754 4128 31760 4140
rect 30984 4100 31760 4128
rect 30984 4088 30990 4100
rect 31754 4088 31760 4100
rect 31812 4088 31818 4140
rect 32140 4137 32168 4168
rect 41248 4168 41460 4196
rect 32125 4131 32183 4137
rect 32125 4097 32137 4131
rect 32171 4097 32183 4131
rect 36170 4128 36176 4140
rect 36131 4100 36176 4128
rect 32125 4091 32183 4097
rect 36170 4088 36176 4100
rect 36228 4088 36234 4140
rect 37826 4128 37832 4140
rect 37787 4100 37832 4128
rect 37826 4088 37832 4100
rect 37884 4088 37890 4140
rect 37921 4131 37979 4137
rect 37921 4097 37933 4131
rect 37967 4128 37979 4131
rect 40497 4131 40555 4137
rect 37967 4100 38424 4128
rect 37967 4097 37979 4100
rect 37921 4091 37979 4097
rect 21008 4032 29132 4060
rect 35342 4020 35348 4072
rect 35400 4060 35406 4072
rect 35400 4032 38148 4060
rect 35400 4020 35406 4032
rect 10686 3992 10692 4004
rect 9140 3964 10692 3992
rect 10686 3952 10692 3964
rect 10744 3952 10750 4004
rect 10778 3952 10784 4004
rect 10836 3992 10842 4004
rect 10836 3964 18368 3992
rect 10836 3952 10842 3964
rect 1394 3884 1400 3936
rect 1452 3924 1458 3936
rect 2041 3927 2099 3933
rect 2041 3924 2053 3927
rect 1452 3896 2053 3924
rect 1452 3884 1458 3896
rect 2041 3893 2053 3896
rect 2087 3893 2099 3927
rect 2041 3887 2099 3893
rect 3605 3927 3663 3933
rect 3605 3893 3617 3927
rect 3651 3924 3663 3927
rect 3786 3924 3792 3936
rect 3651 3896 3792 3924
rect 3651 3893 3663 3896
rect 3605 3887 3663 3893
rect 3786 3884 3792 3896
rect 3844 3884 3850 3936
rect 3970 3884 3976 3936
rect 4028 3924 4034 3936
rect 4249 3927 4307 3933
rect 4249 3924 4261 3927
rect 4028 3896 4261 3924
rect 4028 3884 4034 3896
rect 4249 3893 4261 3896
rect 4295 3893 4307 3927
rect 4890 3924 4896 3936
rect 4851 3896 4896 3924
rect 4249 3887 4307 3893
rect 4890 3884 4896 3896
rect 4948 3884 4954 3936
rect 6454 3884 6460 3936
rect 6512 3924 6518 3936
rect 6641 3927 6699 3933
rect 6641 3924 6653 3927
rect 6512 3896 6653 3924
rect 6512 3884 6518 3896
rect 6641 3893 6653 3896
rect 6687 3893 6699 3927
rect 6641 3887 6699 3893
rect 10318 3884 10324 3936
rect 10376 3924 10382 3936
rect 13262 3924 13268 3936
rect 10376 3896 13268 3924
rect 10376 3884 10382 3896
rect 13262 3884 13268 3896
rect 13320 3884 13326 3936
rect 13909 3927 13967 3933
rect 13909 3893 13921 3927
rect 13955 3924 13967 3927
rect 14274 3924 14280 3936
rect 13955 3896 14280 3924
rect 13955 3893 13967 3896
rect 13909 3887 13967 3893
rect 14274 3884 14280 3896
rect 14332 3884 14338 3936
rect 15102 3884 15108 3936
rect 15160 3924 15166 3936
rect 15289 3927 15347 3933
rect 15289 3924 15301 3927
rect 15160 3896 15301 3924
rect 15160 3884 15166 3896
rect 15289 3893 15301 3896
rect 15335 3893 15347 3927
rect 15289 3887 15347 3893
rect 17954 3884 17960 3936
rect 18012 3924 18018 3936
rect 18233 3927 18291 3933
rect 18233 3924 18245 3927
rect 18012 3896 18245 3924
rect 18012 3884 18018 3896
rect 18233 3893 18245 3896
rect 18279 3893 18291 3927
rect 18340 3924 18368 3964
rect 22554 3952 22560 4004
rect 22612 3992 22618 4004
rect 30926 3992 30932 4004
rect 22612 3964 30932 3992
rect 22612 3952 22618 3964
rect 30926 3952 30932 3964
rect 30984 3952 30990 4004
rect 31110 3952 31116 4004
rect 31168 3992 31174 4004
rect 31168 3964 36584 3992
rect 31168 3952 31174 3964
rect 19978 3924 19984 3936
rect 18340 3896 19984 3924
rect 18233 3887 18291 3893
rect 19978 3884 19984 3896
rect 20036 3884 20042 3936
rect 20073 3927 20131 3933
rect 20073 3893 20085 3927
rect 20119 3924 20131 3927
rect 20254 3924 20260 3936
rect 20119 3896 20260 3924
rect 20119 3893 20131 3896
rect 20073 3887 20131 3893
rect 20254 3884 20260 3896
rect 20312 3884 20318 3936
rect 20898 3924 20904 3936
rect 20859 3896 20904 3924
rect 20898 3884 20904 3896
rect 20956 3884 20962 3936
rect 23385 3927 23443 3933
rect 23385 3893 23397 3927
rect 23431 3924 23443 3927
rect 23566 3924 23572 3936
rect 23431 3896 23572 3924
rect 23431 3893 23443 3896
rect 23385 3887 23443 3893
rect 23566 3884 23572 3896
rect 23624 3884 23630 3936
rect 25958 3884 25964 3936
rect 26016 3924 26022 3936
rect 26145 3927 26203 3933
rect 26145 3924 26157 3927
rect 26016 3896 26157 3924
rect 26016 3884 26022 3896
rect 26145 3893 26157 3896
rect 26191 3893 26203 3927
rect 26145 3887 26203 3893
rect 29730 3884 29736 3936
rect 29788 3924 29794 3936
rect 30009 3927 30067 3933
rect 30009 3924 30021 3927
rect 29788 3896 30021 3924
rect 29788 3884 29794 3896
rect 30009 3893 30021 3896
rect 30055 3893 30067 3927
rect 30009 3887 30067 3893
rect 31021 3927 31079 3933
rect 31021 3893 31033 3927
rect 31067 3924 31079 3927
rect 31386 3924 31392 3936
rect 31067 3896 31392 3924
rect 31067 3893 31079 3896
rect 31021 3887 31079 3893
rect 31386 3884 31392 3896
rect 31444 3884 31450 3936
rect 32217 3927 32275 3933
rect 32217 3893 32229 3927
rect 32263 3924 32275 3927
rect 32398 3924 32404 3936
rect 32263 3896 32404 3924
rect 32263 3893 32275 3896
rect 32217 3887 32275 3893
rect 32398 3884 32404 3896
rect 32456 3884 32462 3936
rect 32950 3924 32956 3936
rect 32911 3896 32956 3924
rect 32950 3884 32956 3896
rect 33008 3884 33014 3936
rect 36265 3927 36323 3933
rect 36265 3893 36277 3927
rect 36311 3924 36323 3927
rect 36446 3924 36452 3936
rect 36311 3896 36452 3924
rect 36311 3893 36323 3896
rect 36265 3887 36323 3893
rect 36446 3884 36452 3896
rect 36504 3884 36510 3936
rect 36556 3924 36584 3964
rect 38010 3924 38016 3936
rect 36556 3896 38016 3924
rect 38010 3884 38016 3896
rect 38068 3884 38074 3936
rect 38120 3924 38148 4032
rect 38396 3992 38424 4100
rect 40497 4097 40509 4131
rect 40543 4128 40555 4131
rect 41248 4128 41276 4168
rect 40543 4100 41276 4128
rect 41325 4131 41383 4137
rect 40543 4097 40555 4100
rect 40497 4091 40555 4097
rect 41325 4097 41337 4131
rect 41371 4097 41383 4131
rect 41432 4128 41460 4168
rect 46750 4156 46756 4208
rect 46808 4196 46814 4208
rect 47949 4199 48007 4205
rect 47949 4196 47961 4199
rect 46808 4168 47961 4196
rect 46808 4156 46814 4168
rect 47949 4165 47961 4168
rect 47995 4165 48007 4199
rect 47949 4159 48007 4165
rect 46382 4128 46388 4140
rect 41432 4100 46388 4128
rect 41325 4091 41383 4097
rect 38654 4060 38660 4072
rect 38615 4032 38660 4060
rect 38654 4020 38660 4032
rect 38712 4020 38718 4072
rect 38841 4063 38899 4069
rect 38841 4029 38853 4063
rect 38887 4029 38899 4063
rect 41340 4060 41368 4091
rect 46382 4088 46388 4100
rect 46440 4088 46446 4140
rect 46845 4131 46903 4137
rect 46845 4097 46857 4131
rect 46891 4128 46903 4131
rect 46934 4128 46940 4140
rect 46891 4100 46940 4128
rect 46891 4097 46903 4100
rect 46845 4091 46903 4097
rect 46934 4088 46940 4100
rect 46992 4128 46998 4140
rect 47486 4128 47492 4140
rect 46992 4100 47492 4128
rect 46992 4088 46998 4100
rect 47486 4088 47492 4100
rect 47544 4088 47550 4140
rect 47210 4060 47216 4072
rect 41340 4032 47216 4060
rect 38841 4023 38899 4029
rect 38856 3992 38884 4023
rect 47210 4020 47216 4032
rect 47268 4020 47274 4072
rect 48133 3995 48191 4001
rect 48133 3992 48145 3995
rect 38396 3964 38884 3992
rect 38948 3964 48145 3992
rect 38948 3924 38976 3964
rect 48133 3961 48145 3964
rect 48179 3961 48191 3995
rect 48133 3955 48191 3961
rect 38120 3896 38976 3924
rect 41417 3927 41475 3933
rect 41417 3893 41429 3927
rect 41463 3924 41475 3927
rect 41598 3924 41604 3936
rect 41463 3896 41604 3924
rect 41463 3893 41475 3896
rect 41417 3887 41475 3893
rect 41598 3884 41604 3896
rect 41656 3884 41662 3936
rect 42426 3884 42432 3936
rect 42484 3924 42490 3936
rect 42613 3927 42671 3933
rect 42613 3924 42625 3927
rect 42484 3896 42625 3924
rect 42484 3884 42490 3896
rect 42613 3893 42625 3896
rect 42659 3893 42671 3927
rect 42613 3887 42671 3893
rect 43990 3884 43996 3936
rect 44048 3924 44054 3936
rect 44269 3927 44327 3933
rect 44269 3924 44281 3927
rect 44048 3896 44281 3924
rect 44048 3884 44054 3896
rect 44269 3893 44281 3896
rect 44315 3893 44327 3927
rect 44910 3924 44916 3936
rect 44871 3896 44916 3924
rect 44269 3887 44327 3893
rect 44910 3884 44916 3896
rect 44968 3884 44974 3936
rect 46474 3884 46480 3936
rect 46532 3924 46538 3936
rect 46937 3927 46995 3933
rect 46937 3924 46949 3927
rect 46532 3896 46949 3924
rect 46532 3884 46538 3896
rect 46937 3893 46949 3896
rect 46983 3893 46995 3927
rect 46937 3887 46995 3893
rect 1104 3834 48852 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 48852 3834
rect 1104 3760 48852 3782
rect 3878 3680 3884 3732
rect 3936 3720 3942 3732
rect 9306 3720 9312 3732
rect 3936 3692 6914 3720
rect 9267 3692 9312 3720
rect 3936 3680 3942 3692
rect 3234 3612 3240 3664
rect 3292 3652 3298 3664
rect 6886 3652 6914 3692
rect 9306 3680 9312 3692
rect 9364 3680 9370 3732
rect 11606 3680 11612 3732
rect 11664 3720 11670 3732
rect 13078 3720 13084 3732
rect 11664 3692 13084 3720
rect 11664 3680 11670 3692
rect 13078 3680 13084 3692
rect 13136 3680 13142 3732
rect 17862 3720 17868 3732
rect 13188 3692 17868 3720
rect 12158 3652 12164 3664
rect 3292 3624 4292 3652
rect 6886 3624 12164 3652
rect 3292 3612 3298 3624
rect 1394 3584 1400 3596
rect 1355 3556 1400 3584
rect 1394 3544 1400 3556
rect 1452 3544 1458 3596
rect 1854 3584 1860 3596
rect 1815 3556 1860 3584
rect 1854 3544 1860 3556
rect 1912 3544 1918 3596
rect 3786 3584 3792 3596
rect 3747 3556 3792 3584
rect 3786 3544 3792 3556
rect 3844 3544 3850 3596
rect 3970 3584 3976 3596
rect 3931 3556 3976 3584
rect 3970 3544 3976 3556
rect 4028 3544 4034 3596
rect 4264 3593 4292 3624
rect 12158 3612 12164 3624
rect 12216 3612 12222 3664
rect 12250 3612 12256 3664
rect 12308 3652 12314 3664
rect 12308 3624 12572 3652
rect 12308 3612 12314 3624
rect 4249 3587 4307 3593
rect 4249 3553 4261 3587
rect 4295 3553 4307 3587
rect 4249 3547 4307 3553
rect 11793 3587 11851 3593
rect 11793 3553 11805 3587
rect 11839 3584 11851 3587
rect 12434 3584 12440 3596
rect 11839 3556 12440 3584
rect 11839 3553 11851 3556
rect 11793 3547 11851 3553
rect 12434 3544 12440 3556
rect 12492 3544 12498 3596
rect 12544 3593 12572 3624
rect 12618 3612 12624 3664
rect 12676 3652 12682 3664
rect 13188 3652 13216 3692
rect 17862 3680 17868 3692
rect 17920 3680 17926 3732
rect 21450 3680 21456 3732
rect 21508 3720 21514 3732
rect 21508 3692 35112 3720
rect 21508 3680 21514 3692
rect 14090 3652 14096 3664
rect 12676 3624 13216 3652
rect 14003 3624 14096 3652
rect 12676 3612 12682 3624
rect 14090 3612 14096 3624
rect 14148 3652 14154 3664
rect 26878 3652 26884 3664
rect 14148 3624 26884 3652
rect 14148 3612 14154 3624
rect 26878 3612 26884 3624
rect 26936 3612 26942 3664
rect 27522 3612 27528 3664
rect 27580 3652 27586 3664
rect 31110 3652 31116 3664
rect 27580 3624 31116 3652
rect 27580 3612 27586 3624
rect 31110 3612 31116 3624
rect 31168 3612 31174 3664
rect 35084 3652 35112 3692
rect 38654 3680 38660 3732
rect 38712 3720 38718 3732
rect 38841 3723 38899 3729
rect 38841 3720 38853 3723
rect 38712 3692 38853 3720
rect 38712 3680 38718 3692
rect 38841 3689 38853 3692
rect 38887 3689 38899 3723
rect 38841 3683 38899 3689
rect 43438 3680 43444 3732
rect 43496 3720 43502 3732
rect 47026 3720 47032 3732
rect 43496 3692 47032 3720
rect 43496 3680 43502 3692
rect 47026 3680 47032 3692
rect 47084 3680 47090 3732
rect 48038 3652 48044 3664
rect 35084 3624 48044 3652
rect 48038 3612 48044 3624
rect 48096 3612 48102 3664
rect 12529 3587 12587 3593
rect 12529 3553 12541 3587
rect 12575 3553 12587 3587
rect 12529 3547 12587 3553
rect 6086 3516 6092 3528
rect 6047 3488 6092 3516
rect 6086 3476 6092 3488
rect 6144 3476 6150 3528
rect 6362 3476 6368 3528
rect 6420 3516 6426 3528
rect 6917 3519 6975 3525
rect 6917 3516 6929 3519
rect 6420 3488 6929 3516
rect 6420 3476 6426 3488
rect 6917 3485 6929 3488
rect 6963 3485 6975 3519
rect 6917 3479 6975 3485
rect 7469 3519 7527 3525
rect 7469 3485 7481 3519
rect 7515 3516 7527 3519
rect 9217 3519 9275 3525
rect 9217 3516 9229 3519
rect 7515 3488 9229 3516
rect 7515 3485 7527 3488
rect 7469 3479 7527 3485
rect 9217 3485 9229 3488
rect 9263 3516 9275 3519
rect 10778 3516 10784 3528
rect 9263 3488 10784 3516
rect 9263 3485 9275 3488
rect 9217 3479 9275 3485
rect 10778 3476 10784 3488
rect 10836 3476 10842 3528
rect 14108 3525 14136 3612
rect 15102 3584 15108 3596
rect 15063 3556 15108 3584
rect 15102 3544 15108 3556
rect 15160 3544 15166 3596
rect 15470 3584 15476 3596
rect 15431 3556 15476 3584
rect 15470 3544 15476 3556
rect 15528 3544 15534 3596
rect 20254 3584 20260 3596
rect 20215 3556 20260 3584
rect 20254 3544 20260 3556
rect 20312 3544 20318 3596
rect 20622 3584 20628 3596
rect 20583 3556 20628 3584
rect 20622 3544 20628 3556
rect 20680 3544 20686 3596
rect 25958 3584 25964 3596
rect 25919 3556 25964 3584
rect 25958 3544 25964 3556
rect 26016 3544 26022 3596
rect 26418 3584 26424 3596
rect 26379 3556 26424 3584
rect 26418 3544 26424 3556
rect 26476 3544 26482 3596
rect 27172 3556 30144 3584
rect 11149 3519 11207 3525
rect 11149 3485 11161 3519
rect 11195 3516 11207 3519
rect 11609 3519 11667 3525
rect 11609 3516 11621 3519
rect 11195 3488 11621 3516
rect 11195 3485 11207 3488
rect 11149 3479 11207 3485
rect 11609 3485 11621 3488
rect 11655 3485 11667 3519
rect 11609 3479 11667 3485
rect 14093 3519 14151 3525
rect 14093 3485 14105 3519
rect 14139 3485 14151 3519
rect 14918 3516 14924 3528
rect 14879 3488 14924 3516
rect 14093 3479 14151 3485
rect 14918 3476 14924 3488
rect 14976 3476 14982 3528
rect 20070 3516 20076 3528
rect 20031 3488 20076 3516
rect 20070 3476 20076 3488
rect 20128 3476 20134 3528
rect 23382 3476 23388 3528
rect 23440 3516 23446 3528
rect 23661 3519 23719 3525
rect 23661 3516 23673 3519
rect 23440 3488 23673 3516
rect 23440 3476 23446 3488
rect 23661 3485 23673 3488
rect 23707 3485 23719 3519
rect 25774 3516 25780 3528
rect 25735 3488 25780 3516
rect 23661 3479 23719 3485
rect 25774 3476 25780 3488
rect 25832 3476 25838 3528
rect 1581 3451 1639 3457
rect 1581 3417 1593 3451
rect 1627 3448 1639 3451
rect 2130 3448 2136 3460
rect 1627 3420 2136 3448
rect 1627 3417 1639 3420
rect 1581 3411 1639 3417
rect 2130 3408 2136 3420
rect 2188 3408 2194 3460
rect 8938 3408 8944 3460
rect 8996 3448 9002 3460
rect 18782 3448 18788 3460
rect 8996 3420 18788 3448
rect 8996 3408 9002 3420
rect 18782 3408 18788 3420
rect 18840 3408 18846 3460
rect 20806 3408 20812 3460
rect 20864 3448 20870 3460
rect 25682 3448 25688 3460
rect 20864 3420 25688 3448
rect 20864 3408 20870 3420
rect 25682 3408 25688 3420
rect 25740 3448 25746 3460
rect 27172 3448 27200 3556
rect 28994 3516 29000 3528
rect 28955 3488 29000 3516
rect 28994 3476 29000 3488
rect 29052 3476 29058 3528
rect 29270 3476 29276 3528
rect 29328 3516 29334 3528
rect 29541 3519 29599 3525
rect 29541 3516 29553 3519
rect 29328 3488 29553 3516
rect 29328 3476 29334 3488
rect 29541 3485 29553 3488
rect 29587 3485 29599 3519
rect 30116 3518 30144 3556
rect 31570 3544 31576 3596
rect 31628 3584 31634 3596
rect 31665 3587 31723 3593
rect 31665 3584 31677 3587
rect 31628 3556 31677 3584
rect 31628 3544 31634 3556
rect 31665 3553 31677 3556
rect 31711 3553 31723 3587
rect 36446 3584 36452 3596
rect 36407 3556 36452 3584
rect 31665 3547 31723 3553
rect 36446 3544 36452 3556
rect 36504 3544 36510 3596
rect 36722 3584 36728 3596
rect 36683 3556 36728 3584
rect 36722 3544 36728 3556
rect 36780 3544 36786 3596
rect 37182 3544 37188 3596
rect 37240 3584 37246 3596
rect 41598 3584 41604 3596
rect 37240 3556 39896 3584
rect 41559 3556 41604 3584
rect 37240 3544 37246 3556
rect 30193 3519 30251 3525
rect 30193 3518 30205 3519
rect 30116 3490 30205 3518
rect 29541 3479 29599 3485
rect 30193 3485 30205 3490
rect 30239 3485 30251 3519
rect 31202 3516 31208 3528
rect 31163 3488 31208 3516
rect 30193 3479 30251 3485
rect 31202 3476 31208 3488
rect 31260 3476 31266 3528
rect 36262 3516 36268 3528
rect 36223 3488 36268 3516
rect 36262 3476 36268 3488
rect 36320 3476 36326 3528
rect 39868 3525 39896 3556
rect 41598 3544 41604 3556
rect 41656 3544 41662 3596
rect 41874 3584 41880 3596
rect 41835 3556 41880 3584
rect 41874 3544 41880 3556
rect 41932 3544 41938 3596
rect 42058 3544 42064 3596
rect 42116 3584 42122 3596
rect 46198 3584 46204 3596
rect 42116 3556 46204 3584
rect 42116 3544 42122 3556
rect 46198 3544 46204 3556
rect 46256 3544 46262 3596
rect 46474 3584 46480 3596
rect 46435 3556 46480 3584
rect 46474 3544 46480 3556
rect 46532 3544 46538 3596
rect 39853 3519 39911 3525
rect 39853 3485 39865 3519
rect 39899 3485 39911 3519
rect 39853 3479 39911 3485
rect 40957 3519 41015 3525
rect 40957 3485 40969 3519
rect 41003 3516 41015 3519
rect 41417 3519 41475 3525
rect 41417 3516 41429 3519
rect 41003 3488 41429 3516
rect 41003 3485 41015 3488
rect 40957 3479 41015 3485
rect 41417 3485 41429 3488
rect 41463 3485 41475 3519
rect 43898 3516 43904 3528
rect 43859 3488 43904 3516
rect 41417 3479 41475 3485
rect 43898 3476 43904 3488
rect 43956 3476 43962 3528
rect 45005 3519 45063 3525
rect 45005 3485 45017 3519
rect 45051 3516 45063 3519
rect 45833 3519 45891 3525
rect 45051 3488 45554 3516
rect 45051 3485 45063 3488
rect 45005 3479 45063 3485
rect 29638 3448 29644 3460
rect 25740 3420 27200 3448
rect 29599 3420 29644 3448
rect 25740 3408 25746 3420
rect 29638 3408 29644 3420
rect 29696 3408 29702 3460
rect 29822 3408 29828 3460
rect 29880 3448 29886 3460
rect 31386 3448 31392 3460
rect 29880 3420 30420 3448
rect 31347 3420 31392 3448
rect 29880 3408 29886 3420
rect 1302 3340 1308 3392
rect 1360 3380 1366 3392
rect 3326 3380 3332 3392
rect 1360 3352 3332 3380
rect 1360 3340 1366 3352
rect 3326 3340 3332 3352
rect 3384 3340 3390 3392
rect 6181 3383 6239 3389
rect 6181 3349 6193 3383
rect 6227 3380 6239 3383
rect 6546 3380 6552 3392
rect 6227 3352 6552 3380
rect 6227 3349 6239 3352
rect 6181 3343 6239 3349
rect 6546 3340 6552 3352
rect 6604 3340 6610 3392
rect 6914 3340 6920 3392
rect 6972 3380 6978 3392
rect 7561 3383 7619 3389
rect 7561 3380 7573 3383
rect 6972 3352 7573 3380
rect 6972 3340 6978 3352
rect 7561 3349 7573 3352
rect 7607 3349 7619 3383
rect 7561 3343 7619 3349
rect 12434 3340 12440 3392
rect 12492 3380 12498 3392
rect 14185 3383 14243 3389
rect 14185 3380 14197 3383
rect 12492 3352 14197 3380
rect 12492 3340 12498 3352
rect 14185 3349 14197 3352
rect 14231 3349 14243 3383
rect 14185 3343 14243 3349
rect 14642 3340 14648 3392
rect 14700 3380 14706 3392
rect 25498 3380 25504 3392
rect 14700 3352 25504 3380
rect 14700 3340 14706 3352
rect 25498 3340 25504 3352
rect 25556 3380 25562 3392
rect 29454 3380 29460 3392
rect 25556 3352 29460 3380
rect 25556 3340 25562 3352
rect 29454 3340 29460 3352
rect 29512 3340 29518 3392
rect 29914 3340 29920 3392
rect 29972 3380 29978 3392
rect 30285 3383 30343 3389
rect 30285 3380 30297 3383
rect 29972 3352 30297 3380
rect 29972 3340 29978 3352
rect 30285 3349 30297 3352
rect 30331 3349 30343 3383
rect 30392 3380 30420 3420
rect 31386 3408 31392 3420
rect 31444 3408 31450 3460
rect 43438 3448 43444 3460
rect 31726 3420 43444 3448
rect 31726 3380 31754 3420
rect 43438 3408 43444 3420
rect 43496 3408 43502 3460
rect 45526 3448 45554 3488
rect 45833 3485 45845 3519
rect 45879 3516 45891 3519
rect 46293 3519 46351 3525
rect 46293 3516 46305 3519
rect 45879 3488 46305 3516
rect 45879 3485 45891 3488
rect 45833 3479 45891 3485
rect 46293 3485 46305 3488
rect 46339 3485 46351 3519
rect 46293 3479 46351 3485
rect 46934 3448 46940 3460
rect 45526 3420 46940 3448
rect 46934 3408 46940 3420
rect 46992 3408 46998 3460
rect 48133 3451 48191 3457
rect 48133 3417 48145 3451
rect 48179 3448 48191 3451
rect 48314 3448 48320 3460
rect 48179 3420 48320 3448
rect 48179 3417 48191 3420
rect 48133 3411 48191 3417
rect 48314 3408 48320 3420
rect 48372 3408 48378 3460
rect 30392 3352 31754 3380
rect 39945 3383 40003 3389
rect 30285 3343 30343 3349
rect 39945 3349 39957 3383
rect 39991 3380 40003 3383
rect 40034 3380 40040 3392
rect 39991 3352 40040 3380
rect 39991 3349 40003 3352
rect 39945 3343 40003 3349
rect 40034 3340 40040 3352
rect 40092 3340 40098 3392
rect 43993 3383 44051 3389
rect 43993 3349 44005 3383
rect 44039 3380 44051 3383
rect 44174 3380 44180 3392
rect 44039 3352 44180 3380
rect 44039 3349 44051 3352
rect 43993 3343 44051 3349
rect 44174 3340 44180 3352
rect 44232 3340 44238 3392
rect 45097 3383 45155 3389
rect 45097 3349 45109 3383
rect 45143 3380 45155 3383
rect 45186 3380 45192 3392
rect 45143 3352 45192 3380
rect 45143 3349 45155 3352
rect 45097 3343 45155 3349
rect 45186 3340 45192 3352
rect 45244 3340 45250 3392
rect 1104 3290 48852 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 48852 3290
rect 1104 3216 48852 3238
rect 2130 3176 2136 3188
rect 2091 3148 2136 3176
rect 2130 3136 2136 3148
rect 2188 3136 2194 3188
rect 2406 3136 2412 3188
rect 2464 3176 2470 3188
rect 22554 3176 22560 3188
rect 2464 3148 22560 3176
rect 2464 3136 2470 3148
rect 22554 3136 22560 3148
rect 22612 3136 22618 3188
rect 22646 3136 22652 3188
rect 22704 3176 22710 3188
rect 22833 3179 22891 3185
rect 22833 3176 22845 3179
rect 22704 3148 22845 3176
rect 22704 3136 22710 3148
rect 22833 3145 22845 3148
rect 22879 3145 22891 3179
rect 22833 3139 22891 3145
rect 23124 3148 23704 3176
rect 4157 3111 4215 3117
rect 4157 3077 4169 3111
rect 4203 3108 4215 3111
rect 4890 3108 4896 3120
rect 4203 3080 4896 3108
rect 4203 3077 4215 3080
rect 4157 3071 4215 3077
rect 4890 3068 4896 3080
rect 4948 3068 4954 3120
rect 6546 3108 6552 3120
rect 6507 3080 6552 3108
rect 6546 3068 6552 3080
rect 6604 3068 6610 3120
rect 10229 3111 10287 3117
rect 10229 3077 10241 3111
rect 10275 3108 10287 3111
rect 17862 3108 17868 3120
rect 10275 3080 17868 3108
rect 10275 3077 10287 3080
rect 10229 3071 10287 3077
rect 17862 3068 17868 3080
rect 17920 3068 17926 3120
rect 18138 3108 18144 3120
rect 18099 3080 18144 3108
rect 18138 3068 18144 3080
rect 18196 3068 18202 3120
rect 19978 3068 19984 3120
rect 20036 3108 20042 3120
rect 20036 3080 20944 3108
rect 20036 3068 20042 3080
rect 1946 3000 1952 3052
rect 2004 3040 2010 3052
rect 2041 3043 2099 3049
rect 2041 3040 2053 3043
rect 2004 3012 2053 3040
rect 2004 3000 2010 3012
rect 2041 3009 2053 3012
rect 2087 3009 2099 3043
rect 6362 3040 6368 3052
rect 6323 3012 6368 3040
rect 2041 3003 2099 3009
rect 2056 2904 2084 3003
rect 6362 3000 6368 3012
rect 6420 3000 6426 3052
rect 8938 3040 8944 3052
rect 8899 3012 8944 3040
rect 8938 3000 8944 3012
rect 8996 3000 9002 3052
rect 9674 3000 9680 3052
rect 9732 3040 9738 3052
rect 10045 3043 10103 3049
rect 10045 3040 10057 3043
rect 9732 3012 10057 3040
rect 9732 3000 9738 3012
rect 10045 3009 10057 3012
rect 10091 3009 10103 3043
rect 10045 3003 10103 3009
rect 12158 3000 12164 3052
rect 12216 3040 12222 3052
rect 12253 3043 12311 3049
rect 12253 3040 12265 3043
rect 12216 3012 12265 3040
rect 12216 3000 12222 3012
rect 12253 3009 12265 3012
rect 12299 3009 12311 3043
rect 12253 3003 12311 3009
rect 14182 3000 14188 3052
rect 14240 3040 14246 3052
rect 14553 3043 14611 3049
rect 14553 3040 14565 3043
rect 14240 3012 14565 3040
rect 14240 3000 14246 3012
rect 14553 3009 14565 3012
rect 14599 3009 14611 3043
rect 14553 3003 14611 3009
rect 14918 3000 14924 3052
rect 14976 3040 14982 3052
rect 15473 3043 15531 3049
rect 15473 3040 15485 3043
rect 14976 3012 15485 3040
rect 14976 3000 14982 3012
rect 15473 3009 15485 3012
rect 15519 3009 15531 3043
rect 17954 3040 17960 3052
rect 17915 3012 17960 3040
rect 15473 3003 15531 3009
rect 17954 3000 17960 3012
rect 18012 3000 18018 3052
rect 20070 3000 20076 3052
rect 20128 3040 20134 3052
rect 20916 3049 20944 3080
rect 20441 3043 20499 3049
rect 20441 3040 20453 3043
rect 20128 3012 20453 3040
rect 20128 3000 20134 3012
rect 20441 3009 20453 3012
rect 20487 3009 20499 3043
rect 20441 3003 20499 3009
rect 20901 3043 20959 3049
rect 20901 3009 20913 3043
rect 20947 3009 20959 3043
rect 20901 3003 20959 3009
rect 22554 3000 22560 3052
rect 22612 3040 22618 3052
rect 22741 3043 22799 3049
rect 22741 3040 22753 3043
rect 22612 3012 22753 3040
rect 22612 3000 22618 3012
rect 22741 3009 22753 3012
rect 22787 3009 22799 3043
rect 22741 3003 22799 3009
rect 3973 2975 4031 2981
rect 3973 2941 3985 2975
rect 4019 2972 4031 2975
rect 4614 2972 4620 2984
rect 4019 2944 4620 2972
rect 4019 2941 4031 2944
rect 3973 2935 4031 2941
rect 4614 2932 4620 2944
rect 4672 2932 4678 2984
rect 5166 2972 5172 2984
rect 5127 2944 5172 2972
rect 5166 2932 5172 2944
rect 5224 2932 5230 2984
rect 6546 2932 6552 2984
rect 6604 2972 6610 2984
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 6604 2944 6837 2972
rect 6604 2932 6610 2944
rect 6825 2941 6837 2944
rect 6871 2941 6883 2975
rect 6825 2935 6883 2941
rect 7742 2932 7748 2984
rect 7800 2972 7806 2984
rect 8665 2975 8723 2981
rect 8665 2972 8677 2975
rect 7800 2944 8677 2972
rect 7800 2932 7806 2944
rect 8665 2941 8677 2944
rect 8711 2941 8723 2975
rect 8665 2935 8723 2941
rect 12176 2928 12388 2956
rect 12434 2932 12440 2984
rect 12492 2972 12498 2984
rect 12894 2972 12900 2984
rect 12492 2944 12537 2972
rect 12855 2944 12900 2972
rect 12492 2932 12498 2944
rect 12894 2932 12900 2944
rect 12952 2932 12958 2984
rect 18138 2932 18144 2984
rect 18196 2972 18202 2984
rect 18417 2975 18475 2981
rect 18417 2972 18429 2975
rect 18196 2944 18429 2972
rect 18196 2932 18202 2944
rect 18417 2941 18429 2944
rect 18463 2941 18475 2975
rect 18417 2935 18475 2941
rect 12176 2904 12204 2928
rect 2056 2876 12204 2904
rect 12360 2904 12388 2928
rect 14642 2904 14648 2916
rect 12360 2876 14648 2904
rect 14642 2864 14648 2876
rect 14700 2864 14706 2916
rect 14737 2907 14795 2913
rect 14737 2873 14749 2907
rect 14783 2904 14795 2907
rect 23124 2904 23152 3148
rect 23566 3108 23572 3120
rect 23527 3080 23572 3108
rect 23566 3068 23572 3080
rect 23624 3068 23630 3120
rect 23676 3108 23704 3148
rect 26142 3136 26148 3188
rect 26200 3176 26206 3188
rect 26973 3179 27031 3185
rect 26973 3176 26985 3179
rect 26200 3148 26985 3176
rect 26200 3136 26206 3148
rect 26973 3145 26985 3148
rect 27019 3145 27031 3179
rect 26973 3139 27031 3145
rect 28902 3136 28908 3188
rect 28960 3176 28966 3188
rect 30834 3176 30840 3188
rect 28960 3148 30840 3176
rect 28960 3136 28966 3148
rect 30834 3136 30840 3148
rect 30892 3136 30898 3188
rect 36170 3136 36176 3188
rect 36228 3176 36234 3188
rect 36228 3148 40356 3176
rect 36228 3136 36234 3148
rect 29914 3108 29920 3120
rect 23676 3080 27292 3108
rect 29875 3080 29920 3108
rect 23382 3040 23388 3052
rect 23343 3012 23388 3040
rect 23382 3000 23388 3012
rect 23440 3000 23446 3052
rect 25774 3000 25780 3052
rect 25832 3040 25838 3052
rect 26053 3043 26111 3049
rect 26053 3040 26065 3043
rect 25832 3012 26065 3040
rect 25832 3000 25838 3012
rect 26053 3009 26065 3012
rect 26099 3009 26111 3043
rect 26053 3003 26111 3009
rect 27157 3043 27215 3049
rect 27157 3009 27169 3043
rect 27203 3009 27215 3043
rect 27157 3003 27215 3009
rect 23842 2972 23848 2984
rect 23803 2944 23848 2972
rect 23842 2932 23848 2944
rect 23900 2932 23906 2984
rect 14783 2876 23152 2904
rect 14783 2873 14795 2876
rect 14737 2867 14795 2873
rect 23198 2864 23204 2916
rect 23256 2904 23262 2916
rect 27172 2904 27200 3003
rect 23256 2876 27200 2904
rect 27264 2904 27292 3080
rect 29914 3068 29920 3080
rect 29972 3068 29978 3120
rect 32398 3108 32404 3120
rect 32359 3080 32404 3108
rect 32398 3068 32404 3080
rect 32456 3068 32462 3120
rect 33042 3068 33048 3120
rect 33100 3108 33106 3120
rect 40218 3108 40224 3120
rect 33100 3080 39804 3108
rect 40179 3080 40224 3108
rect 33100 3068 33106 3080
rect 29730 3040 29736 3052
rect 29691 3012 29736 3040
rect 29730 3000 29736 3012
rect 29788 3000 29794 3052
rect 36262 3000 36268 3052
rect 36320 3040 36326 3052
rect 36541 3043 36599 3049
rect 36541 3040 36553 3043
rect 36320 3012 36553 3040
rect 36320 3000 36326 3012
rect 36541 3009 36553 3012
rect 36587 3009 36599 3043
rect 36541 3003 36599 3009
rect 30282 2972 30288 2984
rect 30243 2944 30288 2972
rect 30282 2932 30288 2944
rect 30340 2932 30346 2984
rect 32217 2975 32275 2981
rect 32217 2941 32229 2975
rect 32263 2972 32275 2975
rect 32950 2972 32956 2984
rect 32263 2944 32956 2972
rect 32263 2941 32275 2944
rect 32217 2935 32275 2941
rect 32950 2932 32956 2944
rect 33008 2932 33014 2984
rect 33413 2975 33471 2981
rect 33413 2941 33425 2975
rect 33459 2972 33471 2975
rect 33459 2944 33548 2972
rect 33459 2941 33471 2944
rect 33413 2935 33471 2941
rect 33520 2916 33548 2944
rect 37734 2932 37740 2984
rect 37792 2972 37798 2984
rect 37792 2944 39712 2972
rect 37792 2932 37798 2944
rect 30742 2904 30748 2916
rect 27264 2876 30748 2904
rect 23256 2864 23262 2876
rect 30742 2864 30748 2876
rect 30800 2864 30806 2916
rect 33502 2864 33508 2916
rect 33560 2864 33566 2916
rect 10962 2796 10968 2848
rect 11020 2836 11026 2848
rect 16574 2836 16580 2848
rect 11020 2808 16580 2836
rect 11020 2796 11026 2808
rect 16574 2796 16580 2808
rect 16632 2796 16638 2848
rect 20993 2839 21051 2845
rect 20993 2805 21005 2839
rect 21039 2836 21051 2839
rect 22002 2836 22008 2848
rect 21039 2808 22008 2836
rect 21039 2805 21051 2808
rect 20993 2799 21051 2805
rect 22002 2796 22008 2808
rect 22060 2796 22066 2848
rect 26878 2796 26884 2848
rect 26936 2836 26942 2848
rect 33410 2836 33416 2848
rect 26936 2808 33416 2836
rect 26936 2796 26942 2808
rect 33410 2796 33416 2808
rect 33468 2796 33474 2848
rect 39574 2836 39580 2848
rect 39535 2808 39580 2836
rect 39574 2796 39580 2808
rect 39632 2796 39638 2848
rect 39684 2836 39712 2944
rect 39776 2904 39804 3080
rect 40218 3068 40224 3080
rect 40276 3068 40282 3120
rect 40328 3108 40356 3148
rect 40402 3136 40408 3188
rect 40460 3176 40466 3188
rect 43898 3176 43904 3188
rect 40460 3148 43904 3176
rect 40460 3136 40466 3148
rect 43898 3136 43904 3148
rect 43956 3136 43962 3188
rect 46106 3136 46112 3188
rect 46164 3176 46170 3188
rect 46477 3179 46535 3185
rect 46477 3176 46489 3179
rect 46164 3148 46489 3176
rect 46164 3136 46170 3148
rect 46477 3145 46489 3148
rect 46523 3145 46535 3179
rect 48038 3176 48044 3188
rect 47999 3148 48044 3176
rect 46477 3139 46535 3145
rect 48038 3136 48044 3148
rect 48096 3136 48102 3188
rect 44174 3108 44180 3120
rect 40328 3080 42748 3108
rect 44135 3080 44180 3108
rect 42429 3043 42487 3049
rect 42429 3009 42441 3043
rect 42475 3009 42487 3043
rect 42429 3003 42487 3009
rect 40037 2975 40095 2981
rect 40037 2941 40049 2975
rect 40083 2972 40095 2975
rect 40494 2972 40500 2984
rect 40083 2944 40500 2972
rect 40083 2941 40095 2944
rect 40037 2935 40095 2941
rect 40494 2932 40500 2944
rect 40552 2932 40558 2984
rect 41230 2972 41236 2984
rect 41191 2944 41236 2972
rect 41230 2932 41236 2944
rect 41288 2932 41294 2984
rect 40402 2904 40408 2916
rect 39776 2876 40408 2904
rect 40402 2864 40408 2876
rect 40460 2864 40466 2916
rect 42444 2904 42472 3003
rect 41386 2876 42472 2904
rect 41386 2836 41414 2876
rect 39684 2808 41414 2836
rect 42521 2839 42579 2845
rect 42521 2805 42533 2839
rect 42567 2836 42579 2839
rect 42610 2836 42616 2848
rect 42567 2808 42616 2836
rect 42567 2805 42579 2808
rect 42521 2799 42579 2805
rect 42610 2796 42616 2808
rect 42668 2796 42674 2848
rect 42720 2836 42748 3080
rect 44174 3068 44180 3080
rect 44232 3068 44238 3120
rect 43162 3000 43168 3052
rect 43220 3040 43226 3052
rect 43257 3043 43315 3049
rect 43257 3040 43269 3043
rect 43220 3012 43269 3040
rect 43220 3000 43226 3012
rect 43257 3009 43269 3012
rect 43303 3009 43315 3043
rect 43990 3040 43996 3052
rect 43951 3012 43996 3040
rect 43257 3003 43315 3009
rect 43990 3000 43996 3012
rect 44048 3000 44054 3052
rect 45738 3000 45744 3052
rect 45796 3040 45802 3052
rect 46293 3043 46351 3049
rect 46293 3040 46305 3043
rect 45796 3012 46305 3040
rect 45796 3000 45802 3012
rect 46293 3009 46305 3012
rect 46339 3009 46351 3043
rect 46293 3003 46351 3009
rect 47857 3043 47915 3049
rect 47857 3009 47869 3043
rect 47903 3040 47915 3043
rect 49602 3040 49608 3052
rect 47903 3012 49608 3040
rect 47903 3009 47915 3012
rect 47857 3003 47915 3009
rect 49602 3000 49608 3012
rect 49660 3000 49666 3052
rect 44450 2972 44456 2984
rect 44411 2944 44456 2972
rect 44450 2932 44456 2944
rect 44508 2932 44514 2984
rect 43438 2904 43444 2916
rect 43399 2876 43444 2904
rect 43438 2864 43444 2876
rect 43496 2864 43502 2916
rect 45646 2836 45652 2848
rect 42720 2808 45652 2836
rect 45646 2796 45652 2808
rect 45704 2796 45710 2848
rect 1104 2746 48852 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 48852 2746
rect 1104 2672 48852 2694
rect 3142 2592 3148 2644
rect 3200 2632 3206 2644
rect 3200 2604 10180 2632
rect 3200 2592 3206 2604
rect 2961 2567 3019 2573
rect 2961 2533 2973 2567
rect 3007 2564 3019 2567
rect 3694 2564 3700 2576
rect 3007 2536 3700 2564
rect 3007 2533 3019 2536
rect 2961 2527 3019 2533
rect 3694 2524 3700 2536
rect 3752 2524 3758 2576
rect 4798 2564 4804 2576
rect 4759 2536 4804 2564
rect 4798 2524 4804 2536
rect 4856 2524 4862 2576
rect 5810 2524 5816 2576
rect 5868 2564 5874 2576
rect 5868 2536 7052 2564
rect 5868 2524 5874 2536
rect 6454 2496 6460 2508
rect 6415 2468 6460 2496
rect 6454 2456 6460 2468
rect 6512 2456 6518 2508
rect 6641 2499 6699 2505
rect 6641 2465 6653 2499
rect 6687 2496 6699 2499
rect 6914 2496 6920 2508
rect 6687 2468 6920 2496
rect 6687 2465 6699 2468
rect 6641 2459 6699 2465
rect 6914 2456 6920 2468
rect 6972 2456 6978 2508
rect 7024 2505 7052 2536
rect 7009 2499 7067 2505
rect 7009 2465 7021 2499
rect 7055 2465 7067 2499
rect 7009 2459 7067 2465
rect 7098 2456 7104 2508
rect 7156 2496 7162 2508
rect 8941 2499 8999 2505
rect 8941 2496 8953 2499
rect 7156 2468 8953 2496
rect 7156 2456 7162 2468
rect 8941 2465 8953 2468
rect 8987 2465 8999 2499
rect 10152 2496 10180 2604
rect 12158 2592 12164 2644
rect 12216 2632 12222 2644
rect 12437 2635 12495 2641
rect 12437 2632 12449 2635
rect 12216 2604 12449 2632
rect 12216 2592 12222 2604
rect 12437 2601 12449 2604
rect 12483 2601 12495 2635
rect 12437 2595 12495 2601
rect 22094 2592 22100 2644
rect 22152 2632 22158 2644
rect 45830 2632 45836 2644
rect 22152 2604 45836 2632
rect 22152 2592 22158 2604
rect 45830 2592 45836 2604
rect 45888 2592 45894 2644
rect 10413 2567 10471 2573
rect 10413 2533 10425 2567
rect 10459 2564 10471 2567
rect 20349 2567 20407 2573
rect 10459 2536 20300 2564
rect 10459 2533 10471 2536
rect 10413 2527 10471 2533
rect 12526 2496 12532 2508
rect 10152 2468 12532 2496
rect 8941 2459 8999 2465
rect 12526 2456 12532 2468
rect 12584 2456 12590 2508
rect 13538 2456 13544 2508
rect 13596 2496 13602 2508
rect 14553 2499 14611 2505
rect 14553 2496 14565 2499
rect 13596 2468 14565 2496
rect 13596 2456 13602 2468
rect 14553 2465 14565 2468
rect 14599 2465 14611 2499
rect 14553 2459 14611 2465
rect 1946 2388 1952 2440
rect 2004 2428 2010 2440
rect 2777 2431 2835 2437
rect 2777 2428 2789 2431
rect 2004 2400 2789 2428
rect 2004 2388 2010 2400
rect 2777 2397 2789 2400
rect 2823 2397 2835 2431
rect 2777 2391 2835 2397
rect 4522 2388 4528 2440
rect 4580 2428 4586 2440
rect 4617 2431 4675 2437
rect 4617 2428 4629 2431
rect 4580 2400 4629 2428
rect 4580 2388 4586 2400
rect 4617 2397 4629 2400
rect 4663 2397 4675 2431
rect 4617 2391 4675 2397
rect 10229 2431 10287 2437
rect 10229 2397 10241 2431
rect 10275 2397 10287 2431
rect 10229 2391 10287 2397
rect 13081 2431 13139 2437
rect 13081 2397 13093 2431
rect 13127 2428 13139 2431
rect 14093 2431 14151 2437
rect 14093 2428 14105 2431
rect 13127 2400 14105 2428
rect 13127 2397 13139 2400
rect 13081 2391 13139 2397
rect 14093 2397 14105 2400
rect 14139 2397 14151 2431
rect 14093 2391 14151 2397
rect 1854 2360 1860 2372
rect 1815 2332 1860 2360
rect 1854 2320 1860 2332
rect 1912 2320 1918 2372
rect 2222 2360 2228 2372
rect 2183 2332 2228 2360
rect 2222 2320 2228 2332
rect 2280 2320 2286 2372
rect 8386 2320 8392 2372
rect 8444 2360 8450 2372
rect 10244 2360 10272 2391
rect 17402 2388 17408 2440
rect 17460 2428 17466 2440
rect 17497 2431 17555 2437
rect 17497 2428 17509 2431
rect 17460 2400 17509 2428
rect 17460 2388 17466 2400
rect 17497 2397 17509 2400
rect 17543 2397 17555 2431
rect 17497 2391 17555 2397
rect 14274 2360 14280 2372
rect 8444 2332 10272 2360
rect 14235 2332 14280 2360
rect 8444 2320 8450 2332
rect 14274 2320 14280 2332
rect 14332 2320 14338 2372
rect 19978 2320 19984 2372
rect 20036 2360 20042 2372
rect 20165 2363 20223 2369
rect 20165 2360 20177 2363
rect 20036 2332 20177 2360
rect 20036 2320 20042 2332
rect 20165 2329 20177 2332
rect 20211 2329 20223 2363
rect 20272 2360 20300 2536
rect 20349 2533 20361 2567
rect 20395 2564 20407 2567
rect 20990 2564 20996 2576
rect 20395 2536 20996 2564
rect 20395 2533 20407 2536
rect 20349 2527 20407 2533
rect 20990 2524 20996 2536
rect 21048 2524 21054 2576
rect 21266 2524 21272 2576
rect 21324 2564 21330 2576
rect 21324 2536 22324 2564
rect 21324 2524 21330 2536
rect 20898 2456 20904 2508
rect 20956 2496 20962 2508
rect 21821 2499 21879 2505
rect 21821 2496 21833 2499
rect 20956 2468 21833 2496
rect 20956 2456 20962 2468
rect 21821 2465 21833 2468
rect 21867 2465 21879 2499
rect 22002 2496 22008 2508
rect 21963 2468 22008 2496
rect 21821 2459 21879 2465
rect 22002 2456 22008 2468
rect 22060 2456 22066 2508
rect 22296 2505 22324 2536
rect 23106 2524 23112 2576
rect 23164 2564 23170 2576
rect 27341 2567 27399 2573
rect 27341 2564 27353 2567
rect 23164 2536 27353 2564
rect 23164 2524 23170 2536
rect 27341 2533 27353 2536
rect 27387 2533 27399 2567
rect 27341 2527 27399 2533
rect 28074 2524 28080 2576
rect 28132 2564 28138 2576
rect 28169 2567 28227 2573
rect 28169 2564 28181 2567
rect 28132 2536 28181 2564
rect 28132 2524 28138 2536
rect 28169 2533 28181 2536
rect 28215 2533 28227 2567
rect 28169 2527 28227 2533
rect 32674 2524 32680 2576
rect 32732 2564 32738 2576
rect 34149 2567 34207 2573
rect 34149 2564 34161 2567
rect 32732 2536 34161 2564
rect 32732 2524 32738 2536
rect 34149 2533 34161 2536
rect 34195 2533 34207 2567
rect 34149 2527 34207 2533
rect 39942 2524 39948 2576
rect 40000 2564 40006 2576
rect 40000 2536 40356 2564
rect 40000 2524 40006 2536
rect 22281 2499 22339 2505
rect 22281 2465 22293 2499
rect 22327 2465 22339 2499
rect 22281 2459 22339 2465
rect 24670 2456 24676 2508
rect 24728 2496 24734 2508
rect 26142 2496 26148 2508
rect 24728 2468 26148 2496
rect 24728 2456 24734 2468
rect 26142 2456 26148 2468
rect 26200 2456 26206 2508
rect 26237 2499 26295 2505
rect 26237 2465 26249 2499
rect 26283 2496 26295 2499
rect 28718 2496 28724 2508
rect 26283 2468 28724 2496
rect 26283 2465 26295 2468
rect 26237 2459 26295 2465
rect 28718 2456 28724 2468
rect 28776 2456 28782 2508
rect 28994 2456 29000 2508
rect 29052 2496 29058 2508
rect 29549 2499 29607 2505
rect 29549 2496 29561 2499
rect 29052 2468 29561 2496
rect 29052 2456 29058 2468
rect 29549 2465 29561 2468
rect 29595 2465 29607 2499
rect 29730 2496 29736 2508
rect 29691 2468 29736 2496
rect 29549 2459 29607 2465
rect 29730 2456 29736 2468
rect 29788 2456 29794 2508
rect 30926 2496 30932 2508
rect 30887 2468 30932 2496
rect 30926 2456 30932 2468
rect 30984 2456 30990 2508
rect 32490 2456 32496 2508
rect 32548 2496 32554 2508
rect 35345 2499 35403 2505
rect 35345 2496 35357 2499
rect 32548 2468 35357 2496
rect 32548 2456 32554 2468
rect 35345 2465 35357 2468
rect 35391 2465 35403 2499
rect 35345 2459 35403 2465
rect 39574 2456 39580 2508
rect 39632 2496 39638 2508
rect 39853 2499 39911 2505
rect 39853 2496 39865 2499
rect 39632 2468 39865 2496
rect 39632 2456 39638 2468
rect 39853 2465 39865 2468
rect 39899 2465 39911 2499
rect 40034 2496 40040 2508
rect 39995 2468 40040 2496
rect 39853 2459 39911 2465
rect 40034 2456 40040 2468
rect 40092 2456 40098 2508
rect 40328 2505 40356 2536
rect 40313 2499 40371 2505
rect 40313 2465 40325 2499
rect 40359 2465 40371 2499
rect 42426 2496 42432 2508
rect 42387 2468 42432 2496
rect 40313 2459 40371 2465
rect 42426 2456 42432 2468
rect 42484 2456 42490 2508
rect 42610 2496 42616 2508
rect 42571 2468 42616 2496
rect 42610 2456 42616 2468
rect 42668 2456 42674 2508
rect 42702 2456 42708 2508
rect 42760 2496 42766 2508
rect 42889 2499 42947 2505
rect 42889 2496 42901 2499
rect 42760 2468 42901 2496
rect 42760 2456 42766 2468
rect 42889 2465 42901 2468
rect 42935 2465 42947 2499
rect 42889 2459 42947 2465
rect 44910 2456 44916 2508
rect 44968 2496 44974 2508
rect 45005 2499 45063 2505
rect 45005 2496 45017 2499
rect 44968 2468 45017 2496
rect 44968 2456 44974 2468
rect 45005 2465 45017 2468
rect 45051 2465 45063 2499
rect 45186 2496 45192 2508
rect 45147 2468 45192 2496
rect 45005 2459 45063 2465
rect 45186 2456 45192 2468
rect 45244 2456 45250 2508
rect 45370 2456 45376 2508
rect 45428 2496 45434 2508
rect 45557 2499 45615 2505
rect 45557 2496 45569 2499
rect 45428 2468 45569 2496
rect 45428 2456 45434 2468
rect 45557 2465 45569 2468
rect 45603 2465 45615 2499
rect 45557 2459 45615 2465
rect 25501 2431 25559 2437
rect 25501 2397 25513 2431
rect 25547 2428 25559 2431
rect 25547 2400 26234 2428
rect 25547 2397 25559 2400
rect 25501 2391 25559 2397
rect 22922 2360 22928 2372
rect 20272 2332 22928 2360
rect 20165 2323 20223 2329
rect 22922 2320 22928 2332
rect 22980 2320 22986 2372
rect 25130 2320 25136 2372
rect 25188 2360 25194 2372
rect 25317 2363 25375 2369
rect 25317 2360 25329 2363
rect 25188 2332 25329 2360
rect 25188 2320 25194 2332
rect 25317 2329 25329 2332
rect 25363 2329 25375 2363
rect 25317 2323 25375 2329
rect 26053 2363 26111 2369
rect 26053 2329 26065 2363
rect 26099 2329 26111 2363
rect 26206 2360 26234 2400
rect 27062 2388 27068 2440
rect 27120 2428 27126 2440
rect 27157 2431 27215 2437
rect 27157 2428 27169 2431
rect 27120 2400 27169 2428
rect 27120 2388 27126 2400
rect 27157 2397 27169 2400
rect 27203 2397 27215 2431
rect 28258 2428 28264 2440
rect 27157 2391 27215 2397
rect 27264 2400 28264 2428
rect 27264 2360 27292 2400
rect 28258 2388 28264 2400
rect 28316 2388 28322 2440
rect 32858 2388 32864 2440
rect 32916 2428 32922 2440
rect 32953 2431 33011 2437
rect 32953 2428 32965 2431
rect 32916 2400 32965 2428
rect 32916 2388 32922 2400
rect 32953 2397 32965 2400
rect 32999 2397 33011 2431
rect 36449 2431 36507 2437
rect 36449 2428 36461 2431
rect 32953 2391 33011 2397
rect 33060 2400 36461 2428
rect 26206 2332 27292 2360
rect 26053 2323 26111 2329
rect 9171 2295 9229 2301
rect 9171 2261 9183 2295
rect 9217 2292 9229 2295
rect 15194 2292 15200 2304
rect 9217 2264 15200 2292
rect 9217 2261 9229 2264
rect 9171 2255 9229 2261
rect 15194 2252 15200 2264
rect 15252 2252 15258 2304
rect 17678 2292 17684 2304
rect 17639 2264 17684 2292
rect 17678 2252 17684 2264
rect 17736 2252 17742 2304
rect 24486 2252 24492 2304
rect 24544 2292 24550 2304
rect 26068 2292 26096 2323
rect 27706 2320 27712 2372
rect 27764 2360 27770 2372
rect 27985 2363 28043 2369
rect 27985 2360 27997 2363
rect 27764 2332 27997 2360
rect 27764 2320 27770 2332
rect 27985 2329 27997 2332
rect 28031 2329 28043 2363
rect 27985 2323 28043 2329
rect 28442 2320 28448 2372
rect 28500 2360 28506 2372
rect 33060 2360 33088 2400
rect 36449 2397 36461 2400
rect 36495 2397 36507 2431
rect 36449 2391 36507 2397
rect 38473 2431 38531 2437
rect 38473 2397 38485 2431
rect 38519 2428 38531 2431
rect 38654 2428 38660 2440
rect 38519 2400 38660 2428
rect 38519 2397 38531 2400
rect 38473 2391 38531 2397
rect 38654 2388 38660 2400
rect 38712 2388 38718 2440
rect 38746 2388 38752 2440
rect 38804 2428 38810 2440
rect 38804 2400 38849 2428
rect 38804 2388 38810 2400
rect 28500 2332 33088 2360
rect 33965 2363 34023 2369
rect 28500 2320 28506 2332
rect 33965 2329 33977 2363
rect 34011 2360 34023 2363
rect 34146 2360 34152 2372
rect 34011 2332 34152 2360
rect 34011 2329 34023 2332
rect 33965 2323 34023 2329
rect 34146 2320 34152 2332
rect 34204 2320 34210 2372
rect 34790 2320 34796 2372
rect 34848 2360 34854 2372
rect 35161 2363 35219 2369
rect 35161 2360 35173 2363
rect 34848 2332 35173 2360
rect 34848 2320 34854 2332
rect 35161 2329 35173 2332
rect 35207 2329 35219 2363
rect 35161 2323 35219 2329
rect 36078 2320 36084 2372
rect 36136 2360 36142 2372
rect 36265 2363 36323 2369
rect 36265 2360 36277 2363
rect 36136 2332 36277 2360
rect 36136 2320 36142 2332
rect 36265 2329 36277 2332
rect 36311 2329 36323 2363
rect 47762 2360 47768 2372
rect 47723 2332 47768 2360
rect 36265 2323 36323 2329
rect 47762 2320 47768 2332
rect 47820 2320 47826 2372
rect 24544 2264 26096 2292
rect 24544 2252 24550 2264
rect 26142 2252 26148 2304
rect 26200 2292 26206 2304
rect 33137 2295 33195 2301
rect 33137 2292 33149 2295
rect 26200 2264 33149 2292
rect 26200 2252 26206 2264
rect 33137 2261 33149 2264
rect 33183 2261 33195 2295
rect 47854 2292 47860 2304
rect 47815 2264 47860 2292
rect 33137 2255 33195 2261
rect 47854 2252 47860 2264
rect 47912 2252 47918 2304
rect 1104 2202 48852 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 48852 2202
rect 1104 2128 48852 2150
rect 24302 1980 24308 2032
rect 24360 2020 24366 2032
rect 47854 2020 47860 2032
rect 24360 1992 47860 2020
rect 24360 1980 24366 1992
rect 47854 1980 47860 1992
rect 47912 1980 47918 2032
rect 22278 1912 22284 1964
rect 22336 1952 22342 1964
rect 38746 1952 38752 1964
rect 22336 1924 38752 1952
rect 22336 1912 22342 1924
rect 38746 1912 38752 1924
rect 38804 1912 38810 1964
rect 17678 1844 17684 1896
rect 17736 1884 17742 1896
rect 31662 1884 31668 1896
rect 17736 1856 31668 1884
rect 17736 1844 17742 1856
rect 31662 1844 31668 1856
rect 31720 1844 31726 1896
<< via1 >>
rect 41420 50192 41472 50244
rect 46848 50192 46900 50244
rect 3424 49716 3476 49768
rect 9220 49716 9272 49768
rect 21272 49716 21324 49768
rect 46756 49716 46808 49768
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 3976 49240 4028 49292
rect 4068 49240 4120 49292
rect 8668 49240 8720 49292
rect 12716 49283 12768 49292
rect 12716 49249 12725 49283
rect 12725 49249 12759 49283
rect 12759 49249 12768 49283
rect 12716 49240 12768 49249
rect 13820 49240 13872 49292
rect 18052 49240 18104 49292
rect 20444 49240 20496 49292
rect 664 49172 716 49224
rect 3240 49172 3292 49224
rect 6460 49172 6512 49224
rect 9864 49215 9916 49224
rect 5448 49104 5500 49156
rect 6644 49104 6696 49156
rect 9864 49181 9873 49215
rect 9873 49181 9907 49215
rect 9907 49181 9916 49215
rect 9864 49172 9916 49181
rect 11612 49172 11664 49224
rect 12992 49215 13044 49224
rect 12992 49181 13001 49215
rect 13001 49181 13035 49215
rect 13035 49181 13044 49215
rect 12992 49172 13044 49181
rect 14372 49215 14424 49224
rect 14372 49181 14381 49215
rect 14381 49181 14415 49215
rect 14415 49181 14424 49215
rect 14372 49172 14424 49181
rect 16580 49172 16632 49224
rect 16672 49172 16724 49224
rect 19340 49215 19392 49224
rect 19340 49181 19349 49215
rect 19349 49181 19383 49215
rect 19383 49181 19392 49215
rect 19340 49172 19392 49181
rect 19984 49172 20036 49224
rect 23848 49308 23900 49360
rect 40040 49308 40092 49360
rect 22560 49283 22612 49292
rect 22560 49249 22569 49283
rect 22569 49249 22603 49283
rect 22603 49249 22612 49283
rect 22560 49240 22612 49249
rect 24768 49240 24820 49292
rect 27620 49283 27672 49292
rect 27620 49249 27629 49283
rect 27629 49249 27663 49283
rect 27663 49249 27672 49283
rect 27620 49240 27672 49249
rect 30564 49240 30616 49292
rect 30932 49283 30984 49292
rect 30932 49249 30941 49283
rect 30941 49249 30975 49283
rect 30975 49249 30984 49283
rect 30932 49240 30984 49249
rect 22008 49215 22060 49224
rect 22008 49181 22017 49215
rect 22017 49181 22051 49215
rect 22051 49181 22060 49215
rect 22008 49172 22060 49181
rect 24400 49215 24452 49224
rect 24400 49181 24409 49215
rect 24409 49181 24443 49215
rect 24443 49181 24452 49215
rect 24400 49172 24452 49181
rect 26976 49215 27028 49224
rect 26976 49181 26985 49215
rect 26985 49181 27019 49215
rect 27019 49181 27028 49215
rect 26976 49172 27028 49181
rect 31944 49172 31996 49224
rect 34888 49172 34940 49224
rect 38108 49215 38160 49224
rect 38108 49181 38117 49215
rect 38117 49181 38151 49215
rect 38151 49181 38160 49215
rect 38108 49172 38160 49181
rect 40592 49240 40644 49292
rect 46664 49240 46716 49292
rect 46848 49283 46900 49292
rect 46848 49249 46857 49283
rect 46857 49249 46891 49283
rect 46891 49249 46900 49283
rect 46848 49240 46900 49249
rect 39764 49172 39816 49224
rect 41972 49172 42024 49224
rect 44088 49172 44140 49224
rect 48964 49172 49016 49224
rect 12164 49147 12216 49156
rect 12164 49113 12173 49147
rect 12173 49113 12207 49147
rect 12207 49113 12216 49147
rect 12164 49104 12216 49113
rect 22192 49147 22244 49156
rect 22192 49113 22201 49147
rect 22201 49113 22235 49147
rect 22235 49113 22244 49147
rect 22192 49104 22244 49113
rect 24584 49147 24636 49156
rect 24584 49113 24593 49147
rect 24593 49113 24627 49147
rect 24627 49113 24636 49147
rect 24584 49104 24636 49113
rect 27160 49147 27212 49156
rect 27160 49113 27169 49147
rect 27169 49113 27203 49147
rect 27203 49113 27212 49147
rect 27160 49104 27212 49113
rect 29920 49147 29972 49156
rect 29920 49113 29929 49147
rect 29929 49113 29963 49147
rect 29963 49113 29972 49147
rect 29920 49104 29972 49113
rect 40040 49147 40092 49156
rect 40040 49113 40049 49147
rect 40049 49113 40083 49147
rect 40083 49113 40092 49147
rect 40040 49104 40092 49113
rect 43720 49104 43772 49156
rect 45376 49147 45428 49156
rect 45376 49113 45385 49147
rect 45385 49113 45419 49147
rect 45419 49113 45428 49147
rect 45376 49104 45428 49113
rect 1676 49036 1728 49088
rect 3148 49079 3200 49088
rect 3148 49045 3157 49079
rect 3157 49045 3191 49079
rect 3191 49045 3200 49079
rect 3148 49036 3200 49045
rect 6920 49079 6972 49088
rect 6920 49045 6929 49079
rect 6929 49045 6963 49079
rect 6963 49045 6972 49079
rect 6920 49036 6972 49045
rect 8944 49036 8996 49088
rect 20168 49036 20220 49088
rect 20352 49036 20404 49088
rect 23480 49036 23532 49088
rect 32128 49079 32180 49088
rect 32128 49045 32137 49079
rect 32137 49045 32171 49079
rect 32171 49045 32180 49079
rect 32128 49036 32180 49045
rect 38292 49079 38344 49088
rect 38292 49045 38301 49079
rect 38301 49045 38335 49079
rect 38335 49045 38344 49079
rect 38292 49036 38344 49045
rect 39212 49079 39264 49088
rect 39212 49045 39221 49079
rect 39221 49045 39255 49079
rect 39255 49045 39264 49079
rect 39212 49036 39264 49045
rect 47952 49036 48004 49088
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 20168 48832 20220 48884
rect 26792 48832 26844 48884
rect 2872 48764 2924 48816
rect 14372 48764 14424 48816
rect 22928 48764 22980 48816
rect 25780 48764 25832 48816
rect 26424 48764 26476 48816
rect 29000 48764 29052 48816
rect 38752 48764 38804 48816
rect 41420 48764 41472 48816
rect 41880 48764 41932 48816
rect 47768 48807 47820 48816
rect 47768 48773 47777 48807
rect 47777 48773 47811 48807
rect 47811 48773 47820 48807
rect 47768 48764 47820 48773
rect 6644 48739 6696 48748
rect 6644 48705 6653 48739
rect 6653 48705 6687 48739
rect 6687 48705 6696 48739
rect 6644 48696 6696 48705
rect 8944 48739 8996 48748
rect 8944 48705 8953 48739
rect 8953 48705 8987 48739
rect 8987 48705 8996 48739
rect 8944 48696 8996 48705
rect 14004 48739 14056 48748
rect 14004 48705 14013 48739
rect 14013 48705 14047 48739
rect 14047 48705 14056 48739
rect 14004 48696 14056 48705
rect 16120 48696 16172 48748
rect 16672 48739 16724 48748
rect 16672 48705 16681 48739
rect 16681 48705 16715 48739
rect 16715 48705 16724 48739
rect 16672 48696 16724 48705
rect 22008 48696 22060 48748
rect 32128 48739 32180 48748
rect 32128 48705 32137 48739
rect 32137 48705 32171 48739
rect 32171 48705 32180 48739
rect 32128 48696 32180 48705
rect 34888 48739 34940 48748
rect 34888 48705 34897 48739
rect 34897 48705 34931 48739
rect 34931 48705 34940 48739
rect 34888 48696 34940 48705
rect 3056 48628 3108 48680
rect 3792 48671 3844 48680
rect 3792 48637 3801 48671
rect 3801 48637 3835 48671
rect 3835 48637 3844 48671
rect 3792 48628 3844 48637
rect 4068 48628 4120 48680
rect 4712 48671 4764 48680
rect 4712 48637 4721 48671
rect 4721 48637 4755 48671
rect 4755 48637 4764 48671
rect 4712 48628 4764 48637
rect 7748 48628 7800 48680
rect 9128 48671 9180 48680
rect 3884 48560 3936 48612
rect 7104 48560 7156 48612
rect 9128 48637 9137 48671
rect 9137 48637 9171 48671
rect 9171 48637 9180 48671
rect 9128 48628 9180 48637
rect 9680 48671 9732 48680
rect 9680 48637 9689 48671
rect 9689 48637 9723 48671
rect 9723 48637 9732 48671
rect 9680 48628 9732 48637
rect 11520 48671 11572 48680
rect 11520 48637 11529 48671
rect 11529 48637 11563 48671
rect 11563 48637 11572 48671
rect 11520 48628 11572 48637
rect 11704 48671 11756 48680
rect 11704 48637 11713 48671
rect 11713 48637 11747 48671
rect 11747 48637 11756 48671
rect 11704 48628 11756 48637
rect 12440 48671 12492 48680
rect 12440 48637 12449 48671
rect 12449 48637 12483 48671
rect 12483 48637 12492 48671
rect 12440 48628 12492 48637
rect 16856 48671 16908 48680
rect 16856 48637 16865 48671
rect 16865 48637 16899 48671
rect 16899 48637 16908 48671
rect 16856 48628 16908 48637
rect 16948 48628 17000 48680
rect 23664 48628 23716 48680
rect 18604 48560 18656 48612
rect 20812 48560 20864 48612
rect 23204 48560 23256 48612
rect 29368 48671 29420 48680
rect 29368 48637 29377 48671
rect 29377 48637 29411 48671
rect 29411 48637 29420 48671
rect 29644 48671 29696 48680
rect 29368 48628 29420 48637
rect 29644 48637 29653 48671
rect 29653 48637 29687 48671
rect 29687 48637 29696 48671
rect 29644 48628 29696 48637
rect 32312 48671 32364 48680
rect 32312 48637 32321 48671
rect 32321 48637 32355 48671
rect 32355 48637 32364 48671
rect 32312 48628 32364 48637
rect 32864 48671 32916 48680
rect 32864 48637 32873 48671
rect 32873 48637 32907 48671
rect 32907 48637 32916 48671
rect 32864 48628 32916 48637
rect 36084 48671 36136 48680
rect 27620 48603 27672 48612
rect 27620 48569 27629 48603
rect 27629 48569 27663 48603
rect 27663 48569 27672 48603
rect 27620 48560 27672 48569
rect 29276 48560 29328 48612
rect 36084 48637 36093 48671
rect 36093 48637 36127 48671
rect 36127 48637 36136 48671
rect 36084 48628 36136 48637
rect 42800 48671 42852 48680
rect 36176 48560 36228 48612
rect 42800 48637 42809 48671
rect 42809 48637 42843 48671
rect 42843 48637 42852 48671
rect 42800 48628 42852 48637
rect 43168 48671 43220 48680
rect 43168 48637 43177 48671
rect 43177 48637 43211 48671
rect 43211 48637 43220 48671
rect 43168 48628 43220 48637
rect 44916 48671 44968 48680
rect 44916 48637 44925 48671
rect 44925 48637 44959 48671
rect 44959 48637 44968 48671
rect 44916 48628 44968 48637
rect 45100 48671 45152 48680
rect 45100 48637 45109 48671
rect 45109 48637 45143 48671
rect 45143 48637 45152 48671
rect 45100 48628 45152 48637
rect 45744 48671 45796 48680
rect 45744 48637 45753 48671
rect 45753 48637 45787 48671
rect 45787 48637 45796 48671
rect 45744 48628 45796 48637
rect 42984 48560 43036 48612
rect 20260 48535 20312 48544
rect 20260 48501 20269 48535
rect 20269 48501 20303 48535
rect 20303 48501 20312 48535
rect 20260 48492 20312 48501
rect 25412 48535 25464 48544
rect 25412 48501 25421 48535
rect 25421 48501 25455 48535
rect 25455 48501 25464 48535
rect 25412 48492 25464 48501
rect 25504 48492 25556 48544
rect 28448 48492 28500 48544
rect 33784 48492 33836 48544
rect 34152 48492 34204 48544
rect 37464 48535 37516 48544
rect 37464 48501 37473 48535
rect 37473 48501 37507 48535
rect 37507 48501 37516 48535
rect 37464 48492 37516 48501
rect 41604 48535 41656 48544
rect 41604 48501 41613 48535
rect 41613 48501 41647 48535
rect 41647 48501 41656 48535
rect 41604 48492 41656 48501
rect 48228 48492 48280 48544
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 9128 48331 9180 48340
rect 9128 48297 9137 48331
rect 9137 48297 9171 48331
rect 9171 48297 9180 48331
rect 9128 48288 9180 48297
rect 11704 48288 11756 48340
rect 29920 48288 29972 48340
rect 38752 48331 38804 48340
rect 38752 48297 38761 48331
rect 38761 48297 38795 48331
rect 38795 48297 38804 48331
rect 38752 48288 38804 48297
rect 20 48220 72 48272
rect 7748 48263 7800 48272
rect 1308 48152 1360 48204
rect 7748 48229 7757 48263
rect 7757 48229 7791 48263
rect 7791 48229 7800 48263
rect 7748 48220 7800 48229
rect 17132 48220 17184 48272
rect 23664 48263 23716 48272
rect 5172 48152 5224 48204
rect 9864 48152 9916 48204
rect 10324 48195 10376 48204
rect 10324 48161 10333 48195
rect 10333 48161 10367 48195
rect 10367 48161 10376 48195
rect 10324 48152 10376 48161
rect 14924 48195 14976 48204
rect 14924 48161 14933 48195
rect 14933 48161 14967 48195
rect 14967 48161 14976 48195
rect 14924 48152 14976 48161
rect 16580 48152 16632 48204
rect 17408 48195 17460 48204
rect 17408 48161 17417 48195
rect 17417 48161 17451 48195
rect 17451 48161 17460 48195
rect 17408 48152 17460 48161
rect 20260 48152 20312 48204
rect 20628 48152 20680 48204
rect 5356 48127 5408 48136
rect 5356 48093 5365 48127
rect 5365 48093 5399 48127
rect 5399 48093 5408 48127
rect 5356 48084 5408 48093
rect 7104 48084 7156 48136
rect 8944 48084 8996 48136
rect 9128 48084 9180 48136
rect 11980 48127 12032 48136
rect 11980 48093 11989 48127
rect 11989 48093 12023 48127
rect 12023 48093 12032 48127
rect 11980 48084 12032 48093
rect 14464 48127 14516 48136
rect 14464 48093 14473 48127
rect 14473 48093 14507 48127
rect 14507 48093 14516 48127
rect 14464 48084 14516 48093
rect 1584 48059 1636 48068
rect 1584 48025 1593 48059
rect 1593 48025 1627 48059
rect 1627 48025 1636 48059
rect 1584 48016 1636 48025
rect 4436 48059 4488 48068
rect 4436 48025 4445 48059
rect 4445 48025 4479 48059
rect 4479 48025 4488 48059
rect 4436 48016 4488 48025
rect 5540 48059 5592 48068
rect 5540 48025 5549 48059
rect 5549 48025 5583 48059
rect 5583 48025 5592 48059
rect 5540 48016 5592 48025
rect 9956 48016 10008 48068
rect 14372 48016 14424 48068
rect 17408 48016 17460 48068
rect 20168 48059 20220 48068
rect 20168 48025 20177 48059
rect 20177 48025 20211 48059
rect 20211 48025 20220 48059
rect 20168 48016 20220 48025
rect 4712 47948 4764 48000
rect 7380 47948 7432 48000
rect 21916 48084 21968 48136
rect 21640 47948 21692 48000
rect 23664 48229 23673 48263
rect 23673 48229 23707 48263
rect 23707 48229 23716 48263
rect 23664 48220 23716 48229
rect 25320 48220 25372 48272
rect 25412 48152 25464 48204
rect 29368 48220 29420 48272
rect 32312 48220 32364 48272
rect 36728 48220 36780 48272
rect 27712 48152 27764 48204
rect 31944 48152 31996 48204
rect 32220 48195 32272 48204
rect 32220 48161 32229 48195
rect 32229 48161 32263 48195
rect 32263 48161 32272 48195
rect 32220 48152 32272 48161
rect 37464 48152 37516 48204
rect 40040 48220 40092 48272
rect 47032 48220 47084 48272
rect 49608 48220 49660 48272
rect 42524 48195 42576 48204
rect 42524 48161 42533 48195
rect 42533 48161 42567 48195
rect 42567 48161 42576 48195
rect 42524 48152 42576 48161
rect 48320 48152 48372 48204
rect 23848 48084 23900 48136
rect 24952 48059 25004 48068
rect 24952 48025 24961 48059
rect 24961 48025 24995 48059
rect 24995 48025 25004 48059
rect 24952 48016 25004 48025
rect 25228 47991 25280 48000
rect 25228 47957 25237 47991
rect 25237 47957 25271 47991
rect 25271 47957 25280 47991
rect 25228 47948 25280 47957
rect 28080 48084 28132 48136
rect 30104 48127 30156 48136
rect 28172 48016 28224 48068
rect 30104 48093 30113 48127
rect 30113 48093 30147 48127
rect 30147 48093 30156 48127
rect 30104 48084 30156 48093
rect 30748 48127 30800 48136
rect 30748 48093 30757 48127
rect 30757 48093 30791 48127
rect 30791 48093 30800 48127
rect 30748 48084 30800 48093
rect 33784 48084 33836 48136
rect 35716 48127 35768 48136
rect 35716 48093 35725 48127
rect 35725 48093 35759 48127
rect 35759 48093 35768 48127
rect 35716 48084 35768 48093
rect 38660 48127 38712 48136
rect 38660 48093 38669 48127
rect 38669 48093 38703 48127
rect 38703 48093 38712 48127
rect 38660 48084 38712 48093
rect 39856 48127 39908 48136
rect 39856 48093 39865 48127
rect 39865 48093 39899 48127
rect 39899 48093 39908 48127
rect 39856 48084 39908 48093
rect 41052 48127 41104 48136
rect 41052 48093 41061 48127
rect 41061 48093 41095 48127
rect 41095 48093 41104 48127
rect 41052 48084 41104 48093
rect 43904 48127 43956 48136
rect 43904 48093 43913 48127
rect 43913 48093 43947 48127
rect 43947 48093 43956 48127
rect 43904 48084 43956 48093
rect 44456 48084 44508 48136
rect 32220 48016 32272 48068
rect 40408 48016 40460 48068
rect 43812 48016 43864 48068
rect 47676 48016 47728 48068
rect 32128 47948 32180 48000
rect 43996 47948 44048 48000
rect 45192 47991 45244 48000
rect 45192 47957 45201 47991
rect 45201 47957 45235 47991
rect 45235 47957 45244 47991
rect 45192 47948 45244 47957
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 1584 47744 1636 47796
rect 3056 47787 3108 47796
rect 3056 47753 3065 47787
rect 3065 47753 3099 47787
rect 3099 47753 3108 47787
rect 3056 47744 3108 47753
rect 5448 47787 5500 47796
rect 5448 47753 5457 47787
rect 5457 47753 5491 47787
rect 5491 47753 5500 47787
rect 5448 47744 5500 47753
rect 7472 47744 7524 47796
rect 8668 47744 8720 47796
rect 9956 47787 10008 47796
rect 9956 47753 9965 47787
rect 9965 47753 9999 47787
rect 9999 47753 10008 47787
rect 9956 47744 10008 47753
rect 16856 47744 16908 47796
rect 17408 47787 17460 47796
rect 17408 47753 17417 47787
rect 17417 47753 17451 47787
rect 17451 47753 17460 47787
rect 17408 47744 17460 47753
rect 20168 47744 20220 47796
rect 22192 47744 22244 47796
rect 24584 47744 24636 47796
rect 24768 47744 24820 47796
rect 30748 47744 30800 47796
rect 32220 47787 32272 47796
rect 32220 47753 32229 47787
rect 32229 47753 32263 47787
rect 32263 47753 32272 47787
rect 32220 47744 32272 47753
rect 36176 47787 36228 47796
rect 2136 47719 2188 47728
rect 2136 47685 2145 47719
rect 2145 47685 2179 47719
rect 2179 47685 2188 47719
rect 2136 47676 2188 47685
rect 3332 47676 3384 47728
rect 3516 47608 3568 47660
rect 3792 47608 3844 47660
rect 4620 47651 4672 47660
rect 4620 47617 4629 47651
rect 4629 47617 4663 47651
rect 4663 47617 4672 47651
rect 4620 47608 4672 47617
rect 7380 47608 7432 47660
rect 8944 47608 8996 47660
rect 11520 47608 11572 47660
rect 14464 47608 14516 47660
rect 16672 47651 16724 47660
rect 16672 47617 16681 47651
rect 16681 47617 16715 47651
rect 16715 47617 16724 47651
rect 16672 47608 16724 47617
rect 17316 47651 17368 47660
rect 17316 47617 17325 47651
rect 17325 47617 17359 47651
rect 17359 47617 17368 47651
rect 17316 47608 17368 47617
rect 20076 47608 20128 47660
rect 2504 47540 2556 47592
rect 7472 47583 7524 47592
rect 4436 47472 4488 47524
rect 5448 47472 5500 47524
rect 7472 47549 7481 47583
rect 7481 47549 7515 47583
rect 7515 47549 7524 47583
rect 7472 47540 7524 47549
rect 9036 47540 9088 47592
rect 9220 47583 9272 47592
rect 9220 47549 9229 47583
rect 9229 47549 9263 47583
rect 9263 47549 9272 47583
rect 9220 47540 9272 47549
rect 11980 47540 12032 47592
rect 17132 47540 17184 47592
rect 17224 47472 17276 47524
rect 24952 47676 25004 47728
rect 24216 47608 24268 47660
rect 25228 47651 25280 47660
rect 25228 47617 25237 47651
rect 25237 47617 25271 47651
rect 25271 47617 25280 47651
rect 25228 47608 25280 47617
rect 22008 47583 22060 47592
rect 22008 47549 22017 47583
rect 22017 47549 22051 47583
rect 22051 47549 22060 47583
rect 22008 47540 22060 47549
rect 25136 47540 25188 47592
rect 26700 47540 26752 47592
rect 26884 47608 26936 47660
rect 27160 47608 27212 47660
rect 28080 47651 28132 47660
rect 28080 47617 28089 47651
rect 28089 47617 28123 47651
rect 28123 47617 28132 47651
rect 28080 47608 28132 47617
rect 27528 47540 27580 47592
rect 28540 47540 28592 47592
rect 1952 47404 2004 47456
rect 4804 47447 4856 47456
rect 4804 47413 4813 47447
rect 4813 47413 4847 47447
rect 4847 47413 4856 47447
rect 4804 47404 4856 47413
rect 25412 47472 25464 47524
rect 28356 47472 28408 47524
rect 24308 47404 24360 47456
rect 29552 47540 29604 47592
rect 30104 47676 30156 47728
rect 36176 47753 36185 47787
rect 36185 47753 36219 47787
rect 36219 47753 36228 47787
rect 36176 47744 36228 47753
rect 40408 47787 40460 47796
rect 40408 47753 40417 47787
rect 40417 47753 40451 47787
rect 40451 47753 40460 47787
rect 40408 47744 40460 47753
rect 42800 47744 42852 47796
rect 45376 47744 45428 47796
rect 46664 47719 46716 47728
rect 46664 47685 46673 47719
rect 46673 47685 46707 47719
rect 46707 47685 46716 47719
rect 46664 47676 46716 47685
rect 47860 47676 47912 47728
rect 30564 47651 30616 47660
rect 30564 47617 30573 47651
rect 30573 47617 30607 47651
rect 30607 47617 30616 47651
rect 30564 47608 30616 47617
rect 31852 47608 31904 47660
rect 32128 47651 32180 47660
rect 32128 47617 32137 47651
rect 32137 47617 32171 47651
rect 32171 47617 32180 47651
rect 32128 47608 32180 47617
rect 33140 47651 33192 47660
rect 33140 47617 33149 47651
rect 33149 47617 33183 47651
rect 33183 47617 33192 47651
rect 33140 47608 33192 47617
rect 33784 47651 33836 47660
rect 33784 47617 33793 47651
rect 33793 47617 33827 47651
rect 33827 47617 33836 47651
rect 33784 47608 33836 47617
rect 36084 47651 36136 47660
rect 36084 47617 36093 47651
rect 36093 47617 36127 47651
rect 36127 47617 36136 47651
rect 36084 47608 36136 47617
rect 39764 47651 39816 47660
rect 39764 47617 39773 47651
rect 39773 47617 39807 47651
rect 39807 47617 39816 47651
rect 39764 47608 39816 47617
rect 40316 47651 40368 47660
rect 40316 47617 40325 47651
rect 40325 47617 40359 47651
rect 40359 47617 40368 47651
rect 40316 47608 40368 47617
rect 41052 47608 41104 47660
rect 41972 47608 42024 47660
rect 43536 47651 43588 47660
rect 34796 47583 34848 47592
rect 34796 47549 34805 47583
rect 34805 47549 34839 47583
rect 34839 47549 34848 47583
rect 34796 47540 34848 47549
rect 43536 47617 43545 47651
rect 43545 47617 43579 47651
rect 43579 47617 43588 47651
rect 43536 47608 43588 47617
rect 44180 47583 44232 47592
rect 44180 47549 44189 47583
rect 44189 47549 44223 47583
rect 44223 47549 44232 47583
rect 44180 47540 44232 47549
rect 44364 47583 44416 47592
rect 44364 47549 44373 47583
rect 44373 47549 44407 47583
rect 44407 47549 44416 47583
rect 44364 47540 44416 47549
rect 45008 47583 45060 47592
rect 45008 47549 45017 47583
rect 45017 47549 45051 47583
rect 45051 47549 45060 47583
rect 45008 47540 45060 47549
rect 47584 47472 47636 47524
rect 47124 47404 47176 47456
rect 47768 47404 47820 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 3976 47243 4028 47252
rect 3976 47209 3985 47243
rect 3985 47209 4019 47243
rect 4019 47209 4028 47243
rect 3976 47200 4028 47209
rect 5540 47243 5592 47252
rect 5540 47209 5549 47243
rect 5549 47209 5583 47243
rect 5583 47209 5592 47243
rect 5540 47200 5592 47209
rect 9036 47243 9088 47252
rect 9036 47209 9045 47243
rect 9045 47209 9079 47243
rect 9079 47209 9088 47243
rect 9036 47200 9088 47209
rect 14372 47243 14424 47252
rect 14372 47209 14381 47243
rect 14381 47209 14415 47243
rect 14415 47209 14424 47243
rect 14372 47200 14424 47209
rect 16672 47200 16724 47252
rect 24308 47200 24360 47252
rect 24400 47200 24452 47252
rect 24860 47200 24912 47252
rect 26148 47200 26200 47252
rect 26700 47200 26752 47252
rect 36084 47200 36136 47252
rect 37188 47200 37240 47252
rect 42984 47243 43036 47252
rect 42984 47209 42993 47243
rect 42993 47209 43027 47243
rect 43027 47209 43036 47243
rect 42984 47200 43036 47209
rect 43812 47243 43864 47252
rect 43812 47209 43821 47243
rect 43821 47209 43855 47243
rect 43855 47209 43864 47243
rect 43812 47200 43864 47209
rect 44364 47243 44416 47252
rect 44364 47209 44373 47243
rect 44373 47209 44407 47243
rect 44407 47209 44416 47243
rect 44364 47200 44416 47209
rect 45100 47200 45152 47252
rect 3608 47132 3660 47184
rect 3884 47132 3936 47184
rect 17316 47132 17368 47184
rect 1860 47107 1912 47116
rect 1860 47073 1869 47107
rect 1869 47073 1903 47107
rect 1903 47073 1912 47107
rect 1860 47064 1912 47073
rect 9128 47064 9180 47116
rect 24768 47064 24820 47116
rect 4896 46996 4948 47048
rect 9404 46996 9456 47048
rect 14280 47039 14332 47048
rect 14280 47005 14289 47039
rect 14289 47005 14323 47039
rect 14323 47005 14332 47039
rect 14280 46996 14332 47005
rect 21732 46996 21784 47048
rect 1584 46971 1636 46980
rect 1584 46937 1593 46971
rect 1593 46937 1627 46971
rect 1627 46937 1636 46971
rect 1584 46928 1636 46937
rect 15476 46928 15528 46980
rect 16580 46928 16632 46980
rect 17224 46928 17276 46980
rect 24860 46996 24912 47048
rect 22008 46928 22060 46980
rect 33140 47064 33192 47116
rect 33692 47064 33744 47116
rect 25228 46996 25280 47048
rect 27528 46996 27580 47048
rect 21916 46903 21968 46912
rect 21916 46869 21925 46903
rect 21925 46869 21959 46903
rect 21959 46869 21968 46903
rect 21916 46860 21968 46869
rect 28264 46996 28316 47048
rect 28540 47039 28592 47048
rect 28540 47005 28549 47039
rect 28549 47005 28583 47039
rect 28583 47005 28592 47039
rect 28540 46996 28592 47005
rect 45560 46996 45612 47048
rect 46296 47039 46348 47048
rect 46296 47005 46305 47039
rect 46305 47005 46339 47039
rect 46339 47005 46348 47039
rect 46296 46996 46348 47005
rect 48136 47039 48188 47048
rect 48136 47005 48145 47039
rect 48145 47005 48179 47039
rect 48179 47005 48188 47039
rect 48136 46996 48188 47005
rect 44548 46928 44600 46980
rect 46480 46971 46532 46980
rect 46480 46937 46489 46971
rect 46489 46937 46523 46971
rect 46523 46937 46532 46971
rect 46480 46928 46532 46937
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 1584 46656 1636 46708
rect 43720 46656 43772 46708
rect 47676 46699 47728 46708
rect 47676 46665 47685 46699
rect 47685 46665 47719 46699
rect 47719 46665 47728 46699
rect 47676 46656 47728 46665
rect 21272 46631 21324 46640
rect 21272 46597 21281 46631
rect 21281 46597 21315 46631
rect 21315 46597 21324 46631
rect 21272 46588 21324 46597
rect 25228 46588 25280 46640
rect 47032 46631 47084 46640
rect 47032 46597 47041 46631
rect 47041 46597 47075 46631
rect 47075 46597 47084 46631
rect 47032 46588 47084 46597
rect 1400 46563 1452 46572
rect 1400 46529 1409 46563
rect 1409 46529 1443 46563
rect 1443 46529 1452 46563
rect 1400 46520 1452 46529
rect 2136 46563 2188 46572
rect 2136 46529 2145 46563
rect 2145 46529 2179 46563
rect 2179 46529 2188 46563
rect 2136 46520 2188 46529
rect 3608 46563 3660 46572
rect 3608 46529 3617 46563
rect 3617 46529 3651 46563
rect 3651 46529 3660 46563
rect 3608 46520 3660 46529
rect 4712 46520 4764 46572
rect 26976 46520 27028 46572
rect 44088 46563 44140 46572
rect 44088 46529 44097 46563
rect 44097 46529 44131 46563
rect 44131 46529 44140 46563
rect 44088 46520 44140 46529
rect 44548 46563 44600 46572
rect 44548 46529 44557 46563
rect 44557 46529 44591 46563
rect 44591 46529 44600 46563
rect 44548 46520 44600 46529
rect 47584 46563 47636 46572
rect 47584 46529 47593 46563
rect 47593 46529 47627 46563
rect 47627 46529 47636 46563
rect 47584 46520 47636 46529
rect 3056 46452 3108 46504
rect 14280 46452 14332 46504
rect 19340 46452 19392 46504
rect 19708 46452 19760 46504
rect 45192 46495 45244 46504
rect 45192 46461 45201 46495
rect 45201 46461 45235 46495
rect 45235 46461 45244 46495
rect 45192 46452 45244 46461
rect 46112 46452 46164 46504
rect 4896 46384 4948 46436
rect 1584 46359 1636 46368
rect 1584 46325 1593 46359
rect 1593 46325 1627 46359
rect 1627 46325 1636 46359
rect 1584 46316 1636 46325
rect 2872 46359 2924 46368
rect 2872 46325 2881 46359
rect 2881 46325 2915 46359
rect 2915 46325 2924 46359
rect 2872 46316 2924 46325
rect 7932 46316 7984 46368
rect 28080 46316 28132 46368
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 19708 46155 19760 46164
rect 19708 46121 19717 46155
rect 19717 46121 19751 46155
rect 19751 46121 19760 46155
rect 19708 46112 19760 46121
rect 44180 46112 44232 46164
rect 44916 46112 44968 46164
rect 2872 45976 2924 46028
rect 2964 46019 3016 46028
rect 2964 45985 2973 46019
rect 2973 45985 3007 46019
rect 3007 45985 3016 46019
rect 25412 46019 25464 46028
rect 2964 45976 3016 45985
rect 25412 45985 25421 46019
rect 25421 45985 25455 46019
rect 25455 45985 25464 46019
rect 25412 45976 25464 45985
rect 48136 46019 48188 46028
rect 48136 45985 48145 46019
rect 48145 45985 48179 46019
rect 48179 45985 48188 46019
rect 48136 45976 48188 45985
rect 20076 45908 20128 45960
rect 25228 45951 25280 45960
rect 25228 45917 25237 45951
rect 25237 45917 25271 45951
rect 25271 45917 25280 45951
rect 25228 45908 25280 45917
rect 45652 45951 45704 45960
rect 45652 45917 45661 45951
rect 45661 45917 45695 45951
rect 45695 45917 45704 45951
rect 45652 45908 45704 45917
rect 45836 45908 45888 45960
rect 2872 45840 2924 45892
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 1860 45543 1912 45552
rect 1860 45509 1869 45543
rect 1869 45509 1903 45543
rect 1903 45509 1912 45543
rect 1860 45500 1912 45509
rect 2872 45475 2924 45484
rect 2872 45441 2881 45475
rect 2881 45441 2915 45475
rect 2915 45441 2924 45475
rect 2872 45432 2924 45441
rect 7932 45475 7984 45484
rect 7932 45441 7941 45475
rect 7941 45441 7975 45475
rect 7975 45441 7984 45475
rect 7932 45432 7984 45441
rect 23756 45475 23808 45484
rect 23756 45441 23765 45475
rect 23765 45441 23799 45475
rect 23799 45441 23808 45475
rect 23756 45432 23808 45441
rect 26148 45432 26200 45484
rect 45192 45432 45244 45484
rect 45836 45432 45888 45484
rect 46112 45500 46164 45552
rect 46480 45500 46532 45552
rect 46204 45475 46256 45484
rect 46204 45441 46213 45475
rect 46213 45441 46247 45475
rect 46247 45441 46256 45475
rect 46204 45432 46256 45441
rect 47584 45475 47636 45484
rect 8116 45407 8168 45416
rect 8116 45373 8125 45407
rect 8125 45373 8159 45407
rect 8159 45373 8168 45407
rect 8116 45364 8168 45373
rect 8392 45407 8444 45416
rect 8392 45373 8401 45407
rect 8401 45373 8435 45407
rect 8435 45373 8444 45407
rect 8392 45364 8444 45373
rect 24124 45364 24176 45416
rect 47584 45441 47593 45475
rect 47593 45441 47627 45475
rect 47627 45441 47636 45475
rect 47584 45432 47636 45441
rect 45744 45296 45796 45348
rect 1492 45228 1544 45280
rect 46480 45228 46532 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 8116 45024 8168 45076
rect 46296 45024 46348 45076
rect 2044 44820 2096 44872
rect 15108 44888 15160 44940
rect 22376 44888 22428 44940
rect 30104 44888 30156 44940
rect 46480 44931 46532 44940
rect 46480 44897 46489 44931
rect 46489 44897 46523 44931
rect 46523 44897 46532 44931
rect 46480 44888 46532 44897
rect 48136 44931 48188 44940
rect 48136 44897 48145 44931
rect 48145 44897 48179 44931
rect 48179 44897 48188 44931
rect 48136 44888 48188 44897
rect 8944 44863 8996 44872
rect 8944 44829 8953 44863
rect 8953 44829 8987 44863
rect 8987 44829 8996 44863
rect 8944 44820 8996 44829
rect 46296 44863 46348 44872
rect 46296 44829 46305 44863
rect 46305 44829 46339 44863
rect 46339 44829 46348 44863
rect 46296 44820 46348 44829
rect 2228 44684 2280 44736
rect 3516 44684 3568 44736
rect 23756 44752 23808 44804
rect 25596 44684 25648 44736
rect 38660 44684 38712 44736
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 2228 44455 2280 44464
rect 2228 44421 2237 44455
rect 2237 44421 2271 44455
rect 2271 44421 2280 44455
rect 2228 44412 2280 44421
rect 2044 44387 2096 44396
rect 2044 44353 2053 44387
rect 2053 44353 2087 44387
rect 2087 44353 2096 44387
rect 2044 44344 2096 44353
rect 23756 44387 23808 44396
rect 23756 44353 23765 44387
rect 23765 44353 23799 44387
rect 23799 44353 23808 44387
rect 23756 44344 23808 44353
rect 46296 44344 46348 44396
rect 2780 44319 2832 44328
rect 2780 44285 2789 44319
rect 2789 44285 2823 44319
rect 2823 44285 2832 44319
rect 2780 44276 2832 44285
rect 23848 44276 23900 44328
rect 24768 44319 24820 44328
rect 24768 44285 24777 44319
rect 24777 44285 24811 44319
rect 24811 44285 24820 44319
rect 24768 44276 24820 44285
rect 47032 44183 47084 44192
rect 47032 44149 47041 44183
rect 47041 44149 47075 44183
rect 47075 44149 47084 44183
rect 47032 44140 47084 44149
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 8944 43868 8996 43920
rect 15108 43800 15160 43852
rect 1860 43775 1912 43784
rect 1860 43741 1869 43775
rect 1869 43741 1903 43775
rect 1903 43741 1912 43775
rect 1860 43732 1912 43741
rect 20168 43732 20220 43784
rect 23756 43732 23808 43784
rect 26884 43732 26936 43784
rect 2320 43664 2372 43716
rect 23572 43664 23624 43716
rect 24952 43664 25004 43716
rect 47032 43800 47084 43852
rect 45836 43664 45888 43716
rect 46940 43664 46992 43716
rect 48136 43707 48188 43716
rect 48136 43673 48145 43707
rect 48145 43673 48179 43707
rect 48179 43673 48188 43707
rect 48136 43664 48188 43673
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 28816 43392 28868 43444
rect 46940 43435 46992 43444
rect 46940 43401 46949 43435
rect 46949 43401 46983 43435
rect 46983 43401 46992 43435
rect 46940 43392 46992 43401
rect 1860 43367 1912 43376
rect 1860 43333 1869 43367
rect 1869 43333 1903 43367
rect 1903 43333 1912 43367
rect 1860 43324 1912 43333
rect 20536 43367 20588 43376
rect 2136 43188 2188 43240
rect 20536 43333 20545 43367
rect 20545 43333 20579 43367
rect 20579 43333 20588 43367
rect 20536 43324 20588 43333
rect 20168 43299 20220 43308
rect 20168 43265 20177 43299
rect 20177 43265 20211 43299
rect 20211 43265 20220 43299
rect 20168 43256 20220 43265
rect 22008 43256 22060 43308
rect 22744 43256 22796 43308
rect 24676 43299 24728 43308
rect 24676 43265 24685 43299
rect 24685 43265 24719 43299
rect 24719 43265 24728 43299
rect 24676 43256 24728 43265
rect 24584 43188 24636 43240
rect 24860 43299 24912 43308
rect 24860 43265 24869 43299
rect 24869 43265 24903 43299
rect 24903 43265 24912 43299
rect 24860 43256 24912 43265
rect 25044 43299 25096 43308
rect 25044 43265 25053 43299
rect 25053 43265 25087 43299
rect 25087 43265 25096 43299
rect 27160 43299 27212 43308
rect 25044 43256 25096 43265
rect 27160 43265 27169 43299
rect 27169 43265 27203 43299
rect 27203 43265 27212 43299
rect 27160 43256 27212 43265
rect 27436 43299 27488 43308
rect 27436 43265 27445 43299
rect 27445 43265 27479 43299
rect 27479 43265 27488 43299
rect 27436 43256 27488 43265
rect 45836 43256 45888 43308
rect 47860 43299 47912 43308
rect 47860 43265 47869 43299
rect 47869 43265 47903 43299
rect 47903 43265 47912 43299
rect 47860 43256 47912 43265
rect 40316 43188 40368 43240
rect 2412 43052 2464 43104
rect 22284 43095 22336 43104
rect 22284 43061 22293 43095
rect 22293 43061 22327 43095
rect 22327 43061 22336 43095
rect 22284 43052 22336 43061
rect 24952 43052 25004 43104
rect 26976 43095 27028 43104
rect 26976 43061 26985 43095
rect 26985 43061 27019 43095
rect 27019 43061 27028 43095
rect 26976 43052 27028 43061
rect 47216 43052 47268 43104
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 20168 42644 20220 42696
rect 21364 42687 21416 42696
rect 21364 42653 21373 42687
rect 21373 42653 21407 42687
rect 21407 42653 21416 42687
rect 21364 42644 21416 42653
rect 24032 42644 24084 42696
rect 24952 42687 25004 42696
rect 24952 42653 24986 42687
rect 24986 42653 25004 42687
rect 24952 42644 25004 42653
rect 25688 42644 25740 42696
rect 26884 42687 26936 42696
rect 26884 42653 26893 42687
rect 26893 42653 26927 42687
rect 26927 42653 26936 42687
rect 26884 42644 26936 42653
rect 26976 42687 27028 42696
rect 26976 42653 26985 42687
rect 26985 42653 27019 42687
rect 27019 42653 27028 42687
rect 26976 42644 27028 42653
rect 27528 42644 27580 42696
rect 27988 42644 28040 42696
rect 29092 42712 29144 42764
rect 28816 42687 28868 42696
rect 28816 42653 28825 42687
rect 28825 42653 28859 42687
rect 28859 42653 28868 42687
rect 28816 42644 28868 42653
rect 29368 42644 29420 42696
rect 29552 42687 29604 42696
rect 29552 42653 29561 42687
rect 29561 42653 29595 42687
rect 29595 42653 29604 42687
rect 29552 42644 29604 42653
rect 20076 42619 20128 42628
rect 20076 42585 20085 42619
rect 20085 42585 20119 42619
rect 20119 42585 20128 42619
rect 20076 42576 20128 42585
rect 21824 42576 21876 42628
rect 23388 42576 23440 42628
rect 22744 42551 22796 42560
rect 22744 42517 22753 42551
rect 22753 42517 22787 42551
rect 22787 42517 22796 42551
rect 22744 42508 22796 42517
rect 24860 42576 24912 42628
rect 27896 42576 27948 42628
rect 47952 42619 48004 42628
rect 47952 42585 47961 42619
rect 47961 42585 47995 42619
rect 47995 42585 48004 42619
rect 47952 42576 48004 42585
rect 26148 42508 26200 42560
rect 26516 42551 26568 42560
rect 26516 42517 26525 42551
rect 26525 42517 26559 42551
rect 26559 42517 26568 42551
rect 26516 42508 26568 42517
rect 27804 42508 27856 42560
rect 30196 42508 30248 42560
rect 48044 42551 48096 42560
rect 48044 42517 48053 42551
rect 48053 42517 48087 42551
rect 48087 42517 48096 42551
rect 48044 42508 48096 42517
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 5448 42304 5500 42356
rect 21824 42347 21876 42356
rect 21824 42313 21833 42347
rect 21833 42313 21867 42347
rect 21867 42313 21876 42347
rect 21824 42304 21876 42313
rect 22100 42304 22152 42356
rect 23388 42304 23440 42356
rect 25688 42347 25740 42356
rect 25688 42313 25697 42347
rect 25697 42313 25731 42347
rect 25731 42313 25740 42347
rect 25688 42304 25740 42313
rect 21732 42168 21784 42220
rect 23848 42236 23900 42288
rect 24676 42236 24728 42288
rect 29184 42304 29236 42356
rect 29368 42304 29420 42356
rect 29644 42304 29696 42356
rect 29920 42304 29972 42356
rect 30840 42304 30892 42356
rect 48044 42304 48096 42356
rect 28816 42236 28868 42288
rect 21456 42100 21508 42152
rect 22284 42211 22336 42220
rect 22284 42177 22293 42211
rect 22293 42177 22327 42211
rect 22327 42177 22336 42211
rect 22284 42168 22336 42177
rect 23940 42168 23992 42220
rect 24032 42168 24084 42220
rect 23664 42100 23716 42152
rect 22744 42032 22796 42084
rect 27804 42211 27856 42220
rect 27804 42177 27813 42211
rect 27813 42177 27847 42211
rect 27847 42177 27856 42211
rect 27804 42168 27856 42177
rect 27988 42211 28040 42220
rect 27988 42177 27997 42211
rect 27997 42177 28031 42211
rect 28031 42177 28040 42211
rect 27988 42168 28040 42177
rect 29920 42168 29972 42220
rect 27712 42032 27764 42084
rect 1400 41964 1452 42016
rect 15752 41964 15804 42016
rect 24952 41964 25004 42016
rect 25964 41964 26016 42016
rect 29092 41964 29144 42016
rect 30196 42100 30248 42152
rect 30288 42007 30340 42016
rect 30288 41973 30297 42007
rect 30297 41973 30331 42007
rect 30331 41973 30340 42007
rect 30288 41964 30340 41973
rect 46296 41964 46348 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 23848 41760 23900 41812
rect 26148 41760 26200 41812
rect 24032 41692 24084 41744
rect 24768 41692 24820 41744
rect 1400 41667 1452 41676
rect 1400 41633 1409 41667
rect 1409 41633 1443 41667
rect 1443 41633 1452 41667
rect 1400 41624 1452 41633
rect 1860 41667 1912 41676
rect 1860 41633 1869 41667
rect 1869 41633 1903 41667
rect 1903 41633 1912 41667
rect 1860 41624 1912 41633
rect 15752 41667 15804 41676
rect 15752 41633 15761 41667
rect 15761 41633 15795 41667
rect 15795 41633 15804 41667
rect 15752 41624 15804 41633
rect 16580 41667 16632 41676
rect 16580 41633 16589 41667
rect 16589 41633 16623 41667
rect 16623 41633 16632 41667
rect 16580 41624 16632 41633
rect 25964 41667 26016 41676
rect 25964 41633 25973 41667
rect 25973 41633 26007 41667
rect 26007 41633 26016 41667
rect 25964 41624 26016 41633
rect 15568 41599 15620 41608
rect 15568 41565 15577 41599
rect 15577 41565 15611 41599
rect 15611 41565 15620 41599
rect 15568 41556 15620 41565
rect 20628 41556 20680 41608
rect 21364 41556 21416 41608
rect 24032 41556 24084 41608
rect 2596 41488 2648 41540
rect 20904 41488 20956 41540
rect 22744 41531 22796 41540
rect 22744 41497 22778 41531
rect 22778 41497 22796 41531
rect 22744 41488 22796 41497
rect 23664 41488 23716 41540
rect 24584 41488 24636 41540
rect 24952 41556 25004 41608
rect 25044 41599 25096 41608
rect 25044 41565 25053 41599
rect 25053 41565 25087 41599
rect 25087 41565 25096 41599
rect 25044 41556 25096 41565
rect 26516 41556 26568 41608
rect 27436 41760 27488 41812
rect 27896 41803 27948 41812
rect 27896 41769 27905 41803
rect 27905 41769 27939 41803
rect 27939 41769 27948 41803
rect 27896 41760 27948 41769
rect 27712 41624 27764 41676
rect 30288 41760 30340 41812
rect 29552 41667 29604 41676
rect 29552 41633 29561 41667
rect 29561 41633 29595 41667
rect 29595 41633 29604 41667
rect 29552 41624 29604 41633
rect 46296 41667 46348 41676
rect 46296 41633 46305 41667
rect 46305 41633 46339 41667
rect 46339 41633 46348 41667
rect 46296 41624 46348 41633
rect 48136 41599 48188 41608
rect 22008 41420 22060 41472
rect 23204 41420 23256 41472
rect 23848 41463 23900 41472
rect 23848 41429 23857 41463
rect 23857 41429 23891 41463
rect 23891 41429 23900 41463
rect 23848 41420 23900 41429
rect 23940 41420 23992 41472
rect 27528 41488 27580 41540
rect 48136 41565 48145 41599
rect 48145 41565 48179 41599
rect 48179 41565 48188 41599
rect 48136 41556 48188 41565
rect 29000 41488 29052 41540
rect 46480 41531 46532 41540
rect 46480 41497 46489 41531
rect 46489 41497 46523 41531
rect 46523 41497 46532 41531
rect 46480 41488 46532 41497
rect 26516 41420 26568 41472
rect 27160 41420 27212 41472
rect 29092 41420 29144 41472
rect 30932 41463 30984 41472
rect 30932 41429 30941 41463
rect 30941 41429 30975 41463
rect 30975 41429 30984 41463
rect 30932 41420 30984 41429
rect 33324 41420 33376 41472
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 2596 41259 2648 41268
rect 2596 41225 2605 41259
rect 2605 41225 2639 41259
rect 2639 41225 2648 41259
rect 2596 41216 2648 41225
rect 1860 41123 1912 41132
rect 1860 41089 1869 41123
rect 1869 41089 1903 41123
rect 1903 41089 1912 41123
rect 1860 41080 1912 41089
rect 2136 41080 2188 41132
rect 15200 41148 15252 41200
rect 15016 41123 15068 41132
rect 15016 41089 15050 41123
rect 15050 41089 15068 41123
rect 20812 41123 20864 41132
rect 15016 41080 15068 41089
rect 20812 41089 20821 41123
rect 20821 41089 20855 41123
rect 20855 41089 20864 41123
rect 20812 41080 20864 41089
rect 22744 41216 22796 41268
rect 24216 41216 24268 41268
rect 29000 41216 29052 41268
rect 29184 41259 29236 41268
rect 29184 41225 29193 41259
rect 29193 41225 29227 41259
rect 29227 41225 29236 41259
rect 29184 41216 29236 41225
rect 46480 41216 46532 41268
rect 21180 41123 21232 41132
rect 21180 41089 21189 41123
rect 21189 41089 21223 41123
rect 21223 41089 21232 41123
rect 21180 41080 21232 41089
rect 22008 41123 22060 41132
rect 21456 41012 21508 41064
rect 20904 40944 20956 40996
rect 1400 40876 1452 40928
rect 15660 40876 15712 40928
rect 22008 41089 22017 41123
rect 22017 41089 22051 41123
rect 22051 41089 22060 41123
rect 22008 41080 22060 41089
rect 22836 41080 22888 41132
rect 23017 41126 23069 41135
rect 23017 41092 23026 41126
rect 23026 41092 23060 41126
rect 23060 41092 23069 41126
rect 23017 41083 23069 41092
rect 25228 41148 25280 41200
rect 26884 41148 26936 41200
rect 23296 41123 23348 41132
rect 23296 41089 23305 41123
rect 23305 41089 23339 41123
rect 23339 41089 23348 41123
rect 23296 41080 23348 41089
rect 23664 41080 23716 41132
rect 23848 41080 23900 41132
rect 23204 41012 23256 41064
rect 23296 40944 23348 40996
rect 27436 40944 27488 40996
rect 29092 41080 29144 41132
rect 30932 41080 30984 41132
rect 32128 41080 32180 41132
rect 46664 41123 46716 41132
rect 46664 41089 46673 41123
rect 46673 41089 46707 41123
rect 46707 41089 46716 41123
rect 46664 41080 46716 41089
rect 47952 41123 48004 41132
rect 47952 41089 47961 41123
rect 47961 41089 47995 41123
rect 47995 41089 48004 41123
rect 47952 41080 48004 41089
rect 29552 41012 29604 41064
rect 30288 41012 30340 41064
rect 32312 41055 32364 41064
rect 32312 41021 32321 41055
rect 32321 41021 32355 41055
rect 32355 41021 32364 41055
rect 32312 41012 32364 41021
rect 22100 40876 22152 40928
rect 22468 40876 22520 40928
rect 23112 40876 23164 40928
rect 25228 40876 25280 40928
rect 33784 40876 33836 40928
rect 47400 40876 47452 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 23296 40672 23348 40724
rect 27344 40672 27396 40724
rect 28816 40604 28868 40656
rect 32220 40672 32272 40724
rect 29184 40468 29236 40520
rect 31116 40511 31168 40520
rect 1860 40443 1912 40452
rect 1860 40409 1869 40443
rect 1869 40409 1903 40443
rect 1903 40409 1912 40443
rect 1860 40400 1912 40409
rect 23388 40400 23440 40452
rect 29828 40400 29880 40452
rect 17132 40332 17184 40384
rect 23664 40332 23716 40384
rect 30748 40400 30800 40452
rect 30840 40332 30892 40384
rect 31116 40477 31125 40511
rect 31125 40477 31159 40511
rect 31159 40477 31168 40511
rect 31116 40468 31168 40477
rect 32404 40536 32456 40588
rect 32956 40536 33008 40588
rect 33324 40511 33376 40520
rect 33324 40477 33333 40511
rect 33333 40477 33367 40511
rect 33367 40477 33376 40511
rect 33324 40468 33376 40477
rect 31760 40400 31812 40452
rect 31668 40375 31720 40384
rect 31668 40341 31677 40375
rect 31677 40341 31711 40375
rect 31711 40341 31720 40375
rect 31668 40332 31720 40341
rect 33784 40400 33836 40452
rect 46480 40443 46532 40452
rect 46480 40409 46489 40443
rect 46489 40409 46523 40443
rect 46523 40409 46532 40443
rect 46480 40400 46532 40409
rect 48136 40443 48188 40452
rect 48136 40409 48145 40443
rect 48145 40409 48179 40443
rect 48179 40409 48188 40443
rect 48136 40400 48188 40409
rect 33416 40332 33468 40384
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 29828 40171 29880 40180
rect 21272 40060 21324 40112
rect 23848 40060 23900 40112
rect 24492 40060 24544 40112
rect 22008 39992 22060 40044
rect 23204 39992 23256 40044
rect 29828 40137 29837 40171
rect 29837 40137 29871 40171
rect 29871 40137 29880 40171
rect 29828 40128 29880 40137
rect 24860 39992 24912 40044
rect 25780 40035 25832 40044
rect 25780 40001 25789 40035
rect 25789 40001 25823 40035
rect 25823 40001 25832 40035
rect 25780 39992 25832 40001
rect 26976 40060 27028 40112
rect 31024 40060 31076 40112
rect 32220 40128 32272 40180
rect 33416 40128 33468 40180
rect 46480 40128 46532 40180
rect 31668 40060 31720 40112
rect 26056 40035 26108 40044
rect 26056 40001 26065 40035
rect 26065 40001 26099 40035
rect 26099 40001 26108 40035
rect 26056 39992 26108 40001
rect 29828 39992 29880 40044
rect 20536 39924 20588 39976
rect 23296 39924 23348 39976
rect 30748 39992 30800 40044
rect 2044 39788 2096 39840
rect 5540 39788 5592 39840
rect 6092 39788 6144 39840
rect 17224 39788 17276 39840
rect 20352 39788 20404 39840
rect 24400 39856 24452 39908
rect 24768 39788 24820 39840
rect 25964 39788 26016 39840
rect 30196 39856 30248 39908
rect 32312 39924 32364 39976
rect 33232 40035 33284 40044
rect 33232 40001 33266 40035
rect 33266 40001 33284 40035
rect 33232 39992 33284 40001
rect 35900 39992 35952 40044
rect 37188 39992 37240 40044
rect 32404 39788 32456 39840
rect 32496 39831 32548 39840
rect 32496 39797 32505 39831
rect 32505 39797 32539 39831
rect 32539 39797 32548 39831
rect 32496 39788 32548 39797
rect 33968 39788 34020 39840
rect 46296 39788 46348 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 17224 39584 17276 39636
rect 23204 39627 23256 39636
rect 21272 39559 21324 39568
rect 21272 39525 21281 39559
rect 21281 39525 21315 39559
rect 21315 39525 21324 39559
rect 21272 39516 21324 39525
rect 23204 39593 23213 39627
rect 23213 39593 23247 39627
rect 23247 39593 23256 39627
rect 23204 39584 23256 39593
rect 23296 39584 23348 39636
rect 31852 39584 31904 39636
rect 32128 39627 32180 39636
rect 32128 39593 32137 39627
rect 32137 39593 32171 39627
rect 32171 39593 32180 39627
rect 32128 39584 32180 39593
rect 25136 39516 25188 39568
rect 32496 39516 32548 39568
rect 5540 39380 5592 39432
rect 20720 39380 20772 39432
rect 21824 39380 21876 39432
rect 22468 39380 22520 39432
rect 23480 39423 23532 39432
rect 23480 39389 23489 39423
rect 23489 39389 23523 39423
rect 23523 39389 23532 39423
rect 23480 39380 23532 39389
rect 19984 39312 20036 39364
rect 23940 39380 23992 39432
rect 24768 39380 24820 39432
rect 25964 39380 26016 39432
rect 26424 39380 26476 39432
rect 27252 39448 27304 39500
rect 30288 39491 30340 39500
rect 24400 39312 24452 39364
rect 2228 39244 2280 39296
rect 22192 39244 22244 39296
rect 23480 39244 23532 39296
rect 23664 39244 23716 39296
rect 24860 39312 24912 39364
rect 24952 39312 25004 39364
rect 27160 39312 27212 39364
rect 24584 39244 24636 39296
rect 27436 39244 27488 39296
rect 27988 39380 28040 39432
rect 30288 39457 30297 39491
rect 30297 39457 30331 39491
rect 30331 39457 30340 39491
rect 30288 39448 30340 39457
rect 32312 39380 32364 39432
rect 33232 39491 33284 39500
rect 33232 39457 33241 39491
rect 33241 39457 33275 39491
rect 33275 39457 33284 39491
rect 33232 39448 33284 39457
rect 33324 39448 33376 39500
rect 46296 39491 46348 39500
rect 32772 39423 32824 39432
rect 32772 39389 32781 39423
rect 32781 39389 32815 39423
rect 32815 39389 32824 39423
rect 33508 39423 33560 39432
rect 32772 39380 32824 39389
rect 33508 39389 33531 39423
rect 33531 39389 33560 39423
rect 33508 39380 33560 39389
rect 46296 39457 46305 39491
rect 46305 39457 46339 39491
rect 46339 39457 46348 39491
rect 46296 39448 46348 39457
rect 48136 39491 48188 39500
rect 48136 39457 48145 39491
rect 48145 39457 48179 39491
rect 48179 39457 48188 39491
rect 48136 39448 48188 39457
rect 33876 39423 33928 39432
rect 28080 39355 28132 39364
rect 28080 39321 28089 39355
rect 28089 39321 28123 39355
rect 28123 39321 28132 39355
rect 28080 39312 28132 39321
rect 28816 39312 28868 39364
rect 30380 39312 30432 39364
rect 33324 39312 33376 39364
rect 33876 39389 33885 39423
rect 33885 39389 33919 39423
rect 33919 39389 33928 39423
rect 33876 39380 33928 39389
rect 35900 39380 35952 39432
rect 33968 39312 34020 39364
rect 34244 39312 34296 39364
rect 35992 39312 36044 39364
rect 46756 39312 46808 39364
rect 30932 39244 30984 39296
rect 31024 39244 31076 39296
rect 31668 39287 31720 39296
rect 31668 39253 31677 39287
rect 31677 39253 31711 39287
rect 31711 39253 31720 39287
rect 31668 39244 31720 39253
rect 33600 39244 33652 39296
rect 37464 39244 37516 39296
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 19984 39040 20036 39092
rect 26056 39040 26108 39092
rect 26424 39083 26476 39092
rect 26424 39049 26433 39083
rect 26433 39049 26467 39083
rect 26467 39049 26476 39083
rect 26424 39040 26476 39049
rect 26976 39083 27028 39092
rect 26976 39049 26985 39083
rect 26985 39049 27019 39083
rect 27019 39049 27028 39083
rect 26976 39040 27028 39049
rect 28080 39040 28132 39092
rect 29092 39040 29144 39092
rect 29644 39083 29696 39092
rect 29644 39049 29653 39083
rect 29653 39049 29687 39083
rect 29687 39049 29696 39083
rect 29644 39040 29696 39049
rect 30380 39083 30432 39092
rect 30380 39049 30389 39083
rect 30389 39049 30423 39083
rect 30423 39049 30432 39083
rect 30380 39040 30432 39049
rect 31852 39040 31904 39092
rect 35992 39083 36044 39092
rect 2228 39015 2280 39024
rect 2228 38981 2237 39015
rect 2237 38981 2271 39015
rect 2271 38981 2280 39015
rect 2228 38972 2280 38981
rect 2044 38947 2096 38956
rect 2044 38913 2053 38947
rect 2053 38913 2087 38947
rect 2087 38913 2096 38947
rect 2044 38904 2096 38913
rect 18604 38904 18656 38956
rect 2780 38879 2832 38888
rect 2780 38845 2789 38879
rect 2789 38845 2823 38879
rect 2823 38845 2832 38879
rect 2780 38836 2832 38845
rect 20352 38947 20404 38956
rect 20352 38913 20361 38947
rect 20361 38913 20395 38947
rect 20395 38913 20404 38947
rect 20352 38904 20404 38913
rect 21916 38904 21968 38956
rect 22100 38947 22152 38956
rect 22100 38913 22134 38947
rect 22134 38913 22152 38947
rect 22100 38904 22152 38913
rect 20628 38836 20680 38888
rect 21824 38879 21876 38888
rect 21824 38845 21833 38879
rect 21833 38845 21867 38879
rect 21867 38845 21876 38879
rect 21824 38836 21876 38845
rect 21272 38700 21324 38752
rect 23388 38904 23440 38956
rect 24768 38904 24820 38956
rect 25688 38904 25740 38956
rect 25872 38904 25924 38956
rect 23756 38836 23808 38888
rect 24676 38836 24728 38888
rect 27436 38947 27488 38956
rect 27436 38913 27445 38947
rect 27445 38913 27479 38947
rect 27479 38913 27488 38947
rect 27436 38904 27488 38913
rect 30380 38904 30432 38956
rect 33324 38972 33376 39024
rect 33600 39015 33652 39024
rect 33600 38981 33609 39015
rect 33609 38981 33643 39015
rect 33643 38981 33652 39015
rect 33600 38972 33652 38981
rect 34244 39015 34296 39024
rect 34244 38981 34253 39015
rect 34253 38981 34287 39015
rect 34287 38981 34296 39015
rect 34244 38972 34296 38981
rect 34336 38972 34388 39024
rect 35992 39049 36001 39083
rect 36001 39049 36035 39083
rect 36035 39049 36044 39083
rect 35992 39040 36044 39049
rect 36084 39040 36136 39092
rect 27988 38836 28040 38888
rect 28908 38836 28960 38888
rect 29828 38879 29880 38888
rect 29828 38845 29837 38879
rect 29837 38845 29871 38879
rect 29871 38845 29880 38879
rect 29828 38836 29880 38845
rect 23480 38700 23532 38752
rect 24584 38700 24636 38752
rect 29276 38768 29328 38820
rect 30840 38947 30892 38956
rect 30840 38913 30849 38947
rect 30849 38913 30883 38947
rect 30883 38913 30892 38947
rect 30840 38904 30892 38913
rect 31300 38904 31352 38956
rect 32772 38904 32824 38956
rect 34428 38904 34480 38956
rect 36176 38972 36228 39024
rect 46756 39083 46808 39092
rect 46756 39049 46765 39083
rect 46765 39049 46799 39083
rect 46799 39049 46808 39083
rect 46756 39040 46808 39049
rect 37464 39015 37516 39024
rect 37464 38981 37473 39015
rect 37473 38981 37507 39015
rect 37507 38981 37516 39015
rect 37464 38972 37516 38981
rect 36636 38947 36688 38956
rect 36636 38913 36645 38947
rect 36645 38913 36679 38947
rect 36679 38913 36688 38947
rect 36636 38904 36688 38913
rect 37280 38947 37332 38956
rect 37280 38913 37289 38947
rect 37289 38913 37323 38947
rect 37323 38913 37332 38947
rect 37280 38904 37332 38913
rect 37372 38904 37424 38956
rect 48136 38947 48188 38956
rect 48136 38913 48145 38947
rect 48145 38913 48179 38947
rect 48179 38913 48188 38947
rect 48136 38904 48188 38913
rect 45928 38836 45980 38888
rect 34428 38700 34480 38752
rect 34520 38700 34572 38752
rect 35716 38700 35768 38752
rect 35808 38700 35860 38752
rect 37280 38700 37332 38752
rect 46756 38700 46808 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 22100 38496 22152 38548
rect 22468 38496 22520 38548
rect 25688 38539 25740 38548
rect 25688 38505 25697 38539
rect 25697 38505 25731 38539
rect 25731 38505 25740 38539
rect 25688 38496 25740 38505
rect 18604 38292 18656 38344
rect 21824 38292 21876 38344
rect 21916 38292 21968 38344
rect 23020 38428 23072 38480
rect 22192 38335 22244 38344
rect 22192 38301 22201 38335
rect 22201 38301 22235 38335
rect 22235 38301 22244 38335
rect 22192 38292 22244 38301
rect 23940 38428 23992 38480
rect 25780 38428 25832 38480
rect 27804 38496 27856 38548
rect 23480 38360 23532 38412
rect 24676 38292 24728 38344
rect 27160 38428 27212 38480
rect 18696 38224 18748 38276
rect 21364 38224 21416 38276
rect 23020 38224 23072 38276
rect 23664 38224 23716 38276
rect 29276 38360 29328 38412
rect 19984 38156 20036 38208
rect 26056 38156 26108 38208
rect 28816 38335 28868 38344
rect 28816 38301 28825 38335
rect 28825 38301 28859 38335
rect 28859 38301 28868 38335
rect 28816 38292 28868 38301
rect 29000 38335 29052 38344
rect 29000 38301 29009 38335
rect 29009 38301 29043 38335
rect 29043 38301 29052 38335
rect 29000 38292 29052 38301
rect 30288 38292 30340 38344
rect 32864 38335 32916 38344
rect 32864 38301 32873 38335
rect 32873 38301 32907 38335
rect 32907 38301 32916 38335
rect 32864 38292 32916 38301
rect 33140 38292 33192 38344
rect 33876 38292 33928 38344
rect 30380 38156 30432 38208
rect 32496 38156 32548 38208
rect 35900 38292 35952 38344
rect 47860 38335 47912 38344
rect 47860 38301 47869 38335
rect 47869 38301 47903 38335
rect 47903 38301 47912 38335
rect 47860 38292 47912 38301
rect 33140 38156 33192 38208
rect 34520 38156 34572 38208
rect 35624 38156 35676 38208
rect 35808 38199 35860 38208
rect 35808 38165 35817 38199
rect 35817 38165 35851 38199
rect 35851 38165 35860 38199
rect 35808 38156 35860 38165
rect 36084 38224 36136 38276
rect 47124 38156 47176 38208
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 18696 37952 18748 38004
rect 22008 37995 22060 38004
rect 22008 37961 22017 37995
rect 22017 37961 22051 37995
rect 22051 37961 22060 37995
rect 22008 37952 22060 37961
rect 25780 37952 25832 38004
rect 27436 37952 27488 38004
rect 28816 37952 28868 38004
rect 36084 37995 36136 38004
rect 36084 37961 36093 37995
rect 36093 37961 36127 37995
rect 36127 37961 36136 37995
rect 36084 37952 36136 37961
rect 1860 37859 1912 37868
rect 1860 37825 1869 37859
rect 1869 37825 1903 37859
rect 1903 37825 1912 37859
rect 1860 37816 1912 37825
rect 18880 37859 18932 37868
rect 18880 37825 18889 37859
rect 18889 37825 18923 37859
rect 18923 37825 18932 37859
rect 18880 37816 18932 37825
rect 19800 37884 19852 37936
rect 19984 37884 20036 37936
rect 24584 37884 24636 37936
rect 24676 37884 24728 37936
rect 26240 37884 26292 37936
rect 2596 37680 2648 37732
rect 20352 37816 20404 37868
rect 20536 37816 20588 37868
rect 21364 37816 21416 37868
rect 26424 37816 26476 37868
rect 27344 37816 27396 37868
rect 28080 37816 28132 37868
rect 29092 37884 29144 37936
rect 29736 37816 29788 37868
rect 30288 37816 30340 37868
rect 31760 37816 31812 37868
rect 32496 37816 32548 37868
rect 23940 37791 23992 37800
rect 23940 37757 23949 37791
rect 23949 37757 23983 37791
rect 23983 37757 23992 37791
rect 23940 37748 23992 37757
rect 27528 37748 27580 37800
rect 29828 37748 29880 37800
rect 36176 37748 36228 37800
rect 19616 37680 19668 37732
rect 20536 37680 20588 37732
rect 35808 37680 35860 37732
rect 36728 37859 36780 37868
rect 36728 37825 36737 37859
rect 36737 37825 36771 37859
rect 36771 37825 36780 37859
rect 36728 37816 36780 37825
rect 46756 37816 46808 37868
rect 21180 37612 21232 37664
rect 26332 37612 26384 37664
rect 32680 37612 32732 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 21916 37408 21968 37460
rect 29000 37408 29052 37460
rect 31300 37408 31352 37460
rect 32864 37408 32916 37460
rect 19616 37340 19668 37392
rect 21548 37383 21600 37392
rect 21548 37349 21557 37383
rect 21557 37349 21591 37383
rect 21591 37349 21600 37383
rect 21548 37340 21600 37349
rect 29276 37340 29328 37392
rect 19432 37204 19484 37256
rect 29092 37272 29144 37324
rect 29828 37272 29880 37324
rect 1860 37179 1912 37188
rect 1860 37145 1869 37179
rect 1869 37145 1903 37179
rect 1903 37145 1912 37179
rect 1860 37136 1912 37145
rect 19248 37111 19300 37120
rect 19248 37077 19257 37111
rect 19257 37077 19291 37111
rect 19291 37077 19300 37111
rect 19248 37068 19300 37077
rect 19800 37204 19852 37256
rect 19984 37136 20036 37188
rect 21824 37204 21876 37256
rect 23940 37204 23992 37256
rect 24768 37204 24820 37256
rect 26700 37247 26752 37256
rect 26700 37213 26709 37247
rect 26709 37213 26743 37247
rect 26743 37213 26752 37247
rect 26700 37204 26752 37213
rect 27344 37204 27396 37256
rect 32404 37340 32456 37392
rect 36176 37340 36228 37392
rect 33324 37272 33376 37324
rect 32404 37247 32456 37256
rect 21364 37179 21416 37188
rect 20812 37068 20864 37120
rect 21364 37145 21373 37179
rect 21373 37145 21407 37179
rect 21407 37145 21416 37179
rect 21364 37136 21416 37145
rect 22652 37179 22704 37188
rect 22652 37145 22661 37179
rect 22661 37145 22695 37179
rect 22695 37145 22704 37179
rect 22652 37136 22704 37145
rect 23296 37136 23348 37188
rect 24584 37179 24636 37188
rect 24584 37145 24593 37179
rect 24593 37145 24627 37179
rect 24627 37145 24636 37179
rect 24584 37136 24636 37145
rect 21548 37068 21600 37120
rect 22928 37068 22980 37120
rect 24400 37068 24452 37120
rect 25780 37136 25832 37188
rect 26056 37179 26108 37188
rect 24860 37068 24912 37120
rect 26056 37145 26065 37179
rect 26065 37145 26099 37179
rect 26099 37145 26108 37179
rect 26056 37136 26108 37145
rect 26332 37136 26384 37188
rect 26976 37179 27028 37188
rect 26976 37145 27010 37179
rect 27010 37145 27028 37179
rect 26976 37136 27028 37145
rect 27988 37136 28040 37188
rect 29000 37136 29052 37188
rect 29736 37179 29788 37188
rect 29736 37145 29745 37179
rect 29745 37145 29779 37179
rect 29779 37145 29788 37179
rect 29736 37136 29788 37145
rect 27436 37068 27488 37120
rect 28080 37111 28132 37120
rect 28080 37077 28089 37111
rect 28089 37077 28123 37111
rect 28123 37077 28132 37111
rect 28080 37068 28132 37077
rect 28540 37068 28592 37120
rect 29368 37068 29420 37120
rect 32404 37213 32413 37247
rect 32413 37213 32447 37247
rect 32447 37213 32456 37247
rect 32404 37204 32456 37213
rect 32680 37247 32732 37256
rect 32680 37213 32689 37247
rect 32689 37213 32723 37247
rect 32723 37213 32732 37247
rect 32680 37204 32732 37213
rect 30748 37111 30800 37120
rect 30748 37077 30757 37111
rect 30757 37077 30791 37111
rect 30791 37077 30800 37111
rect 30748 37068 30800 37077
rect 33232 37136 33284 37188
rect 33600 37247 33652 37256
rect 33600 37213 33609 37247
rect 33609 37213 33643 37247
rect 33643 37213 33652 37247
rect 33600 37204 33652 37213
rect 33876 37204 33928 37256
rect 36084 37247 36136 37256
rect 36084 37213 36093 37247
rect 36093 37213 36127 37247
rect 36127 37213 36136 37247
rect 36084 37204 36136 37213
rect 40684 37272 40736 37324
rect 46848 37272 46900 37324
rect 36636 37204 36688 37256
rect 35532 37136 35584 37188
rect 33140 37111 33192 37120
rect 33140 37077 33149 37111
rect 33149 37077 33183 37111
rect 33183 37077 33192 37111
rect 33140 37068 33192 37077
rect 35716 37068 35768 37120
rect 35992 37068 36044 37120
rect 36360 37136 36412 37188
rect 42800 37204 42852 37256
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 17408 36864 17460 36916
rect 24400 36864 24452 36916
rect 24584 36864 24636 36916
rect 19248 36796 19300 36848
rect 20352 36796 20404 36848
rect 22652 36796 22704 36848
rect 18604 36771 18656 36780
rect 18604 36737 18613 36771
rect 18613 36737 18647 36771
rect 18647 36737 18656 36771
rect 18604 36728 18656 36737
rect 20812 36703 20864 36712
rect 20812 36669 20821 36703
rect 20821 36669 20855 36703
rect 20855 36669 20864 36703
rect 20812 36660 20864 36669
rect 22468 36728 22520 36780
rect 23940 36796 23992 36848
rect 24768 36796 24820 36848
rect 24400 36728 24452 36780
rect 26700 36864 26752 36916
rect 26976 36839 27028 36848
rect 26976 36805 26985 36839
rect 26985 36805 27019 36839
rect 27019 36805 27028 36839
rect 26976 36796 27028 36805
rect 27068 36796 27120 36848
rect 21824 36660 21876 36712
rect 26884 36660 26936 36712
rect 27436 36771 27488 36780
rect 27436 36737 27445 36771
rect 27445 36737 27479 36771
rect 27479 36737 27488 36771
rect 27988 36796 28040 36848
rect 28172 36839 28224 36848
rect 28172 36805 28181 36839
rect 28181 36805 28215 36839
rect 28215 36805 28224 36839
rect 28172 36796 28224 36805
rect 33600 36864 33652 36916
rect 35992 36907 36044 36916
rect 35992 36873 36001 36907
rect 36001 36873 36035 36907
rect 36035 36873 36044 36907
rect 35992 36864 36044 36873
rect 27436 36728 27488 36737
rect 28816 36728 28868 36780
rect 29368 36771 29420 36780
rect 29368 36737 29382 36771
rect 29382 36737 29416 36771
rect 29416 36737 29420 36771
rect 29368 36728 29420 36737
rect 29552 36771 29604 36780
rect 29552 36737 29561 36771
rect 29561 36737 29595 36771
rect 29595 36737 29604 36771
rect 33140 36796 33192 36848
rect 35532 36796 35584 36848
rect 37004 36796 37056 36848
rect 29552 36728 29604 36737
rect 30104 36728 30156 36780
rect 31392 36728 31444 36780
rect 31944 36728 31996 36780
rect 32312 36728 32364 36780
rect 32404 36728 32456 36780
rect 33232 36771 33284 36780
rect 33232 36737 33241 36771
rect 33241 36737 33275 36771
rect 33275 36737 33284 36771
rect 33232 36728 33284 36737
rect 33324 36771 33376 36780
rect 33324 36737 33333 36771
rect 33333 36737 33367 36771
rect 33367 36737 33376 36771
rect 35624 36771 35676 36780
rect 33324 36728 33376 36737
rect 35624 36737 35633 36771
rect 35633 36737 35667 36771
rect 35667 36737 35676 36771
rect 35624 36728 35676 36737
rect 31760 36660 31812 36712
rect 33232 36592 33284 36644
rect 23204 36524 23256 36576
rect 23296 36567 23348 36576
rect 23296 36533 23305 36567
rect 23305 36533 23339 36567
rect 23339 36533 23348 36567
rect 23296 36524 23348 36533
rect 28816 36524 28868 36576
rect 30748 36524 30800 36576
rect 33324 36524 33376 36576
rect 46296 36524 46348 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 20536 36320 20588 36372
rect 22468 36363 22520 36372
rect 21548 36252 21600 36304
rect 22468 36329 22477 36363
rect 22477 36329 22511 36363
rect 22511 36329 22520 36363
rect 22468 36320 22520 36329
rect 22744 36320 22796 36372
rect 23296 36320 23348 36372
rect 24400 36363 24452 36372
rect 24400 36329 24409 36363
rect 24409 36329 24443 36363
rect 24443 36329 24452 36363
rect 24400 36320 24452 36329
rect 26056 36320 26108 36372
rect 28080 36320 28132 36372
rect 28172 36320 28224 36372
rect 2044 36116 2096 36168
rect 16672 36116 16724 36168
rect 20444 36184 20496 36236
rect 23020 36252 23072 36304
rect 23204 36252 23256 36304
rect 22744 36159 22796 36168
rect 19156 36048 19208 36100
rect 22744 36125 22753 36159
rect 22753 36125 22787 36159
rect 22787 36125 22796 36159
rect 22744 36116 22796 36125
rect 2964 36023 3016 36032
rect 2964 35989 2973 36023
rect 2973 35989 3007 36023
rect 3007 35989 3016 36023
rect 2964 35980 3016 35989
rect 19248 36023 19300 36032
rect 19248 35989 19257 36023
rect 19257 35989 19291 36023
rect 19291 35989 19300 36023
rect 19248 35980 19300 35989
rect 20812 36048 20864 36100
rect 21640 36048 21692 36100
rect 21916 35980 21968 36032
rect 22928 36159 22980 36168
rect 22928 36125 22937 36159
rect 22937 36125 22971 36159
rect 22971 36125 22980 36159
rect 22928 36116 22980 36125
rect 24676 36159 24728 36168
rect 24676 36125 24685 36159
rect 24685 36125 24719 36159
rect 24719 36125 24728 36159
rect 24676 36116 24728 36125
rect 23020 36048 23072 36100
rect 24860 36159 24912 36168
rect 24860 36125 24869 36159
rect 24869 36125 24903 36159
rect 24903 36125 24912 36159
rect 24860 36116 24912 36125
rect 29552 36252 29604 36304
rect 27252 36227 27304 36236
rect 27252 36193 27261 36227
rect 27261 36193 27295 36227
rect 27295 36193 27304 36227
rect 27252 36184 27304 36193
rect 27528 36184 27580 36236
rect 27988 36184 28040 36236
rect 24952 36048 25004 36100
rect 27068 36116 27120 36168
rect 28356 36116 28408 36168
rect 30012 36159 30064 36168
rect 30012 36125 30026 36159
rect 30026 36125 30060 36159
rect 30060 36125 30064 36159
rect 30012 36116 30064 36125
rect 30564 36116 30616 36168
rect 33232 36320 33284 36372
rect 34704 36320 34756 36372
rect 31760 36252 31812 36304
rect 35900 36320 35952 36372
rect 37004 36363 37056 36372
rect 37004 36329 37013 36363
rect 37013 36329 37047 36363
rect 37047 36329 37056 36363
rect 37004 36320 37056 36329
rect 46296 36227 46348 36236
rect 46296 36193 46305 36227
rect 46305 36193 46339 36227
rect 46339 36193 46348 36227
rect 46296 36184 46348 36193
rect 48136 36227 48188 36236
rect 48136 36193 48145 36227
rect 48145 36193 48179 36227
rect 48179 36193 48188 36227
rect 48136 36184 48188 36193
rect 35716 36116 35768 36168
rect 26240 36048 26292 36100
rect 26608 35980 26660 36032
rect 28172 36091 28224 36100
rect 28172 36057 28181 36091
rect 28181 36057 28215 36091
rect 28215 36057 28224 36091
rect 28172 36048 28224 36057
rect 30104 36048 30156 36100
rect 30748 36091 30800 36100
rect 30748 36057 30757 36091
rect 30757 36057 30791 36091
rect 30791 36057 30800 36091
rect 30748 36048 30800 36057
rect 47676 36048 47728 36100
rect 29828 35980 29880 36032
rect 30196 35980 30248 36032
rect 33324 35980 33376 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 20812 35819 20864 35828
rect 2964 35708 3016 35760
rect 19248 35708 19300 35760
rect 20812 35785 20821 35819
rect 20821 35785 20855 35819
rect 20855 35785 20864 35819
rect 20812 35776 20864 35785
rect 27988 35776 28040 35828
rect 28356 35819 28408 35828
rect 28356 35785 28365 35819
rect 28365 35785 28399 35819
rect 28399 35785 28408 35819
rect 28356 35776 28408 35785
rect 26424 35708 26476 35760
rect 26608 35708 26660 35760
rect 29920 35776 29972 35828
rect 30104 35708 30156 35760
rect 2044 35683 2096 35692
rect 2044 35649 2053 35683
rect 2053 35649 2087 35683
rect 2087 35649 2096 35683
rect 2044 35640 2096 35649
rect 11704 35640 11756 35692
rect 19432 35640 19484 35692
rect 20444 35683 20496 35692
rect 20444 35649 20453 35683
rect 20453 35649 20487 35683
rect 20487 35649 20496 35683
rect 20444 35640 20496 35649
rect 21456 35640 21508 35692
rect 26700 35640 26752 35692
rect 2780 35615 2832 35624
rect 2780 35581 2789 35615
rect 2789 35581 2823 35615
rect 2823 35581 2832 35615
rect 2780 35572 2832 35581
rect 18604 35615 18656 35624
rect 18604 35581 18613 35615
rect 18613 35581 18647 35615
rect 18647 35581 18656 35615
rect 18604 35572 18656 35581
rect 26240 35572 26292 35624
rect 26884 35572 26936 35624
rect 28172 35572 28224 35624
rect 29736 35640 29788 35692
rect 31300 35751 31352 35760
rect 31300 35717 31309 35751
rect 31309 35717 31343 35751
rect 31343 35717 31352 35751
rect 31300 35708 31352 35717
rect 31392 35708 31444 35760
rect 22836 35504 22888 35556
rect 28908 35504 28960 35556
rect 31484 35640 31536 35692
rect 47860 35683 47912 35692
rect 30196 35572 30248 35624
rect 30472 35615 30524 35624
rect 30472 35581 30481 35615
rect 30481 35581 30515 35615
rect 30515 35581 30524 35615
rect 30472 35572 30524 35581
rect 32036 35572 32088 35624
rect 30564 35504 30616 35556
rect 32588 35504 32640 35556
rect 47860 35649 47869 35683
rect 47869 35649 47903 35683
rect 47903 35649 47912 35683
rect 47860 35640 47912 35649
rect 1584 35436 1636 35488
rect 2596 35436 2648 35488
rect 15844 35436 15896 35488
rect 20812 35436 20864 35488
rect 21548 35436 21600 35488
rect 22008 35479 22060 35488
rect 22008 35445 22017 35479
rect 22017 35445 22051 35479
rect 22051 35445 22060 35479
rect 22008 35436 22060 35445
rect 32128 35479 32180 35488
rect 32128 35445 32137 35479
rect 32137 35445 32171 35479
rect 32171 35445 32180 35479
rect 32128 35436 32180 35445
rect 46296 35436 46348 35488
rect 47032 35479 47084 35488
rect 47032 35445 47041 35479
rect 47041 35445 47075 35479
rect 47075 35445 47084 35479
rect 47032 35436 47084 35445
rect 48044 35479 48096 35488
rect 48044 35445 48053 35479
rect 48053 35445 48087 35479
rect 48087 35445 48096 35479
rect 48044 35436 48096 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 17776 35232 17828 35284
rect 5356 35164 5408 35216
rect 15844 35164 15896 35216
rect 11704 35096 11756 35148
rect 20812 35232 20864 35284
rect 27528 35232 27580 35284
rect 29368 35164 29420 35216
rect 21456 35139 21508 35148
rect 21456 35105 21465 35139
rect 21465 35105 21499 35139
rect 21499 35105 21508 35139
rect 21456 35096 21508 35105
rect 28172 35096 28224 35148
rect 1400 35071 1452 35080
rect 1400 35037 1409 35071
rect 1409 35037 1443 35071
rect 1443 35037 1452 35071
rect 1400 35028 1452 35037
rect 15200 35028 15252 35080
rect 18604 35028 18656 35080
rect 19156 35028 19208 35080
rect 19984 35028 20036 35080
rect 21640 35028 21692 35080
rect 22560 35028 22612 35080
rect 23480 35071 23532 35080
rect 23480 35037 23489 35071
rect 23489 35037 23523 35071
rect 23523 35037 23532 35071
rect 23480 35028 23532 35037
rect 23848 35028 23900 35080
rect 18696 34892 18748 34944
rect 22652 34960 22704 35012
rect 26240 35028 26292 35080
rect 32036 35232 32088 35284
rect 31760 35096 31812 35148
rect 46296 35139 46348 35148
rect 46296 35105 46305 35139
rect 46305 35105 46339 35139
rect 46339 35105 46348 35139
rect 46296 35096 46348 35105
rect 48136 35139 48188 35148
rect 48136 35105 48145 35139
rect 48145 35105 48179 35139
rect 48179 35105 48188 35139
rect 48136 35096 48188 35105
rect 26332 34960 26384 35012
rect 26976 34960 27028 35012
rect 32128 35028 32180 35080
rect 45560 35028 45612 35080
rect 28724 34960 28776 35012
rect 29644 34960 29696 35012
rect 29828 35003 29880 35012
rect 29828 34969 29862 35003
rect 29862 34969 29880 35003
rect 29828 34960 29880 34969
rect 31576 35003 31628 35012
rect 31576 34969 31585 35003
rect 31585 34969 31619 35003
rect 31619 34969 31628 35003
rect 31576 34960 31628 34969
rect 32036 34960 32088 35012
rect 20628 34935 20680 34944
rect 20628 34901 20637 34935
rect 20637 34901 20671 34935
rect 20671 34901 20680 34935
rect 20628 34892 20680 34901
rect 23204 34892 23256 34944
rect 29552 34892 29604 34944
rect 29920 34892 29972 34944
rect 33232 34892 33284 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 12992 34688 13044 34740
rect 18696 34731 18748 34740
rect 15844 34663 15896 34672
rect 15844 34629 15853 34663
rect 15853 34629 15887 34663
rect 15887 34629 15896 34663
rect 15844 34620 15896 34629
rect 2044 34595 2096 34604
rect 2044 34561 2053 34595
rect 2053 34561 2087 34595
rect 2087 34561 2096 34595
rect 2044 34552 2096 34561
rect 3056 34552 3108 34604
rect 15200 34552 15252 34604
rect 17684 34552 17736 34604
rect 18696 34697 18705 34731
rect 18705 34697 18739 34731
rect 18739 34697 18748 34731
rect 18696 34688 18748 34697
rect 19064 34688 19116 34740
rect 19248 34620 19300 34672
rect 22284 34688 22336 34740
rect 23204 34688 23256 34740
rect 31484 34688 31536 34740
rect 31576 34688 31628 34740
rect 47676 34731 47728 34740
rect 47676 34697 47685 34731
rect 47685 34697 47719 34731
rect 47719 34697 47728 34731
rect 47676 34688 47728 34697
rect 20628 34620 20680 34672
rect 1768 34484 1820 34536
rect 14464 34527 14516 34536
rect 14464 34493 14473 34527
rect 14473 34493 14507 34527
rect 14507 34493 14516 34527
rect 14464 34484 14516 34493
rect 16580 34484 16632 34536
rect 19432 34552 19484 34604
rect 20444 34552 20496 34604
rect 22100 34595 22152 34604
rect 22100 34561 22134 34595
rect 22134 34561 22152 34595
rect 17776 34416 17828 34468
rect 22100 34552 22152 34561
rect 21824 34527 21876 34536
rect 21824 34493 21833 34527
rect 21833 34493 21867 34527
rect 21867 34493 21876 34527
rect 21824 34484 21876 34493
rect 23940 34595 23992 34604
rect 23940 34561 23949 34595
rect 23949 34561 23983 34595
rect 23983 34561 23992 34595
rect 23940 34552 23992 34561
rect 24216 34595 24268 34604
rect 24216 34561 24250 34595
rect 24250 34561 24268 34595
rect 26240 34595 26292 34604
rect 24216 34552 24268 34561
rect 26240 34561 26249 34595
rect 26249 34561 26283 34595
rect 26283 34561 26292 34595
rect 26240 34552 26292 34561
rect 26516 34620 26568 34672
rect 28540 34595 28592 34604
rect 28540 34561 28549 34595
rect 28549 34561 28583 34595
rect 28583 34561 28592 34595
rect 28540 34552 28592 34561
rect 30748 34620 30800 34672
rect 33232 34620 33284 34672
rect 39856 34620 39908 34672
rect 28172 34484 28224 34536
rect 28908 34484 28960 34536
rect 29644 34552 29696 34604
rect 46112 34595 46164 34604
rect 46112 34561 46121 34595
rect 46121 34561 46155 34595
rect 46155 34561 46164 34595
rect 46112 34552 46164 34561
rect 46572 34552 46624 34604
rect 47584 34595 47636 34604
rect 47584 34561 47593 34595
rect 47593 34561 47627 34595
rect 47627 34561 47636 34595
rect 47584 34552 47636 34561
rect 1400 34348 1452 34400
rect 2136 34391 2188 34400
rect 2136 34357 2145 34391
rect 2145 34357 2179 34391
rect 2179 34357 2188 34391
rect 2136 34348 2188 34357
rect 17500 34348 17552 34400
rect 21272 34391 21324 34400
rect 21272 34357 21281 34391
rect 21281 34357 21315 34391
rect 21315 34357 21324 34391
rect 21272 34348 21324 34357
rect 32220 34484 32272 34536
rect 33324 34484 33376 34536
rect 33508 34484 33560 34536
rect 46848 34527 46900 34536
rect 46848 34493 46857 34527
rect 46857 34493 46891 34527
rect 46891 34493 46900 34527
rect 46848 34484 46900 34493
rect 47676 34484 47728 34536
rect 48044 34484 48096 34536
rect 30564 34416 30616 34468
rect 23112 34348 23164 34400
rect 25688 34348 25740 34400
rect 30472 34348 30524 34400
rect 46480 34348 46532 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 17684 34187 17736 34196
rect 1400 34051 1452 34060
rect 1400 34017 1409 34051
rect 1409 34017 1443 34051
rect 1443 34017 1452 34051
rect 1400 34008 1452 34017
rect 2136 34008 2188 34060
rect 2780 34051 2832 34060
rect 2780 34017 2789 34051
rect 2789 34017 2823 34051
rect 2823 34017 2832 34051
rect 2780 34008 2832 34017
rect 17684 34153 17693 34187
rect 17693 34153 17727 34187
rect 17727 34153 17736 34187
rect 17684 34144 17736 34153
rect 22100 34144 22152 34196
rect 22192 34144 22244 34196
rect 23020 34144 23072 34196
rect 24216 34144 24268 34196
rect 30472 34144 30524 34196
rect 18144 34076 18196 34128
rect 19984 34119 20036 34128
rect 19984 34085 19993 34119
rect 19993 34085 20027 34119
rect 20027 34085 20036 34119
rect 19984 34076 20036 34085
rect 21916 34076 21968 34128
rect 11888 33915 11940 33924
rect 11888 33881 11897 33915
rect 11897 33881 11931 33915
rect 11931 33881 11940 33915
rect 11888 33872 11940 33881
rect 9864 33804 9916 33856
rect 15200 34008 15252 34060
rect 21272 34008 21324 34060
rect 16672 33872 16724 33924
rect 16580 33804 16632 33856
rect 21732 33983 21784 33992
rect 17500 33872 17552 33924
rect 20904 33872 20956 33924
rect 17868 33847 17920 33856
rect 17868 33813 17877 33847
rect 17877 33813 17911 33847
rect 17911 33813 17920 33847
rect 17868 33804 17920 33813
rect 21732 33949 21741 33983
rect 21741 33949 21775 33983
rect 21775 33949 21784 33983
rect 21732 33940 21784 33949
rect 22284 34008 22336 34060
rect 22560 33983 22612 33992
rect 22560 33949 22569 33983
rect 22569 33949 22603 33983
rect 22603 33949 22612 33983
rect 22560 33940 22612 33949
rect 23112 33940 23164 33992
rect 24768 34076 24820 34128
rect 23940 33940 23992 33992
rect 25044 33983 25096 33992
rect 25044 33949 25053 33983
rect 25053 33949 25087 33983
rect 25087 33949 25096 33983
rect 25044 33940 25096 33949
rect 25688 34076 25740 34128
rect 26884 34008 26936 34060
rect 27712 33940 27764 33992
rect 28172 33983 28224 33992
rect 28172 33949 28181 33983
rect 28181 33949 28215 33983
rect 28215 33949 28224 33983
rect 31484 34076 31536 34128
rect 31668 34008 31720 34060
rect 33508 34008 33560 34060
rect 47032 34076 47084 34128
rect 46480 34051 46532 34060
rect 46480 34017 46489 34051
rect 46489 34017 46523 34051
rect 46523 34017 46532 34051
rect 46480 34008 46532 34017
rect 48136 34051 48188 34060
rect 48136 34017 48145 34051
rect 48145 34017 48179 34051
rect 48179 34017 48188 34051
rect 48136 34008 48188 34017
rect 28172 33940 28224 33949
rect 22652 33804 22704 33856
rect 27436 33872 27488 33924
rect 29644 33915 29696 33924
rect 29644 33881 29653 33915
rect 29653 33881 29687 33915
rect 29687 33881 29696 33915
rect 29644 33872 29696 33881
rect 31576 33983 31628 33992
rect 31576 33949 31585 33983
rect 31585 33949 31619 33983
rect 31619 33949 31628 33983
rect 31576 33940 31628 33949
rect 32496 33940 32548 33992
rect 34428 33940 34480 33992
rect 25688 33804 25740 33856
rect 27160 33804 27212 33856
rect 29920 33804 29972 33856
rect 33324 33872 33376 33924
rect 33876 33915 33928 33924
rect 33876 33881 33885 33915
rect 33885 33881 33919 33915
rect 33919 33881 33928 33915
rect 33876 33872 33928 33881
rect 32036 33804 32088 33856
rect 32128 33804 32180 33856
rect 33140 33804 33192 33856
rect 33784 33847 33836 33856
rect 33784 33813 33793 33847
rect 33793 33813 33827 33847
rect 33827 33813 33836 33847
rect 33784 33804 33836 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 11888 33643 11940 33652
rect 11888 33609 11897 33643
rect 11897 33609 11931 33643
rect 11931 33609 11940 33643
rect 11888 33600 11940 33609
rect 14464 33600 14516 33652
rect 16764 33600 16816 33652
rect 23112 33600 23164 33652
rect 27436 33643 27488 33652
rect 1768 33507 1820 33516
rect 1768 33473 1777 33507
rect 1777 33473 1811 33507
rect 1811 33473 1820 33507
rect 1768 33464 1820 33473
rect 11704 33464 11756 33516
rect 16028 33532 16080 33584
rect 22284 33532 22336 33584
rect 27436 33609 27445 33643
rect 27445 33609 27479 33643
rect 27479 33609 27488 33643
rect 27436 33600 27488 33609
rect 28356 33600 28408 33652
rect 29644 33600 29696 33652
rect 30380 33643 30432 33652
rect 30380 33609 30389 33643
rect 30389 33609 30423 33643
rect 30423 33609 30432 33643
rect 30380 33600 30432 33609
rect 31576 33600 31628 33652
rect 33784 33600 33836 33652
rect 1952 33439 2004 33448
rect 1952 33405 1961 33439
rect 1961 33405 1995 33439
rect 1995 33405 2004 33439
rect 1952 33396 2004 33405
rect 2780 33439 2832 33448
rect 2780 33405 2789 33439
rect 2789 33405 2823 33439
rect 2823 33405 2832 33439
rect 2780 33396 2832 33405
rect 15752 33464 15804 33516
rect 16580 33464 16632 33516
rect 15936 33439 15988 33448
rect 15936 33405 15945 33439
rect 15945 33405 15979 33439
rect 15979 33405 15988 33439
rect 15936 33396 15988 33405
rect 17868 33464 17920 33516
rect 19432 33464 19484 33516
rect 23112 33507 23164 33516
rect 23112 33473 23123 33507
rect 23123 33473 23157 33507
rect 23157 33473 23164 33507
rect 24492 33532 24544 33584
rect 25044 33532 25096 33584
rect 26424 33532 26476 33584
rect 27712 33532 27764 33584
rect 32128 33575 32180 33584
rect 32128 33541 32137 33575
rect 32137 33541 32171 33575
rect 32171 33541 32180 33575
rect 32128 33532 32180 33541
rect 23112 33464 23164 33473
rect 17500 33439 17552 33448
rect 15292 33328 15344 33380
rect 17500 33405 17509 33439
rect 17509 33405 17543 33439
rect 17543 33405 17552 33439
rect 17500 33396 17552 33405
rect 18052 33396 18104 33448
rect 25780 33464 25832 33516
rect 27988 33464 28040 33516
rect 28172 33464 28224 33516
rect 28816 33464 28868 33516
rect 31392 33464 31444 33516
rect 32036 33464 32088 33516
rect 32496 33464 32548 33516
rect 33048 33507 33100 33516
rect 33048 33473 33057 33507
rect 33057 33473 33091 33507
rect 33091 33473 33100 33507
rect 33048 33464 33100 33473
rect 33324 33507 33376 33516
rect 33324 33473 33358 33507
rect 33358 33473 33376 33507
rect 33324 33464 33376 33473
rect 23388 33396 23440 33448
rect 28080 33439 28132 33448
rect 28080 33405 28089 33439
rect 28089 33405 28123 33439
rect 28123 33405 28132 33439
rect 28080 33396 28132 33405
rect 30472 33439 30524 33448
rect 30472 33405 30481 33439
rect 30481 33405 30515 33439
rect 30515 33405 30524 33439
rect 30472 33396 30524 33405
rect 34244 33396 34296 33448
rect 42800 33396 42852 33448
rect 46204 33439 46256 33448
rect 46204 33405 46213 33439
rect 46213 33405 46247 33439
rect 46247 33405 46256 33439
rect 46204 33396 46256 33405
rect 16672 33371 16724 33380
rect 16672 33337 16681 33371
rect 16681 33337 16715 33371
rect 16715 33337 16724 33371
rect 16672 33328 16724 33337
rect 26884 33328 26936 33380
rect 34428 33371 34480 33380
rect 34428 33337 34437 33371
rect 34437 33337 34471 33371
rect 34471 33337 34480 33371
rect 34428 33328 34480 33337
rect 2596 33260 2648 33312
rect 2780 33260 2832 33312
rect 11704 33260 11756 33312
rect 20536 33260 20588 33312
rect 24308 33260 24360 33312
rect 47768 33303 47820 33312
rect 47768 33269 47777 33303
rect 47777 33269 47811 33303
rect 47811 33269 47820 33303
rect 47768 33260 47820 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 1952 33056 2004 33108
rect 2596 33056 2648 33108
rect 23756 33099 23808 33108
rect 16028 32988 16080 33040
rect 23756 33065 23765 33099
rect 23765 33065 23799 33099
rect 23799 33065 23808 33099
rect 23756 33056 23808 33065
rect 28540 33056 28592 33108
rect 9036 32920 9088 32972
rect 2044 32784 2096 32836
rect 15936 32852 15988 32904
rect 18328 32895 18380 32904
rect 18328 32861 18337 32895
rect 18337 32861 18371 32895
rect 18371 32861 18380 32895
rect 18328 32852 18380 32861
rect 18512 32895 18564 32904
rect 18512 32861 18526 32895
rect 18526 32861 18560 32895
rect 18560 32861 18564 32895
rect 18512 32852 18564 32861
rect 19064 32852 19116 32904
rect 24124 32988 24176 33040
rect 19248 32963 19300 32972
rect 19248 32929 19257 32963
rect 19257 32929 19291 32963
rect 19291 32929 19300 32963
rect 19248 32920 19300 32929
rect 27068 32895 27120 32904
rect 27068 32861 27077 32895
rect 27077 32861 27111 32895
rect 27111 32861 27120 32895
rect 27068 32852 27120 32861
rect 27160 32852 27212 32904
rect 27620 32852 27672 32904
rect 30380 33056 30432 33108
rect 31392 33099 31444 33108
rect 31392 33065 31401 33099
rect 31401 33065 31435 33099
rect 31435 33065 31444 33099
rect 31392 33056 31444 33065
rect 34244 33056 34296 33108
rect 31484 32920 31536 32972
rect 31760 32852 31812 32904
rect 32220 32895 32272 32904
rect 32220 32861 32229 32895
rect 32229 32861 32263 32895
rect 32263 32861 32272 32895
rect 32220 32852 32272 32861
rect 47768 32920 47820 32972
rect 48044 32963 48096 32972
rect 48044 32929 48053 32963
rect 48053 32929 48087 32963
rect 48087 32929 48096 32963
rect 48044 32920 48096 32929
rect 32588 32895 32640 32904
rect 32588 32861 32597 32895
rect 32597 32861 32631 32895
rect 32631 32861 32640 32895
rect 32588 32852 32640 32861
rect 33140 32852 33192 32904
rect 23388 32784 23440 32836
rect 23848 32784 23900 32836
rect 29368 32784 29420 32836
rect 32496 32784 32548 32836
rect 46848 32784 46900 32836
rect 19156 32716 19208 32768
rect 20628 32759 20680 32768
rect 20628 32725 20637 32759
rect 20637 32725 20671 32759
rect 20671 32725 20680 32759
rect 20628 32716 20680 32725
rect 24768 32716 24820 32768
rect 25780 32759 25832 32768
rect 25780 32725 25789 32759
rect 25789 32725 25823 32759
rect 25823 32725 25832 32759
rect 25780 32716 25832 32725
rect 27988 32716 28040 32768
rect 28816 32716 28868 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 2688 32444 2740 32496
rect 2044 32419 2096 32428
rect 2044 32385 2053 32419
rect 2053 32385 2087 32419
rect 2087 32385 2096 32419
rect 2044 32376 2096 32385
rect 15200 32444 15252 32496
rect 15936 32512 15988 32564
rect 16764 32555 16816 32564
rect 16764 32521 16773 32555
rect 16773 32521 16807 32555
rect 16807 32521 16816 32555
rect 16764 32512 16816 32521
rect 18512 32512 18564 32564
rect 14096 32376 14148 32428
rect 15384 32419 15436 32428
rect 15384 32385 15393 32419
rect 15393 32385 15427 32419
rect 15427 32385 15436 32419
rect 15384 32376 15436 32385
rect 16856 32419 16908 32428
rect 2964 32308 3016 32360
rect 3056 32351 3108 32360
rect 3056 32317 3065 32351
rect 3065 32317 3099 32351
rect 3099 32317 3108 32351
rect 3056 32308 3108 32317
rect 15568 32308 15620 32360
rect 16856 32385 16865 32419
rect 16865 32385 16899 32419
rect 16899 32385 16908 32419
rect 16856 32376 16908 32385
rect 19156 32419 19208 32428
rect 19156 32385 19165 32419
rect 19165 32385 19199 32419
rect 19199 32385 19208 32419
rect 19156 32376 19208 32385
rect 19432 32419 19484 32428
rect 18052 32308 18104 32360
rect 18696 32308 18748 32360
rect 19432 32385 19441 32419
rect 19441 32385 19475 32419
rect 19475 32385 19484 32419
rect 19432 32376 19484 32385
rect 20628 32444 20680 32496
rect 21548 32444 21600 32496
rect 19892 32419 19944 32428
rect 19892 32385 19901 32419
rect 19901 32385 19935 32419
rect 19935 32385 19944 32419
rect 22652 32512 22704 32564
rect 23020 32512 23072 32564
rect 23848 32555 23900 32564
rect 23848 32521 23857 32555
rect 23857 32521 23891 32555
rect 23891 32521 23900 32555
rect 23848 32512 23900 32521
rect 24124 32512 24176 32564
rect 27620 32512 27672 32564
rect 28080 32512 28132 32564
rect 28540 32512 28592 32564
rect 29368 32555 29420 32564
rect 29368 32521 29377 32555
rect 29377 32521 29411 32555
rect 29411 32521 29420 32555
rect 29368 32512 29420 32521
rect 29736 32512 29788 32564
rect 29920 32512 29972 32564
rect 21732 32444 21784 32496
rect 23756 32444 23808 32496
rect 19892 32376 19944 32385
rect 21916 32376 21968 32428
rect 22560 32376 22612 32428
rect 23020 32419 23072 32428
rect 23020 32385 23029 32419
rect 23029 32385 23063 32419
rect 23063 32385 23072 32419
rect 23020 32376 23072 32385
rect 23204 32419 23256 32428
rect 23204 32385 23213 32419
rect 23213 32385 23247 32419
rect 23247 32385 23256 32419
rect 23204 32376 23256 32385
rect 22468 32351 22520 32360
rect 22468 32317 22477 32351
rect 22477 32317 22511 32351
rect 22511 32317 22520 32351
rect 22468 32308 22520 32317
rect 22836 32308 22888 32360
rect 25780 32444 25832 32496
rect 12164 32172 12216 32224
rect 22376 32240 22428 32292
rect 24308 32419 24360 32428
rect 24308 32385 24317 32419
rect 24317 32385 24351 32419
rect 24351 32385 24360 32419
rect 24308 32376 24360 32385
rect 24492 32419 24544 32428
rect 24492 32385 24501 32419
rect 24501 32385 24535 32419
rect 24535 32385 24544 32419
rect 24492 32376 24544 32385
rect 26424 32376 26476 32428
rect 27344 32419 27396 32428
rect 27344 32385 27353 32419
rect 27353 32385 27387 32419
rect 27387 32385 27396 32419
rect 27344 32376 27396 32385
rect 27712 32419 27764 32428
rect 26884 32308 26936 32360
rect 27712 32385 27721 32419
rect 27721 32385 27755 32419
rect 27755 32385 27764 32419
rect 27712 32376 27764 32385
rect 28356 32308 28408 32360
rect 28724 32419 28776 32428
rect 28724 32385 28733 32419
rect 28733 32385 28767 32419
rect 28767 32385 28776 32419
rect 28724 32376 28776 32385
rect 30748 32444 30800 32496
rect 47676 32419 47728 32428
rect 47676 32385 47685 32419
rect 47685 32385 47719 32419
rect 47719 32385 47728 32419
rect 47676 32376 47728 32385
rect 30196 32308 30248 32360
rect 47492 32308 47544 32360
rect 24308 32240 24360 32292
rect 25780 32240 25832 32292
rect 39212 32240 39264 32292
rect 15200 32172 15252 32224
rect 15476 32215 15528 32224
rect 15476 32181 15485 32215
rect 15485 32181 15519 32215
rect 15519 32181 15528 32215
rect 15476 32172 15528 32181
rect 18788 32215 18840 32224
rect 18788 32181 18797 32215
rect 18797 32181 18831 32215
rect 18831 32181 18840 32215
rect 18788 32172 18840 32181
rect 18880 32172 18932 32224
rect 19892 32172 19944 32224
rect 20904 32215 20956 32224
rect 20904 32181 20913 32215
rect 20913 32181 20947 32215
rect 20947 32181 20956 32215
rect 20904 32172 20956 32181
rect 23756 32172 23808 32224
rect 26148 32172 26200 32224
rect 26884 32172 26936 32224
rect 27620 32172 27672 32224
rect 28172 32172 28224 32224
rect 28724 32172 28776 32224
rect 29460 32172 29512 32224
rect 30288 32172 30340 32224
rect 31760 32172 31812 32224
rect 33048 32172 33100 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 2596 31968 2648 32020
rect 2964 32011 3016 32020
rect 2964 31977 2973 32011
rect 2973 31977 3007 32011
rect 3007 31977 3016 32011
rect 2964 31968 3016 31977
rect 14096 32011 14148 32020
rect 14096 31977 14105 32011
rect 14105 31977 14139 32011
rect 14139 31977 14148 32011
rect 14096 31968 14148 31977
rect 17408 32011 17460 32020
rect 17408 31977 17417 32011
rect 17417 31977 17451 32011
rect 17451 31977 17460 32011
rect 17408 31968 17460 31977
rect 18696 32011 18748 32020
rect 18696 31977 18705 32011
rect 18705 31977 18739 32011
rect 18739 31977 18748 32011
rect 18696 31968 18748 31977
rect 1400 31807 1452 31816
rect 1400 31773 1409 31807
rect 1409 31773 1443 31807
rect 1443 31773 1452 31807
rect 1400 31764 1452 31773
rect 1952 31764 2004 31816
rect 12164 31764 12216 31816
rect 12256 31739 12308 31748
rect 12256 31705 12265 31739
rect 12265 31705 12299 31739
rect 12299 31705 12308 31739
rect 12256 31696 12308 31705
rect 13176 31832 13228 31884
rect 15292 31900 15344 31952
rect 23940 31968 23992 32020
rect 25688 31968 25740 32020
rect 29644 31968 29696 32020
rect 15200 31832 15252 31884
rect 14556 31807 14608 31816
rect 14556 31773 14565 31807
rect 14565 31773 14599 31807
rect 14599 31773 14608 31807
rect 14556 31764 14608 31773
rect 17132 31764 17184 31816
rect 18052 31764 18104 31816
rect 22928 31900 22980 31952
rect 19248 31875 19300 31884
rect 19248 31841 19257 31875
rect 19257 31841 19291 31875
rect 19291 31841 19300 31875
rect 19248 31832 19300 31841
rect 21824 31832 21876 31884
rect 18788 31764 18840 31816
rect 21916 31764 21968 31816
rect 11520 31628 11572 31680
rect 15844 31696 15896 31748
rect 18880 31696 18932 31748
rect 12624 31671 12676 31680
rect 12624 31637 12633 31671
rect 12633 31637 12667 31671
rect 12667 31637 12676 31671
rect 12624 31628 12676 31637
rect 15568 31628 15620 31680
rect 19432 31628 19484 31680
rect 21272 31628 21324 31680
rect 21456 31628 21508 31680
rect 22560 31801 22612 31810
rect 22560 31767 22569 31801
rect 22569 31767 22603 31801
rect 22603 31767 22612 31801
rect 22744 31807 22796 31816
rect 22560 31758 22612 31767
rect 22744 31773 22753 31807
rect 22753 31773 22787 31807
rect 22787 31773 22796 31807
rect 22744 31764 22796 31773
rect 23480 31807 23532 31816
rect 23480 31773 23489 31807
rect 23489 31773 23523 31807
rect 23523 31773 23532 31807
rect 23480 31764 23532 31773
rect 22836 31696 22888 31748
rect 23756 31764 23808 31816
rect 29552 31900 29604 31952
rect 28540 31832 28592 31884
rect 28908 31832 28960 31884
rect 26884 31764 26936 31816
rect 22376 31628 22428 31680
rect 22468 31628 22520 31680
rect 22744 31628 22796 31680
rect 27528 31696 27580 31748
rect 29368 31696 29420 31748
rect 29644 31764 29696 31816
rect 31760 31943 31812 31952
rect 31760 31909 31769 31943
rect 31769 31909 31803 31943
rect 31803 31909 31812 31943
rect 31760 31900 31812 31909
rect 30288 31832 30340 31884
rect 30196 31807 30248 31816
rect 30196 31773 30205 31807
rect 30205 31773 30239 31807
rect 30239 31773 30248 31807
rect 30196 31764 30248 31773
rect 45928 31832 45980 31884
rect 32496 31764 32548 31816
rect 26240 31628 26292 31680
rect 27436 31628 27488 31680
rect 29828 31628 29880 31680
rect 30380 31696 30432 31748
rect 30748 31696 30800 31748
rect 32404 31696 32456 31748
rect 32772 31807 32824 31816
rect 32772 31773 32781 31807
rect 32781 31773 32815 31807
rect 32815 31773 32824 31807
rect 32772 31764 32824 31773
rect 33508 31764 33560 31816
rect 47308 31807 47360 31816
rect 47308 31773 47317 31807
rect 47317 31773 47351 31807
rect 47351 31773 47360 31807
rect 47308 31764 47360 31773
rect 33324 31628 33376 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 4804 31424 4856 31476
rect 13176 31467 13228 31476
rect 1952 31331 2004 31340
rect 1952 31297 1961 31331
rect 1961 31297 1995 31331
rect 1995 31297 2004 31331
rect 1952 31288 2004 31297
rect 2872 31220 2924 31272
rect 3056 31263 3108 31272
rect 3056 31229 3065 31263
rect 3065 31229 3099 31263
rect 3099 31229 3108 31263
rect 3056 31220 3108 31229
rect 8484 31220 8536 31272
rect 11520 31356 11572 31408
rect 10324 31288 10376 31340
rect 11888 31288 11940 31340
rect 13176 31433 13185 31467
rect 13185 31433 13219 31467
rect 13219 31433 13228 31467
rect 13176 31424 13228 31433
rect 14096 31424 14148 31476
rect 15384 31424 15436 31476
rect 15936 31424 15988 31476
rect 16856 31424 16908 31476
rect 18880 31424 18932 31476
rect 12256 31356 12308 31408
rect 14372 31356 14424 31408
rect 15292 31356 15344 31408
rect 16212 31356 16264 31408
rect 21548 31424 21600 31476
rect 23940 31399 23992 31408
rect 13360 31288 13412 31340
rect 15568 31288 15620 31340
rect 15752 31288 15804 31340
rect 16120 31331 16172 31340
rect 16120 31297 16129 31331
rect 16129 31297 16163 31331
rect 16163 31297 16172 31331
rect 16120 31288 16172 31297
rect 15384 31263 15436 31272
rect 15384 31229 15393 31263
rect 15393 31229 15427 31263
rect 15427 31229 15436 31263
rect 15384 31220 15436 31229
rect 18052 31288 18104 31340
rect 20812 31288 20864 31340
rect 14556 31152 14608 31204
rect 15844 31195 15896 31204
rect 15844 31161 15853 31195
rect 15853 31161 15887 31195
rect 15887 31161 15896 31195
rect 15844 31152 15896 31161
rect 15936 31152 15988 31204
rect 20352 31220 20404 31272
rect 20076 31152 20128 31204
rect 21088 31331 21140 31340
rect 21088 31297 21097 31331
rect 21097 31297 21131 31331
rect 21131 31297 21140 31331
rect 21272 31331 21324 31340
rect 21088 31288 21140 31297
rect 21272 31297 21281 31331
rect 21281 31297 21315 31331
rect 21315 31297 21324 31331
rect 21272 31288 21324 31297
rect 23940 31365 23974 31399
rect 23974 31365 23992 31399
rect 23940 31356 23992 31365
rect 28632 31424 28684 31476
rect 30380 31424 30432 31476
rect 30840 31424 30892 31476
rect 32772 31424 32824 31476
rect 32496 31356 32548 31408
rect 33324 31399 33376 31408
rect 33324 31365 33358 31399
rect 33358 31365 33376 31399
rect 33324 31356 33376 31365
rect 22928 31288 22980 31340
rect 26148 31331 26200 31340
rect 26148 31297 26157 31331
rect 26157 31297 26191 31331
rect 26191 31297 26200 31331
rect 26148 31288 26200 31297
rect 26240 31331 26292 31340
rect 26240 31297 26249 31331
rect 26249 31297 26283 31331
rect 26283 31297 26292 31331
rect 26240 31288 26292 31297
rect 27712 31288 27764 31340
rect 28264 31288 28316 31340
rect 28540 31288 28592 31340
rect 28724 31288 28776 31340
rect 30012 31288 30064 31340
rect 30748 31288 30800 31340
rect 31944 31288 31996 31340
rect 32220 31331 32272 31340
rect 21456 31152 21508 31204
rect 26976 31220 27028 31272
rect 27252 31263 27304 31272
rect 27252 31229 27261 31263
rect 27261 31229 27295 31263
rect 27295 31229 27304 31263
rect 27252 31220 27304 31229
rect 27528 31263 27580 31272
rect 27528 31229 27537 31263
rect 27537 31229 27571 31263
rect 27571 31229 27580 31263
rect 27528 31220 27580 31229
rect 30840 31263 30892 31272
rect 25044 31195 25096 31204
rect 10140 31084 10192 31136
rect 15476 31084 15528 31136
rect 18420 31084 18472 31136
rect 20904 31084 20956 31136
rect 21824 31084 21876 31136
rect 25044 31161 25053 31195
rect 25053 31161 25087 31195
rect 25087 31161 25096 31195
rect 25044 31152 25096 31161
rect 27344 31152 27396 31204
rect 28908 31152 28960 31204
rect 30840 31229 30849 31263
rect 30849 31229 30883 31263
rect 30883 31229 30892 31263
rect 30840 31220 30892 31229
rect 32220 31297 32229 31331
rect 32229 31297 32263 31331
rect 32263 31297 32272 31331
rect 32220 31288 32272 31297
rect 33048 31331 33100 31340
rect 33048 31297 33057 31331
rect 33057 31297 33091 31331
rect 33091 31297 33100 31331
rect 33048 31288 33100 31297
rect 25780 31127 25832 31136
rect 25780 31093 25789 31127
rect 25789 31093 25823 31127
rect 25823 31093 25832 31127
rect 25780 31084 25832 31093
rect 28172 31084 28224 31136
rect 33416 31084 33468 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 2872 30923 2924 30932
rect 2872 30889 2881 30923
rect 2881 30889 2915 30923
rect 2915 30889 2924 30923
rect 2872 30880 2924 30889
rect 10324 30880 10376 30932
rect 11888 30880 11940 30932
rect 16120 30880 16172 30932
rect 21088 30880 21140 30932
rect 22560 30923 22612 30932
rect 22560 30889 22569 30923
rect 22569 30889 22603 30923
rect 22603 30889 22612 30923
rect 22560 30880 22612 30889
rect 23664 30880 23716 30932
rect 28356 30880 28408 30932
rect 32220 30880 32272 30932
rect 1768 30676 1820 30728
rect 12164 30812 12216 30864
rect 13268 30812 13320 30864
rect 19524 30812 19576 30864
rect 10416 30676 10468 30728
rect 10784 30719 10836 30728
rect 10784 30685 10793 30719
rect 10793 30685 10827 30719
rect 10827 30685 10836 30719
rect 10784 30676 10836 30685
rect 9680 30608 9732 30660
rect 10048 30608 10100 30660
rect 10876 30540 10928 30592
rect 11152 30676 11204 30728
rect 13360 30744 13412 30796
rect 12440 30719 12492 30728
rect 12440 30685 12449 30719
rect 12449 30685 12483 30719
rect 12483 30685 12492 30719
rect 12440 30676 12492 30685
rect 13268 30719 13320 30728
rect 13268 30685 13277 30719
rect 13277 30685 13311 30719
rect 13311 30685 13320 30719
rect 13268 30676 13320 30685
rect 14096 30719 14148 30728
rect 14096 30685 14105 30719
rect 14105 30685 14139 30719
rect 14139 30685 14148 30719
rect 14096 30676 14148 30685
rect 15476 30676 15528 30728
rect 21456 30812 21508 30864
rect 23112 30744 23164 30796
rect 27528 30812 27580 30864
rect 20352 30719 20404 30728
rect 12624 30608 12676 30660
rect 15936 30651 15988 30660
rect 15936 30617 15945 30651
rect 15945 30617 15979 30651
rect 15979 30617 15988 30651
rect 15936 30608 15988 30617
rect 17408 30608 17460 30660
rect 19432 30608 19484 30660
rect 20352 30685 20361 30719
rect 20361 30685 20395 30719
rect 20395 30685 20404 30719
rect 20352 30676 20404 30685
rect 20536 30651 20588 30660
rect 20536 30617 20545 30651
rect 20545 30617 20579 30651
rect 20579 30617 20588 30651
rect 20536 30608 20588 30617
rect 22652 30676 22704 30728
rect 22744 30676 22796 30728
rect 23664 30676 23716 30728
rect 27068 30676 27120 30728
rect 27528 30676 27580 30728
rect 28172 30719 28224 30728
rect 28172 30685 28181 30719
rect 28181 30685 28215 30719
rect 28215 30685 28224 30719
rect 28172 30676 28224 30685
rect 30840 30744 30892 30796
rect 29736 30719 29788 30728
rect 29736 30685 29745 30719
rect 29745 30685 29779 30719
rect 29779 30685 29788 30719
rect 29736 30676 29788 30685
rect 29828 30676 29880 30728
rect 31944 30676 31996 30728
rect 33232 30676 33284 30728
rect 20720 30608 20772 30660
rect 20812 30608 20864 30660
rect 21272 30608 21324 30660
rect 21548 30651 21600 30660
rect 21548 30617 21557 30651
rect 21557 30617 21591 30651
rect 21591 30617 21600 30651
rect 21548 30608 21600 30617
rect 25044 30608 25096 30660
rect 25780 30608 25832 30660
rect 12440 30540 12492 30592
rect 17592 30540 17644 30592
rect 19340 30540 19392 30592
rect 20076 30540 20128 30592
rect 23572 30540 23624 30592
rect 27160 30540 27212 30592
rect 27436 30540 27488 30592
rect 30012 30540 30064 30592
rect 32956 30608 33008 30660
rect 33140 30540 33192 30592
rect 33416 30540 33468 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 15936 30336 15988 30388
rect 9680 30268 9732 30320
rect 12256 30268 12308 30320
rect 17132 30268 17184 30320
rect 18420 30311 18472 30320
rect 18420 30277 18429 30311
rect 18429 30277 18463 30311
rect 18463 30277 18472 30311
rect 18420 30268 18472 30277
rect 19340 30311 19392 30320
rect 19340 30277 19374 30311
rect 19374 30277 19392 30311
rect 19340 30268 19392 30277
rect 23112 30268 23164 30320
rect 27528 30336 27580 30388
rect 29736 30336 29788 30388
rect 29460 30311 29512 30320
rect 1768 30243 1820 30252
rect 1768 30209 1777 30243
rect 1777 30209 1811 30243
rect 1811 30209 1820 30243
rect 1768 30200 1820 30209
rect 4804 30243 4856 30252
rect 4804 30209 4813 30243
rect 4813 30209 4847 30243
rect 4847 30209 4856 30243
rect 4804 30200 4856 30209
rect 10232 30200 10284 30252
rect 10600 30243 10652 30252
rect 10600 30209 10609 30243
rect 10609 30209 10643 30243
rect 10643 30209 10652 30243
rect 10600 30200 10652 30209
rect 10784 30200 10836 30252
rect 16028 30200 16080 30252
rect 16304 30200 16356 30252
rect 2136 30132 2188 30184
rect 2780 30175 2832 30184
rect 2780 30141 2789 30175
rect 2789 30141 2823 30175
rect 2823 30141 2832 30175
rect 2780 30132 2832 30141
rect 7748 30132 7800 30184
rect 8484 30175 8536 30184
rect 8484 30141 8493 30175
rect 8493 30141 8527 30175
rect 8527 30141 8536 30175
rect 8484 30132 8536 30141
rect 17776 30200 17828 30252
rect 4068 30064 4120 30116
rect 12440 30064 12492 30116
rect 17776 30064 17828 30116
rect 18604 30107 18656 30116
rect 18604 30073 18613 30107
rect 18613 30073 18647 30107
rect 18647 30073 18656 30107
rect 18604 30064 18656 30073
rect 10600 29996 10652 30048
rect 10692 29996 10744 30048
rect 21364 30200 21416 30252
rect 27344 30200 27396 30252
rect 27620 30200 27672 30252
rect 29460 30277 29469 30311
rect 29469 30277 29503 30311
rect 29503 30277 29512 30311
rect 29460 30268 29512 30277
rect 45468 30336 45520 30388
rect 27528 30175 27580 30184
rect 27528 30141 27537 30175
rect 27537 30141 27571 30175
rect 27571 30141 27580 30175
rect 27528 30132 27580 30141
rect 20076 29996 20128 30048
rect 20536 30064 20588 30116
rect 32956 30243 33008 30252
rect 32956 30209 32965 30243
rect 32965 30209 32999 30243
rect 32999 30209 33008 30243
rect 32956 30200 33008 30209
rect 33508 30200 33560 30252
rect 47952 30243 48004 30252
rect 47952 30209 47961 30243
rect 47961 30209 47995 30243
rect 47995 30209 48004 30243
rect 47952 30200 48004 30209
rect 33048 30132 33100 30184
rect 33600 30175 33652 30184
rect 33600 30141 33609 30175
rect 33609 30141 33643 30175
rect 33643 30141 33652 30175
rect 33600 30132 33652 30141
rect 20628 29996 20680 30048
rect 22008 29996 22060 30048
rect 25596 29996 25648 30048
rect 32404 30064 32456 30116
rect 32864 30064 32916 30116
rect 28724 29996 28776 30048
rect 34612 29996 34664 30048
rect 48044 30039 48096 30048
rect 48044 30005 48053 30039
rect 48053 30005 48087 30039
rect 48087 30005 48096 30039
rect 48044 29996 48096 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 2136 29835 2188 29844
rect 2136 29801 2145 29835
rect 2145 29801 2179 29835
rect 2179 29801 2188 29835
rect 2136 29792 2188 29801
rect 10232 29835 10284 29844
rect 10232 29801 10241 29835
rect 10241 29801 10275 29835
rect 10275 29801 10284 29835
rect 10232 29792 10284 29801
rect 10508 29792 10560 29844
rect 2688 29724 2740 29776
rect 20352 29792 20404 29844
rect 20904 29792 20956 29844
rect 32404 29792 32456 29844
rect 33140 29792 33192 29844
rect 13728 29724 13780 29776
rect 1768 29588 1820 29640
rect 9128 29631 9180 29640
rect 9128 29597 9137 29631
rect 9137 29597 9171 29631
rect 9171 29597 9180 29631
rect 9128 29588 9180 29597
rect 10508 29631 10560 29640
rect 10508 29597 10517 29631
rect 10517 29597 10551 29631
rect 10551 29597 10560 29631
rect 10508 29588 10560 29597
rect 10784 29656 10836 29708
rect 12440 29699 12492 29708
rect 12440 29665 12449 29699
rect 12449 29665 12483 29699
rect 12483 29665 12492 29699
rect 16304 29699 16356 29708
rect 12440 29656 12492 29665
rect 16304 29665 16313 29699
rect 16313 29665 16347 29699
rect 16347 29665 16356 29699
rect 16304 29656 16356 29665
rect 17224 29656 17276 29708
rect 22008 29656 22060 29708
rect 10692 29631 10744 29640
rect 10692 29597 10701 29631
rect 10701 29597 10735 29631
rect 10735 29597 10744 29631
rect 10692 29588 10744 29597
rect 10876 29631 10928 29640
rect 10876 29597 10885 29631
rect 10885 29597 10919 29631
rect 10919 29597 10928 29631
rect 10876 29588 10928 29597
rect 14372 29631 14424 29640
rect 11704 29520 11756 29572
rect 12256 29563 12308 29572
rect 12256 29529 12265 29563
rect 12265 29529 12299 29563
rect 12299 29529 12308 29563
rect 12256 29520 12308 29529
rect 14372 29597 14381 29631
rect 14381 29597 14415 29631
rect 14415 29597 14424 29631
rect 14372 29588 14424 29597
rect 15384 29588 15436 29640
rect 16028 29588 16080 29640
rect 17776 29588 17828 29640
rect 18604 29588 18656 29640
rect 20720 29631 20772 29640
rect 20720 29597 20729 29631
rect 20729 29597 20763 29631
rect 20763 29597 20772 29631
rect 20720 29588 20772 29597
rect 20904 29631 20956 29640
rect 20904 29597 20913 29631
rect 20913 29597 20947 29631
rect 20947 29597 20956 29631
rect 20904 29588 20956 29597
rect 1952 29452 2004 29504
rect 8944 29495 8996 29504
rect 8944 29461 8953 29495
rect 8953 29461 8987 29495
rect 8987 29461 8996 29495
rect 8944 29452 8996 29461
rect 10232 29452 10284 29504
rect 10416 29452 10468 29504
rect 13636 29452 13688 29504
rect 14372 29452 14424 29504
rect 14556 29495 14608 29504
rect 14556 29461 14565 29495
rect 14565 29461 14599 29495
rect 14599 29461 14608 29495
rect 14556 29452 14608 29461
rect 16764 29452 16816 29504
rect 19340 29520 19392 29572
rect 23112 29656 23164 29708
rect 23480 29588 23532 29640
rect 48044 29724 48096 29776
rect 24952 29656 25004 29708
rect 27252 29656 27304 29708
rect 32680 29656 32732 29708
rect 24860 29631 24912 29640
rect 24860 29597 24869 29631
rect 24869 29597 24903 29631
rect 24903 29597 24912 29631
rect 24860 29588 24912 29597
rect 25136 29588 25188 29640
rect 25596 29631 25648 29640
rect 25596 29597 25605 29631
rect 25605 29597 25639 29631
rect 25639 29597 25648 29631
rect 25596 29588 25648 29597
rect 28172 29588 28224 29640
rect 28908 29588 28960 29640
rect 33784 29656 33836 29708
rect 33968 29699 34020 29708
rect 33968 29665 33977 29699
rect 33977 29665 34011 29699
rect 34011 29665 34020 29699
rect 38016 29699 38068 29708
rect 33968 29656 34020 29665
rect 38016 29665 38025 29699
rect 38025 29665 38059 29699
rect 38059 29665 38068 29699
rect 38016 29656 38068 29665
rect 18328 29495 18380 29504
rect 18328 29461 18337 29495
rect 18337 29461 18371 29495
rect 18371 29461 18380 29495
rect 18328 29452 18380 29461
rect 20076 29452 20128 29504
rect 20812 29452 20864 29504
rect 28356 29520 28408 29572
rect 31208 29563 31260 29572
rect 31208 29529 31217 29563
rect 31217 29529 31251 29563
rect 31251 29529 31260 29563
rect 31208 29520 31260 29529
rect 33324 29520 33376 29572
rect 36452 29520 36504 29572
rect 22928 29452 22980 29504
rect 24400 29495 24452 29504
rect 24400 29461 24409 29495
rect 24409 29461 24443 29495
rect 24443 29461 24452 29495
rect 24400 29452 24452 29461
rect 24584 29452 24636 29504
rect 24768 29452 24820 29504
rect 25044 29452 25096 29504
rect 31484 29452 31536 29504
rect 33048 29452 33100 29504
rect 34612 29452 34664 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 1952 29223 2004 29232
rect 1952 29189 1961 29223
rect 1961 29189 1995 29223
rect 1995 29189 2004 29223
rect 1952 29180 2004 29189
rect 8944 29180 8996 29232
rect 10232 29248 10284 29300
rect 13728 29291 13780 29300
rect 13728 29257 13737 29291
rect 13737 29257 13771 29291
rect 13771 29257 13780 29291
rect 13728 29248 13780 29257
rect 18144 29248 18196 29300
rect 19340 29248 19392 29300
rect 24860 29248 24912 29300
rect 9864 29223 9916 29232
rect 9864 29189 9889 29223
rect 9889 29189 9916 29223
rect 15476 29223 15528 29232
rect 9864 29180 9916 29189
rect 15476 29189 15485 29223
rect 15485 29189 15519 29223
rect 15519 29189 15528 29223
rect 15476 29180 15528 29189
rect 1768 29155 1820 29164
rect 1768 29121 1777 29155
rect 1777 29121 1811 29155
rect 1811 29121 1820 29155
rect 1768 29112 1820 29121
rect 4068 29112 4120 29164
rect 11520 29155 11572 29164
rect 11520 29121 11529 29155
rect 11529 29121 11563 29155
rect 11563 29121 11572 29155
rect 11520 29112 11572 29121
rect 11612 29112 11664 29164
rect 12900 29112 12952 29164
rect 13636 29155 13688 29164
rect 13636 29121 13645 29155
rect 13645 29121 13679 29155
rect 13679 29121 13688 29155
rect 13636 29112 13688 29121
rect 14372 29155 14424 29164
rect 14372 29121 14381 29155
rect 14381 29121 14415 29155
rect 14415 29121 14424 29155
rect 14372 29112 14424 29121
rect 15752 29155 15804 29164
rect 15752 29121 15761 29155
rect 15761 29121 15795 29155
rect 15795 29121 15804 29155
rect 15752 29112 15804 29121
rect 16580 29180 16632 29232
rect 16948 29155 17000 29164
rect 16948 29121 16982 29155
rect 16982 29121 17000 29155
rect 3332 29087 3384 29096
rect 3332 29053 3341 29087
rect 3341 29053 3375 29087
rect 3375 29053 3384 29087
rect 3332 29044 3384 29053
rect 7748 29044 7800 29096
rect 9680 29044 9732 29096
rect 16028 29044 16080 29096
rect 8852 28976 8904 29028
rect 1400 28908 1452 28960
rect 9772 28908 9824 28960
rect 10508 28908 10560 28960
rect 12532 28908 12584 28960
rect 13360 28908 13412 28960
rect 15660 28908 15712 28960
rect 16028 28908 16080 28960
rect 16948 29112 17000 29121
rect 20076 29180 20128 29232
rect 24400 29180 24452 29232
rect 18604 29112 18656 29164
rect 20352 29112 20404 29164
rect 20812 29155 20864 29164
rect 20812 29121 20821 29155
rect 20821 29121 20855 29155
rect 20855 29121 20864 29155
rect 20812 29112 20864 29121
rect 20996 29155 21048 29164
rect 20996 29121 21005 29155
rect 21005 29121 21039 29155
rect 21039 29121 21048 29155
rect 20996 29112 21048 29121
rect 22008 29112 22060 29164
rect 22189 29158 22241 29167
rect 22189 29124 22198 29158
rect 22198 29124 22232 29158
rect 22232 29124 22241 29158
rect 22189 29115 22241 29124
rect 22284 29155 22336 29164
rect 22284 29121 22298 29155
rect 22298 29121 22332 29155
rect 22332 29121 22336 29155
rect 22284 29112 22336 29121
rect 22560 29112 22612 29164
rect 22928 29112 22980 29164
rect 27620 29180 27672 29232
rect 28080 29180 28132 29232
rect 28356 29248 28408 29300
rect 32680 29248 32732 29300
rect 36452 29291 36504 29300
rect 36452 29257 36461 29291
rect 36461 29257 36495 29291
rect 36495 29257 36504 29291
rect 36452 29248 36504 29257
rect 47308 29248 47360 29300
rect 47492 29248 47544 29300
rect 27344 29155 27396 29164
rect 27344 29121 27353 29155
rect 27353 29121 27387 29155
rect 27387 29121 27396 29155
rect 27344 29112 27396 29121
rect 27988 29155 28040 29164
rect 27988 29121 27997 29155
rect 27997 29121 28031 29155
rect 28031 29121 28040 29155
rect 27988 29112 28040 29121
rect 30196 29180 30248 29232
rect 32496 29223 32548 29232
rect 32496 29189 32505 29223
rect 32505 29189 32539 29223
rect 32539 29189 32548 29223
rect 32496 29180 32548 29189
rect 33048 29180 33100 29232
rect 24492 29087 24544 29096
rect 17316 28908 17368 28960
rect 18052 28908 18104 28960
rect 21180 28976 21232 29028
rect 20352 28951 20404 28960
rect 20352 28917 20361 28951
rect 20361 28917 20395 28951
rect 20395 28917 20404 28951
rect 20352 28908 20404 28917
rect 24492 29053 24501 29087
rect 24501 29053 24535 29087
rect 24535 29053 24544 29087
rect 24492 29044 24544 29053
rect 22100 28976 22152 29028
rect 28172 28976 28224 29028
rect 28356 29019 28408 29028
rect 28356 28985 28365 29019
rect 28365 28985 28399 29019
rect 28399 28985 28408 29019
rect 28356 28976 28408 28985
rect 21456 28908 21508 28960
rect 24860 28908 24912 28960
rect 28080 28908 28132 28960
rect 30748 28951 30800 28960
rect 30748 28917 30757 28951
rect 30757 28917 30791 28951
rect 30791 28917 30800 28951
rect 30748 28908 30800 28917
rect 31116 28976 31168 29028
rect 31760 29112 31812 29164
rect 32404 29112 32456 29164
rect 32864 29155 32916 29164
rect 32864 29121 32873 29155
rect 32873 29121 32907 29155
rect 32907 29121 32916 29155
rect 32864 29112 32916 29121
rect 33508 29112 33560 29164
rect 33600 29112 33652 29164
rect 33784 29112 33836 29164
rect 36360 29155 36412 29164
rect 36360 29121 36369 29155
rect 36369 29121 36403 29155
rect 36403 29121 36412 29155
rect 36360 29112 36412 29121
rect 46296 29112 46348 29164
rect 32496 29044 32548 29096
rect 47492 29044 47544 29096
rect 47768 29044 47820 29096
rect 35532 28976 35584 29028
rect 47676 28951 47728 28960
rect 47676 28917 47685 28951
rect 47685 28917 47719 28951
rect 47719 28917 47728 28951
rect 47676 28908 47728 28917
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 8300 28704 8352 28756
rect 9128 28704 9180 28756
rect 11612 28704 11664 28756
rect 15660 28747 15712 28756
rect 15660 28713 15669 28747
rect 15669 28713 15703 28747
rect 15703 28713 15712 28747
rect 15660 28704 15712 28713
rect 8852 28636 8904 28688
rect 1400 28611 1452 28620
rect 1400 28577 1409 28611
rect 1409 28577 1443 28611
rect 1443 28577 1452 28611
rect 1400 28568 1452 28577
rect 2780 28611 2832 28620
rect 2780 28577 2789 28611
rect 2789 28577 2823 28611
rect 2823 28577 2832 28611
rect 2780 28568 2832 28577
rect 2320 28432 2372 28484
rect 9772 28611 9824 28620
rect 9772 28577 9781 28611
rect 9781 28577 9815 28611
rect 9815 28577 9824 28611
rect 9772 28568 9824 28577
rect 13360 28568 13412 28620
rect 14004 28568 14056 28620
rect 18604 28704 18656 28756
rect 20904 28704 20956 28756
rect 27988 28704 28040 28756
rect 31208 28704 31260 28756
rect 33324 28704 33376 28756
rect 17776 28636 17828 28688
rect 10232 28500 10284 28552
rect 11520 28543 11572 28552
rect 11520 28509 11529 28543
rect 11529 28509 11563 28543
rect 11563 28509 11572 28543
rect 11520 28500 11572 28509
rect 12256 28543 12308 28552
rect 12256 28509 12265 28543
rect 12265 28509 12299 28543
rect 12299 28509 12308 28543
rect 12256 28500 12308 28509
rect 10968 28432 11020 28484
rect 12532 28500 12584 28552
rect 14280 28543 14332 28552
rect 12716 28432 12768 28484
rect 12992 28432 13044 28484
rect 14280 28509 14289 28543
rect 14289 28509 14323 28543
rect 14323 28509 14332 28543
rect 14280 28500 14332 28509
rect 15752 28500 15804 28552
rect 18328 28568 18380 28620
rect 21824 28611 21876 28620
rect 21824 28577 21833 28611
rect 21833 28577 21867 28611
rect 21867 28577 21876 28611
rect 21824 28568 21876 28577
rect 24492 28568 24544 28620
rect 28724 28611 28776 28620
rect 28724 28577 28733 28611
rect 28733 28577 28767 28611
rect 28767 28577 28776 28611
rect 28724 28568 28776 28577
rect 31392 28568 31444 28620
rect 33968 28611 34020 28620
rect 33968 28577 33977 28611
rect 33977 28577 34011 28611
rect 34011 28577 34020 28611
rect 33968 28568 34020 28577
rect 47676 28568 47728 28620
rect 48136 28611 48188 28620
rect 48136 28577 48145 28611
rect 48145 28577 48179 28611
rect 48179 28577 48188 28611
rect 48136 28568 48188 28577
rect 18052 28543 18104 28552
rect 14648 28432 14700 28484
rect 14740 28432 14792 28484
rect 18052 28509 18061 28543
rect 18061 28509 18095 28543
rect 18095 28509 18104 28543
rect 18052 28500 18104 28509
rect 20076 28500 20128 28552
rect 22100 28543 22152 28552
rect 22100 28509 22134 28543
rect 22134 28509 22152 28543
rect 22100 28500 22152 28509
rect 27620 28500 27672 28552
rect 28816 28500 28868 28552
rect 33784 28500 33836 28552
rect 34428 28500 34480 28552
rect 20352 28432 20404 28484
rect 24584 28432 24636 28484
rect 32588 28432 32640 28484
rect 47676 28432 47728 28484
rect 9956 28364 10008 28416
rect 11980 28407 12032 28416
rect 11980 28373 11989 28407
rect 11989 28373 12023 28407
rect 12023 28373 12032 28407
rect 11980 28364 12032 28373
rect 12440 28364 12492 28416
rect 23480 28364 23532 28416
rect 26056 28407 26108 28416
rect 26056 28373 26065 28407
rect 26065 28373 26099 28407
rect 26099 28373 26108 28407
rect 26056 28364 26108 28373
rect 27436 28407 27488 28416
rect 27436 28373 27445 28407
rect 27445 28373 27479 28407
rect 27479 28373 27488 28407
rect 27436 28364 27488 28373
rect 28632 28407 28684 28416
rect 28632 28373 28641 28407
rect 28641 28373 28675 28407
rect 28675 28373 28684 28407
rect 28632 28364 28684 28373
rect 29828 28407 29880 28416
rect 29828 28373 29837 28407
rect 29837 28373 29871 28407
rect 29871 28373 29880 28407
rect 29828 28364 29880 28373
rect 31576 28364 31628 28416
rect 35532 28364 35584 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 2320 28203 2372 28212
rect 2320 28169 2329 28203
rect 2329 28169 2363 28203
rect 2363 28169 2372 28203
rect 2320 28160 2372 28169
rect 8300 28160 8352 28212
rect 11520 28160 11572 28212
rect 12256 28160 12308 28212
rect 12992 28203 13044 28212
rect 12992 28169 13001 28203
rect 13001 28169 13035 28203
rect 13035 28169 13044 28203
rect 12992 28160 13044 28169
rect 14372 28160 14424 28212
rect 14648 28203 14700 28212
rect 14648 28169 14657 28203
rect 14657 28169 14691 28203
rect 14691 28169 14700 28203
rect 14648 28160 14700 28169
rect 16580 28160 16632 28212
rect 22284 28160 22336 28212
rect 24584 28160 24636 28212
rect 33784 28160 33836 28212
rect 11888 28092 11940 28144
rect 3516 28024 3568 28076
rect 8300 28024 8352 28076
rect 9772 28024 9824 28076
rect 9864 28024 9916 28076
rect 9312 27956 9364 28008
rect 12716 28024 12768 28076
rect 12992 28024 13044 28076
rect 14096 28092 14148 28144
rect 16764 28092 16816 28144
rect 18144 28092 18196 28144
rect 20996 28092 21048 28144
rect 14004 28067 14056 28076
rect 14004 28033 14013 28067
rect 14013 28033 14047 28067
rect 14047 28033 14056 28067
rect 14004 28024 14056 28033
rect 22192 28067 22244 28076
rect 12164 27956 12216 28008
rect 22192 28033 22201 28067
rect 22201 28033 22235 28067
rect 22235 28033 22244 28067
rect 22192 28024 22244 28033
rect 22284 28067 22336 28076
rect 22284 28033 22293 28067
rect 22293 28033 22327 28067
rect 22327 28033 22336 28067
rect 22560 28092 22612 28144
rect 22284 28024 22336 28033
rect 22928 28067 22980 28076
rect 22928 28033 22937 28067
rect 22937 28033 22971 28067
rect 22971 28033 22980 28067
rect 22928 28024 22980 28033
rect 23480 28024 23532 28076
rect 24400 28024 24452 28076
rect 24860 28067 24912 28076
rect 24860 28033 24869 28067
rect 24869 28033 24903 28067
rect 24903 28033 24912 28067
rect 24860 28024 24912 28033
rect 24952 28067 25004 28076
rect 24952 28033 24961 28067
rect 24961 28033 24995 28067
rect 24995 28033 25004 28067
rect 24952 28024 25004 28033
rect 25136 28067 25188 28076
rect 25136 28033 25145 28067
rect 25145 28033 25179 28067
rect 25179 28033 25188 28067
rect 25136 28024 25188 28033
rect 27620 28024 27672 28076
rect 32496 28092 32548 28144
rect 30748 28024 30800 28076
rect 31944 28024 31996 28076
rect 47952 28067 48004 28076
rect 47952 28033 47961 28067
rect 47961 28033 47995 28067
rect 47995 28033 48004 28067
rect 47952 28024 48004 28033
rect 22836 27956 22888 28008
rect 27528 27956 27580 28008
rect 32496 27999 32548 28008
rect 12532 27888 12584 27940
rect 20260 27888 20312 27940
rect 25780 27888 25832 27940
rect 7288 27820 7340 27872
rect 8760 27863 8812 27872
rect 8760 27829 8769 27863
rect 8769 27829 8803 27863
rect 8803 27829 8812 27863
rect 8760 27820 8812 27829
rect 9680 27820 9732 27872
rect 11980 27863 12032 27872
rect 11980 27829 11989 27863
rect 11989 27829 12023 27863
rect 12023 27829 12032 27863
rect 11980 27820 12032 27829
rect 22100 27820 22152 27872
rect 32496 27965 32505 27999
rect 32505 27965 32539 27999
rect 32539 27965 32548 27999
rect 32496 27956 32548 27965
rect 27896 27820 27948 27872
rect 28632 27820 28684 27872
rect 31576 27863 31628 27872
rect 31576 27829 31585 27863
rect 31585 27829 31619 27863
rect 31619 27829 31628 27863
rect 31576 27820 31628 27829
rect 32404 27820 32456 27872
rect 32772 27820 32824 27872
rect 44180 27820 44232 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 9864 27659 9916 27668
rect 9864 27625 9873 27659
rect 9873 27625 9907 27659
rect 9907 27625 9916 27659
rect 9864 27616 9916 27625
rect 12716 27659 12768 27668
rect 12716 27625 12725 27659
rect 12725 27625 12759 27659
rect 12759 27625 12768 27659
rect 12716 27616 12768 27625
rect 24952 27659 25004 27668
rect 24952 27625 24961 27659
rect 24961 27625 24995 27659
rect 24995 27625 25004 27659
rect 24952 27616 25004 27625
rect 10968 27548 11020 27600
rect 12900 27591 12952 27600
rect 9036 27480 9088 27532
rect 1400 27412 1452 27464
rect 2044 27455 2096 27464
rect 2044 27421 2053 27455
rect 2053 27421 2087 27455
rect 2087 27421 2096 27455
rect 2044 27412 2096 27421
rect 2320 27412 2372 27464
rect 1768 27344 1820 27396
rect 7748 27412 7800 27464
rect 7288 27387 7340 27396
rect 7288 27353 7322 27387
rect 7322 27353 7340 27387
rect 7288 27344 7340 27353
rect 9956 27412 10008 27464
rect 10876 27412 10928 27464
rect 10416 27344 10468 27396
rect 10968 27344 11020 27396
rect 1952 27276 2004 27328
rect 9312 27276 9364 27328
rect 10692 27319 10744 27328
rect 10692 27285 10701 27319
rect 10701 27285 10735 27319
rect 10735 27285 10744 27319
rect 10692 27276 10744 27285
rect 12900 27557 12909 27591
rect 12909 27557 12943 27591
rect 12943 27557 12952 27591
rect 12900 27548 12952 27557
rect 14280 27548 14332 27600
rect 17132 27548 17184 27600
rect 26056 27548 26108 27600
rect 27620 27548 27672 27600
rect 27712 27548 27764 27600
rect 30196 27591 30248 27600
rect 12532 27523 12584 27532
rect 12532 27489 12541 27523
rect 12541 27489 12575 27523
rect 12575 27489 12584 27523
rect 12532 27480 12584 27489
rect 17592 27480 17644 27532
rect 21824 27480 21876 27532
rect 16764 27412 16816 27464
rect 17868 27412 17920 27464
rect 20168 27412 20220 27464
rect 23480 27480 23532 27532
rect 24492 27412 24544 27464
rect 28356 27480 28408 27532
rect 27988 27412 28040 27464
rect 29828 27455 29880 27464
rect 29828 27421 29837 27455
rect 29837 27421 29871 27455
rect 29871 27421 29880 27455
rect 29828 27412 29880 27421
rect 30196 27557 30205 27591
rect 30205 27557 30239 27591
rect 30239 27557 30248 27591
rect 30196 27548 30248 27557
rect 31944 27548 31996 27600
rect 47676 27591 47728 27600
rect 47676 27557 47685 27591
rect 47685 27557 47719 27591
rect 47719 27557 47728 27591
rect 47676 27548 47728 27557
rect 12624 27344 12676 27396
rect 14740 27344 14792 27396
rect 19432 27344 19484 27396
rect 19524 27344 19576 27396
rect 20812 27387 20864 27396
rect 20812 27353 20821 27387
rect 20821 27353 20855 27387
rect 20855 27353 20864 27387
rect 20812 27344 20864 27353
rect 22100 27344 22152 27396
rect 22928 27344 22980 27396
rect 26056 27344 26108 27396
rect 28908 27344 28960 27396
rect 31484 27412 31536 27464
rect 31760 27412 31812 27464
rect 32312 27412 32364 27464
rect 12808 27276 12860 27328
rect 17040 27276 17092 27328
rect 17776 27276 17828 27328
rect 18236 27276 18288 27328
rect 23480 27276 23532 27328
rect 31116 27276 31168 27328
rect 32864 27276 32916 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 8760 27072 8812 27124
rect 11888 27072 11940 27124
rect 12808 27072 12860 27124
rect 1952 27047 2004 27056
rect 1952 27013 1961 27047
rect 1961 27013 1995 27047
rect 1995 27013 2004 27047
rect 1952 27004 2004 27013
rect 8392 27004 8444 27056
rect 10324 27004 10376 27056
rect 11980 27047 12032 27056
rect 11980 27013 11989 27047
rect 11989 27013 12023 27047
rect 12023 27013 12032 27047
rect 11980 27004 12032 27013
rect 12992 27004 13044 27056
rect 1768 26979 1820 26988
rect 1768 26945 1777 26979
rect 1777 26945 1811 26979
rect 1811 26945 1820 26979
rect 1768 26936 1820 26945
rect 9864 26936 9916 26988
rect 10416 26979 10468 26988
rect 10416 26945 10425 26979
rect 10425 26945 10459 26979
rect 10459 26945 10468 26979
rect 10416 26936 10468 26945
rect 2780 26911 2832 26920
rect 2780 26877 2789 26911
rect 2789 26877 2823 26911
rect 2823 26877 2832 26911
rect 2780 26868 2832 26877
rect 8300 26800 8352 26852
rect 9680 26868 9732 26920
rect 10140 26911 10192 26920
rect 10140 26877 10149 26911
rect 10149 26877 10183 26911
rect 10183 26877 10192 26911
rect 10140 26868 10192 26877
rect 10692 26800 10744 26852
rect 13360 26800 13412 26852
rect 14188 26979 14240 26988
rect 14188 26945 14197 26979
rect 14197 26945 14231 26979
rect 14231 26945 14240 26979
rect 14372 26979 14424 26988
rect 14188 26936 14240 26945
rect 14372 26945 14381 26979
rect 14381 26945 14415 26979
rect 14415 26945 14424 26979
rect 14372 26936 14424 26945
rect 17776 27004 17828 27056
rect 17020 26979 17072 26988
rect 17020 26945 17046 26979
rect 17046 26945 17072 26979
rect 17020 26936 17072 26945
rect 15476 26868 15528 26920
rect 17316 26979 17368 26988
rect 17316 26945 17325 26979
rect 17325 26945 17359 26979
rect 17359 26945 17368 26979
rect 17316 26936 17368 26945
rect 17592 26936 17644 26988
rect 20536 27004 20588 27056
rect 18236 26979 18288 26988
rect 18236 26945 18245 26979
rect 18245 26945 18279 26979
rect 18279 26945 18288 26979
rect 18236 26936 18288 26945
rect 18512 26936 18564 26988
rect 17224 26800 17276 26852
rect 17868 26868 17920 26920
rect 20168 26936 20220 26988
rect 18512 26800 18564 26852
rect 20260 26800 20312 26852
rect 22284 27072 22336 27124
rect 23940 27072 23992 27124
rect 24216 27072 24268 27124
rect 25044 27072 25096 27124
rect 27712 27072 27764 27124
rect 31116 27072 31168 27124
rect 24124 27004 24176 27056
rect 23848 26936 23900 26988
rect 24216 26936 24268 26988
rect 24768 26936 24820 26988
rect 28908 27004 28960 27056
rect 32404 27004 32456 27056
rect 25596 26936 25648 26988
rect 26056 26979 26108 26988
rect 26056 26945 26065 26979
rect 26065 26945 26099 26979
rect 26099 26945 26108 26979
rect 26056 26936 26108 26945
rect 26516 26936 26568 26988
rect 23480 26868 23532 26920
rect 27988 26979 28040 26988
rect 27988 26945 27997 26979
rect 27997 26945 28031 26979
rect 28031 26945 28040 26979
rect 27988 26936 28040 26945
rect 28540 26936 28592 26988
rect 31208 26979 31260 26988
rect 31208 26945 31217 26979
rect 31217 26945 31251 26979
rect 31251 26945 31260 26979
rect 31208 26936 31260 26945
rect 32864 26979 32916 26988
rect 32864 26945 32873 26979
rect 32873 26945 32907 26979
rect 32907 26945 32916 26979
rect 32864 26936 32916 26945
rect 36452 27004 36504 27056
rect 33232 26979 33284 26988
rect 31760 26868 31812 26920
rect 33232 26945 33241 26979
rect 33241 26945 33275 26979
rect 33275 26945 33284 26979
rect 33232 26936 33284 26945
rect 35716 26936 35768 26988
rect 35348 26868 35400 26920
rect 9680 26775 9732 26784
rect 9680 26741 9689 26775
rect 9689 26741 9723 26775
rect 9723 26741 9732 26775
rect 9680 26732 9732 26741
rect 14464 26732 14516 26784
rect 16672 26775 16724 26784
rect 16672 26741 16681 26775
rect 16681 26741 16715 26775
rect 16715 26741 16724 26775
rect 16672 26732 16724 26741
rect 18236 26732 18288 26784
rect 18328 26732 18380 26784
rect 24676 26775 24728 26784
rect 24676 26741 24685 26775
rect 24685 26741 24719 26775
rect 24719 26741 24728 26775
rect 24676 26732 24728 26741
rect 25044 26732 25096 26784
rect 25596 26732 25648 26784
rect 27988 26732 28040 26784
rect 30564 26732 30616 26784
rect 32864 26732 32916 26784
rect 35624 26732 35676 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 11428 26571 11480 26580
rect 11428 26537 11437 26571
rect 11437 26537 11471 26571
rect 11471 26537 11480 26571
rect 11428 26528 11480 26537
rect 14372 26528 14424 26580
rect 1308 26460 1360 26512
rect 1584 26460 1636 26512
rect 10140 26460 10192 26512
rect 10784 26460 10836 26512
rect 10876 26460 10928 26512
rect 1400 26435 1452 26444
rect 1400 26401 1409 26435
rect 1409 26401 1443 26435
rect 1443 26401 1452 26435
rect 1400 26392 1452 26401
rect 2780 26435 2832 26444
rect 2780 26401 2789 26435
rect 2789 26401 2823 26435
rect 2823 26401 2832 26435
rect 17132 26528 17184 26580
rect 26056 26528 26108 26580
rect 28540 26528 28592 26580
rect 31208 26528 31260 26580
rect 37280 26528 37332 26580
rect 20536 26460 20588 26512
rect 2780 26392 2832 26401
rect 24492 26392 24544 26444
rect 27160 26435 27212 26444
rect 27160 26401 27169 26435
rect 27169 26401 27203 26435
rect 27203 26401 27212 26435
rect 27160 26392 27212 26401
rect 29000 26460 29052 26512
rect 30012 26435 30064 26444
rect 30012 26401 30021 26435
rect 30021 26401 30055 26435
rect 30055 26401 30064 26435
rect 30012 26392 30064 26401
rect 7748 26324 7800 26376
rect 12164 26367 12216 26376
rect 12164 26333 12173 26367
rect 12173 26333 12207 26367
rect 12207 26333 12216 26367
rect 12164 26324 12216 26333
rect 12532 26324 12584 26376
rect 13360 26367 13412 26376
rect 13360 26333 13369 26367
rect 13369 26333 13403 26367
rect 13403 26333 13412 26367
rect 13360 26324 13412 26333
rect 1584 26299 1636 26308
rect 1584 26265 1593 26299
rect 1593 26265 1627 26299
rect 1627 26265 1636 26299
rect 1584 26256 1636 26265
rect 9220 26299 9272 26308
rect 9220 26265 9254 26299
rect 9254 26265 9272 26299
rect 9220 26256 9272 26265
rect 10968 26188 11020 26240
rect 11796 26256 11848 26308
rect 13176 26256 13228 26308
rect 14280 26324 14332 26376
rect 14464 26367 14516 26376
rect 14464 26333 14498 26367
rect 14498 26333 14516 26367
rect 14464 26324 14516 26333
rect 16672 26324 16724 26376
rect 20076 26324 20128 26376
rect 24676 26324 24728 26376
rect 33968 26392 34020 26444
rect 31392 26324 31444 26376
rect 32772 26367 32824 26376
rect 32772 26333 32781 26367
rect 32781 26333 32815 26367
rect 32815 26333 32824 26367
rect 32772 26324 32824 26333
rect 32864 26324 32916 26376
rect 34704 26324 34756 26376
rect 15292 26256 15344 26308
rect 17960 26256 18012 26308
rect 31116 26299 31168 26308
rect 31116 26265 31125 26299
rect 31125 26265 31159 26299
rect 31159 26265 31168 26299
rect 31116 26256 31168 26265
rect 33784 26256 33836 26308
rect 35256 26324 35308 26376
rect 35624 26324 35676 26376
rect 37372 26256 37424 26308
rect 46020 26256 46072 26308
rect 47952 26299 48004 26308
rect 47952 26265 47961 26299
rect 47961 26265 47995 26299
rect 47995 26265 48004 26299
rect 47952 26256 48004 26265
rect 48136 26299 48188 26308
rect 48136 26265 48145 26299
rect 48145 26265 48179 26299
rect 48179 26265 48188 26299
rect 48136 26256 48188 26265
rect 12256 26188 12308 26240
rect 12532 26231 12584 26240
rect 12532 26197 12541 26231
rect 12541 26197 12575 26231
rect 12575 26197 12584 26231
rect 12532 26188 12584 26197
rect 15568 26231 15620 26240
rect 15568 26197 15577 26231
rect 15577 26197 15611 26231
rect 15611 26197 15620 26231
rect 15568 26188 15620 26197
rect 18052 26188 18104 26240
rect 18788 26188 18840 26240
rect 22284 26188 22336 26240
rect 23940 26188 23992 26240
rect 26240 26231 26292 26240
rect 26240 26197 26249 26231
rect 26249 26197 26283 26231
rect 26283 26197 26292 26231
rect 26240 26188 26292 26197
rect 29276 26188 29328 26240
rect 34704 26231 34756 26240
rect 34704 26197 34713 26231
rect 34713 26197 34747 26231
rect 34747 26197 34756 26231
rect 34704 26188 34756 26197
rect 36544 26188 36596 26240
rect 46572 26188 46624 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 1584 25984 1636 26036
rect 9220 25984 9272 26036
rect 10324 26027 10376 26036
rect 10324 25993 10333 26027
rect 10333 25993 10367 26027
rect 10367 25993 10376 26027
rect 10324 25984 10376 25993
rect 12256 25984 12308 26036
rect 12716 25984 12768 26036
rect 13728 25984 13780 26036
rect 15292 26027 15344 26036
rect 15292 25993 15301 26027
rect 15301 25993 15335 26027
rect 15335 25993 15344 26027
rect 15292 25984 15344 25993
rect 17224 25984 17276 26036
rect 19432 25984 19484 26036
rect 20168 25984 20220 26036
rect 21824 25984 21876 26036
rect 25872 25984 25924 26036
rect 28264 25984 28316 26036
rect 29276 26027 29328 26036
rect 29276 25993 29285 26027
rect 29285 25993 29319 26027
rect 29319 25993 29328 26027
rect 29276 25984 29328 25993
rect 11980 25916 12032 25968
rect 12440 25916 12492 25968
rect 22284 25916 22336 25968
rect 24492 25916 24544 25968
rect 1400 25891 1452 25900
rect 1400 25857 1409 25891
rect 1409 25857 1443 25891
rect 1443 25857 1452 25891
rect 1400 25848 1452 25857
rect 1768 25848 1820 25900
rect 7104 25891 7156 25900
rect 7104 25857 7113 25891
rect 7113 25857 7147 25891
rect 7147 25857 7156 25891
rect 7104 25848 7156 25857
rect 9680 25848 9732 25900
rect 10876 25848 10928 25900
rect 12808 25891 12860 25900
rect 12808 25857 12817 25891
rect 12817 25857 12851 25891
rect 12851 25857 12860 25891
rect 12808 25848 12860 25857
rect 14096 25848 14148 25900
rect 15568 25848 15620 25900
rect 15752 25891 15804 25900
rect 15752 25857 15761 25891
rect 15761 25857 15795 25891
rect 15795 25857 15804 25891
rect 15752 25848 15804 25857
rect 16764 25848 16816 25900
rect 18052 25848 18104 25900
rect 18236 25848 18288 25900
rect 12440 25780 12492 25832
rect 14832 25780 14884 25832
rect 15660 25780 15712 25832
rect 17132 25780 17184 25832
rect 11704 25755 11756 25764
rect 11704 25721 11713 25755
rect 11713 25721 11747 25755
rect 11747 25721 11756 25755
rect 11704 25712 11756 25721
rect 1584 25687 1636 25696
rect 1584 25653 1593 25687
rect 1593 25653 1627 25687
rect 1627 25653 1636 25687
rect 1584 25644 1636 25653
rect 6736 25644 6788 25696
rect 10324 25687 10376 25696
rect 10324 25653 10333 25687
rect 10333 25653 10367 25687
rect 10367 25653 10376 25687
rect 10324 25644 10376 25653
rect 10508 25687 10560 25696
rect 10508 25653 10517 25687
rect 10517 25653 10551 25687
rect 10551 25653 10560 25687
rect 10508 25644 10560 25653
rect 12532 25712 12584 25764
rect 19984 25780 20036 25832
rect 20444 25780 20496 25832
rect 22468 25891 22520 25900
rect 22468 25857 22477 25891
rect 22477 25857 22511 25891
rect 22511 25857 22520 25891
rect 23480 25891 23532 25900
rect 22468 25848 22520 25857
rect 23480 25857 23489 25891
rect 23489 25857 23523 25891
rect 23523 25857 23532 25891
rect 23480 25848 23532 25857
rect 28632 25916 28684 25968
rect 32956 25984 33008 26036
rect 33232 25984 33284 26036
rect 29552 25916 29604 25968
rect 33968 25959 34020 25968
rect 33968 25925 33977 25959
rect 33977 25925 34011 25959
rect 34011 25925 34020 25959
rect 33968 25916 34020 25925
rect 36544 25984 36596 26036
rect 37372 26027 37424 26036
rect 37372 25993 37381 26027
rect 37381 25993 37415 26027
rect 37415 25993 37424 26027
rect 37372 25984 37424 25993
rect 25872 25848 25924 25900
rect 26056 25848 26108 25900
rect 26884 25848 26936 25900
rect 27988 25848 28040 25900
rect 31392 25848 31444 25900
rect 33048 25891 33100 25900
rect 33048 25857 33057 25891
rect 33057 25857 33091 25891
rect 33091 25857 33100 25891
rect 33048 25848 33100 25857
rect 34704 25916 34756 25968
rect 26240 25780 26292 25832
rect 27896 25823 27948 25832
rect 27896 25789 27905 25823
rect 27905 25789 27939 25823
rect 27939 25789 27948 25823
rect 27896 25780 27948 25789
rect 30932 25823 30984 25832
rect 30932 25789 30941 25823
rect 30941 25789 30975 25823
rect 30975 25789 30984 25823
rect 37280 25891 37332 25900
rect 30932 25780 30984 25789
rect 20168 25712 20220 25764
rect 12624 25644 12676 25696
rect 13176 25644 13228 25696
rect 14280 25644 14332 25696
rect 14556 25644 14608 25696
rect 20352 25644 20404 25696
rect 27712 25712 27764 25764
rect 31116 25712 31168 25764
rect 37280 25857 37289 25891
rect 37289 25857 37323 25891
rect 37323 25857 37332 25891
rect 37280 25848 37332 25857
rect 34704 25780 34756 25832
rect 36452 25712 36504 25764
rect 37372 25712 37424 25764
rect 45652 25712 45704 25764
rect 24860 25687 24912 25696
rect 24860 25653 24869 25687
rect 24869 25653 24903 25687
rect 24903 25653 24912 25687
rect 24860 25644 24912 25653
rect 27620 25644 27672 25696
rect 28816 25644 28868 25696
rect 32588 25644 32640 25696
rect 33048 25644 33100 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 7104 25440 7156 25492
rect 10324 25440 10376 25492
rect 11980 25440 12032 25492
rect 12900 25440 12952 25492
rect 17040 25440 17092 25492
rect 26056 25440 26108 25492
rect 27620 25440 27672 25492
rect 27712 25440 27764 25492
rect 30012 25440 30064 25492
rect 6736 25347 6788 25356
rect 6736 25313 6745 25347
rect 6745 25313 6779 25347
rect 6779 25313 6788 25347
rect 6736 25304 6788 25313
rect 8116 25347 8168 25356
rect 8116 25313 8125 25347
rect 8125 25313 8159 25347
rect 8159 25313 8168 25347
rect 8116 25304 8168 25313
rect 17960 25304 18012 25356
rect 19432 25304 19484 25356
rect 20352 25347 20404 25356
rect 20352 25313 20361 25347
rect 20361 25313 20395 25347
rect 20395 25313 20404 25347
rect 20352 25304 20404 25313
rect 21548 25347 21600 25356
rect 21548 25313 21557 25347
rect 21557 25313 21591 25347
rect 21591 25313 21600 25347
rect 21548 25304 21600 25313
rect 10508 25236 10560 25288
rect 10968 25236 11020 25288
rect 11428 25236 11480 25288
rect 11796 25236 11848 25288
rect 12900 25236 12952 25288
rect 13360 25236 13412 25288
rect 14096 25279 14148 25288
rect 14096 25245 14105 25279
rect 14105 25245 14139 25279
rect 14139 25245 14148 25279
rect 14096 25236 14148 25245
rect 14280 25279 14332 25288
rect 14280 25245 14289 25279
rect 14289 25245 14323 25279
rect 14323 25245 14332 25279
rect 14280 25236 14332 25245
rect 8944 25143 8996 25152
rect 8944 25109 8953 25143
rect 8953 25109 8987 25143
rect 8987 25109 8996 25143
rect 8944 25100 8996 25109
rect 12808 25168 12860 25220
rect 13728 25168 13780 25220
rect 17776 25168 17828 25220
rect 18328 25279 18380 25288
rect 18328 25245 18337 25279
rect 18337 25245 18371 25279
rect 18371 25245 18380 25279
rect 18328 25236 18380 25245
rect 30932 25372 30984 25424
rect 34612 25372 34664 25424
rect 34888 25372 34940 25424
rect 22468 25304 22520 25356
rect 23848 25304 23900 25356
rect 25872 25304 25924 25356
rect 24860 25236 24912 25288
rect 26884 25236 26936 25288
rect 20628 25168 20680 25220
rect 21824 25168 21876 25220
rect 24492 25168 24544 25220
rect 28356 25236 28408 25288
rect 28632 25279 28684 25288
rect 28632 25245 28655 25279
rect 28655 25245 28684 25279
rect 28632 25236 28684 25245
rect 29276 25304 29328 25356
rect 30564 25347 30616 25356
rect 30564 25313 30573 25347
rect 30573 25313 30607 25347
rect 30607 25313 30616 25347
rect 30564 25304 30616 25313
rect 31760 25347 31812 25356
rect 31760 25313 31769 25347
rect 31769 25313 31803 25347
rect 31803 25313 31812 25347
rect 31760 25304 31812 25313
rect 30380 25279 30432 25288
rect 30380 25245 30389 25279
rect 30389 25245 30423 25279
rect 30423 25245 30432 25279
rect 30380 25236 30432 25245
rect 32772 25236 32824 25288
rect 34704 25236 34756 25288
rect 34796 25236 34848 25288
rect 35532 25304 35584 25356
rect 36452 25304 36504 25356
rect 35164 25279 35216 25288
rect 35164 25245 35173 25279
rect 35173 25245 35207 25279
rect 35207 25245 35216 25279
rect 35164 25236 35216 25245
rect 35900 25236 35952 25288
rect 37280 25236 37332 25288
rect 47860 25279 47912 25288
rect 47860 25245 47869 25279
rect 47869 25245 47903 25279
rect 47903 25245 47912 25279
rect 47860 25236 47912 25245
rect 29368 25168 29420 25220
rect 11704 25100 11756 25152
rect 12900 25143 12952 25152
rect 12900 25109 12909 25143
rect 12909 25109 12943 25143
rect 12943 25109 12952 25143
rect 12900 25100 12952 25109
rect 13820 25100 13872 25152
rect 17040 25100 17092 25152
rect 21640 25100 21692 25152
rect 27160 25100 27212 25152
rect 27344 25100 27396 25152
rect 29460 25100 29512 25152
rect 29644 25168 29696 25220
rect 31116 25168 31168 25220
rect 33324 25168 33376 25220
rect 34612 25168 34664 25220
rect 48504 25168 48556 25220
rect 30380 25100 30432 25152
rect 34520 25100 34572 25152
rect 35624 25100 35676 25152
rect 39948 25100 40000 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 9404 24896 9456 24948
rect 29552 24896 29604 24948
rect 30380 24896 30432 24948
rect 31392 24939 31444 24948
rect 31392 24905 31401 24939
rect 31401 24905 31435 24939
rect 31435 24905 31444 24939
rect 31392 24896 31444 24905
rect 14832 24871 14884 24880
rect 14832 24837 14841 24871
rect 14841 24837 14875 24871
rect 14875 24837 14884 24871
rect 14832 24828 14884 24837
rect 22100 24871 22152 24880
rect 22100 24837 22134 24871
rect 22134 24837 22152 24871
rect 22100 24828 22152 24837
rect 7748 24803 7800 24812
rect 7748 24769 7757 24803
rect 7757 24769 7791 24803
rect 7791 24769 7800 24803
rect 7748 24760 7800 24769
rect 8944 24760 8996 24812
rect 10784 24760 10836 24812
rect 14188 24760 14240 24812
rect 15016 24760 15068 24812
rect 10600 24692 10652 24744
rect 15752 24692 15804 24744
rect 21824 24735 21876 24744
rect 21824 24701 21833 24735
rect 21833 24701 21867 24735
rect 21867 24701 21876 24735
rect 21824 24692 21876 24701
rect 25872 24760 25924 24812
rect 26884 24760 26936 24812
rect 11796 24624 11848 24676
rect 20628 24624 20680 24676
rect 26240 24692 26292 24744
rect 27712 24828 27764 24880
rect 27344 24803 27396 24812
rect 27344 24769 27353 24803
rect 27353 24769 27387 24803
rect 27387 24769 27396 24803
rect 28264 24828 28316 24880
rect 33784 24896 33836 24948
rect 35164 24896 35216 24948
rect 27344 24760 27396 24769
rect 28632 24760 28684 24812
rect 35624 24871 35676 24880
rect 35624 24837 35658 24871
rect 35658 24837 35676 24871
rect 35624 24828 35676 24837
rect 29000 24760 29052 24812
rect 29460 24760 29512 24812
rect 30012 24760 30064 24812
rect 24400 24624 24452 24676
rect 9128 24599 9180 24608
rect 9128 24565 9137 24599
rect 9137 24565 9171 24599
rect 9171 24565 9180 24599
rect 9128 24556 9180 24565
rect 10232 24599 10284 24608
rect 10232 24565 10241 24599
rect 10241 24565 10275 24599
rect 10275 24565 10284 24599
rect 10232 24556 10284 24565
rect 10324 24556 10376 24608
rect 11888 24556 11940 24608
rect 14096 24556 14148 24608
rect 26056 24599 26108 24608
rect 26056 24565 26065 24599
rect 26065 24565 26099 24599
rect 26099 24565 26108 24599
rect 26056 24556 26108 24565
rect 26332 24624 26384 24676
rect 27804 24692 27856 24744
rect 27896 24692 27948 24744
rect 30380 24692 30432 24744
rect 34244 24735 34296 24744
rect 34244 24701 34253 24735
rect 34253 24701 34287 24735
rect 34287 24701 34296 24735
rect 34244 24692 34296 24701
rect 34704 24692 34756 24744
rect 37280 24760 37332 24812
rect 47308 24760 47360 24812
rect 47584 24803 47636 24812
rect 47584 24769 47593 24803
rect 47593 24769 47627 24803
rect 47627 24769 47636 24803
rect 47584 24760 47636 24769
rect 28908 24624 28960 24676
rect 27804 24556 27856 24608
rect 28080 24556 28132 24608
rect 28540 24556 28592 24608
rect 33048 24556 33100 24608
rect 33232 24556 33284 24608
rect 36728 24599 36780 24608
rect 36728 24565 36737 24599
rect 36737 24565 36771 24599
rect 36771 24565 36780 24599
rect 36728 24556 36780 24565
rect 37648 24556 37700 24608
rect 38200 24599 38252 24608
rect 38200 24565 38209 24599
rect 38209 24565 38243 24599
rect 38243 24565 38252 24599
rect 38200 24556 38252 24565
rect 46296 24556 46348 24608
rect 47676 24599 47728 24608
rect 47676 24565 47685 24599
rect 47685 24565 47719 24599
rect 47719 24565 47728 24599
rect 47676 24556 47728 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 9312 24327 9364 24336
rect 9312 24293 9321 24327
rect 9321 24293 9355 24327
rect 9355 24293 9364 24327
rect 9312 24284 9364 24293
rect 10232 24259 10284 24268
rect 10232 24225 10241 24259
rect 10241 24225 10275 24259
rect 10275 24225 10284 24259
rect 10232 24216 10284 24225
rect 10508 24216 10560 24268
rect 10968 24216 11020 24268
rect 11152 24327 11204 24336
rect 11152 24293 11161 24327
rect 11161 24293 11195 24327
rect 11195 24293 11204 24327
rect 11152 24284 11204 24293
rect 11244 24216 11296 24268
rect 11796 24259 11848 24268
rect 11796 24225 11805 24259
rect 11805 24225 11839 24259
rect 11839 24225 11848 24259
rect 11796 24216 11848 24225
rect 12900 24352 12952 24404
rect 22744 24352 22796 24404
rect 23388 24395 23440 24404
rect 23388 24361 23397 24395
rect 23397 24361 23431 24395
rect 23431 24361 23440 24395
rect 23388 24352 23440 24361
rect 13820 24216 13872 24268
rect 14188 24216 14240 24268
rect 8852 24148 8904 24200
rect 10140 24191 10192 24200
rect 10140 24157 10149 24191
rect 10149 24157 10183 24191
rect 10183 24157 10192 24191
rect 10140 24148 10192 24157
rect 10324 24191 10376 24200
rect 10324 24157 10333 24191
rect 10333 24157 10367 24191
rect 10367 24157 10376 24191
rect 10324 24148 10376 24157
rect 10876 24148 10928 24200
rect 11888 24191 11940 24200
rect 11888 24157 11897 24191
rect 11897 24157 11931 24191
rect 11931 24157 11940 24191
rect 11888 24148 11940 24157
rect 12900 24191 12952 24200
rect 12900 24157 12909 24191
rect 12909 24157 12943 24191
rect 12943 24157 12952 24191
rect 12900 24148 12952 24157
rect 13912 24148 13964 24200
rect 14096 24191 14148 24200
rect 14096 24157 14105 24191
rect 14105 24157 14139 24191
rect 14139 24157 14148 24191
rect 14096 24148 14148 24157
rect 1860 24123 1912 24132
rect 1860 24089 1869 24123
rect 1869 24089 1903 24123
rect 1903 24089 1912 24123
rect 1860 24080 1912 24089
rect 2688 24080 2740 24132
rect 9128 24080 9180 24132
rect 10968 24123 11020 24132
rect 10968 24089 10977 24123
rect 10977 24089 11011 24123
rect 11011 24089 11020 24123
rect 10968 24080 11020 24089
rect 11428 24080 11480 24132
rect 9404 24012 9456 24064
rect 11704 24012 11756 24064
rect 11888 24012 11940 24064
rect 14832 24148 14884 24200
rect 15292 24191 15344 24200
rect 15292 24157 15301 24191
rect 15301 24157 15335 24191
rect 15335 24157 15344 24191
rect 15292 24148 15344 24157
rect 14924 24080 14976 24132
rect 17316 24148 17368 24200
rect 18696 24191 18748 24200
rect 16672 24080 16724 24132
rect 18236 24080 18288 24132
rect 18696 24157 18705 24191
rect 18705 24157 18739 24191
rect 18739 24157 18748 24191
rect 18696 24148 18748 24157
rect 19984 24148 20036 24200
rect 20260 24148 20312 24200
rect 19432 24080 19484 24132
rect 20352 24080 20404 24132
rect 20628 24123 20680 24132
rect 20628 24089 20637 24123
rect 20637 24089 20671 24123
rect 20671 24089 20680 24123
rect 20628 24080 20680 24089
rect 22100 24123 22152 24132
rect 22100 24089 22109 24123
rect 22109 24089 22143 24123
rect 22143 24089 22152 24123
rect 24768 24148 24820 24200
rect 26332 24284 26384 24336
rect 29368 24352 29420 24404
rect 30104 24395 30156 24404
rect 30104 24361 30113 24395
rect 30113 24361 30147 24395
rect 30147 24361 30156 24395
rect 30104 24352 30156 24361
rect 30656 24352 30708 24404
rect 31852 24352 31904 24404
rect 33324 24395 33376 24404
rect 33324 24361 33333 24395
rect 33333 24361 33367 24395
rect 33367 24361 33376 24395
rect 33324 24352 33376 24361
rect 33508 24352 33560 24404
rect 34244 24352 34296 24404
rect 35532 24352 35584 24404
rect 35900 24395 35952 24404
rect 35900 24361 35909 24395
rect 35909 24361 35943 24395
rect 35943 24361 35952 24395
rect 35900 24352 35952 24361
rect 48044 24352 48096 24404
rect 36452 24284 36504 24336
rect 45008 24284 45060 24336
rect 26148 24148 26200 24200
rect 27896 24148 27948 24200
rect 22100 24080 22152 24089
rect 14832 24055 14884 24064
rect 14832 24021 14841 24055
rect 14841 24021 14875 24055
rect 14875 24021 14884 24055
rect 14832 24012 14884 24021
rect 15568 24012 15620 24064
rect 17408 24055 17460 24064
rect 17408 24021 17417 24055
rect 17417 24021 17451 24055
rect 17451 24021 17460 24055
rect 17408 24012 17460 24021
rect 18052 24055 18104 24064
rect 18052 24021 18061 24055
rect 18061 24021 18095 24055
rect 18095 24021 18104 24055
rect 18052 24012 18104 24021
rect 21180 24012 21232 24064
rect 24860 24012 24912 24064
rect 25504 24012 25556 24064
rect 26056 24012 26108 24064
rect 26792 24012 26844 24064
rect 27068 24080 27120 24132
rect 27528 24012 27580 24064
rect 28724 24191 28776 24200
rect 28724 24157 28733 24191
rect 28733 24157 28767 24191
rect 28767 24157 28776 24191
rect 28724 24148 28776 24157
rect 28908 24216 28960 24268
rect 31300 24216 31352 24268
rect 31576 24216 31628 24268
rect 37648 24259 37700 24268
rect 28908 24080 28960 24132
rect 31392 24080 31444 24132
rect 32864 24148 32916 24200
rect 37648 24225 37657 24259
rect 37657 24225 37691 24259
rect 37691 24225 37700 24259
rect 37648 24216 37700 24225
rect 46296 24259 46348 24268
rect 46296 24225 46305 24259
rect 46305 24225 46339 24259
rect 46339 24225 46348 24259
rect 46296 24216 46348 24225
rect 47676 24216 47728 24268
rect 48136 24259 48188 24268
rect 48136 24225 48145 24259
rect 48145 24225 48179 24259
rect 48179 24225 48188 24259
rect 48136 24216 48188 24225
rect 33784 24191 33836 24200
rect 33784 24157 33793 24191
rect 33793 24157 33827 24191
rect 33827 24157 33836 24191
rect 33784 24148 33836 24157
rect 36728 24148 36780 24200
rect 33232 24080 33284 24132
rect 28632 24055 28684 24064
rect 28632 24021 28641 24055
rect 28641 24021 28675 24055
rect 28675 24021 28684 24055
rect 28632 24012 28684 24021
rect 30104 24012 30156 24064
rect 34520 24080 34572 24132
rect 34888 24123 34940 24132
rect 34888 24089 34897 24123
rect 34897 24089 34931 24123
rect 34931 24089 34940 24123
rect 35716 24123 35768 24132
rect 34888 24080 34940 24089
rect 35716 24089 35725 24123
rect 35725 24089 35759 24123
rect 35759 24089 35768 24123
rect 35716 24080 35768 24089
rect 35992 24080 36044 24132
rect 39304 24123 39356 24132
rect 39304 24089 39313 24123
rect 39313 24089 39347 24123
rect 39347 24089 39356 24123
rect 39304 24080 39356 24089
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 8852 23851 8904 23860
rect 8852 23817 8861 23851
rect 8861 23817 8895 23851
rect 8895 23817 8904 23851
rect 8852 23808 8904 23817
rect 12900 23808 12952 23860
rect 13820 23808 13872 23860
rect 14832 23808 14884 23860
rect 16672 23851 16724 23860
rect 16672 23817 16681 23851
rect 16681 23817 16715 23851
rect 16715 23817 16724 23851
rect 16672 23808 16724 23817
rect 1492 23740 1544 23792
rect 9220 23672 9272 23724
rect 9404 23672 9456 23724
rect 10416 23715 10468 23724
rect 10416 23681 10425 23715
rect 10425 23681 10459 23715
rect 10459 23681 10468 23715
rect 10600 23715 10652 23724
rect 10416 23672 10468 23681
rect 10600 23681 10609 23715
rect 10609 23681 10643 23715
rect 10643 23681 10652 23715
rect 10600 23672 10652 23681
rect 10784 23715 10836 23724
rect 10784 23681 10793 23715
rect 10793 23681 10827 23715
rect 10827 23681 10836 23715
rect 10784 23672 10836 23681
rect 10876 23672 10928 23724
rect 11704 23715 11756 23724
rect 11704 23681 11713 23715
rect 11713 23681 11747 23715
rect 11747 23681 11756 23715
rect 11704 23672 11756 23681
rect 10508 23647 10560 23656
rect 10508 23613 10517 23647
rect 10517 23613 10551 23647
rect 10551 23613 10560 23647
rect 10508 23604 10560 23613
rect 10968 23604 11020 23656
rect 2044 23511 2096 23520
rect 2044 23477 2053 23511
rect 2053 23477 2087 23511
rect 2087 23477 2096 23511
rect 2044 23468 2096 23477
rect 9312 23468 9364 23520
rect 10140 23468 10192 23520
rect 10324 23468 10376 23520
rect 10416 23468 10468 23520
rect 12624 23715 12676 23724
rect 12624 23681 12633 23715
rect 12633 23681 12667 23715
rect 12667 23681 12676 23715
rect 12624 23672 12676 23681
rect 14280 23740 14332 23792
rect 14648 23740 14700 23792
rect 14924 23783 14976 23792
rect 14924 23749 14933 23783
rect 14933 23749 14967 23783
rect 14967 23749 14976 23783
rect 14924 23740 14976 23749
rect 15568 23783 15620 23792
rect 15568 23749 15577 23783
rect 15577 23749 15611 23783
rect 15611 23749 15620 23783
rect 15568 23740 15620 23749
rect 18236 23808 18288 23860
rect 20260 23808 20312 23860
rect 20812 23808 20864 23860
rect 27804 23851 27856 23860
rect 14096 23715 14148 23724
rect 14096 23681 14105 23715
rect 14105 23681 14139 23715
rect 14139 23681 14148 23715
rect 14096 23672 14148 23681
rect 15292 23672 15344 23724
rect 18052 23740 18104 23792
rect 17132 23715 17184 23724
rect 17132 23681 17141 23715
rect 17141 23681 17175 23715
rect 17175 23681 17184 23715
rect 17132 23672 17184 23681
rect 18144 23672 18196 23724
rect 18696 23740 18748 23792
rect 17868 23604 17920 23656
rect 17316 23536 17368 23588
rect 20904 23536 20956 23588
rect 21272 23715 21324 23724
rect 21272 23681 21281 23715
rect 21281 23681 21315 23715
rect 21315 23681 21324 23715
rect 21272 23672 21324 23681
rect 21824 23672 21876 23724
rect 23480 23740 23532 23792
rect 24492 23672 24544 23724
rect 24860 23740 24912 23792
rect 25504 23740 25556 23792
rect 27804 23817 27813 23851
rect 27813 23817 27847 23851
rect 27847 23817 27856 23851
rect 27804 23808 27856 23817
rect 27896 23808 27948 23860
rect 28908 23808 28960 23860
rect 29644 23851 29696 23860
rect 29644 23817 29653 23851
rect 29653 23817 29687 23851
rect 29687 23817 29696 23851
rect 29644 23808 29696 23817
rect 31576 23808 31628 23860
rect 33784 23740 33836 23792
rect 35348 23740 35400 23792
rect 47492 23740 47544 23792
rect 47952 23783 48004 23792
rect 47952 23749 47961 23783
rect 47961 23749 47995 23783
rect 47995 23749 48004 23783
rect 47952 23740 48004 23749
rect 21180 23604 21232 23656
rect 24124 23604 24176 23656
rect 25044 23672 25096 23724
rect 25596 23715 25648 23724
rect 25596 23681 25605 23715
rect 25605 23681 25639 23715
rect 25639 23681 25648 23715
rect 25596 23672 25648 23681
rect 27528 23672 27580 23724
rect 29000 23672 29052 23724
rect 30012 23672 30064 23724
rect 30656 23672 30708 23724
rect 31668 23672 31720 23724
rect 32128 23715 32180 23724
rect 32128 23681 32137 23715
rect 32137 23681 32171 23715
rect 32171 23681 32180 23715
rect 32128 23672 32180 23681
rect 32220 23672 32272 23724
rect 33048 23672 33100 23724
rect 34520 23672 34572 23724
rect 34612 23672 34664 23724
rect 34949 23721 35001 23724
rect 34796 23681 34818 23708
rect 34818 23681 34848 23708
rect 34949 23687 34952 23721
rect 34952 23687 35001 23721
rect 34796 23656 34848 23681
rect 34949 23672 35001 23687
rect 25504 23604 25556 23656
rect 28632 23604 28684 23656
rect 23572 23536 23624 23588
rect 24492 23536 24544 23588
rect 27712 23536 27764 23588
rect 28264 23536 28316 23588
rect 12440 23511 12492 23520
rect 12440 23477 12449 23511
rect 12449 23477 12483 23511
rect 12483 23477 12492 23511
rect 12440 23468 12492 23477
rect 14372 23468 14424 23520
rect 15936 23511 15988 23520
rect 15936 23477 15945 23511
rect 15945 23477 15979 23511
rect 15979 23477 15988 23511
rect 15936 23468 15988 23477
rect 19524 23468 19576 23520
rect 20720 23468 20772 23520
rect 24768 23468 24820 23520
rect 25872 23468 25924 23520
rect 30380 23604 30432 23656
rect 30472 23604 30524 23656
rect 30748 23647 30800 23656
rect 30748 23613 30757 23647
rect 30757 23613 30791 23647
rect 30791 23613 30800 23647
rect 30748 23604 30800 23613
rect 32588 23604 32640 23656
rect 35624 23672 35676 23724
rect 35992 23672 36044 23724
rect 36728 23672 36780 23724
rect 29920 23536 29972 23588
rect 33784 23536 33836 23588
rect 35348 23536 35400 23588
rect 38200 23604 38252 23656
rect 43444 23604 43496 23656
rect 36084 23536 36136 23588
rect 46664 23536 46716 23588
rect 30564 23468 30616 23520
rect 30748 23468 30800 23520
rect 31024 23511 31076 23520
rect 31024 23477 31033 23511
rect 31033 23477 31067 23511
rect 31067 23477 31076 23511
rect 31024 23468 31076 23477
rect 34796 23468 34848 23520
rect 35532 23468 35584 23520
rect 45560 23468 45612 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 1584 23264 1636 23316
rect 11704 23196 11756 23248
rect 2044 23128 2096 23180
rect 2780 23171 2832 23180
rect 2780 23137 2789 23171
rect 2789 23137 2823 23171
rect 2823 23137 2832 23171
rect 10324 23171 10376 23180
rect 2780 23128 2832 23137
rect 10324 23137 10333 23171
rect 10333 23137 10367 23171
rect 10367 23137 10376 23171
rect 10324 23128 10376 23137
rect 11888 23128 11940 23180
rect 13268 23128 13320 23180
rect 15660 23171 15712 23180
rect 10784 23060 10836 23112
rect 12992 23060 13044 23112
rect 13084 23060 13136 23112
rect 15660 23137 15669 23171
rect 15669 23137 15703 23171
rect 15703 23137 15712 23171
rect 15660 23128 15712 23137
rect 16580 23128 16632 23180
rect 14280 23060 14332 23112
rect 14740 23060 14792 23112
rect 2596 22992 2648 23044
rect 12440 22992 12492 23044
rect 6920 22924 6972 22976
rect 14464 22924 14516 22976
rect 16580 22992 16632 23044
rect 17132 23196 17184 23248
rect 19432 23196 19484 23248
rect 25596 23264 25648 23316
rect 25872 23264 25924 23316
rect 27068 23264 27120 23316
rect 31116 23264 31168 23316
rect 29368 23196 29420 23248
rect 29460 23196 29512 23248
rect 44180 23264 44232 23316
rect 32956 23196 33008 23248
rect 33692 23196 33744 23248
rect 17224 23128 17276 23180
rect 16856 23060 16908 23112
rect 17316 23103 17368 23112
rect 17316 23069 17325 23103
rect 17325 23069 17359 23103
rect 17359 23069 17368 23103
rect 17316 23060 17368 23069
rect 23480 23128 23532 23180
rect 17868 23060 17920 23112
rect 22376 23060 22428 23112
rect 23940 23060 23992 23112
rect 29644 23128 29696 23180
rect 26792 23103 26844 23112
rect 26792 23069 26801 23103
rect 26801 23069 26835 23103
rect 26835 23069 26844 23103
rect 26792 23060 26844 23069
rect 27068 23060 27120 23112
rect 27436 23060 27488 23112
rect 28080 23060 28132 23112
rect 28632 23060 28684 23112
rect 33968 23128 34020 23180
rect 34704 23171 34756 23180
rect 34704 23137 34713 23171
rect 34713 23137 34747 23171
rect 34747 23137 34756 23171
rect 34704 23128 34756 23137
rect 19156 22992 19208 23044
rect 19340 22992 19392 23044
rect 19432 23035 19484 23044
rect 19432 23001 19441 23035
rect 19441 23001 19475 23035
rect 19475 23001 19484 23035
rect 20720 23035 20772 23044
rect 19432 22992 19484 23001
rect 20720 23001 20754 23035
rect 20754 23001 20772 23035
rect 20720 22992 20772 23001
rect 20812 22992 20864 23044
rect 24952 22992 25004 23044
rect 27896 22992 27948 23044
rect 29368 22992 29420 23044
rect 30564 23060 30616 23112
rect 32128 23060 32180 23112
rect 32312 23060 32364 23112
rect 33048 23060 33100 23112
rect 17960 22924 18012 22976
rect 18052 22924 18104 22976
rect 20628 22924 20680 22976
rect 23664 22967 23716 22976
rect 23664 22933 23673 22967
rect 23673 22933 23707 22967
rect 23707 22933 23716 22967
rect 23664 22924 23716 22933
rect 25780 22924 25832 22976
rect 30288 22924 30340 22976
rect 30472 22992 30524 23044
rect 30932 22924 30984 22976
rect 31116 22992 31168 23044
rect 38292 23060 38344 23112
rect 48136 23103 48188 23112
rect 48136 23069 48145 23103
rect 48145 23069 48179 23103
rect 48179 23069 48188 23103
rect 48136 23060 48188 23069
rect 34520 22992 34572 23044
rect 32956 22924 33008 22976
rect 33048 22924 33100 22976
rect 35900 22924 35952 22976
rect 46112 22924 46164 22976
rect 47584 22924 47636 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 2596 22763 2648 22772
rect 2596 22729 2605 22763
rect 2605 22729 2639 22763
rect 2639 22729 2648 22763
rect 2596 22720 2648 22729
rect 10600 22720 10652 22772
rect 13820 22720 13872 22772
rect 14280 22720 14332 22772
rect 14464 22763 14516 22772
rect 14464 22729 14473 22763
rect 14473 22729 14507 22763
rect 14507 22729 14516 22763
rect 14464 22720 14516 22729
rect 17224 22720 17276 22772
rect 17960 22720 18012 22772
rect 23940 22720 23992 22772
rect 24124 22720 24176 22772
rect 25228 22720 25280 22772
rect 26700 22720 26752 22772
rect 30840 22720 30892 22772
rect 33140 22720 33192 22772
rect 36360 22720 36412 22772
rect 13084 22652 13136 22704
rect 13268 22695 13320 22704
rect 13268 22661 13277 22695
rect 13277 22661 13311 22695
rect 13311 22661 13320 22695
rect 13268 22652 13320 22661
rect 1860 22627 1912 22636
rect 1860 22593 1869 22627
rect 1869 22593 1903 22627
rect 1903 22593 1912 22627
rect 1860 22584 1912 22593
rect 2504 22627 2556 22636
rect 2504 22593 2513 22627
rect 2513 22593 2547 22627
rect 2547 22593 2556 22627
rect 2504 22584 2556 22593
rect 9496 22584 9548 22636
rect 10784 22584 10836 22636
rect 14096 22652 14148 22704
rect 14372 22695 14424 22704
rect 14372 22661 14381 22695
rect 14381 22661 14415 22695
rect 14415 22661 14424 22695
rect 14372 22652 14424 22661
rect 15936 22652 15988 22704
rect 14464 22584 14516 22636
rect 18236 22627 18288 22636
rect 18236 22593 18245 22627
rect 18245 22593 18279 22627
rect 18279 22593 18288 22627
rect 18236 22584 18288 22593
rect 18328 22627 18380 22636
rect 18328 22593 18337 22627
rect 18337 22593 18371 22627
rect 18371 22593 18380 22627
rect 18328 22584 18380 22593
rect 20720 22652 20772 22704
rect 9956 22559 10008 22568
rect 9956 22525 9965 22559
rect 9965 22525 9999 22559
rect 9999 22525 10008 22559
rect 9956 22516 10008 22525
rect 10416 22516 10468 22568
rect 10968 22559 11020 22568
rect 10968 22525 10977 22559
rect 10977 22525 11011 22559
rect 11011 22525 11020 22559
rect 10968 22516 11020 22525
rect 13728 22516 13780 22568
rect 19892 22584 19944 22636
rect 9772 22380 9824 22432
rect 10416 22380 10468 22432
rect 14280 22448 14332 22500
rect 14832 22448 14884 22500
rect 14924 22448 14976 22500
rect 17960 22448 18012 22500
rect 18144 22448 18196 22500
rect 20076 22516 20128 22568
rect 21088 22627 21140 22636
rect 21088 22593 21102 22627
rect 21102 22593 21136 22627
rect 21136 22593 21140 22627
rect 21088 22584 21140 22593
rect 21272 22627 21324 22636
rect 21272 22593 21281 22627
rect 21281 22593 21315 22627
rect 21315 22593 21324 22627
rect 21272 22584 21324 22593
rect 18420 22448 18472 22500
rect 19432 22448 19484 22500
rect 20904 22448 20956 22500
rect 13820 22380 13872 22432
rect 13912 22380 13964 22432
rect 16028 22380 16080 22432
rect 20812 22380 20864 22432
rect 24768 22652 24820 22704
rect 26148 22652 26200 22704
rect 30748 22652 30800 22704
rect 31116 22652 31168 22704
rect 24400 22627 24452 22636
rect 24400 22593 24409 22627
rect 24409 22593 24443 22627
rect 24443 22593 24452 22627
rect 24400 22584 24452 22593
rect 25228 22627 25280 22636
rect 24768 22516 24820 22568
rect 25228 22593 25237 22627
rect 25237 22593 25271 22627
rect 25271 22593 25280 22627
rect 25228 22584 25280 22593
rect 25504 22584 25556 22636
rect 25872 22627 25924 22636
rect 25872 22593 25881 22627
rect 25881 22593 25915 22627
rect 25915 22593 25924 22627
rect 25872 22584 25924 22593
rect 29460 22627 29512 22636
rect 29460 22593 29469 22627
rect 29469 22593 29503 22627
rect 29503 22593 29512 22627
rect 29460 22584 29512 22593
rect 29644 22584 29696 22636
rect 30840 22584 30892 22636
rect 31484 22584 31536 22636
rect 32128 22584 32180 22636
rect 33600 22652 33652 22704
rect 47124 22652 47176 22704
rect 47400 22652 47452 22704
rect 33140 22584 33192 22636
rect 35716 22627 35768 22636
rect 35716 22593 35725 22627
rect 35725 22593 35759 22627
rect 35759 22593 35768 22627
rect 35716 22584 35768 22593
rect 35900 22627 35952 22636
rect 35900 22593 35909 22627
rect 35909 22593 35943 22627
rect 35943 22593 35952 22627
rect 35900 22584 35952 22593
rect 36084 22584 36136 22636
rect 47584 22627 47636 22636
rect 47584 22593 47593 22627
rect 47593 22593 47627 22627
rect 47627 22593 47636 22627
rect 47584 22584 47636 22593
rect 25136 22516 25188 22568
rect 29552 22559 29604 22568
rect 29552 22525 29561 22559
rect 29561 22525 29595 22559
rect 29595 22525 29604 22559
rect 29552 22516 29604 22525
rect 31576 22516 31628 22568
rect 33600 22559 33652 22568
rect 24952 22491 25004 22500
rect 24952 22457 24961 22491
rect 24961 22457 24995 22491
rect 24995 22457 25004 22491
rect 24952 22448 25004 22457
rect 25228 22448 25280 22500
rect 26148 22380 26200 22432
rect 29368 22380 29420 22432
rect 31392 22448 31444 22500
rect 33600 22525 33609 22559
rect 33609 22525 33643 22559
rect 33643 22525 33652 22559
rect 33600 22516 33652 22525
rect 42064 22516 42116 22568
rect 35624 22448 35676 22500
rect 36268 22448 36320 22500
rect 34612 22380 34664 22432
rect 47676 22423 47728 22432
rect 47676 22389 47685 22423
rect 47685 22389 47719 22423
rect 47719 22389 47728 22423
rect 47676 22380 47728 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 4804 22176 4856 22228
rect 9496 22108 9548 22160
rect 15292 22108 15344 22160
rect 18328 22176 18380 22228
rect 18512 22108 18564 22160
rect 20076 22151 20128 22160
rect 20076 22117 20085 22151
rect 20085 22117 20119 22151
rect 20119 22117 20128 22151
rect 20076 22108 20128 22117
rect 21088 22176 21140 22228
rect 29460 22176 29512 22228
rect 29736 22219 29788 22228
rect 29736 22185 29745 22219
rect 29745 22185 29779 22219
rect 29779 22185 29788 22219
rect 29736 22176 29788 22185
rect 26700 22108 26752 22160
rect 26884 22108 26936 22160
rect 30196 22219 30248 22228
rect 30196 22185 30205 22219
rect 30205 22185 30239 22219
rect 30239 22185 30248 22219
rect 30840 22219 30892 22228
rect 30196 22176 30248 22185
rect 30840 22185 30849 22219
rect 30849 22185 30883 22219
rect 30883 22185 30892 22219
rect 30840 22176 30892 22185
rect 31484 22176 31536 22228
rect 46940 22176 46992 22228
rect 47860 22219 47912 22228
rect 47860 22185 47869 22219
rect 47869 22185 47903 22219
rect 47903 22185 47912 22219
rect 47860 22176 47912 22185
rect 7840 22040 7892 22092
rect 8024 21972 8076 22024
rect 9956 22015 10008 22024
rect 9956 21981 9965 22015
rect 9965 21981 9999 22015
rect 9999 21981 10008 22015
rect 9956 21972 10008 21981
rect 14096 21972 14148 22024
rect 14556 22040 14608 22092
rect 17224 22040 17276 22092
rect 2320 21836 2372 21888
rect 7196 21836 7248 21888
rect 7288 21836 7340 21888
rect 9956 21879 10008 21888
rect 9956 21845 9965 21879
rect 9965 21845 9999 21879
rect 9999 21845 10008 21879
rect 9956 21836 10008 21845
rect 10140 21904 10192 21956
rect 10968 21904 11020 21956
rect 14464 21947 14516 21956
rect 14464 21913 14473 21947
rect 14473 21913 14507 21947
rect 14507 21913 14516 21947
rect 14464 21904 14516 21913
rect 16672 21972 16724 22024
rect 17960 22015 18012 22024
rect 17592 21904 17644 21956
rect 17960 21981 17969 22015
rect 17969 21981 18003 22015
rect 18003 21981 18012 22015
rect 17960 21972 18012 21981
rect 19432 21972 19484 22024
rect 20628 21972 20680 22024
rect 20996 21972 21048 22024
rect 24860 21972 24912 22024
rect 25136 22015 25188 22024
rect 25136 21981 25145 22015
rect 25145 21981 25179 22015
rect 25179 21981 25188 22015
rect 25136 21972 25188 21981
rect 19340 21904 19392 21956
rect 20352 21904 20404 21956
rect 22192 21904 22244 21956
rect 22284 21904 22336 21956
rect 25320 21904 25372 21956
rect 26332 22040 26384 22092
rect 28540 22040 28592 22092
rect 28724 22040 28776 22092
rect 29644 22040 29696 22092
rect 30932 22083 30984 22092
rect 25504 22015 25556 22024
rect 25504 21981 25513 22015
rect 25513 21981 25547 22015
rect 25547 21981 25556 22015
rect 26240 22015 26292 22024
rect 25504 21972 25556 21981
rect 26240 21981 26249 22015
rect 26249 21981 26283 22015
rect 26283 21981 26292 22015
rect 26240 21972 26292 21981
rect 26424 22015 26476 22024
rect 26424 21981 26433 22015
rect 26433 21981 26467 22015
rect 26467 21981 26476 22015
rect 26424 21972 26476 21981
rect 26240 21836 26292 21888
rect 26424 21879 26476 21888
rect 26424 21845 26433 21879
rect 26433 21845 26467 21879
rect 26467 21845 26476 21879
rect 26424 21836 26476 21845
rect 26516 21836 26568 21888
rect 27804 21972 27856 22024
rect 28816 22015 28868 22024
rect 27252 21836 27304 21888
rect 28816 21981 28825 22015
rect 28825 21981 28859 22015
rect 28859 21981 28868 22015
rect 28816 21972 28868 21981
rect 28264 21904 28316 21956
rect 29736 21972 29788 22024
rect 30932 22049 30941 22083
rect 30941 22049 30975 22083
rect 30975 22049 30984 22083
rect 30932 22040 30984 22049
rect 32864 22040 32916 22092
rect 29184 21904 29236 21956
rect 29460 21904 29512 21956
rect 30012 22015 30064 22024
rect 30012 21981 30021 22015
rect 30021 21981 30055 22015
rect 30055 21981 30064 22015
rect 30012 21972 30064 21981
rect 31392 21972 31444 22024
rect 32128 21972 32180 22024
rect 33416 21972 33468 22024
rect 36268 22108 36320 22160
rect 47400 22083 47452 22092
rect 33968 22015 34020 22024
rect 33968 21981 33977 22015
rect 33977 21981 34011 22015
rect 34011 21981 34020 22015
rect 33968 21972 34020 21981
rect 34612 21972 34664 22024
rect 34704 21972 34756 22024
rect 29092 21836 29144 21888
rect 29920 21836 29972 21888
rect 31208 21904 31260 21956
rect 31300 21904 31352 21956
rect 32680 21904 32732 21956
rect 34520 21904 34572 21956
rect 34796 21904 34848 21956
rect 47400 22049 47409 22083
rect 47409 22049 47443 22083
rect 47443 22049 47452 22083
rect 47400 22040 47452 22049
rect 36268 21972 36320 22024
rect 47584 21972 47636 22024
rect 47860 22015 47912 22024
rect 47860 21981 47869 22015
rect 47869 21981 47903 22015
rect 47903 21981 47912 22015
rect 47860 21972 47912 21981
rect 37372 21904 37424 21956
rect 40776 21904 40828 21956
rect 36176 21836 36228 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 2688 21632 2740 21684
rect 14556 21632 14608 21684
rect 14832 21632 14884 21684
rect 15660 21632 15712 21684
rect 19340 21632 19392 21684
rect 20352 21632 20404 21684
rect 20628 21632 20680 21684
rect 2412 21564 2464 21616
rect 7104 21564 7156 21616
rect 7196 21564 7248 21616
rect 17224 21564 17276 21616
rect 17408 21564 17460 21616
rect 22284 21564 22336 21616
rect 22376 21564 22428 21616
rect 2228 21496 2280 21548
rect 7288 21539 7340 21548
rect 7288 21505 7297 21539
rect 7297 21505 7331 21539
rect 7331 21505 7340 21539
rect 7288 21496 7340 21505
rect 9956 21496 10008 21548
rect 10232 21496 10284 21548
rect 13820 21496 13872 21548
rect 14188 21539 14240 21548
rect 14188 21505 14197 21539
rect 14197 21505 14231 21539
rect 14231 21505 14240 21539
rect 14188 21496 14240 21505
rect 14464 21539 14516 21548
rect 14464 21505 14473 21539
rect 14473 21505 14507 21539
rect 14507 21505 14516 21539
rect 14464 21496 14516 21505
rect 15384 21539 15436 21548
rect 15384 21505 15393 21539
rect 15393 21505 15427 21539
rect 15427 21505 15436 21539
rect 15384 21496 15436 21505
rect 16488 21496 16540 21548
rect 20168 21539 20220 21548
rect 7472 21471 7524 21480
rect 7472 21437 7481 21471
rect 7481 21437 7515 21471
rect 7515 21437 7524 21471
rect 7472 21428 7524 21437
rect 3424 21360 3476 21412
rect 12164 21428 12216 21480
rect 13084 21471 13136 21480
rect 13084 21437 13093 21471
rect 13093 21437 13127 21471
rect 13127 21437 13136 21471
rect 13084 21428 13136 21437
rect 14648 21428 14700 21480
rect 15292 21471 15344 21480
rect 15292 21437 15301 21471
rect 15301 21437 15335 21471
rect 15335 21437 15344 21471
rect 15292 21428 15344 21437
rect 20168 21505 20177 21539
rect 20177 21505 20211 21539
rect 20211 21505 20220 21539
rect 20168 21496 20220 21505
rect 20812 21428 20864 21480
rect 21272 21496 21324 21548
rect 22560 21496 22612 21548
rect 23112 21564 23164 21616
rect 22376 21428 22428 21480
rect 11612 21360 11664 21412
rect 25228 21632 25280 21684
rect 26056 21632 26108 21684
rect 26240 21632 26292 21684
rect 29828 21675 29880 21684
rect 24860 21564 24912 21616
rect 26424 21564 26476 21616
rect 26884 21564 26936 21616
rect 24952 21539 25004 21548
rect 24952 21505 24961 21539
rect 24961 21505 24995 21539
rect 24995 21505 25004 21539
rect 24952 21496 25004 21505
rect 26056 21539 26108 21548
rect 26056 21505 26065 21539
rect 26065 21505 26099 21539
rect 26099 21505 26108 21539
rect 26056 21496 26108 21505
rect 26148 21539 26200 21548
rect 26148 21505 26157 21539
rect 26157 21505 26191 21539
rect 26191 21505 26200 21539
rect 27252 21539 27304 21548
rect 26148 21496 26200 21505
rect 27252 21505 27261 21539
rect 27261 21505 27295 21539
rect 27295 21505 27304 21539
rect 27252 21496 27304 21505
rect 28172 21496 28224 21548
rect 28448 21564 28500 21616
rect 28724 21564 28776 21616
rect 29828 21641 29837 21675
rect 29837 21641 29871 21675
rect 29871 21641 29880 21675
rect 29828 21632 29880 21641
rect 31300 21632 31352 21684
rect 31576 21675 31628 21684
rect 31576 21641 31585 21675
rect 31585 21641 31619 21675
rect 31619 21641 31628 21675
rect 31576 21632 31628 21641
rect 31944 21632 31996 21684
rect 32312 21632 32364 21684
rect 32588 21675 32640 21684
rect 32588 21641 32597 21675
rect 32597 21641 32631 21675
rect 32631 21641 32640 21675
rect 32588 21632 32640 21641
rect 33600 21632 33652 21684
rect 36268 21632 36320 21684
rect 37372 21675 37424 21684
rect 37372 21641 37381 21675
rect 37381 21641 37415 21675
rect 37415 21641 37424 21675
rect 37372 21632 37424 21641
rect 26332 21428 26384 21480
rect 26424 21428 26476 21480
rect 27344 21428 27396 21480
rect 27620 21428 27672 21480
rect 28540 21539 28592 21548
rect 28540 21505 28549 21539
rect 28549 21505 28583 21539
rect 28583 21505 28592 21539
rect 29368 21539 29420 21548
rect 28540 21496 28592 21505
rect 29368 21505 29377 21539
rect 29377 21505 29411 21539
rect 29411 21505 29420 21539
rect 29368 21496 29420 21505
rect 30012 21564 30064 21616
rect 47860 21632 47912 21684
rect 47952 21607 48004 21616
rect 47952 21573 47961 21607
rect 47961 21573 47995 21607
rect 47995 21573 48004 21607
rect 47952 21564 48004 21573
rect 30748 21496 30800 21548
rect 31944 21496 31996 21548
rect 12256 21292 12308 21344
rect 14096 21292 14148 21344
rect 15384 21292 15436 21344
rect 16764 21292 16816 21344
rect 18236 21292 18288 21344
rect 20352 21335 20404 21344
rect 20352 21301 20361 21335
rect 20361 21301 20395 21335
rect 20395 21301 20404 21335
rect 20352 21292 20404 21301
rect 20720 21292 20772 21344
rect 22928 21292 22980 21344
rect 23020 21292 23072 21344
rect 23664 21292 23716 21344
rect 26976 21360 27028 21412
rect 29460 21428 29512 21480
rect 27344 21292 27396 21344
rect 28264 21335 28316 21344
rect 28264 21301 28273 21335
rect 28273 21301 28307 21335
rect 28307 21301 28316 21335
rect 28264 21292 28316 21301
rect 28908 21292 28960 21344
rect 30932 21428 30984 21480
rect 32036 21428 32088 21480
rect 32496 21496 32548 21548
rect 32956 21496 33008 21548
rect 36360 21496 36412 21548
rect 37280 21539 37332 21548
rect 37280 21505 37289 21539
rect 37289 21505 37323 21539
rect 37323 21505 37332 21539
rect 37280 21496 37332 21505
rect 32312 21471 32364 21480
rect 32312 21437 32321 21471
rect 32321 21437 32355 21471
rect 32355 21437 32364 21471
rect 32312 21428 32364 21437
rect 33416 21428 33468 21480
rect 33876 21471 33928 21480
rect 33876 21437 33885 21471
rect 33885 21437 33919 21471
rect 33919 21437 33928 21471
rect 33876 21428 33928 21437
rect 45468 21428 45520 21480
rect 29184 21292 29236 21344
rect 29276 21292 29328 21344
rect 29460 21292 29512 21344
rect 30932 21292 30984 21344
rect 48228 21360 48280 21412
rect 31760 21292 31812 21344
rect 32772 21292 32824 21344
rect 39948 21292 40000 21344
rect 48044 21335 48096 21344
rect 48044 21301 48053 21335
rect 48053 21301 48087 21335
rect 48087 21301 48096 21335
rect 48044 21292 48096 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 7472 21088 7524 21140
rect 12164 21131 12216 21140
rect 12164 21097 12173 21131
rect 12173 21097 12207 21131
rect 12207 21097 12216 21131
rect 12164 21088 12216 21097
rect 12256 21088 12308 21140
rect 20628 21088 20680 21140
rect 20812 21088 20864 21140
rect 21272 21088 21324 21140
rect 22376 21088 22428 21140
rect 22560 21088 22612 21140
rect 23664 21088 23716 21140
rect 25780 21088 25832 21140
rect 27436 21131 27488 21140
rect 27436 21097 27445 21131
rect 27445 21097 27479 21131
rect 27479 21097 27488 21131
rect 27436 21088 27488 21097
rect 27528 21088 27580 21140
rect 28448 21088 28500 21140
rect 28816 21131 28868 21140
rect 28816 21097 28825 21131
rect 28825 21097 28859 21131
rect 28859 21097 28868 21131
rect 28816 21088 28868 21097
rect 1400 21020 1452 21072
rect 11612 21020 11664 21072
rect 13452 21020 13504 21072
rect 13544 21020 13596 21072
rect 16672 21020 16724 21072
rect 6828 20884 6880 20936
rect 12808 20952 12860 21004
rect 3976 20816 4028 20868
rect 11612 20816 11664 20868
rect 12348 20884 12400 20936
rect 16856 20995 16908 21004
rect 16856 20961 16865 20995
rect 16865 20961 16899 20995
rect 16899 20961 16908 20995
rect 16856 20952 16908 20961
rect 26700 21020 26752 21072
rect 31024 21088 31076 21140
rect 36176 21088 36228 21140
rect 13544 20927 13596 20936
rect 13544 20893 13547 20927
rect 13547 20893 13581 20927
rect 13581 20893 13596 20927
rect 13544 20884 13596 20893
rect 17408 20884 17460 20936
rect 17592 20884 17644 20936
rect 22376 20952 22428 21004
rect 20168 20884 20220 20936
rect 20996 20927 21048 20936
rect 20996 20893 21005 20927
rect 21005 20893 21039 20927
rect 21039 20893 21048 20927
rect 20996 20884 21048 20893
rect 21272 20927 21324 20936
rect 21272 20893 21281 20927
rect 21281 20893 21315 20927
rect 21315 20893 21324 20927
rect 21272 20884 21324 20893
rect 4068 20748 4120 20800
rect 5540 20748 5592 20800
rect 12900 20791 12952 20800
rect 12900 20757 12909 20791
rect 12909 20757 12943 20791
rect 12943 20757 12952 20791
rect 12900 20748 12952 20757
rect 14096 20859 14148 20868
rect 14096 20825 14105 20859
rect 14105 20825 14139 20859
rect 14139 20825 14148 20859
rect 14096 20816 14148 20825
rect 14372 20816 14424 20868
rect 13452 20748 13504 20800
rect 16764 20816 16816 20868
rect 17500 20816 17552 20868
rect 14556 20748 14608 20800
rect 22560 20816 22612 20868
rect 17776 20748 17828 20800
rect 18328 20748 18380 20800
rect 20996 20748 21048 20800
rect 21364 20748 21416 20800
rect 22928 20927 22980 20936
rect 22928 20893 22937 20927
rect 22937 20893 22971 20927
rect 22971 20893 22980 20927
rect 22928 20884 22980 20893
rect 25044 20884 25096 20936
rect 25780 20884 25832 20936
rect 26884 20995 26936 21004
rect 26884 20961 26893 20995
rect 26893 20961 26927 20995
rect 26927 20961 26936 20995
rect 27620 20995 27672 21004
rect 26884 20952 26936 20961
rect 26148 20884 26200 20936
rect 27620 20961 27629 20995
rect 27629 20961 27663 20995
rect 27663 20961 27672 20995
rect 27620 20952 27672 20961
rect 28724 20952 28776 21004
rect 29092 20952 29144 21004
rect 31576 21020 31628 21072
rect 48044 21020 48096 21072
rect 30656 20952 30708 21004
rect 36084 20995 36136 21004
rect 36084 20961 36093 20995
rect 36093 20961 36127 20995
rect 36127 20961 36136 20995
rect 36084 20952 36136 20961
rect 36268 20995 36320 21004
rect 36268 20961 36277 20995
rect 36277 20961 36311 20995
rect 36311 20961 36320 20995
rect 36268 20952 36320 20961
rect 36360 20952 36412 21004
rect 37832 20952 37884 21004
rect 27804 20884 27856 20936
rect 28172 20884 28224 20936
rect 28540 20884 28592 20936
rect 28816 20884 28868 20936
rect 31392 20927 31444 20936
rect 31392 20893 31401 20927
rect 31401 20893 31435 20927
rect 31435 20893 31444 20927
rect 31392 20884 31444 20893
rect 31668 20884 31720 20936
rect 33232 20884 33284 20936
rect 26240 20816 26292 20868
rect 27252 20816 27304 20868
rect 27896 20791 27948 20800
rect 27896 20757 27905 20791
rect 27905 20757 27939 20791
rect 27939 20757 27948 20791
rect 27896 20748 27948 20757
rect 28908 20816 28960 20868
rect 31208 20859 31260 20868
rect 31208 20825 31217 20859
rect 31217 20825 31251 20859
rect 31251 20825 31260 20859
rect 31208 20816 31260 20825
rect 31760 20816 31812 20868
rect 32036 20816 32088 20868
rect 37924 20859 37976 20868
rect 37924 20825 37933 20859
rect 37933 20825 37967 20859
rect 37967 20825 37976 20859
rect 37924 20816 37976 20825
rect 47676 20816 47728 20868
rect 29920 20748 29972 20800
rect 30012 20791 30064 20800
rect 30012 20757 30021 20791
rect 30021 20757 30055 20791
rect 30055 20757 30064 20791
rect 30012 20748 30064 20757
rect 31116 20748 31168 20800
rect 33692 20748 33744 20800
rect 37464 20748 37516 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 7932 20544 7984 20596
rect 17132 20544 17184 20596
rect 17500 20587 17552 20596
rect 17500 20553 17509 20587
rect 17509 20553 17543 20587
rect 17543 20553 17552 20587
rect 17500 20544 17552 20553
rect 17868 20544 17920 20596
rect 17960 20544 18012 20596
rect 41604 20544 41656 20596
rect 12900 20476 12952 20528
rect 19340 20476 19392 20528
rect 20352 20476 20404 20528
rect 10508 20408 10560 20460
rect 11704 20451 11756 20460
rect 11704 20417 11713 20451
rect 11713 20417 11747 20451
rect 11747 20417 11756 20451
rect 11704 20408 11756 20417
rect 12992 20408 13044 20460
rect 15752 20451 15804 20460
rect 15752 20417 15761 20451
rect 15761 20417 15795 20451
rect 15795 20417 15804 20451
rect 15752 20408 15804 20417
rect 8760 20383 8812 20392
rect 8760 20349 8769 20383
rect 8769 20349 8803 20383
rect 8803 20349 8812 20383
rect 8760 20340 8812 20349
rect 8944 20383 8996 20392
rect 8944 20349 8953 20383
rect 8953 20349 8987 20383
rect 8987 20349 8996 20383
rect 8944 20340 8996 20349
rect 10416 20383 10468 20392
rect 10416 20349 10425 20383
rect 10425 20349 10459 20383
rect 10459 20349 10468 20383
rect 10416 20340 10468 20349
rect 15936 20451 15988 20460
rect 15936 20417 15945 20451
rect 15945 20417 15979 20451
rect 15979 20417 15988 20451
rect 15936 20408 15988 20417
rect 17316 20408 17368 20460
rect 4896 20247 4948 20256
rect 4896 20213 4905 20247
rect 4905 20213 4939 20247
rect 4939 20213 4948 20247
rect 4896 20204 4948 20213
rect 11980 20204 12032 20256
rect 12808 20204 12860 20256
rect 14464 20247 14516 20256
rect 14464 20213 14473 20247
rect 14473 20213 14507 20247
rect 14507 20213 14516 20247
rect 14464 20204 14516 20213
rect 15476 20247 15528 20256
rect 15476 20213 15485 20247
rect 15485 20213 15519 20247
rect 15519 20213 15528 20247
rect 15476 20204 15528 20213
rect 18144 20451 18196 20460
rect 18144 20417 18153 20451
rect 18153 20417 18187 20451
rect 18187 20417 18196 20451
rect 18144 20408 18196 20417
rect 19248 20408 19300 20460
rect 19616 20408 19668 20460
rect 21732 20408 21784 20460
rect 21916 20408 21968 20460
rect 23020 20476 23072 20528
rect 23112 20476 23164 20528
rect 25136 20476 25188 20528
rect 27896 20476 27948 20528
rect 23848 20451 23900 20460
rect 18052 20340 18104 20392
rect 19432 20340 19484 20392
rect 23848 20417 23857 20451
rect 23857 20417 23891 20451
rect 23891 20417 23900 20451
rect 23848 20408 23900 20417
rect 28264 20408 28316 20460
rect 28908 20451 28960 20460
rect 28908 20417 28917 20451
rect 28917 20417 28951 20451
rect 28951 20417 28960 20451
rect 28908 20408 28960 20417
rect 30840 20519 30892 20528
rect 30840 20485 30849 20519
rect 30849 20485 30883 20519
rect 30883 20485 30892 20519
rect 30840 20476 30892 20485
rect 31392 20476 31444 20528
rect 31944 20476 31996 20528
rect 32496 20476 32548 20528
rect 33692 20519 33744 20528
rect 33692 20485 33701 20519
rect 33701 20485 33735 20519
rect 33735 20485 33744 20519
rect 33692 20476 33744 20485
rect 37464 20519 37516 20528
rect 37464 20485 37473 20519
rect 37473 20485 37507 20519
rect 37507 20485 37516 20519
rect 37464 20476 37516 20485
rect 39028 20476 39080 20528
rect 23756 20340 23808 20392
rect 24032 20383 24084 20392
rect 24032 20349 24041 20383
rect 24041 20349 24075 20383
rect 24075 20349 24084 20383
rect 24032 20340 24084 20349
rect 24952 20340 25004 20392
rect 28816 20383 28868 20392
rect 28816 20349 28825 20383
rect 28825 20349 28859 20383
rect 28859 20349 28868 20383
rect 28816 20340 28868 20349
rect 17224 20204 17276 20256
rect 17868 20204 17920 20256
rect 21088 20204 21140 20256
rect 22008 20272 22060 20324
rect 22560 20272 22612 20324
rect 29092 20315 29144 20324
rect 22192 20204 22244 20256
rect 22376 20204 22428 20256
rect 22928 20204 22980 20256
rect 27804 20204 27856 20256
rect 29092 20281 29101 20315
rect 29101 20281 29135 20315
rect 29135 20281 29144 20315
rect 29092 20272 29144 20281
rect 29276 20272 29328 20324
rect 30932 20408 30984 20460
rect 33232 20408 33284 20460
rect 45836 20408 45888 20460
rect 47492 20408 47544 20460
rect 31484 20340 31536 20392
rect 33784 20340 33836 20392
rect 34060 20383 34112 20392
rect 34060 20349 34069 20383
rect 34069 20349 34103 20383
rect 34103 20349 34112 20383
rect 34060 20340 34112 20349
rect 30380 20272 30432 20324
rect 31392 20272 31444 20324
rect 36544 20272 36596 20324
rect 46112 20272 46164 20324
rect 29460 20204 29512 20256
rect 30196 20204 30248 20256
rect 30748 20204 30800 20256
rect 33324 20204 33376 20256
rect 46480 20204 46532 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 8944 20000 8996 20052
rect 11704 20043 11756 20052
rect 11704 20009 11713 20043
rect 11713 20009 11747 20043
rect 11747 20009 11756 20043
rect 11704 20000 11756 20009
rect 15936 20000 15988 20052
rect 16672 20000 16724 20052
rect 18052 20000 18104 20052
rect 19616 20000 19668 20052
rect 4896 19907 4948 19916
rect 4896 19873 4905 19907
rect 4905 19873 4939 19907
rect 4939 19873 4948 19907
rect 4896 19864 4948 19873
rect 5540 19907 5592 19916
rect 5540 19873 5549 19907
rect 5549 19873 5583 19907
rect 5583 19873 5592 19907
rect 5540 19864 5592 19873
rect 8024 19864 8076 19916
rect 1768 19796 1820 19848
rect 9404 19796 9456 19848
rect 9588 19839 9640 19848
rect 9588 19805 9597 19839
rect 9597 19805 9631 19839
rect 9631 19805 9640 19839
rect 9588 19796 9640 19805
rect 9680 19839 9732 19848
rect 9680 19805 9689 19839
rect 9689 19805 9723 19839
rect 9723 19805 9732 19839
rect 9680 19796 9732 19805
rect 10232 19796 10284 19848
rect 10416 19796 10468 19848
rect 15200 19932 15252 19984
rect 17132 19932 17184 19984
rect 24032 20000 24084 20052
rect 28264 20000 28316 20052
rect 29368 20000 29420 20052
rect 30380 20043 30432 20052
rect 30380 20009 30389 20043
rect 30389 20009 30423 20043
rect 30423 20009 30432 20043
rect 30380 20000 30432 20009
rect 30564 20043 30616 20052
rect 30564 20009 30573 20043
rect 30573 20009 30607 20043
rect 30607 20009 30616 20043
rect 30564 20000 30616 20009
rect 30840 20000 30892 20052
rect 33876 20043 33928 20052
rect 16212 19864 16264 19916
rect 21732 19932 21784 19984
rect 22008 19932 22060 19984
rect 12992 19796 13044 19848
rect 15936 19796 15988 19848
rect 19340 19796 19392 19848
rect 9220 19703 9272 19712
rect 9220 19669 9229 19703
rect 9229 19669 9263 19703
rect 9263 19669 9272 19703
rect 9220 19660 9272 19669
rect 11520 19728 11572 19780
rect 14372 19771 14424 19780
rect 14372 19737 14381 19771
rect 14381 19737 14415 19771
rect 14415 19737 14424 19771
rect 14372 19728 14424 19737
rect 14556 19771 14608 19780
rect 14556 19737 14565 19771
rect 14565 19737 14599 19771
rect 14599 19737 14608 19771
rect 14556 19728 14608 19737
rect 15476 19771 15528 19780
rect 15476 19737 15510 19771
rect 15510 19737 15528 19771
rect 15476 19728 15528 19737
rect 16856 19771 16908 19780
rect 16856 19737 16865 19771
rect 16865 19737 16899 19771
rect 16899 19737 16908 19771
rect 16856 19728 16908 19737
rect 16948 19728 17000 19780
rect 10968 19660 11020 19712
rect 15108 19660 15160 19712
rect 17500 19771 17552 19780
rect 17500 19737 17509 19771
rect 17509 19737 17543 19771
rect 17543 19737 17552 19771
rect 17500 19728 17552 19737
rect 17776 19728 17828 19780
rect 18604 19771 18656 19780
rect 18604 19737 18613 19771
rect 18613 19737 18647 19771
rect 18647 19737 18656 19771
rect 18604 19728 18656 19737
rect 21088 19728 21140 19780
rect 21640 19839 21692 19848
rect 21640 19805 21649 19839
rect 21649 19805 21683 19839
rect 21683 19805 21692 19839
rect 21640 19796 21692 19805
rect 21732 19796 21784 19848
rect 31392 19932 31444 19984
rect 33876 20009 33885 20043
rect 33885 20009 33919 20043
rect 33919 20009 33928 20043
rect 33876 20000 33928 20009
rect 36544 19932 36596 19984
rect 26240 19796 26292 19848
rect 27712 19864 27764 19916
rect 28540 19907 28592 19916
rect 28540 19873 28549 19907
rect 28549 19873 28583 19907
rect 28583 19873 28592 19907
rect 28540 19864 28592 19873
rect 30196 19907 30248 19916
rect 30196 19873 30205 19907
rect 30205 19873 30239 19907
rect 30239 19873 30248 19907
rect 30196 19864 30248 19873
rect 30656 19864 30708 19916
rect 32312 19864 32364 19916
rect 46480 19907 46532 19916
rect 46480 19873 46489 19907
rect 46489 19873 46523 19907
rect 46523 19873 46532 19907
rect 46480 19864 46532 19873
rect 27344 19839 27396 19848
rect 27344 19805 27353 19839
rect 27353 19805 27387 19839
rect 27387 19805 27396 19839
rect 28448 19839 28500 19848
rect 27344 19796 27396 19805
rect 28448 19805 28457 19839
rect 28457 19805 28491 19839
rect 28491 19805 28500 19839
rect 28448 19796 28500 19805
rect 28816 19796 28868 19848
rect 29000 19796 29052 19848
rect 30288 19796 30340 19848
rect 33232 19796 33284 19848
rect 21824 19728 21876 19780
rect 19156 19660 19208 19712
rect 20812 19660 20864 19712
rect 20996 19660 21048 19712
rect 22284 19660 22336 19712
rect 23848 19728 23900 19780
rect 32128 19728 32180 19780
rect 47676 19728 47728 19780
rect 48136 19771 48188 19780
rect 48136 19737 48145 19771
rect 48145 19737 48179 19771
rect 48179 19737 48188 19771
rect 48136 19728 48188 19737
rect 23940 19660 23992 19712
rect 26976 19660 27028 19712
rect 27804 19660 27856 19712
rect 31760 19660 31812 19712
rect 32588 19660 32640 19712
rect 35624 19660 35676 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 8760 19456 8812 19508
rect 4068 19388 4120 19440
rect 1768 19363 1820 19372
rect 1768 19329 1777 19363
rect 1777 19329 1811 19363
rect 1811 19329 1820 19363
rect 1768 19320 1820 19329
rect 8024 19363 8076 19372
rect 8024 19329 8033 19363
rect 8033 19329 8067 19363
rect 8067 19329 8076 19363
rect 8024 19320 8076 19329
rect 9220 19388 9272 19440
rect 9680 19456 9732 19508
rect 11520 19499 11572 19508
rect 11520 19465 11529 19499
rect 11529 19465 11563 19499
rect 11563 19465 11572 19499
rect 11520 19456 11572 19465
rect 14096 19456 14148 19508
rect 14372 19456 14424 19508
rect 14188 19388 14240 19440
rect 14556 19388 14608 19440
rect 16856 19456 16908 19508
rect 9772 19320 9824 19372
rect 10508 19320 10560 19372
rect 11796 19363 11848 19372
rect 11796 19329 11805 19363
rect 11805 19329 11839 19363
rect 11839 19329 11848 19363
rect 11796 19320 11848 19329
rect 1952 19295 2004 19304
rect 1952 19261 1961 19295
rect 1961 19261 1995 19295
rect 1995 19261 2004 19295
rect 1952 19252 2004 19261
rect 2228 19295 2280 19304
rect 2228 19261 2237 19295
rect 2237 19261 2271 19295
rect 2271 19261 2280 19295
rect 2228 19252 2280 19261
rect 11980 19363 12032 19372
rect 11980 19329 11989 19363
rect 11989 19329 12023 19363
rect 12023 19329 12032 19363
rect 11980 19320 12032 19329
rect 12164 19363 12216 19372
rect 12164 19329 12173 19363
rect 12173 19329 12207 19363
rect 12207 19329 12216 19363
rect 12164 19320 12216 19329
rect 13544 19320 13596 19372
rect 14372 19320 14424 19372
rect 15108 19363 15160 19372
rect 15108 19329 15117 19363
rect 15117 19329 15151 19363
rect 15151 19329 15160 19363
rect 15108 19320 15160 19329
rect 16948 19388 17000 19440
rect 20996 19456 21048 19508
rect 21916 19456 21968 19508
rect 24768 19499 24820 19508
rect 24768 19465 24777 19499
rect 24777 19465 24811 19499
rect 24811 19465 24820 19499
rect 24768 19456 24820 19465
rect 19340 19388 19392 19440
rect 20812 19388 20864 19440
rect 16488 19320 16540 19372
rect 17500 19320 17552 19372
rect 18144 19320 18196 19372
rect 21088 19363 21140 19372
rect 12256 19252 12308 19304
rect 13820 19295 13872 19304
rect 13820 19261 13829 19295
rect 13829 19261 13863 19295
rect 13863 19261 13872 19295
rect 13820 19252 13872 19261
rect 15292 19252 15344 19304
rect 15384 19295 15436 19304
rect 15384 19261 15393 19295
rect 15393 19261 15427 19295
rect 15427 19261 15436 19295
rect 15384 19252 15436 19261
rect 19340 19252 19392 19304
rect 21088 19329 21097 19363
rect 21097 19329 21131 19363
rect 21131 19329 21140 19363
rect 21088 19320 21140 19329
rect 21732 19388 21784 19440
rect 22192 19388 22244 19440
rect 47768 19456 47820 19508
rect 21824 19363 21876 19372
rect 21824 19329 21833 19363
rect 21833 19329 21867 19363
rect 21867 19329 21876 19363
rect 21824 19320 21876 19329
rect 22008 19320 22060 19372
rect 22468 19320 22520 19372
rect 22928 19320 22980 19372
rect 25044 19320 25096 19372
rect 26976 19431 27028 19440
rect 26976 19397 26985 19431
rect 26985 19397 27019 19431
rect 27019 19397 27028 19431
rect 26976 19388 27028 19397
rect 27160 19431 27212 19440
rect 27160 19397 27169 19431
rect 27169 19397 27203 19431
rect 27203 19397 27212 19431
rect 27160 19388 27212 19397
rect 28448 19388 28500 19440
rect 28908 19388 28960 19440
rect 32128 19363 32180 19372
rect 32128 19329 32137 19363
rect 32137 19329 32171 19363
rect 32171 19329 32180 19363
rect 32128 19320 32180 19329
rect 16120 19184 16172 19236
rect 22192 19184 22244 19236
rect 13544 19116 13596 19168
rect 17316 19159 17368 19168
rect 17316 19125 17325 19159
rect 17325 19125 17359 19159
rect 17359 19125 17368 19159
rect 17316 19116 17368 19125
rect 17500 19116 17552 19168
rect 19432 19116 19484 19168
rect 19800 19159 19852 19168
rect 19800 19125 19809 19159
rect 19809 19125 19843 19159
rect 19843 19125 19852 19159
rect 19800 19116 19852 19125
rect 22008 19159 22060 19168
rect 22008 19125 22017 19159
rect 22017 19125 22051 19159
rect 22051 19125 22060 19159
rect 22008 19116 22060 19125
rect 23112 19116 23164 19168
rect 23572 19116 23624 19168
rect 26240 19252 26292 19304
rect 27068 19252 27120 19304
rect 27620 19184 27672 19236
rect 33140 19388 33192 19440
rect 33324 19431 33376 19440
rect 33324 19397 33333 19431
rect 33333 19397 33367 19431
rect 33367 19397 33376 19431
rect 33324 19388 33376 19397
rect 36636 19320 36688 19372
rect 47860 19363 47912 19372
rect 47860 19329 47869 19363
rect 47869 19329 47903 19363
rect 47903 19329 47912 19363
rect 47860 19320 47912 19329
rect 33600 19252 33652 19304
rect 34152 19295 34204 19304
rect 34152 19261 34161 19295
rect 34161 19261 34195 19295
rect 34195 19261 34204 19295
rect 34152 19252 34204 19261
rect 24584 19116 24636 19168
rect 36544 19159 36596 19168
rect 36544 19125 36553 19159
rect 36553 19125 36587 19159
rect 36587 19125 36596 19159
rect 36544 19116 36596 19125
rect 37464 19116 37516 19168
rect 48044 19159 48096 19168
rect 48044 19125 48053 19159
rect 48053 19125 48087 19159
rect 48087 19125 48096 19159
rect 48044 19116 48096 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 1952 18912 2004 18964
rect 2044 18844 2096 18896
rect 2412 18708 2464 18760
rect 4988 18708 5040 18760
rect 9312 18751 9364 18760
rect 9312 18717 9321 18751
rect 9321 18717 9355 18751
rect 9355 18717 9364 18751
rect 9312 18708 9364 18717
rect 9588 18776 9640 18828
rect 9496 18751 9548 18760
rect 9496 18717 9505 18751
rect 9505 18717 9539 18751
rect 9539 18717 9548 18751
rect 9496 18708 9548 18717
rect 10232 18708 10284 18760
rect 3976 18640 4028 18692
rect 12808 18776 12860 18828
rect 11888 18708 11940 18760
rect 12164 18708 12216 18760
rect 9036 18615 9088 18624
rect 9036 18581 9045 18615
rect 9045 18581 9079 18615
rect 9079 18581 9088 18615
rect 9036 18572 9088 18581
rect 11336 18615 11388 18624
rect 11336 18581 11345 18615
rect 11345 18581 11379 18615
rect 11379 18581 11388 18615
rect 11336 18572 11388 18581
rect 12256 18640 12308 18692
rect 13544 18751 13596 18760
rect 13544 18717 13553 18751
rect 13553 18717 13587 18751
rect 13587 18717 13596 18751
rect 13544 18708 13596 18717
rect 13820 18708 13872 18760
rect 14740 18708 14792 18760
rect 16120 18751 16172 18760
rect 16120 18717 16129 18751
rect 16129 18717 16163 18751
rect 16163 18717 16172 18751
rect 16120 18708 16172 18717
rect 14096 18683 14148 18692
rect 14096 18649 14105 18683
rect 14105 18649 14139 18683
rect 14139 18649 14148 18683
rect 14096 18640 14148 18649
rect 12900 18615 12952 18624
rect 12900 18581 12909 18615
rect 12909 18581 12943 18615
rect 12943 18581 12952 18615
rect 12900 18572 12952 18581
rect 15752 18572 15804 18624
rect 19800 18708 19852 18760
rect 20812 18912 20864 18964
rect 21732 18912 21784 18964
rect 22928 18912 22980 18964
rect 33416 18912 33468 18964
rect 47676 18955 47728 18964
rect 47676 18921 47685 18955
rect 47685 18921 47719 18955
rect 47719 18921 47728 18955
rect 47676 18912 47728 18921
rect 19984 18844 20036 18896
rect 20628 18844 20680 18896
rect 16856 18640 16908 18692
rect 20352 18708 20404 18760
rect 20996 18708 21048 18760
rect 22376 18776 22428 18828
rect 21732 18751 21784 18760
rect 21732 18717 21741 18751
rect 21741 18717 21775 18751
rect 21775 18717 21784 18751
rect 21732 18708 21784 18717
rect 22560 18751 22612 18760
rect 22560 18717 22569 18751
rect 22569 18717 22603 18751
rect 22603 18717 22612 18751
rect 22560 18708 22612 18717
rect 25044 18819 25096 18828
rect 25044 18785 25053 18819
rect 25053 18785 25087 18819
rect 25087 18785 25096 18819
rect 25044 18776 25096 18785
rect 24032 18708 24084 18760
rect 19340 18572 19392 18624
rect 20168 18572 20220 18624
rect 21088 18640 21140 18692
rect 23940 18640 23992 18692
rect 34704 18776 34756 18828
rect 36544 18819 36596 18828
rect 36544 18785 36553 18819
rect 36553 18785 36587 18819
rect 36587 18785 36596 18819
rect 36544 18776 36596 18785
rect 24584 18640 24636 18692
rect 26332 18708 26384 18760
rect 26792 18751 26844 18760
rect 26792 18717 26801 18751
rect 26801 18717 26835 18751
rect 26835 18717 26844 18751
rect 26792 18708 26844 18717
rect 26976 18708 27028 18760
rect 27528 18708 27580 18760
rect 28172 18708 28224 18760
rect 27896 18640 27948 18692
rect 28724 18640 28776 18692
rect 29644 18640 29696 18692
rect 35624 18708 35676 18760
rect 32220 18683 32272 18692
rect 32220 18649 32254 18683
rect 32254 18649 32272 18683
rect 32220 18640 32272 18649
rect 33140 18640 33192 18692
rect 36084 18640 36136 18692
rect 46388 18640 46440 18692
rect 20812 18572 20864 18624
rect 21272 18572 21324 18624
rect 21640 18615 21692 18624
rect 21640 18581 21649 18615
rect 21649 18581 21683 18615
rect 21683 18581 21692 18615
rect 21640 18572 21692 18581
rect 22928 18572 22980 18624
rect 23664 18572 23716 18624
rect 23848 18572 23900 18624
rect 24952 18572 25004 18624
rect 27436 18572 27488 18624
rect 29552 18615 29604 18624
rect 29552 18581 29561 18615
rect 29561 18581 29595 18615
rect 29595 18581 29604 18615
rect 29552 18572 29604 18581
rect 34520 18572 34572 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 9496 18368 9548 18420
rect 11888 18411 11940 18420
rect 11888 18377 11897 18411
rect 11897 18377 11931 18411
rect 11931 18377 11940 18411
rect 11888 18368 11940 18377
rect 14372 18411 14424 18420
rect 14372 18377 14381 18411
rect 14381 18377 14415 18411
rect 14415 18377 14424 18411
rect 14372 18368 14424 18377
rect 15936 18411 15988 18420
rect 15936 18377 15945 18411
rect 15945 18377 15979 18411
rect 15979 18377 15988 18411
rect 15936 18368 15988 18377
rect 16856 18411 16908 18420
rect 16856 18377 16865 18411
rect 16865 18377 16899 18411
rect 16899 18377 16908 18411
rect 16856 18368 16908 18377
rect 17224 18368 17276 18420
rect 22560 18368 22612 18420
rect 26056 18411 26108 18420
rect 26056 18377 26065 18411
rect 26065 18377 26099 18411
rect 26099 18377 26108 18411
rect 26056 18368 26108 18377
rect 26240 18368 26292 18420
rect 28172 18411 28224 18420
rect 28172 18377 28181 18411
rect 28181 18377 28215 18411
rect 28215 18377 28224 18411
rect 28172 18368 28224 18377
rect 8024 18300 8076 18352
rect 2136 18232 2188 18284
rect 6828 18275 6880 18284
rect 6828 18241 6837 18275
rect 6837 18241 6871 18275
rect 6871 18241 6880 18275
rect 6828 18232 6880 18241
rect 7472 18275 7524 18284
rect 7472 18241 7481 18275
rect 7481 18241 7515 18275
rect 7515 18241 7524 18275
rect 7472 18232 7524 18241
rect 9036 18232 9088 18284
rect 10140 18300 10192 18352
rect 12900 18300 12952 18352
rect 21640 18300 21692 18352
rect 22192 18300 22244 18352
rect 29552 18300 29604 18352
rect 32220 18368 32272 18420
rect 35624 18411 35676 18420
rect 1584 18028 1636 18080
rect 2872 18071 2924 18080
rect 2872 18037 2881 18071
rect 2881 18037 2915 18071
rect 2915 18037 2924 18071
rect 2872 18028 2924 18037
rect 4068 18028 4120 18080
rect 6828 18028 6880 18080
rect 6920 18071 6972 18080
rect 6920 18037 6929 18071
rect 6929 18037 6963 18071
rect 6963 18037 6972 18071
rect 6920 18028 6972 18037
rect 8208 18028 8260 18080
rect 9404 18071 9456 18080
rect 9404 18037 9413 18071
rect 9413 18037 9447 18071
rect 9447 18037 9456 18071
rect 9404 18028 9456 18037
rect 9588 18096 9640 18148
rect 9864 18275 9916 18284
rect 9864 18241 9873 18275
rect 9873 18241 9907 18275
rect 9907 18241 9916 18275
rect 9864 18232 9916 18241
rect 10232 18232 10284 18284
rect 10508 18275 10560 18284
rect 10508 18241 10517 18275
rect 10517 18241 10551 18275
rect 10551 18241 10560 18275
rect 10508 18232 10560 18241
rect 11704 18275 11756 18284
rect 11704 18241 11713 18275
rect 11713 18241 11747 18275
rect 11747 18241 11756 18275
rect 11704 18232 11756 18241
rect 12992 18275 13044 18284
rect 12992 18241 13001 18275
rect 13001 18241 13035 18275
rect 13035 18241 13044 18275
rect 12992 18232 13044 18241
rect 17040 18232 17092 18284
rect 17500 18275 17552 18284
rect 17500 18241 17509 18275
rect 17509 18241 17543 18275
rect 17543 18241 17552 18275
rect 17500 18232 17552 18241
rect 19984 18232 20036 18284
rect 20168 18275 20220 18284
rect 20168 18241 20202 18275
rect 20202 18241 20220 18275
rect 20168 18232 20220 18241
rect 18144 18096 18196 18148
rect 20168 18028 20220 18080
rect 20536 18028 20588 18080
rect 21088 18028 21140 18080
rect 21272 18071 21324 18080
rect 21272 18037 21281 18071
rect 21281 18037 21315 18071
rect 21315 18037 21324 18071
rect 21272 18028 21324 18037
rect 23664 18164 23716 18216
rect 23940 18275 23992 18284
rect 23940 18241 23949 18275
rect 23949 18241 23983 18275
rect 23983 18241 23992 18275
rect 23940 18232 23992 18241
rect 24216 18232 24268 18284
rect 25044 18275 25096 18284
rect 25044 18241 25053 18275
rect 25053 18241 25087 18275
rect 25087 18241 25096 18275
rect 25044 18232 25096 18241
rect 25320 18232 25372 18284
rect 25872 18232 25924 18284
rect 26148 18207 26200 18216
rect 23848 18096 23900 18148
rect 24032 18096 24084 18148
rect 26148 18173 26157 18207
rect 26157 18173 26191 18207
rect 26191 18173 26200 18207
rect 26148 18164 26200 18173
rect 26332 18207 26384 18216
rect 26332 18173 26341 18207
rect 26341 18173 26375 18207
rect 26375 18173 26384 18207
rect 26332 18164 26384 18173
rect 26700 18164 26752 18216
rect 27252 18275 27304 18284
rect 27252 18241 27258 18275
rect 27258 18241 27292 18275
rect 27292 18241 27304 18275
rect 27252 18232 27304 18241
rect 27712 18207 27764 18216
rect 27712 18173 27721 18207
rect 27721 18173 27755 18207
rect 27755 18173 27764 18207
rect 27712 18164 27764 18173
rect 28172 18232 28224 18284
rect 28356 18232 28408 18284
rect 25780 18096 25832 18148
rect 28724 18207 28776 18216
rect 28724 18173 28733 18207
rect 28733 18173 28767 18207
rect 28767 18173 28776 18207
rect 28724 18164 28776 18173
rect 24584 18028 24636 18080
rect 25596 18028 25648 18080
rect 27436 18028 27488 18080
rect 27988 18028 28040 18080
rect 28724 18028 28776 18080
rect 30840 18232 30892 18284
rect 35624 18377 35633 18411
rect 35633 18377 35667 18411
rect 35667 18377 35676 18411
rect 35624 18368 35676 18377
rect 36636 18300 36688 18352
rect 37464 18343 37516 18352
rect 37464 18309 37473 18343
rect 37473 18309 37507 18343
rect 37507 18309 37516 18343
rect 37464 18300 37516 18309
rect 40132 18300 40184 18352
rect 32772 18275 32824 18284
rect 32772 18241 32781 18275
rect 32781 18241 32815 18275
rect 32815 18241 32824 18275
rect 32772 18232 32824 18241
rect 33140 18232 33192 18284
rect 33416 18275 33468 18284
rect 33416 18241 33425 18275
rect 33425 18241 33459 18275
rect 33459 18241 33468 18275
rect 33416 18232 33468 18241
rect 34796 18232 34848 18284
rect 36084 18275 36136 18284
rect 36084 18241 36093 18275
rect 36093 18241 36127 18275
rect 36127 18241 36136 18275
rect 36084 18232 36136 18241
rect 36176 18232 36228 18284
rect 33692 18164 33744 18216
rect 32496 18096 32548 18148
rect 29552 18028 29604 18080
rect 34612 18028 34664 18080
rect 35348 18028 35400 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 9956 17824 10008 17876
rect 2872 17756 2924 17808
rect 1584 17731 1636 17740
rect 1584 17697 1593 17731
rect 1593 17697 1627 17731
rect 1627 17697 1636 17731
rect 1584 17688 1636 17697
rect 2780 17731 2832 17740
rect 2780 17697 2789 17731
rect 2789 17697 2823 17731
rect 2823 17697 2832 17731
rect 7472 17756 7524 17808
rect 17868 17824 17920 17876
rect 18144 17799 18196 17808
rect 2780 17688 2832 17697
rect 6828 17688 6880 17740
rect 15752 17731 15804 17740
rect 15752 17697 15761 17731
rect 15761 17697 15795 17731
rect 15795 17697 15804 17731
rect 15752 17688 15804 17697
rect 18144 17765 18153 17799
rect 18153 17765 18187 17799
rect 18187 17765 18196 17799
rect 18144 17756 18196 17765
rect 25228 17824 25280 17876
rect 25596 17867 25648 17876
rect 25596 17833 25605 17867
rect 25605 17833 25639 17867
rect 25639 17833 25648 17867
rect 25596 17824 25648 17833
rect 26240 17867 26292 17876
rect 26240 17833 26249 17867
rect 26249 17833 26283 17867
rect 26283 17833 26292 17867
rect 26240 17824 26292 17833
rect 26424 17824 26476 17876
rect 29920 17824 29972 17876
rect 34796 17824 34848 17876
rect 36176 17867 36228 17876
rect 36176 17833 36185 17867
rect 36185 17833 36219 17867
rect 36219 17833 36228 17867
rect 36176 17824 36228 17833
rect 26332 17756 26384 17808
rect 24584 17731 24636 17740
rect 12440 17620 12492 17672
rect 12992 17620 13044 17672
rect 15568 17663 15620 17672
rect 15568 17629 15577 17663
rect 15577 17629 15611 17663
rect 15611 17629 15620 17663
rect 15568 17620 15620 17629
rect 6920 17552 6972 17604
rect 9404 17552 9456 17604
rect 11336 17552 11388 17604
rect 15200 17552 15252 17604
rect 17960 17595 18012 17604
rect 17960 17561 17969 17595
rect 17969 17561 18003 17595
rect 18003 17561 18012 17595
rect 17960 17552 18012 17561
rect 19340 17620 19392 17672
rect 24584 17697 24593 17731
rect 24593 17697 24627 17731
rect 24627 17697 24636 17731
rect 24584 17688 24636 17697
rect 24860 17620 24912 17672
rect 25044 17620 25096 17672
rect 25504 17663 25556 17672
rect 25504 17629 25513 17663
rect 25513 17629 25547 17663
rect 25547 17629 25556 17663
rect 25504 17620 25556 17629
rect 25872 17688 25924 17740
rect 26700 17756 26752 17808
rect 27344 17756 27396 17808
rect 27712 17688 27764 17740
rect 27804 17688 27856 17740
rect 26240 17620 26292 17672
rect 26424 17663 26476 17672
rect 26424 17629 26433 17663
rect 26433 17629 26467 17663
rect 26467 17629 26476 17663
rect 26424 17620 26476 17629
rect 26792 17620 26844 17672
rect 27068 17620 27120 17672
rect 28632 17620 28684 17672
rect 29552 17663 29604 17672
rect 29552 17629 29561 17663
rect 29561 17629 29595 17663
rect 29595 17629 29604 17663
rect 29552 17620 29604 17629
rect 32496 17688 32548 17740
rect 34428 17756 34480 17808
rect 31668 17620 31720 17672
rect 31760 17620 31812 17672
rect 31944 17620 31996 17672
rect 34520 17688 34572 17740
rect 35900 17688 35952 17740
rect 39120 17731 39172 17740
rect 39120 17697 39129 17731
rect 39129 17697 39163 17731
rect 39163 17697 39172 17731
rect 39120 17688 39172 17697
rect 33692 17620 33744 17672
rect 34612 17620 34664 17672
rect 36636 17663 36688 17672
rect 36636 17629 36645 17663
rect 36645 17629 36679 17663
rect 36679 17629 36688 17663
rect 36636 17620 36688 17629
rect 47124 17620 47176 17672
rect 9588 17484 9640 17536
rect 11520 17484 11572 17536
rect 11704 17484 11756 17536
rect 15108 17527 15160 17536
rect 15108 17493 15117 17527
rect 15117 17493 15151 17527
rect 15151 17493 15160 17527
rect 15108 17484 15160 17493
rect 19432 17484 19484 17536
rect 20076 17552 20128 17604
rect 20812 17552 20864 17604
rect 24492 17595 24544 17604
rect 24492 17561 24501 17595
rect 24501 17561 24535 17595
rect 24535 17561 24544 17595
rect 24492 17552 24544 17561
rect 26884 17552 26936 17604
rect 26976 17552 27028 17604
rect 29460 17552 29512 17604
rect 29828 17595 29880 17604
rect 29828 17561 29840 17595
rect 29840 17561 29880 17595
rect 29828 17552 29880 17561
rect 29920 17552 29972 17604
rect 19984 17484 20036 17536
rect 21732 17527 21784 17536
rect 21732 17493 21741 17527
rect 21741 17493 21775 17527
rect 21775 17493 21784 17527
rect 21732 17484 21784 17493
rect 24124 17484 24176 17536
rect 24584 17484 24636 17536
rect 24860 17484 24912 17536
rect 25228 17484 25280 17536
rect 27988 17484 28040 17536
rect 30932 17527 30984 17536
rect 30932 17493 30941 17527
rect 30941 17493 30975 17527
rect 30975 17493 30984 17527
rect 30932 17484 30984 17493
rect 33968 17552 34020 17604
rect 46848 17484 46900 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 23388 17280 23440 17332
rect 1860 17187 1912 17196
rect 1860 17153 1869 17187
rect 1869 17153 1903 17187
rect 1903 17153 1912 17187
rect 1860 17144 1912 17153
rect 9588 17187 9640 17196
rect 9588 17153 9597 17187
rect 9597 17153 9631 17187
rect 9631 17153 9640 17187
rect 9588 17144 9640 17153
rect 9864 17212 9916 17264
rect 20812 17255 20864 17264
rect 10508 17144 10560 17196
rect 3700 17076 3752 17128
rect 12992 17144 13044 17196
rect 14648 17144 14700 17196
rect 16856 17144 16908 17196
rect 20352 17187 20404 17196
rect 16672 17076 16724 17128
rect 19892 17076 19944 17128
rect 20352 17153 20361 17187
rect 20361 17153 20395 17187
rect 20395 17153 20404 17187
rect 20352 17144 20404 17153
rect 20812 17221 20821 17255
rect 20821 17221 20855 17255
rect 20855 17221 20864 17255
rect 20812 17212 20864 17221
rect 21732 17212 21784 17264
rect 23480 17255 23532 17264
rect 23480 17221 23489 17255
rect 23489 17221 23523 17255
rect 23523 17221 23532 17255
rect 23664 17280 23716 17332
rect 23940 17280 23992 17332
rect 24124 17280 24176 17332
rect 24400 17280 24452 17332
rect 24492 17280 24544 17332
rect 25872 17323 25924 17332
rect 25872 17289 25881 17323
rect 25881 17289 25915 17323
rect 25915 17289 25924 17323
rect 25872 17280 25924 17289
rect 27252 17323 27304 17332
rect 27252 17289 27261 17323
rect 27261 17289 27295 17323
rect 27295 17289 27304 17323
rect 27252 17280 27304 17289
rect 27712 17323 27764 17332
rect 27712 17289 27721 17323
rect 27721 17289 27755 17323
rect 27755 17289 27764 17323
rect 27712 17280 27764 17289
rect 27988 17280 28040 17332
rect 29828 17280 29880 17332
rect 33968 17280 34020 17332
rect 23480 17212 23532 17221
rect 23020 17144 23072 17196
rect 23388 17187 23440 17196
rect 23388 17153 23395 17187
rect 23395 17153 23440 17187
rect 23388 17144 23440 17153
rect 29000 17212 29052 17264
rect 35348 17280 35400 17332
rect 25504 17187 25556 17196
rect 25504 17153 25513 17187
rect 25513 17153 25547 17187
rect 25547 17153 25556 17187
rect 25504 17144 25556 17153
rect 25596 17144 25648 17196
rect 15568 17008 15620 17060
rect 20076 17008 20128 17060
rect 20812 17008 20864 17060
rect 25136 17076 25188 17128
rect 26424 17144 26476 17196
rect 26976 17187 27028 17196
rect 26976 17153 26985 17187
rect 26985 17153 27019 17187
rect 27019 17153 27028 17187
rect 26976 17144 27028 17153
rect 27068 17187 27120 17196
rect 27068 17153 27077 17187
rect 27077 17153 27111 17187
rect 27111 17153 27120 17187
rect 27068 17144 27120 17153
rect 27528 17144 27580 17196
rect 28908 17187 28960 17196
rect 18328 16940 18380 16992
rect 25228 17008 25280 17060
rect 23848 16983 23900 16992
rect 23848 16949 23857 16983
rect 23857 16949 23891 16983
rect 23891 16949 23900 16983
rect 23848 16940 23900 16949
rect 24216 16940 24268 16992
rect 25780 17051 25832 17060
rect 25780 17017 25789 17051
rect 25789 17017 25823 17051
rect 25823 17017 25832 17051
rect 28632 17076 28684 17128
rect 28908 17153 28917 17187
rect 28917 17153 28951 17187
rect 28951 17153 28960 17187
rect 28908 17144 28960 17153
rect 29092 17185 29144 17196
rect 29092 17151 29101 17185
rect 29101 17151 29135 17185
rect 29135 17151 29144 17185
rect 29460 17187 29512 17196
rect 29092 17144 29144 17151
rect 29460 17153 29469 17187
rect 29469 17153 29503 17187
rect 29503 17153 29512 17187
rect 29460 17144 29512 17153
rect 31944 17144 31996 17196
rect 32312 17187 32364 17196
rect 32312 17153 32321 17187
rect 32321 17153 32355 17187
rect 32355 17153 32364 17187
rect 32312 17144 32364 17153
rect 29000 17076 29052 17128
rect 25780 17008 25832 17017
rect 27988 17008 28040 17060
rect 29644 17076 29696 17128
rect 31668 17076 31720 17128
rect 34520 17187 34572 17196
rect 34520 17153 34529 17187
rect 34529 17153 34563 17187
rect 34563 17153 34572 17187
rect 35256 17187 35308 17196
rect 34520 17144 34572 17153
rect 35256 17153 35265 17187
rect 35265 17153 35299 17187
rect 35299 17153 35308 17187
rect 35256 17144 35308 17153
rect 34428 17076 34480 17128
rect 35624 17187 35676 17196
rect 35624 17153 35633 17187
rect 35633 17153 35667 17187
rect 35667 17153 35676 17187
rect 36084 17187 36136 17196
rect 35624 17144 35676 17153
rect 36084 17153 36093 17187
rect 36093 17153 36127 17187
rect 36127 17153 36136 17187
rect 36084 17144 36136 17153
rect 36268 17187 36320 17196
rect 36268 17153 36277 17187
rect 36277 17153 36311 17187
rect 36311 17153 36320 17187
rect 36268 17144 36320 17153
rect 36636 17144 36688 17196
rect 30932 17008 30984 17060
rect 26332 16940 26384 16992
rect 31024 16940 31076 16992
rect 31300 16940 31352 16992
rect 33140 16940 33192 16992
rect 34796 16940 34848 16992
rect 37372 16983 37424 16992
rect 37372 16949 37381 16983
rect 37381 16949 37415 16983
rect 37415 16949 37424 16983
rect 37372 16940 37424 16949
rect 46480 16940 46532 16992
rect 47768 16983 47820 16992
rect 47768 16949 47777 16983
rect 47777 16949 47811 16983
rect 47811 16949 47820 16983
rect 47768 16940 47820 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 14648 16736 14700 16788
rect 16856 16779 16908 16788
rect 2044 16532 2096 16584
rect 12072 16668 12124 16720
rect 11612 16532 11664 16584
rect 14832 16668 14884 16720
rect 14740 16600 14792 16652
rect 13728 16532 13780 16584
rect 15108 16532 15160 16584
rect 10140 16507 10192 16516
rect 10140 16473 10149 16507
rect 10149 16473 10183 16507
rect 10183 16473 10192 16507
rect 10140 16464 10192 16473
rect 15384 16532 15436 16584
rect 16856 16745 16865 16779
rect 16865 16745 16899 16779
rect 16899 16745 16908 16779
rect 16856 16736 16908 16745
rect 17960 16736 18012 16788
rect 18512 16736 18564 16788
rect 19432 16736 19484 16788
rect 20812 16736 20864 16788
rect 24216 16736 24268 16788
rect 24400 16779 24452 16788
rect 24400 16745 24409 16779
rect 24409 16745 24443 16779
rect 24443 16745 24452 16779
rect 24400 16736 24452 16745
rect 28908 16736 28960 16788
rect 16396 16600 16448 16652
rect 2228 16396 2280 16448
rect 15200 16396 15252 16448
rect 15660 16439 15712 16448
rect 15660 16405 15669 16439
rect 15669 16405 15703 16439
rect 15703 16405 15712 16439
rect 15660 16396 15712 16405
rect 16396 16464 16448 16516
rect 17316 16575 17368 16584
rect 17316 16541 17325 16575
rect 17325 16541 17359 16575
rect 17359 16541 17368 16575
rect 25228 16668 25280 16720
rect 35900 16736 35952 16788
rect 36268 16736 36320 16788
rect 19248 16643 19300 16652
rect 19248 16609 19257 16643
rect 19257 16609 19291 16643
rect 19291 16609 19300 16643
rect 19248 16600 19300 16609
rect 22468 16643 22520 16652
rect 22468 16609 22477 16643
rect 22477 16609 22511 16643
rect 22511 16609 22520 16643
rect 22468 16600 22520 16609
rect 27988 16600 28040 16652
rect 31300 16600 31352 16652
rect 17316 16532 17368 16541
rect 17868 16532 17920 16584
rect 19340 16464 19392 16516
rect 19064 16396 19116 16448
rect 19892 16464 19944 16516
rect 20076 16464 20128 16516
rect 23848 16532 23900 16584
rect 24860 16532 24912 16584
rect 26884 16575 26936 16584
rect 26884 16541 26893 16575
rect 26893 16541 26927 16575
rect 26927 16541 26936 16575
rect 26884 16532 26936 16541
rect 27068 16532 27120 16584
rect 27620 16532 27672 16584
rect 28908 16532 28960 16584
rect 32496 16600 32548 16652
rect 34704 16643 34756 16652
rect 34704 16609 34713 16643
rect 34713 16609 34747 16643
rect 34747 16609 34756 16643
rect 34704 16600 34756 16609
rect 38568 16643 38620 16652
rect 38568 16609 38577 16643
rect 38577 16609 38611 16643
rect 38611 16609 38620 16643
rect 38568 16600 38620 16609
rect 47768 16668 47820 16720
rect 46480 16643 46532 16652
rect 46480 16609 46489 16643
rect 46489 16609 46523 16643
rect 46523 16609 46532 16643
rect 46480 16600 46532 16609
rect 48136 16643 48188 16652
rect 48136 16609 48145 16643
rect 48145 16609 48179 16643
rect 48179 16609 48188 16643
rect 48136 16600 48188 16609
rect 23940 16464 23992 16516
rect 24216 16464 24268 16516
rect 24400 16507 24452 16516
rect 24400 16473 24409 16507
rect 24409 16473 24443 16507
rect 24443 16473 24452 16507
rect 24400 16464 24452 16473
rect 24492 16464 24544 16516
rect 23112 16396 23164 16448
rect 23664 16396 23716 16448
rect 25504 16396 25556 16448
rect 26148 16396 26200 16448
rect 27160 16396 27212 16448
rect 31944 16439 31996 16448
rect 31944 16405 31953 16439
rect 31953 16405 31987 16439
rect 31987 16405 31996 16439
rect 31944 16396 31996 16405
rect 32772 16532 32824 16584
rect 32864 16532 32916 16584
rect 34796 16532 34848 16584
rect 33140 16464 33192 16516
rect 37372 16464 37424 16516
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 10140 16235 10192 16244
rect 10140 16201 10149 16235
rect 10149 16201 10183 16235
rect 10183 16201 10192 16235
rect 10140 16192 10192 16201
rect 13728 16235 13780 16244
rect 13728 16201 13737 16235
rect 13737 16201 13771 16235
rect 13771 16201 13780 16235
rect 13728 16192 13780 16201
rect 17316 16192 17368 16244
rect 17868 16235 17920 16244
rect 17868 16201 17877 16235
rect 17877 16201 17911 16235
rect 17911 16201 17920 16235
rect 17868 16192 17920 16201
rect 19064 16192 19116 16244
rect 2228 16167 2280 16176
rect 2228 16133 2237 16167
rect 2237 16133 2271 16167
rect 2271 16133 2280 16167
rect 2228 16124 2280 16133
rect 2044 16099 2096 16108
rect 2044 16065 2053 16099
rect 2053 16065 2087 16099
rect 2087 16065 2096 16099
rect 2044 16056 2096 16065
rect 9680 16056 9732 16108
rect 12440 16124 12492 16176
rect 15660 16124 15712 16176
rect 18328 16124 18380 16176
rect 14464 16099 14516 16108
rect 14464 16065 14473 16099
rect 14473 16065 14507 16099
rect 14507 16065 14516 16099
rect 14464 16056 14516 16065
rect 14832 16056 14884 16108
rect 16396 16056 16448 16108
rect 17316 16056 17368 16108
rect 17868 16056 17920 16108
rect 18420 16056 18472 16108
rect 20076 16192 20128 16244
rect 20904 16235 20956 16244
rect 20904 16201 20913 16235
rect 20913 16201 20947 16235
rect 20947 16201 20956 16235
rect 20904 16192 20956 16201
rect 21272 16192 21324 16244
rect 23756 16192 23808 16244
rect 19984 16124 20036 16176
rect 24952 16124 25004 16176
rect 19524 16056 19576 16108
rect 20352 16056 20404 16108
rect 20720 16099 20772 16108
rect 20720 16065 20729 16099
rect 20729 16065 20763 16099
rect 20763 16065 20772 16099
rect 20720 16056 20772 16065
rect 22284 16056 22336 16108
rect 24768 16056 24820 16108
rect 2780 16031 2832 16040
rect 2780 15997 2789 16031
rect 2789 15997 2823 16031
rect 2823 15997 2832 16031
rect 14188 16031 14240 16040
rect 2780 15988 2832 15997
rect 14188 15997 14197 16031
rect 14197 15997 14231 16031
rect 14231 15997 14240 16031
rect 14188 15988 14240 15997
rect 20076 15988 20128 16040
rect 21456 15988 21508 16040
rect 24492 16031 24544 16040
rect 24492 15997 24501 16031
rect 24501 15997 24535 16031
rect 24535 15997 24544 16031
rect 24492 15988 24544 15997
rect 26700 16192 26752 16244
rect 31024 16192 31076 16244
rect 30380 16124 30432 16176
rect 31944 16124 31996 16176
rect 27252 16099 27304 16108
rect 27252 16065 27261 16099
rect 27261 16065 27295 16099
rect 27295 16065 27304 16099
rect 27252 16056 27304 16065
rect 28356 16099 28408 16108
rect 28356 16065 28365 16099
rect 28365 16065 28399 16099
rect 28399 16065 28408 16099
rect 28356 16056 28408 16065
rect 29000 16099 29052 16108
rect 29000 16065 29009 16099
rect 29009 16065 29043 16099
rect 29043 16065 29052 16099
rect 29000 16056 29052 16065
rect 29092 16056 29144 16108
rect 29552 16099 29604 16108
rect 29552 16065 29561 16099
rect 29561 16065 29595 16099
rect 29595 16065 29604 16099
rect 29552 16056 29604 16065
rect 30840 16056 30892 16108
rect 32956 16056 33008 16108
rect 47584 16099 47636 16108
rect 47584 16065 47593 16099
rect 47593 16065 47627 16099
rect 47627 16065 47636 16099
rect 47584 16056 47636 16065
rect 17868 15920 17920 15972
rect 24860 15920 24912 15972
rect 29644 15988 29696 16040
rect 30472 15920 30524 15972
rect 24768 15852 24820 15904
rect 25044 15852 25096 15904
rect 27344 15895 27396 15904
rect 27344 15861 27353 15895
rect 27353 15861 27387 15895
rect 27387 15861 27396 15895
rect 27344 15852 27396 15861
rect 27896 15852 27948 15904
rect 29736 15895 29788 15904
rect 29736 15861 29745 15895
rect 29745 15861 29779 15895
rect 29779 15861 29788 15895
rect 29736 15852 29788 15861
rect 29828 15852 29880 15904
rect 32864 15852 32916 15904
rect 47032 15895 47084 15904
rect 47032 15861 47041 15895
rect 47041 15861 47075 15895
rect 47075 15861 47084 15895
rect 47032 15852 47084 15861
rect 47676 15895 47728 15904
rect 47676 15861 47685 15895
rect 47685 15861 47719 15895
rect 47719 15861 47728 15895
rect 47676 15852 47728 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 15200 15691 15252 15700
rect 15200 15657 15209 15691
rect 15209 15657 15243 15691
rect 15243 15657 15252 15691
rect 15200 15648 15252 15657
rect 17316 15648 17368 15700
rect 20352 15648 20404 15700
rect 1676 15580 1728 15632
rect 24952 15648 25004 15700
rect 27344 15648 27396 15700
rect 27988 15648 28040 15700
rect 30012 15648 30064 15700
rect 9588 15512 9640 15564
rect 10968 15555 11020 15564
rect 10968 15521 10977 15555
rect 10977 15521 11011 15555
rect 11011 15521 11020 15555
rect 10968 15512 11020 15521
rect 11520 15555 11572 15564
rect 11520 15521 11529 15555
rect 11529 15521 11563 15555
rect 11563 15521 11572 15555
rect 11520 15512 11572 15521
rect 9404 15419 9456 15428
rect 9404 15385 9413 15419
rect 9413 15385 9447 15419
rect 9447 15385 9456 15419
rect 9404 15376 9456 15385
rect 11704 15419 11756 15428
rect 11704 15385 11713 15419
rect 11713 15385 11747 15419
rect 11747 15385 11756 15419
rect 11704 15376 11756 15385
rect 13268 15376 13320 15428
rect 10232 15308 10284 15360
rect 14280 15444 14332 15496
rect 14464 15447 14470 15474
rect 14470 15447 14504 15474
rect 14504 15447 14516 15474
rect 14464 15422 14516 15447
rect 14648 15444 14700 15496
rect 16396 15512 16448 15564
rect 15292 15444 15344 15496
rect 16488 15487 16540 15496
rect 16488 15453 16497 15487
rect 16497 15453 16531 15487
rect 16531 15453 16540 15487
rect 16488 15444 16540 15453
rect 20720 15512 20772 15564
rect 19524 15487 19576 15496
rect 19524 15453 19533 15487
rect 19533 15453 19567 15487
rect 19567 15453 19576 15487
rect 19524 15444 19576 15453
rect 26148 15580 26200 15632
rect 28632 15580 28684 15632
rect 24124 15512 24176 15564
rect 17316 15419 17368 15428
rect 17316 15385 17325 15419
rect 17325 15385 17359 15419
rect 17359 15385 17368 15419
rect 17316 15376 17368 15385
rect 17500 15419 17552 15428
rect 17500 15385 17509 15419
rect 17509 15385 17543 15419
rect 17543 15385 17552 15419
rect 17500 15376 17552 15385
rect 17868 15376 17920 15428
rect 20904 15447 20910 15474
rect 20910 15447 20944 15474
rect 20944 15447 20956 15474
rect 20904 15422 20956 15447
rect 21916 15444 21968 15496
rect 23664 15444 23716 15496
rect 24768 15444 24820 15496
rect 21548 15376 21600 15428
rect 21824 15419 21876 15428
rect 21824 15385 21833 15419
rect 21833 15385 21867 15419
rect 21867 15385 21876 15419
rect 21824 15376 21876 15385
rect 24492 15376 24544 15428
rect 24952 15487 25004 15496
rect 24952 15453 24961 15487
rect 24961 15453 24995 15487
rect 24995 15453 25004 15487
rect 27528 15512 27580 15564
rect 29460 15512 29512 15564
rect 29736 15512 29788 15564
rect 24952 15444 25004 15453
rect 26516 15444 26568 15496
rect 26884 15487 26936 15496
rect 26884 15453 26893 15487
rect 26893 15453 26927 15487
rect 26927 15453 26936 15487
rect 26884 15444 26936 15453
rect 27068 15444 27120 15496
rect 29828 15487 29880 15496
rect 27804 15376 27856 15428
rect 29828 15453 29837 15487
rect 29837 15453 29871 15487
rect 29871 15453 29880 15487
rect 29828 15444 29880 15453
rect 30380 15444 30432 15496
rect 47124 15580 47176 15632
rect 47676 15512 47728 15564
rect 48136 15555 48188 15564
rect 48136 15521 48145 15555
rect 48145 15521 48179 15555
rect 48179 15521 48188 15555
rect 48136 15512 48188 15521
rect 34520 15444 34572 15496
rect 29552 15376 29604 15428
rect 31024 15376 31076 15428
rect 32956 15376 33008 15428
rect 36544 15376 36596 15428
rect 14096 15351 14148 15360
rect 14096 15317 14105 15351
rect 14105 15317 14139 15351
rect 14139 15317 14148 15351
rect 14096 15308 14148 15317
rect 16948 15308 17000 15360
rect 17224 15308 17276 15360
rect 20904 15308 20956 15360
rect 22008 15351 22060 15360
rect 22008 15317 22017 15351
rect 22017 15317 22051 15351
rect 22051 15317 22060 15351
rect 22008 15308 22060 15317
rect 24400 15351 24452 15360
rect 24400 15317 24409 15351
rect 24409 15317 24443 15351
rect 24443 15317 24452 15351
rect 24400 15308 24452 15317
rect 26424 15351 26476 15360
rect 26424 15317 26433 15351
rect 26433 15317 26467 15351
rect 26467 15317 26476 15351
rect 26424 15308 26476 15317
rect 26516 15308 26568 15360
rect 27252 15308 27304 15360
rect 30472 15308 30524 15360
rect 32772 15308 32824 15360
rect 33140 15308 33192 15360
rect 35624 15308 35676 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 9404 15104 9456 15156
rect 11704 15104 11756 15156
rect 13728 15104 13780 15156
rect 7932 15036 7984 15088
rect 9680 14968 9732 15020
rect 14280 15036 14332 15088
rect 14648 15104 14700 15156
rect 17500 15104 17552 15156
rect 21548 15104 21600 15156
rect 25504 15104 25556 15156
rect 26240 15104 26292 15156
rect 27160 15104 27212 15156
rect 27528 15147 27580 15156
rect 16948 15079 17000 15088
rect 16948 15045 16982 15079
rect 16982 15045 17000 15079
rect 16948 15036 17000 15045
rect 14096 14968 14148 15020
rect 16672 15011 16724 15020
rect 16672 14977 16681 15011
rect 16681 14977 16715 15011
rect 16715 14977 16724 15011
rect 16672 14968 16724 14977
rect 17960 14968 18012 15020
rect 18604 14968 18656 15020
rect 19432 14968 19484 15020
rect 19892 15011 19944 15020
rect 19892 14977 19901 15011
rect 19901 14977 19935 15011
rect 19935 14977 19944 15011
rect 19892 14968 19944 14977
rect 19984 14968 20036 15020
rect 21916 14968 21968 15020
rect 27068 15036 27120 15088
rect 27528 15113 27537 15147
rect 27537 15113 27571 15147
rect 27571 15113 27580 15147
rect 27528 15104 27580 15113
rect 27804 15104 27856 15156
rect 28908 15104 28960 15156
rect 28724 15036 28776 15088
rect 22192 14968 22244 15020
rect 22284 14968 22336 15020
rect 26056 15011 26108 15020
rect 26056 14977 26065 15011
rect 26065 14977 26099 15011
rect 26099 14977 26108 15011
rect 26056 14968 26108 14977
rect 26424 14968 26476 15020
rect 26608 14968 26660 15020
rect 27804 14968 27856 15020
rect 15200 14900 15252 14952
rect 20996 14900 21048 14952
rect 26240 14943 26292 14952
rect 21824 14832 21876 14884
rect 13728 14807 13780 14816
rect 13728 14773 13737 14807
rect 13737 14773 13771 14807
rect 13771 14773 13780 14807
rect 13728 14764 13780 14773
rect 18604 14807 18656 14816
rect 18604 14773 18613 14807
rect 18613 14773 18647 14807
rect 18647 14773 18656 14807
rect 18604 14764 18656 14773
rect 22468 14832 22520 14884
rect 26240 14909 26249 14943
rect 26249 14909 26283 14943
rect 26283 14909 26292 14943
rect 26240 14900 26292 14909
rect 26332 14943 26384 14952
rect 26332 14909 26341 14943
rect 26341 14909 26375 14943
rect 26375 14909 26384 14943
rect 26332 14900 26384 14909
rect 26516 14900 26568 14952
rect 29184 14968 29236 15020
rect 30840 15104 30892 15156
rect 30932 15147 30984 15156
rect 30932 15113 30941 15147
rect 30941 15113 30975 15147
rect 30975 15113 30984 15147
rect 30932 15104 30984 15113
rect 31116 15104 31168 15156
rect 30472 15079 30524 15088
rect 30472 15045 30481 15079
rect 30481 15045 30515 15079
rect 30515 15045 30524 15079
rect 30472 15036 30524 15045
rect 47952 15104 48004 15156
rect 28632 14900 28684 14952
rect 29092 14900 29144 14952
rect 47860 15036 47912 15088
rect 29552 14943 29604 14952
rect 29552 14909 29561 14943
rect 29561 14909 29595 14943
rect 29595 14909 29604 14943
rect 29552 14900 29604 14909
rect 29644 14943 29696 14952
rect 29644 14909 29653 14943
rect 29653 14909 29687 14943
rect 29687 14909 29696 14943
rect 29644 14900 29696 14909
rect 25136 14764 25188 14816
rect 29736 14832 29788 14884
rect 26792 14764 26844 14816
rect 26976 14764 27028 14816
rect 27620 14764 27672 14816
rect 29276 14764 29328 14816
rect 30656 14968 30708 15020
rect 32496 14968 32548 15020
rect 30288 14900 30340 14952
rect 31668 14900 31720 14952
rect 32220 14900 32272 14952
rect 32588 14900 32640 14952
rect 32312 14832 32364 14884
rect 30104 14764 30156 14816
rect 30380 14764 30432 14816
rect 32496 14764 32548 14816
rect 33140 14968 33192 15020
rect 35440 15011 35492 15020
rect 35440 14977 35474 15011
rect 35474 14977 35492 15011
rect 35440 14968 35492 14977
rect 43536 14968 43588 15020
rect 47584 14968 47636 15020
rect 47952 15011 48004 15020
rect 47952 14977 47961 15011
rect 47961 14977 47995 15011
rect 47995 14977 48004 15011
rect 47952 14968 48004 14977
rect 34612 14900 34664 14952
rect 36544 14807 36596 14816
rect 36544 14773 36553 14807
rect 36553 14773 36587 14807
rect 36587 14773 36596 14807
rect 36544 14764 36596 14773
rect 46480 14764 46532 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 19340 14560 19392 14612
rect 3148 14492 3200 14544
rect 9680 14424 9732 14476
rect 12532 14424 12584 14476
rect 17960 14424 18012 14476
rect 14924 14399 14976 14408
rect 14924 14365 14933 14399
rect 14933 14365 14967 14399
rect 14967 14365 14976 14399
rect 14924 14356 14976 14365
rect 18512 14399 18564 14408
rect 18512 14365 18521 14399
rect 18521 14365 18555 14399
rect 18555 14365 18564 14399
rect 18512 14356 18564 14365
rect 19984 14492 20036 14544
rect 22192 14535 22244 14544
rect 22192 14501 22201 14535
rect 22201 14501 22235 14535
rect 22235 14501 22244 14535
rect 22192 14492 22244 14501
rect 19892 14424 19944 14476
rect 20352 14399 20404 14408
rect 15200 14288 15252 14340
rect 18696 14331 18748 14340
rect 18696 14297 18705 14331
rect 18705 14297 18739 14331
rect 18739 14297 18748 14331
rect 18696 14288 18748 14297
rect 12624 14220 12676 14272
rect 14096 14220 14148 14272
rect 20352 14365 20361 14399
rect 20361 14365 20395 14399
rect 20395 14365 20404 14399
rect 20352 14356 20404 14365
rect 20904 14356 20956 14408
rect 22744 14399 22796 14408
rect 22744 14365 22753 14399
rect 22753 14365 22787 14399
rect 22787 14365 22796 14399
rect 22744 14356 22796 14365
rect 22008 14288 22060 14340
rect 23020 14560 23072 14612
rect 23480 14492 23532 14544
rect 24768 14492 24820 14544
rect 26516 14492 26568 14544
rect 29000 14560 29052 14612
rect 29552 14560 29604 14612
rect 30656 14560 30708 14612
rect 35440 14560 35492 14612
rect 35532 14560 35584 14612
rect 30012 14492 30064 14544
rect 31944 14492 31996 14544
rect 32680 14492 32732 14544
rect 23388 14356 23440 14408
rect 29828 14424 29880 14476
rect 27620 14356 27672 14408
rect 27896 14399 27948 14408
rect 27896 14365 27905 14399
rect 27905 14365 27939 14399
rect 27939 14365 27948 14399
rect 27896 14356 27948 14365
rect 27988 14356 28040 14408
rect 26148 14288 26200 14340
rect 26976 14331 27028 14340
rect 26976 14297 26985 14331
rect 26985 14297 27019 14331
rect 27019 14297 27028 14331
rect 26976 14288 27028 14297
rect 28908 14356 28960 14408
rect 30012 14399 30064 14408
rect 30012 14365 30021 14399
rect 30021 14365 30055 14399
rect 30055 14365 30064 14399
rect 30012 14356 30064 14365
rect 30104 14356 30156 14408
rect 30564 14356 30616 14408
rect 34704 14492 34756 14544
rect 34796 14424 34848 14476
rect 33140 14399 33192 14408
rect 28724 14288 28776 14340
rect 32588 14288 32640 14340
rect 33140 14365 33149 14399
rect 33149 14365 33183 14399
rect 33183 14365 33192 14399
rect 33140 14356 33192 14365
rect 33784 14399 33836 14408
rect 33784 14365 33793 14399
rect 33793 14365 33827 14399
rect 33827 14365 33836 14399
rect 33784 14356 33836 14365
rect 35348 14356 35400 14408
rect 35532 14399 35584 14408
rect 35532 14365 35541 14399
rect 35541 14365 35575 14399
rect 35575 14365 35584 14399
rect 35532 14356 35584 14365
rect 35624 14399 35676 14408
rect 35624 14365 35633 14399
rect 35633 14365 35667 14399
rect 35667 14365 35676 14399
rect 47032 14492 47084 14544
rect 46480 14467 46532 14476
rect 46480 14433 46489 14467
rect 46489 14433 46523 14467
rect 46523 14433 46532 14467
rect 46480 14424 46532 14433
rect 35624 14356 35676 14365
rect 20996 14220 21048 14272
rect 22836 14263 22888 14272
rect 22836 14229 22845 14263
rect 22845 14229 22879 14263
rect 22879 14229 22888 14263
rect 22836 14220 22888 14229
rect 25136 14220 25188 14272
rect 26608 14220 26660 14272
rect 27068 14263 27120 14272
rect 27068 14229 27083 14263
rect 27083 14229 27117 14263
rect 27117 14229 27120 14263
rect 27068 14220 27120 14229
rect 27804 14220 27856 14272
rect 27896 14220 27948 14272
rect 30932 14220 30984 14272
rect 32680 14220 32732 14272
rect 32772 14220 32824 14272
rect 35716 14288 35768 14340
rect 36728 14399 36780 14408
rect 36728 14365 36737 14399
rect 36737 14365 36771 14399
rect 36771 14365 36780 14399
rect 36728 14356 36780 14365
rect 36912 14399 36964 14408
rect 36912 14365 36921 14399
rect 36921 14365 36955 14399
rect 36955 14365 36964 14399
rect 36912 14356 36964 14365
rect 36268 14263 36320 14272
rect 36268 14229 36277 14263
rect 36277 14229 36311 14263
rect 36311 14229 36320 14263
rect 36268 14220 36320 14229
rect 47216 14288 47268 14340
rect 48136 14331 48188 14340
rect 48136 14297 48145 14331
rect 48145 14297 48179 14331
rect 48179 14297 48188 14331
rect 48136 14288 48188 14297
rect 36912 14220 36964 14272
rect 37004 14220 37056 14272
rect 43996 14220 44048 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 20 13948 72 14000
rect 1676 13880 1728 13932
rect 2136 13880 2188 13932
rect 8116 13923 8168 13932
rect 8116 13889 8125 13923
rect 8125 13889 8159 13923
rect 8159 13889 8168 13923
rect 8116 13880 8168 13889
rect 8300 13855 8352 13864
rect 8300 13821 8309 13855
rect 8309 13821 8343 13855
rect 8343 13821 8352 13855
rect 8300 13812 8352 13821
rect 13728 14016 13780 14068
rect 16672 14016 16724 14068
rect 20996 14016 21048 14068
rect 21916 14016 21968 14068
rect 23020 14016 23072 14068
rect 25504 14059 25556 14068
rect 25504 14025 25513 14059
rect 25513 14025 25547 14059
rect 25547 14025 25556 14059
rect 25504 14016 25556 14025
rect 26148 14059 26200 14068
rect 26148 14025 26157 14059
rect 26157 14025 26191 14059
rect 26191 14025 26200 14059
rect 26148 14016 26200 14025
rect 27068 14016 27120 14068
rect 27896 14016 27948 14068
rect 28356 14016 28408 14068
rect 28908 14016 28960 14068
rect 32312 14016 32364 14068
rect 12624 13991 12676 14000
rect 12624 13957 12633 13991
rect 12633 13957 12667 13991
rect 12667 13957 12676 13991
rect 12624 13948 12676 13957
rect 13176 13948 13228 14000
rect 18696 13948 18748 14000
rect 21364 13948 21416 14000
rect 22836 13948 22888 14000
rect 32772 14016 32824 14068
rect 33784 14016 33836 14068
rect 47860 14016 47912 14068
rect 14924 13923 14976 13932
rect 14924 13889 14933 13923
rect 14933 13889 14967 13923
rect 14967 13889 14976 13923
rect 14924 13880 14976 13889
rect 15476 13880 15528 13932
rect 17500 13880 17552 13932
rect 20628 13880 20680 13932
rect 23388 13923 23440 13932
rect 23388 13889 23397 13923
rect 23397 13889 23431 13923
rect 23431 13889 23440 13923
rect 23388 13880 23440 13889
rect 24400 13880 24452 13932
rect 26516 13880 26568 13932
rect 27528 13923 27580 13932
rect 27528 13889 27537 13923
rect 27537 13889 27571 13923
rect 27571 13889 27580 13923
rect 27528 13880 27580 13889
rect 27804 13923 27856 13932
rect 27804 13889 27813 13923
rect 27813 13889 27847 13923
rect 27847 13889 27856 13923
rect 27804 13880 27856 13889
rect 28724 13880 28776 13932
rect 29276 13923 29328 13932
rect 29276 13889 29285 13923
rect 29285 13889 29319 13923
rect 29319 13889 29328 13923
rect 29276 13880 29328 13889
rect 29552 13880 29604 13932
rect 32956 13948 33008 14000
rect 34612 13948 34664 14000
rect 34796 13948 34848 14000
rect 4068 13744 4120 13796
rect 15200 13812 15252 13864
rect 18604 13812 18656 13864
rect 19432 13855 19484 13864
rect 19432 13821 19441 13855
rect 19441 13821 19475 13855
rect 19475 13821 19484 13855
rect 19432 13812 19484 13821
rect 24768 13812 24820 13864
rect 26884 13812 26936 13864
rect 27988 13812 28040 13864
rect 29460 13855 29512 13864
rect 29460 13821 29469 13855
rect 29469 13821 29503 13855
rect 29503 13821 29512 13855
rect 29460 13812 29512 13821
rect 1584 13676 1636 13728
rect 2872 13719 2924 13728
rect 2872 13685 2881 13719
rect 2881 13685 2915 13719
rect 2915 13685 2924 13719
rect 2872 13676 2924 13685
rect 15016 13719 15068 13728
rect 15016 13685 15025 13719
rect 15025 13685 15059 13719
rect 15059 13685 15068 13719
rect 15016 13676 15068 13685
rect 19708 13676 19760 13728
rect 20076 13676 20128 13728
rect 25228 13676 25280 13728
rect 27528 13719 27580 13728
rect 27528 13685 27537 13719
rect 27537 13685 27571 13719
rect 27571 13685 27580 13719
rect 27528 13676 27580 13685
rect 29000 13744 29052 13796
rect 31208 13744 31260 13796
rect 31576 13744 31628 13796
rect 32404 13812 32456 13864
rect 32680 13880 32732 13932
rect 36268 13948 36320 14000
rect 47860 13923 47912 13932
rect 47860 13889 47869 13923
rect 47869 13889 47903 13923
rect 47903 13889 47912 13923
rect 47860 13880 47912 13889
rect 32128 13744 32180 13796
rect 32312 13744 32364 13796
rect 33600 13676 33652 13728
rect 34704 13676 34756 13728
rect 36360 13676 36412 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 8300 13515 8352 13524
rect 8300 13481 8309 13515
rect 8309 13481 8343 13515
rect 8343 13481 8352 13515
rect 8300 13472 8352 13481
rect 15568 13472 15620 13524
rect 2872 13404 2924 13456
rect 1584 13379 1636 13388
rect 1584 13345 1593 13379
rect 1593 13345 1627 13379
rect 1627 13345 1636 13379
rect 1584 13336 1636 13345
rect 2780 13379 2832 13388
rect 2780 13345 2789 13379
rect 2789 13345 2823 13379
rect 2823 13345 2832 13379
rect 2780 13336 2832 13345
rect 14280 13336 14332 13388
rect 7932 13268 7984 13320
rect 8116 13268 8168 13320
rect 15200 13268 15252 13320
rect 23572 13472 23624 13524
rect 26332 13472 26384 13524
rect 27160 13472 27212 13524
rect 27620 13472 27672 13524
rect 29460 13472 29512 13524
rect 29920 13472 29972 13524
rect 27896 13404 27948 13456
rect 18604 13336 18656 13388
rect 23940 13336 23992 13388
rect 27712 13336 27764 13388
rect 30380 13336 30432 13388
rect 15016 13200 15068 13252
rect 17224 13243 17276 13252
rect 17224 13209 17233 13243
rect 17233 13209 17267 13243
rect 17267 13209 17276 13243
rect 17224 13200 17276 13209
rect 18328 13311 18380 13320
rect 18328 13277 18337 13311
rect 18337 13277 18371 13311
rect 18371 13277 18380 13311
rect 18328 13268 18380 13277
rect 18512 13311 18564 13320
rect 18512 13277 18521 13311
rect 18521 13277 18555 13311
rect 18555 13277 18564 13311
rect 19708 13311 19760 13320
rect 18512 13268 18564 13277
rect 19708 13277 19717 13311
rect 19717 13277 19751 13311
rect 19751 13277 19760 13311
rect 19708 13268 19760 13277
rect 20720 13268 20772 13320
rect 23020 13268 23072 13320
rect 25228 13311 25280 13320
rect 25228 13277 25237 13311
rect 25237 13277 25271 13311
rect 25271 13277 25280 13311
rect 25228 13268 25280 13277
rect 26608 13268 26660 13320
rect 26884 13268 26936 13320
rect 29000 13268 29052 13320
rect 29736 13311 29788 13320
rect 29736 13277 29745 13311
rect 29745 13277 29779 13311
rect 29779 13277 29788 13311
rect 29736 13268 29788 13277
rect 25136 13200 25188 13252
rect 17868 13175 17920 13184
rect 17868 13141 17877 13175
rect 17877 13141 17911 13175
rect 17911 13141 17920 13175
rect 17868 13132 17920 13141
rect 20260 13132 20312 13184
rect 23756 13132 23808 13184
rect 25044 13132 25096 13184
rect 29460 13200 29512 13252
rect 29644 13132 29696 13184
rect 30012 13268 30064 13320
rect 30564 13268 30616 13320
rect 33600 13472 33652 13524
rect 36728 13472 36780 13524
rect 30840 13447 30892 13456
rect 30840 13413 30849 13447
rect 30849 13413 30883 13447
rect 30883 13413 30892 13447
rect 30840 13404 30892 13413
rect 35532 13404 35584 13456
rect 32404 13379 32456 13388
rect 32404 13345 32413 13379
rect 32413 13345 32447 13379
rect 32447 13345 32456 13379
rect 32404 13336 32456 13345
rect 30932 13311 30984 13320
rect 30932 13277 30941 13311
rect 30941 13277 30975 13311
rect 30975 13277 30984 13311
rect 30932 13268 30984 13277
rect 31760 13311 31812 13320
rect 31760 13277 31769 13311
rect 31769 13277 31803 13311
rect 31803 13277 31812 13311
rect 31760 13268 31812 13277
rect 32496 13268 32548 13320
rect 35348 13311 35400 13320
rect 35348 13277 35357 13311
rect 35357 13277 35391 13311
rect 35391 13277 35400 13311
rect 35348 13268 35400 13277
rect 35532 13311 35584 13320
rect 35532 13277 35541 13311
rect 35541 13277 35575 13311
rect 35575 13277 35584 13311
rect 35716 13311 35768 13320
rect 35532 13268 35584 13277
rect 35716 13277 35725 13311
rect 35725 13277 35759 13311
rect 35759 13277 35768 13311
rect 35716 13268 35768 13277
rect 36360 13311 36412 13320
rect 36360 13277 36369 13311
rect 36369 13277 36403 13311
rect 36403 13277 36412 13311
rect 36360 13268 36412 13277
rect 34520 13200 34572 13252
rect 30012 13132 30064 13184
rect 30196 13132 30248 13184
rect 32496 13132 32548 13184
rect 35072 13175 35124 13184
rect 35072 13141 35081 13175
rect 35081 13141 35115 13175
rect 35115 13141 35124 13175
rect 35072 13132 35124 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 19340 12928 19392 12980
rect 19984 12971 20036 12980
rect 19984 12937 19993 12971
rect 19993 12937 20027 12971
rect 20027 12937 20036 12971
rect 19984 12928 20036 12937
rect 23572 12928 23624 12980
rect 15292 12860 15344 12912
rect 3976 12792 4028 12844
rect 14096 12835 14148 12844
rect 14096 12801 14105 12835
rect 14105 12801 14139 12835
rect 14139 12801 14148 12835
rect 14096 12792 14148 12801
rect 16672 12835 16724 12844
rect 16672 12801 16681 12835
rect 16681 12801 16715 12835
rect 16715 12801 16724 12835
rect 16672 12792 16724 12801
rect 17868 12860 17920 12912
rect 18696 12860 18748 12912
rect 20996 12860 21048 12912
rect 21364 12860 21416 12912
rect 23756 12860 23808 12912
rect 23572 12792 23624 12844
rect 24492 12835 24544 12844
rect 24492 12801 24501 12835
rect 24501 12801 24535 12835
rect 24535 12801 24544 12835
rect 24492 12792 24544 12801
rect 27252 12928 27304 12980
rect 29092 12928 29144 12980
rect 30012 12928 30064 12980
rect 26792 12860 26844 12912
rect 29736 12860 29788 12912
rect 35072 12860 35124 12912
rect 1400 12767 1452 12776
rect 1400 12733 1409 12767
rect 1409 12733 1443 12767
rect 1443 12733 1452 12767
rect 1400 12724 1452 12733
rect 14280 12767 14332 12776
rect 14280 12733 14289 12767
rect 14289 12733 14323 12767
rect 14323 12733 14332 12767
rect 14280 12724 14332 12733
rect 12440 12656 12492 12708
rect 19156 12724 19208 12776
rect 23756 12767 23808 12776
rect 23756 12733 23765 12767
rect 23765 12733 23799 12767
rect 23799 12733 23808 12767
rect 23756 12724 23808 12733
rect 23940 12767 23992 12776
rect 23940 12733 23949 12767
rect 23949 12733 23983 12767
rect 23983 12733 23992 12767
rect 23940 12724 23992 12733
rect 18052 12631 18104 12640
rect 18052 12597 18061 12631
rect 18061 12597 18095 12631
rect 18095 12597 18104 12631
rect 18052 12588 18104 12597
rect 19248 12588 19300 12640
rect 20076 12588 20128 12640
rect 23480 12588 23532 12640
rect 25136 12792 25188 12844
rect 27712 12792 27764 12844
rect 29276 12792 29328 12844
rect 30380 12792 30432 12844
rect 31300 12792 31352 12844
rect 32404 12835 32456 12844
rect 32404 12801 32413 12835
rect 32413 12801 32447 12835
rect 32447 12801 32456 12835
rect 32404 12792 32456 12801
rect 32772 12792 32824 12844
rect 34796 12792 34848 12844
rect 26332 12724 26384 12776
rect 28356 12724 28408 12776
rect 29460 12767 29512 12776
rect 29460 12733 29469 12767
rect 29469 12733 29503 12767
rect 29503 12733 29512 12767
rect 29460 12724 29512 12733
rect 25136 12656 25188 12708
rect 31760 12724 31812 12776
rect 26792 12588 26844 12640
rect 27252 12588 27304 12640
rect 27988 12588 28040 12640
rect 36360 12631 36412 12640
rect 36360 12597 36369 12631
rect 36369 12597 36403 12631
rect 36403 12597 36412 12631
rect 36360 12588 36412 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 14280 12427 14332 12436
rect 14280 12393 14289 12427
rect 14289 12393 14323 12427
rect 14323 12393 14332 12427
rect 14280 12384 14332 12393
rect 18328 12384 18380 12436
rect 18880 12384 18932 12436
rect 20720 12384 20772 12436
rect 24492 12384 24544 12436
rect 26700 12384 26752 12436
rect 31300 12427 31352 12436
rect 31300 12393 31309 12427
rect 31309 12393 31343 12427
rect 31343 12393 31352 12427
rect 31300 12384 31352 12393
rect 35532 12384 35584 12436
rect 40776 12384 40828 12436
rect 46848 12384 46900 12436
rect 18052 12248 18104 12300
rect 20260 12291 20312 12300
rect 20260 12257 20269 12291
rect 20269 12257 20303 12291
rect 20303 12257 20312 12291
rect 20260 12248 20312 12257
rect 26884 12248 26936 12300
rect 29920 12291 29972 12300
rect 29920 12257 29929 12291
rect 29929 12257 29963 12291
rect 29963 12257 29972 12291
rect 29920 12248 29972 12257
rect 33416 12248 33468 12300
rect 20076 12223 20128 12232
rect 20076 12189 20085 12223
rect 20085 12189 20119 12223
rect 20119 12189 20128 12223
rect 20076 12180 20128 12189
rect 23480 12223 23532 12232
rect 23480 12189 23489 12223
rect 23489 12189 23523 12223
rect 23523 12189 23532 12223
rect 23480 12180 23532 12189
rect 23664 12223 23716 12232
rect 23664 12189 23673 12223
rect 23673 12189 23707 12223
rect 23707 12189 23716 12223
rect 23664 12180 23716 12189
rect 26700 12223 26752 12232
rect 26700 12189 26709 12223
rect 26709 12189 26743 12223
rect 26743 12189 26752 12223
rect 26700 12180 26752 12189
rect 27528 12180 27580 12232
rect 17868 12155 17920 12164
rect 17868 12121 17877 12155
rect 17877 12121 17911 12155
rect 17911 12121 17920 12155
rect 17868 12112 17920 12121
rect 19156 12112 19208 12164
rect 19524 12112 19576 12164
rect 20260 12112 20312 12164
rect 21916 12155 21968 12164
rect 21916 12121 21925 12155
rect 21925 12121 21959 12155
rect 21959 12121 21968 12155
rect 21916 12112 21968 12121
rect 26884 12112 26936 12164
rect 27712 12112 27764 12164
rect 29368 12180 29420 12232
rect 30012 12180 30064 12232
rect 30196 12223 30248 12232
rect 30196 12189 30230 12223
rect 30230 12189 30248 12223
rect 30196 12180 30248 12189
rect 34520 12180 34572 12232
rect 36360 12180 36412 12232
rect 18236 12044 18288 12096
rect 19984 12044 20036 12096
rect 28264 12044 28316 12096
rect 28540 12044 28592 12096
rect 29644 12044 29696 12096
rect 32588 12044 32640 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 20076 11840 20128 11892
rect 17224 11704 17276 11756
rect 19248 11704 19300 11756
rect 19892 11704 19944 11756
rect 20536 11840 20588 11892
rect 21916 11840 21968 11892
rect 46756 11840 46808 11892
rect 23480 11772 23532 11824
rect 24768 11772 24820 11824
rect 20536 11747 20588 11756
rect 20536 11713 20545 11747
rect 20545 11713 20579 11747
rect 20579 11713 20588 11747
rect 20536 11704 20588 11713
rect 20996 11704 21048 11756
rect 25964 11747 26016 11756
rect 16672 11636 16724 11688
rect 17040 11636 17092 11688
rect 20628 11636 20680 11688
rect 20720 11636 20772 11688
rect 22192 11636 22244 11688
rect 25964 11713 25973 11747
rect 25973 11713 26007 11747
rect 26007 11713 26016 11747
rect 25964 11704 26016 11713
rect 28908 11772 28960 11824
rect 27528 11704 27580 11756
rect 28448 11747 28500 11756
rect 28448 11713 28457 11747
rect 28457 11713 28491 11747
rect 28491 11713 28500 11747
rect 28448 11704 28500 11713
rect 28632 11747 28684 11756
rect 28632 11713 28641 11747
rect 28641 11713 28675 11747
rect 28675 11713 28684 11747
rect 28632 11704 28684 11713
rect 29828 11704 29880 11756
rect 26424 11636 26476 11688
rect 28264 11636 28316 11688
rect 29644 11679 29696 11688
rect 29644 11645 29653 11679
rect 29653 11645 29687 11679
rect 29687 11645 29696 11679
rect 29644 11636 29696 11645
rect 26884 11568 26936 11620
rect 29000 11568 29052 11620
rect 18420 11500 18472 11552
rect 20904 11500 20956 11552
rect 25504 11500 25556 11552
rect 27160 11543 27212 11552
rect 27160 11509 27169 11543
rect 27169 11509 27203 11543
rect 27203 11509 27212 11543
rect 27160 11500 27212 11509
rect 27620 11500 27672 11552
rect 27896 11543 27948 11552
rect 27896 11509 27905 11543
rect 27905 11509 27939 11543
rect 27939 11509 27948 11543
rect 27896 11500 27948 11509
rect 30012 11500 30064 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 17960 11296 18012 11348
rect 18880 11296 18932 11348
rect 19248 11339 19300 11348
rect 19248 11305 19257 11339
rect 19257 11305 19291 11339
rect 19291 11305 19300 11339
rect 19248 11296 19300 11305
rect 18604 11228 18656 11280
rect 1768 11092 1820 11144
rect 17132 11092 17184 11144
rect 18236 11092 18288 11144
rect 25136 11296 25188 11348
rect 25964 11296 26016 11348
rect 28448 11296 28500 11348
rect 29920 11296 29972 11348
rect 19984 11160 20036 11212
rect 20076 11160 20128 11212
rect 20444 11160 20496 11212
rect 1860 11067 1912 11076
rect 1860 11033 1869 11067
rect 1869 11033 1903 11067
rect 1903 11033 1912 11067
rect 1860 11024 1912 11033
rect 1952 11024 2004 11076
rect 19432 11024 19484 11076
rect 18512 10956 18564 11008
rect 18880 10956 18932 11008
rect 20168 11092 20220 11144
rect 20904 11135 20956 11144
rect 20904 11101 20913 11135
rect 20913 11101 20947 11135
rect 20947 11101 20956 11135
rect 20904 11092 20956 11101
rect 23848 11228 23900 11280
rect 24216 11228 24268 11280
rect 28264 11271 28316 11280
rect 22192 11092 22244 11144
rect 21456 11024 21508 11076
rect 22376 11024 22428 11076
rect 23480 11135 23532 11144
rect 23480 11101 23489 11135
rect 23489 11101 23523 11135
rect 23523 11101 23532 11135
rect 23480 11092 23532 11101
rect 23848 11092 23900 11144
rect 24400 11135 24452 11144
rect 24400 11101 24409 11135
rect 24409 11101 24443 11135
rect 24443 11101 24452 11135
rect 24400 11092 24452 11101
rect 28264 11237 28273 11271
rect 28273 11237 28307 11271
rect 28307 11237 28316 11271
rect 28264 11228 28316 11237
rect 27528 11160 27580 11212
rect 32588 11228 32640 11280
rect 33140 11228 33192 11280
rect 25228 11135 25280 11144
rect 25228 11101 25237 11135
rect 25237 11101 25271 11135
rect 25271 11101 25280 11135
rect 25228 11092 25280 11101
rect 25504 11135 25556 11144
rect 25504 11101 25538 11135
rect 25538 11101 25556 11135
rect 25504 11092 25556 11101
rect 27988 11092 28040 11144
rect 28264 11092 28316 11144
rect 28724 11092 28776 11144
rect 30012 11135 30064 11144
rect 30012 11101 30021 11135
rect 30021 11101 30055 11135
rect 30055 11101 30064 11135
rect 30012 11092 30064 11101
rect 33048 11160 33100 11212
rect 20444 10999 20496 11008
rect 20444 10965 20453 10999
rect 20453 10965 20487 10999
rect 20487 10965 20496 10999
rect 20444 10956 20496 10965
rect 22284 10956 22336 11008
rect 24032 11024 24084 11076
rect 26976 11024 27028 11076
rect 27528 11067 27580 11076
rect 27528 11033 27537 11067
rect 27537 11033 27571 11067
rect 27571 11033 27580 11067
rect 27528 11024 27580 11033
rect 27896 11024 27948 11076
rect 28540 11024 28592 11076
rect 29920 11024 29972 11076
rect 23664 10956 23716 11008
rect 23848 10999 23900 11008
rect 23848 10965 23857 10999
rect 23857 10965 23891 10999
rect 23891 10965 23900 10999
rect 23848 10956 23900 10965
rect 26332 10956 26384 11008
rect 27252 10956 27304 11008
rect 27712 10999 27764 11008
rect 27712 10965 27721 10999
rect 27721 10965 27755 10999
rect 27755 10965 27764 10999
rect 27712 10956 27764 10965
rect 28724 10999 28776 11008
rect 28724 10965 28733 10999
rect 28733 10965 28767 10999
rect 28767 10965 28776 10999
rect 28724 10956 28776 10965
rect 30012 10956 30064 11008
rect 32404 11092 32456 11144
rect 32956 11092 33008 11144
rect 33140 11092 33192 11144
rect 47216 11135 47268 11144
rect 47216 11101 47225 11135
rect 47225 11101 47259 11135
rect 47259 11101 47268 11135
rect 47216 11092 47268 11101
rect 48044 11135 48096 11144
rect 48044 11101 48053 11135
rect 48053 11101 48087 11135
rect 48087 11101 48096 11135
rect 48044 11092 48096 11101
rect 33416 11024 33468 11076
rect 32588 10956 32640 11008
rect 33784 10956 33836 11008
rect 47308 10999 47360 11008
rect 47308 10965 47317 10999
rect 47317 10965 47351 10999
rect 47351 10965 47360 10999
rect 47308 10956 47360 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 20628 10752 20680 10804
rect 2136 10659 2188 10668
rect 2136 10625 2145 10659
rect 2145 10625 2179 10659
rect 2179 10625 2188 10659
rect 2136 10616 2188 10625
rect 20444 10684 20496 10736
rect 18788 10659 18840 10668
rect 18788 10625 18797 10659
rect 18797 10625 18831 10659
rect 18831 10625 18840 10659
rect 18788 10616 18840 10625
rect 19064 10616 19116 10668
rect 19340 10616 19392 10668
rect 23480 10684 23532 10736
rect 25228 10684 25280 10736
rect 18604 10480 18656 10532
rect 20628 10480 20680 10532
rect 22008 10480 22060 10532
rect 22284 10659 22336 10668
rect 22284 10625 22293 10659
rect 22293 10625 22327 10659
rect 22327 10625 22336 10659
rect 22284 10616 22336 10625
rect 22468 10659 22520 10668
rect 22468 10625 22477 10659
rect 22477 10625 22511 10659
rect 22511 10625 22520 10659
rect 23020 10659 23072 10668
rect 22468 10616 22520 10625
rect 22284 10480 22336 10532
rect 1400 10412 1452 10464
rect 2228 10455 2280 10464
rect 2228 10421 2237 10455
rect 2237 10421 2271 10455
rect 2271 10421 2280 10455
rect 2228 10412 2280 10421
rect 2964 10455 3016 10464
rect 2964 10421 2973 10455
rect 2973 10421 3007 10455
rect 3007 10421 3016 10455
rect 2964 10412 3016 10421
rect 18328 10455 18380 10464
rect 18328 10421 18337 10455
rect 18337 10421 18371 10455
rect 18371 10421 18380 10455
rect 18328 10412 18380 10421
rect 18420 10412 18472 10464
rect 19064 10412 19116 10464
rect 21824 10455 21876 10464
rect 21824 10421 21833 10455
rect 21833 10421 21867 10455
rect 21867 10421 21876 10455
rect 21824 10412 21876 10421
rect 23020 10625 23029 10659
rect 23029 10625 23063 10659
rect 23063 10625 23072 10659
rect 23020 10616 23072 10625
rect 23848 10616 23900 10668
rect 24860 10659 24912 10668
rect 24860 10625 24869 10659
rect 24869 10625 24903 10659
rect 24903 10625 24912 10659
rect 24860 10616 24912 10625
rect 25504 10616 25556 10668
rect 24952 10548 25004 10600
rect 23388 10412 23440 10464
rect 23664 10412 23716 10464
rect 24492 10412 24544 10464
rect 26240 10752 26292 10804
rect 26424 10795 26476 10804
rect 26424 10761 26433 10795
rect 26433 10761 26467 10795
rect 26467 10761 26476 10795
rect 26424 10752 26476 10761
rect 27160 10752 27212 10804
rect 28632 10752 28684 10804
rect 32404 10752 32456 10804
rect 32496 10752 32548 10804
rect 32588 10752 32640 10804
rect 25872 10659 25924 10668
rect 25872 10625 25881 10659
rect 25881 10625 25915 10659
rect 25915 10625 25924 10659
rect 26700 10684 26752 10736
rect 25872 10616 25924 10625
rect 26240 10659 26292 10668
rect 26240 10625 26249 10659
rect 26249 10625 26283 10659
rect 26283 10625 26292 10659
rect 26240 10616 26292 10625
rect 26976 10659 27028 10668
rect 26976 10625 26985 10659
rect 26985 10625 27019 10659
rect 27019 10625 27028 10659
rect 26976 10616 27028 10625
rect 27988 10616 28040 10668
rect 32772 10659 32824 10668
rect 32772 10625 32781 10659
rect 32781 10625 32815 10659
rect 32815 10625 32824 10659
rect 32772 10616 32824 10625
rect 26792 10548 26844 10600
rect 47952 10684 48004 10736
rect 33416 10616 33468 10668
rect 40684 10616 40736 10668
rect 47768 10659 47820 10668
rect 47768 10625 47777 10659
rect 47777 10625 47811 10659
rect 47811 10625 47820 10659
rect 47768 10616 47820 10625
rect 33784 10591 33836 10600
rect 33784 10557 33793 10591
rect 33793 10557 33827 10591
rect 33827 10557 33836 10591
rect 33784 10548 33836 10557
rect 30012 10480 30064 10532
rect 27804 10455 27856 10464
rect 27804 10421 27813 10455
rect 27813 10421 27847 10455
rect 27847 10421 27856 10455
rect 27804 10412 27856 10421
rect 27896 10412 27948 10464
rect 32496 10412 32548 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 18788 10208 18840 10260
rect 22376 10251 22428 10260
rect 22376 10217 22385 10251
rect 22385 10217 22419 10251
rect 22419 10217 22428 10251
rect 22376 10208 22428 10217
rect 25228 10208 25280 10260
rect 27712 10208 27764 10260
rect 25412 10140 25464 10192
rect 25596 10140 25648 10192
rect 27436 10140 27488 10192
rect 1400 10115 1452 10124
rect 1400 10081 1409 10115
rect 1409 10081 1443 10115
rect 1443 10081 1452 10115
rect 1400 10072 1452 10081
rect 2228 10072 2280 10124
rect 2780 10115 2832 10124
rect 2780 10081 2789 10115
rect 2789 10081 2823 10115
rect 2823 10081 2832 10115
rect 2780 10072 2832 10081
rect 17040 10115 17092 10124
rect 17040 10081 17049 10115
rect 17049 10081 17083 10115
rect 17083 10081 17092 10115
rect 17040 10072 17092 10081
rect 19340 10072 19392 10124
rect 23664 10072 23716 10124
rect 24124 10072 24176 10124
rect 24952 10072 25004 10124
rect 18328 10004 18380 10056
rect 20444 10004 20496 10056
rect 21824 10004 21876 10056
rect 22008 10004 22060 10056
rect 26240 10072 26292 10124
rect 28724 10208 28776 10260
rect 33416 10208 33468 10260
rect 28908 10072 28960 10124
rect 29460 10072 29512 10124
rect 48044 10140 48096 10192
rect 47308 10072 47360 10124
rect 48136 10115 48188 10124
rect 48136 10081 48145 10115
rect 48145 10081 48179 10115
rect 48179 10081 48188 10115
rect 48136 10072 48188 10081
rect 27160 10004 27212 10056
rect 27804 10004 27856 10056
rect 28080 10004 28132 10056
rect 29920 10047 29972 10056
rect 19248 9979 19300 9988
rect 19248 9945 19257 9979
rect 19257 9945 19291 9979
rect 19291 9945 19300 9979
rect 19248 9936 19300 9945
rect 18420 9911 18472 9920
rect 18420 9877 18429 9911
rect 18429 9877 18463 9911
rect 18463 9877 18472 9911
rect 22284 9936 22336 9988
rect 23848 9936 23900 9988
rect 24032 9936 24084 9988
rect 24584 9936 24636 9988
rect 26792 9979 26844 9988
rect 18420 9868 18472 9877
rect 23296 9868 23348 9920
rect 24768 9868 24820 9920
rect 25136 9911 25188 9920
rect 25136 9877 25145 9911
rect 25145 9877 25179 9911
rect 25179 9877 25188 9911
rect 25136 9868 25188 9877
rect 26792 9945 26801 9979
rect 26801 9945 26835 9979
rect 26835 9945 26844 9979
rect 26792 9936 26844 9945
rect 26976 9979 27028 9988
rect 26976 9945 26985 9979
rect 26985 9945 27019 9979
rect 27019 9945 27028 9979
rect 27620 9979 27672 9988
rect 26976 9936 27028 9945
rect 27620 9945 27629 9979
rect 27629 9945 27663 9979
rect 27663 9945 27672 9979
rect 27620 9936 27672 9945
rect 27712 9936 27764 9988
rect 29920 10013 29929 10047
rect 29929 10013 29963 10047
rect 29963 10013 29972 10047
rect 29920 10004 29972 10013
rect 30012 10004 30064 10056
rect 32496 10004 32548 10056
rect 27896 9868 27948 9920
rect 29828 9868 29880 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 24860 9707 24912 9716
rect 24860 9673 24869 9707
rect 24869 9673 24903 9707
rect 24903 9673 24912 9707
rect 24860 9664 24912 9673
rect 29920 9664 29972 9716
rect 2964 9596 3016 9648
rect 3424 9596 3476 9648
rect 12440 9596 12492 9648
rect 18420 9596 18472 9648
rect 23756 9596 23808 9648
rect 23204 9571 23256 9580
rect 23204 9537 23213 9571
rect 23213 9537 23247 9571
rect 23247 9537 23256 9571
rect 23204 9528 23256 9537
rect 1952 9503 2004 9512
rect 1952 9469 1961 9503
rect 1961 9469 1995 9503
rect 1995 9469 2004 9503
rect 1952 9460 2004 9469
rect 2780 9503 2832 9512
rect 2780 9469 2789 9503
rect 2789 9469 2823 9503
rect 2823 9469 2832 9503
rect 2780 9460 2832 9469
rect 17776 9503 17828 9512
rect 17776 9469 17785 9503
rect 17785 9469 17819 9503
rect 17819 9469 17828 9503
rect 17776 9460 17828 9469
rect 18236 9503 18288 9512
rect 18236 9469 18245 9503
rect 18245 9469 18279 9503
rect 18279 9469 18288 9503
rect 23296 9503 23348 9512
rect 18236 9460 18288 9469
rect 23296 9469 23305 9503
rect 23305 9469 23339 9503
rect 23339 9469 23348 9503
rect 23296 9460 23348 9469
rect 24400 9596 24452 9648
rect 24768 9596 24820 9648
rect 25412 9596 25464 9648
rect 32128 9664 32180 9716
rect 24492 9571 24544 9580
rect 24492 9537 24501 9571
rect 24501 9537 24535 9571
rect 24535 9537 24544 9571
rect 24492 9528 24544 9537
rect 24584 9528 24636 9580
rect 24860 9528 24912 9580
rect 27160 9528 27212 9580
rect 27988 9571 28040 9580
rect 27988 9537 27997 9571
rect 27997 9537 28031 9571
rect 28031 9537 28040 9571
rect 27988 9528 28040 9537
rect 28540 9528 28592 9580
rect 36544 9596 36596 9648
rect 24400 9460 24452 9512
rect 25136 9460 25188 9512
rect 25412 9503 25464 9512
rect 25412 9469 25421 9503
rect 25421 9469 25455 9503
rect 25455 9469 25464 9503
rect 25412 9460 25464 9469
rect 664 9324 716 9376
rect 29000 9392 29052 9444
rect 29460 9460 29512 9512
rect 29920 9571 29972 9580
rect 29920 9537 29929 9571
rect 29929 9537 29963 9571
rect 29963 9537 29972 9571
rect 29920 9528 29972 9537
rect 30104 9571 30156 9580
rect 30104 9537 30113 9571
rect 30113 9537 30147 9571
rect 30147 9537 30156 9571
rect 30288 9571 30340 9580
rect 30104 9528 30156 9537
rect 30288 9537 30297 9571
rect 30297 9537 30331 9571
rect 30331 9537 30340 9571
rect 30288 9528 30340 9537
rect 31392 9571 31444 9580
rect 30196 9503 30248 9512
rect 30196 9469 30205 9503
rect 30205 9469 30239 9503
rect 30239 9469 30248 9503
rect 30196 9460 30248 9469
rect 31392 9537 31401 9571
rect 31401 9537 31435 9571
rect 31435 9537 31444 9571
rect 31392 9528 31444 9537
rect 32404 9460 32456 9512
rect 32864 9460 32916 9512
rect 33140 9503 33192 9512
rect 33140 9469 33149 9503
rect 33149 9469 33183 9503
rect 33183 9469 33192 9503
rect 33140 9460 33192 9469
rect 30840 9392 30892 9444
rect 32680 9392 32732 9444
rect 16580 9324 16632 9376
rect 18236 9324 18288 9376
rect 24400 9367 24452 9376
rect 24400 9333 24409 9367
rect 24409 9333 24443 9367
rect 24443 9333 24452 9367
rect 24400 9324 24452 9333
rect 24492 9324 24544 9376
rect 26792 9324 26844 9376
rect 26976 9324 27028 9376
rect 28540 9324 28592 9376
rect 30656 9367 30708 9376
rect 30656 9333 30665 9367
rect 30665 9333 30699 9367
rect 30699 9333 30708 9367
rect 30656 9324 30708 9333
rect 31392 9324 31444 9376
rect 33232 9324 33284 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 17776 9120 17828 9172
rect 23204 9120 23256 9172
rect 24400 9120 24452 9172
rect 27896 9163 27948 9172
rect 24768 9052 24820 9104
rect 23572 8984 23624 9036
rect 24492 8984 24544 9036
rect 27896 9129 27905 9163
rect 27905 9129 27939 9163
rect 27939 9129 27948 9163
rect 27896 9120 27948 9129
rect 28080 9163 28132 9172
rect 28080 9129 28089 9163
rect 28089 9129 28123 9163
rect 28123 9129 28132 9163
rect 28080 9120 28132 9129
rect 30196 9120 30248 9172
rect 32220 9120 32272 9172
rect 32680 9120 32732 9172
rect 39304 9120 39356 9172
rect 46848 9120 46900 9172
rect 29920 9052 29972 9104
rect 31484 9052 31536 9104
rect 17960 8959 18012 8968
rect 17960 8925 17969 8959
rect 17969 8925 18003 8959
rect 18003 8925 18012 8959
rect 17960 8916 18012 8925
rect 23296 8916 23348 8968
rect 23572 8848 23624 8900
rect 23756 8848 23808 8900
rect 25412 8916 25464 8968
rect 26976 8959 27028 8968
rect 26976 8925 26985 8959
rect 26985 8925 27019 8959
rect 27019 8925 27028 8959
rect 26976 8916 27028 8925
rect 25872 8780 25924 8832
rect 27712 8916 27764 8968
rect 28540 8959 28592 8968
rect 28540 8925 28549 8959
rect 28549 8925 28583 8959
rect 28583 8925 28592 8959
rect 28540 8916 28592 8925
rect 29552 8916 29604 8968
rect 30012 8959 30064 8968
rect 30012 8925 30021 8959
rect 30021 8925 30055 8959
rect 30055 8925 30064 8959
rect 30012 8916 30064 8925
rect 30656 8916 30708 8968
rect 32128 8916 32180 8968
rect 32588 8959 32640 8968
rect 32588 8925 32597 8959
rect 32597 8925 32631 8959
rect 32631 8925 32640 8959
rect 32588 8916 32640 8925
rect 33140 8984 33192 9036
rect 33232 8984 33284 9036
rect 33416 8959 33468 8968
rect 33416 8925 33425 8959
rect 33425 8925 33459 8959
rect 33459 8925 33468 8959
rect 33416 8916 33468 8925
rect 27804 8848 27856 8900
rect 27988 8848 28040 8900
rect 28632 8848 28684 8900
rect 29460 8848 29512 8900
rect 30104 8848 30156 8900
rect 31944 8848 31996 8900
rect 28908 8823 28960 8832
rect 28908 8789 28917 8823
rect 28917 8789 28951 8823
rect 28951 8789 28960 8823
rect 28908 8780 28960 8789
rect 32220 8823 32272 8832
rect 32220 8789 32229 8823
rect 32229 8789 32263 8823
rect 32263 8789 32272 8823
rect 32220 8780 32272 8789
rect 32772 8848 32824 8900
rect 47952 8891 48004 8900
rect 47952 8857 47961 8891
rect 47961 8857 47995 8891
rect 47995 8857 48004 8891
rect 47952 8848 48004 8857
rect 46480 8780 46532 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 18420 8508 18472 8560
rect 23756 8576 23808 8628
rect 24768 8576 24820 8628
rect 27436 8576 27488 8628
rect 24216 8508 24268 8560
rect 27160 8508 27212 8560
rect 28264 8508 28316 8560
rect 28632 8576 28684 8628
rect 30196 8508 30248 8560
rect 32220 8508 32272 8560
rect 1860 8483 1912 8492
rect 1860 8449 1869 8483
rect 1869 8449 1903 8483
rect 1903 8449 1912 8483
rect 1860 8440 1912 8449
rect 18328 8372 18380 8424
rect 18788 8440 18840 8492
rect 18880 8483 18932 8492
rect 18880 8449 18889 8483
rect 18889 8449 18923 8483
rect 18923 8449 18932 8483
rect 19340 8483 19392 8492
rect 18880 8440 18932 8449
rect 19340 8449 19349 8483
rect 19349 8449 19383 8483
rect 19383 8449 19392 8483
rect 19340 8440 19392 8449
rect 23664 8483 23716 8492
rect 23664 8449 23673 8483
rect 23673 8449 23707 8483
rect 23707 8449 23716 8483
rect 23664 8440 23716 8449
rect 17684 8304 17736 8356
rect 18788 8304 18840 8356
rect 20720 8347 20772 8356
rect 20720 8313 20729 8347
rect 20729 8313 20763 8347
rect 20763 8313 20772 8347
rect 20720 8304 20772 8313
rect 24400 8440 24452 8492
rect 27896 8440 27948 8492
rect 26056 8372 26108 8424
rect 27620 8372 27672 8424
rect 29552 8440 29604 8492
rect 47860 8483 47912 8492
rect 47860 8449 47869 8483
rect 47869 8449 47903 8483
rect 47903 8449 47912 8483
rect 47860 8440 47912 8449
rect 28080 8304 28132 8356
rect 29644 8372 29696 8424
rect 29828 8304 29880 8356
rect 35808 8304 35860 8356
rect 19616 8236 19668 8288
rect 24400 8236 24452 8288
rect 27620 8279 27672 8288
rect 27620 8245 27629 8279
rect 27629 8245 27663 8279
rect 27663 8245 27672 8279
rect 27620 8236 27672 8245
rect 27804 8236 27856 8288
rect 28908 8236 28960 8288
rect 33784 8279 33836 8288
rect 33784 8245 33793 8279
rect 33793 8245 33827 8279
rect 33827 8245 33836 8279
rect 33784 8236 33836 8245
rect 47032 8279 47084 8288
rect 47032 8245 47041 8279
rect 47041 8245 47075 8279
rect 47075 8245 47084 8279
rect 47032 8236 47084 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 18972 8032 19024 8084
rect 19616 8075 19668 8084
rect 19616 8041 19625 8075
rect 19625 8041 19659 8075
rect 19659 8041 19668 8075
rect 19616 8032 19668 8041
rect 20720 8032 20772 8084
rect 1860 7803 1912 7812
rect 1860 7769 1869 7803
rect 1869 7769 1903 7803
rect 1903 7769 1912 7803
rect 1860 7760 1912 7769
rect 18052 7828 18104 7880
rect 17684 7692 17736 7744
rect 18420 7831 18442 7858
rect 18442 7831 18472 7858
rect 18420 7806 18472 7831
rect 20352 7896 20404 7948
rect 24584 7964 24636 8016
rect 24124 7896 24176 7948
rect 27528 8032 27580 8084
rect 33140 8032 33192 8084
rect 19248 7871 19300 7880
rect 19248 7837 19257 7871
rect 19257 7837 19291 7871
rect 19291 7837 19300 7871
rect 19248 7828 19300 7837
rect 20720 7828 20772 7880
rect 24400 7871 24452 7880
rect 24400 7837 24409 7871
rect 24409 7837 24443 7871
rect 24443 7837 24452 7871
rect 24400 7828 24452 7837
rect 24492 7828 24544 7880
rect 18788 7760 18840 7812
rect 19064 7760 19116 7812
rect 20996 7803 21048 7812
rect 20996 7769 21005 7803
rect 21005 7769 21039 7803
rect 21039 7769 21048 7803
rect 20996 7760 21048 7769
rect 22836 7760 22888 7812
rect 20260 7692 20312 7744
rect 21088 7692 21140 7744
rect 21640 7692 21692 7744
rect 23664 7692 23716 7744
rect 25136 7735 25188 7744
rect 25136 7701 25145 7735
rect 25145 7701 25179 7735
rect 25179 7701 25188 7735
rect 25136 7692 25188 7701
rect 28080 7896 28132 7948
rect 29552 7896 29604 7948
rect 47032 7896 47084 7948
rect 27988 7871 28040 7880
rect 27988 7837 27997 7871
rect 27997 7837 28031 7871
rect 28031 7837 28040 7871
rect 27988 7828 28040 7837
rect 33232 7871 33284 7880
rect 33232 7837 33241 7871
rect 33241 7837 33275 7871
rect 33275 7837 33284 7871
rect 33232 7828 33284 7837
rect 33784 7828 33836 7880
rect 25320 7760 25372 7812
rect 27528 7803 27580 7812
rect 27528 7769 27537 7803
rect 27537 7769 27571 7803
rect 27571 7769 27580 7803
rect 27528 7760 27580 7769
rect 30932 7760 30984 7812
rect 32220 7760 32272 7812
rect 32956 7760 33008 7812
rect 46480 7803 46532 7812
rect 46480 7769 46489 7803
rect 46489 7769 46523 7803
rect 46523 7769 46532 7803
rect 46480 7760 46532 7769
rect 48136 7803 48188 7812
rect 48136 7769 48145 7803
rect 48145 7769 48179 7803
rect 48179 7769 48188 7803
rect 48136 7760 48188 7769
rect 26148 7692 26200 7744
rect 27804 7692 27856 7744
rect 29368 7692 29420 7744
rect 32588 7735 32640 7744
rect 32588 7701 32597 7735
rect 32597 7701 32631 7735
rect 32631 7701 32640 7735
rect 32588 7692 32640 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 18052 7488 18104 7540
rect 18236 7488 18288 7540
rect 19432 7488 19484 7540
rect 20996 7531 21048 7540
rect 19340 7420 19392 7472
rect 20260 7463 20312 7472
rect 20260 7429 20269 7463
rect 20269 7429 20303 7463
rect 20303 7429 20312 7463
rect 20260 7420 20312 7429
rect 20996 7497 21005 7531
rect 21005 7497 21039 7531
rect 21039 7497 21048 7531
rect 20996 7488 21048 7497
rect 24584 7488 24636 7540
rect 25136 7420 25188 7472
rect 17684 7352 17736 7404
rect 20904 7395 20956 7404
rect 20904 7361 20913 7395
rect 20913 7361 20947 7395
rect 20947 7361 20956 7395
rect 20904 7352 20956 7361
rect 23480 7395 23532 7404
rect 23480 7361 23489 7395
rect 23489 7361 23523 7395
rect 23523 7361 23532 7395
rect 23480 7352 23532 7361
rect 28264 7488 28316 7540
rect 30932 7531 30984 7540
rect 30932 7497 30941 7531
rect 30941 7497 30975 7531
rect 30975 7497 30984 7531
rect 30932 7488 30984 7497
rect 31576 7488 31628 7540
rect 32772 7488 32824 7540
rect 26056 7395 26108 7404
rect 22192 7284 22244 7336
rect 26056 7361 26065 7395
rect 26065 7361 26099 7395
rect 26099 7361 26108 7395
rect 26056 7352 26108 7361
rect 26240 7352 26292 7404
rect 28540 7395 28592 7404
rect 28540 7361 28549 7395
rect 28549 7361 28583 7395
rect 28583 7361 28592 7395
rect 28540 7352 28592 7361
rect 29368 7395 29420 7404
rect 26148 7327 26200 7336
rect 18788 7216 18840 7268
rect 26148 7293 26157 7327
rect 26157 7293 26191 7327
rect 26191 7293 26200 7327
rect 26148 7284 26200 7293
rect 27436 7327 27488 7336
rect 2044 7191 2096 7200
rect 2044 7157 2053 7191
rect 2053 7157 2087 7191
rect 2087 7157 2096 7191
rect 2044 7148 2096 7157
rect 21088 7148 21140 7200
rect 24124 7148 24176 7200
rect 27068 7216 27120 7268
rect 27436 7293 27445 7327
rect 27445 7293 27479 7327
rect 27479 7293 27488 7327
rect 27436 7284 27488 7293
rect 29368 7361 29377 7395
rect 29377 7361 29411 7395
rect 29411 7361 29420 7395
rect 29368 7352 29420 7361
rect 29460 7352 29512 7404
rect 32496 7420 32548 7472
rect 29644 7327 29696 7336
rect 29644 7293 29653 7327
rect 29653 7293 29687 7327
rect 29687 7293 29696 7327
rect 29644 7284 29696 7293
rect 27804 7216 27856 7268
rect 26148 7148 26200 7200
rect 27620 7148 27672 7200
rect 28540 7148 28592 7200
rect 31576 7395 31628 7404
rect 31576 7361 31585 7395
rect 31585 7361 31619 7395
rect 31619 7361 31628 7395
rect 31576 7352 31628 7361
rect 32956 7488 33008 7540
rect 33416 7420 33468 7472
rect 32496 7284 32548 7336
rect 33232 7284 33284 7336
rect 29920 7216 29972 7268
rect 30104 7191 30156 7200
rect 30104 7157 30113 7191
rect 30113 7157 30147 7191
rect 30147 7157 30156 7191
rect 30104 7148 30156 7157
rect 31852 7148 31904 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 20904 6944 20956 6996
rect 29276 6944 29328 6996
rect 24492 6876 24544 6928
rect 29368 6876 29420 6928
rect 2044 6808 2096 6860
rect 2228 6808 2280 6860
rect 2412 6808 2464 6860
rect 2780 6851 2832 6860
rect 2780 6817 2789 6851
rect 2789 6817 2823 6851
rect 2823 6817 2832 6851
rect 2780 6808 2832 6817
rect 19340 6808 19392 6860
rect 20260 6851 20312 6860
rect 20260 6817 20269 6851
rect 20269 6817 20303 6851
rect 20303 6817 20312 6851
rect 20260 6808 20312 6817
rect 26332 6808 26384 6860
rect 17960 6740 18012 6792
rect 26240 6783 26292 6792
rect 2228 6672 2280 6724
rect 20628 6672 20680 6724
rect 18328 6604 18380 6656
rect 20352 6604 20404 6656
rect 26240 6749 26249 6783
rect 26249 6749 26283 6783
rect 26283 6749 26292 6783
rect 26240 6740 26292 6749
rect 27068 6783 27120 6792
rect 27068 6749 27077 6783
rect 27077 6749 27111 6783
rect 27111 6749 27120 6783
rect 27068 6740 27120 6749
rect 27160 6783 27212 6792
rect 27160 6749 27169 6783
rect 27169 6749 27203 6783
rect 27203 6749 27212 6783
rect 27160 6740 27212 6749
rect 22192 6672 22244 6724
rect 24768 6672 24820 6724
rect 28724 6808 28776 6860
rect 31852 6851 31904 6860
rect 31852 6817 31861 6851
rect 31861 6817 31895 6851
rect 31895 6817 31904 6851
rect 31852 6808 31904 6817
rect 32128 6851 32180 6860
rect 32128 6817 32137 6851
rect 32137 6817 32171 6851
rect 32171 6817 32180 6851
rect 32128 6808 32180 6817
rect 27436 6783 27488 6792
rect 27436 6749 27445 6783
rect 27445 6749 27479 6783
rect 27479 6749 27488 6783
rect 27436 6740 27488 6749
rect 28908 6740 28960 6792
rect 29552 6783 29604 6792
rect 29552 6749 29561 6783
rect 29561 6749 29595 6783
rect 29595 6749 29604 6783
rect 29552 6740 29604 6749
rect 30104 6740 30156 6792
rect 23204 6604 23256 6656
rect 28540 6672 28592 6724
rect 32588 6672 32640 6724
rect 27712 6604 27764 6656
rect 29644 6604 29696 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 2228 6443 2280 6452
rect 2228 6409 2237 6443
rect 2237 6409 2271 6443
rect 2271 6409 2280 6443
rect 2228 6400 2280 6409
rect 18328 6375 18380 6384
rect 18328 6341 18337 6375
rect 18337 6341 18371 6375
rect 18371 6341 18380 6375
rect 18328 6332 18380 6341
rect 2136 6307 2188 6316
rect 2136 6273 2145 6307
rect 2145 6273 2179 6307
rect 2179 6273 2188 6307
rect 2136 6264 2188 6273
rect 18144 6307 18196 6316
rect 18144 6273 18153 6307
rect 18153 6273 18187 6307
rect 18187 6273 18196 6307
rect 18144 6264 18196 6273
rect 28908 6400 28960 6452
rect 22284 6332 22336 6384
rect 22468 6332 22520 6384
rect 19432 6128 19484 6180
rect 15200 6060 15252 6112
rect 21272 6264 21324 6316
rect 21824 6307 21876 6316
rect 21824 6273 21833 6307
rect 21833 6273 21867 6307
rect 21867 6273 21876 6307
rect 21824 6264 21876 6273
rect 21916 6264 21968 6316
rect 22192 6196 22244 6248
rect 23204 6307 23256 6316
rect 23204 6273 23213 6307
rect 23213 6273 23247 6307
rect 23247 6273 23256 6307
rect 23204 6264 23256 6273
rect 23388 6307 23440 6316
rect 23388 6273 23397 6307
rect 23397 6273 23431 6307
rect 23431 6273 23440 6307
rect 29552 6332 29604 6384
rect 23388 6264 23440 6273
rect 27712 6307 27764 6316
rect 27712 6273 27746 6307
rect 27746 6273 27764 6307
rect 27712 6264 27764 6273
rect 26148 6196 26200 6248
rect 22836 6128 22888 6180
rect 20536 6060 20588 6112
rect 23664 6060 23716 6112
rect 46848 6400 46900 6452
rect 32220 6332 32272 6384
rect 32496 6375 32548 6384
rect 32496 6341 32505 6375
rect 32505 6341 32539 6375
rect 32539 6341 32548 6375
rect 32496 6332 32548 6341
rect 32588 6264 32640 6316
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 3424 5856 3476 5908
rect 32128 5856 32180 5908
rect 21640 5831 21692 5840
rect 21640 5797 21649 5831
rect 21649 5797 21683 5831
rect 21683 5797 21692 5831
rect 21640 5788 21692 5797
rect 20260 5763 20312 5772
rect 20260 5729 20269 5763
rect 20269 5729 20303 5763
rect 20303 5729 20312 5763
rect 20260 5720 20312 5729
rect 2320 5652 2372 5704
rect 2964 5695 3016 5704
rect 2964 5661 2973 5695
rect 2973 5661 3007 5695
rect 3007 5661 3016 5695
rect 2964 5652 3016 5661
rect 20076 5652 20128 5704
rect 20536 5695 20588 5704
rect 20536 5661 20570 5695
rect 20570 5661 20588 5695
rect 20536 5652 20588 5661
rect 23480 5652 23532 5704
rect 47860 5695 47912 5704
rect 47860 5661 47869 5695
rect 47869 5661 47903 5695
rect 47903 5661 47912 5695
rect 47860 5652 47912 5661
rect 4804 5584 4856 5636
rect 1584 5516 1636 5568
rect 3884 5559 3936 5568
rect 3884 5525 3893 5559
rect 3893 5525 3927 5559
rect 3927 5525 3936 5559
rect 3884 5516 3936 5525
rect 19340 5559 19392 5568
rect 19340 5525 19349 5559
rect 19349 5525 19383 5559
rect 19383 5525 19392 5559
rect 19340 5516 19392 5525
rect 22192 5584 22244 5636
rect 32036 5584 32088 5636
rect 33048 5584 33100 5636
rect 23848 5559 23900 5568
rect 23848 5525 23857 5559
rect 23857 5525 23891 5559
rect 23891 5525 23900 5559
rect 23848 5516 23900 5525
rect 28632 5516 28684 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 2964 5312 3016 5364
rect 3424 5312 3476 5364
rect 10968 5312 11020 5364
rect 20628 5355 20680 5364
rect 20628 5321 20637 5355
rect 20637 5321 20671 5355
rect 20671 5321 20680 5355
rect 20628 5312 20680 5321
rect 22192 5312 22244 5364
rect 24768 5355 24820 5364
rect 24768 5321 24777 5355
rect 24777 5321 24811 5355
rect 24811 5321 24820 5355
rect 24768 5312 24820 5321
rect 38568 5312 38620 5364
rect 46848 5312 46900 5364
rect 3884 5244 3936 5296
rect 19340 5244 19392 5296
rect 46756 5244 46808 5296
rect 2780 5151 2832 5160
rect 2780 5117 2789 5151
rect 2789 5117 2823 5151
rect 2823 5117 2832 5151
rect 2780 5108 2832 5117
rect 18696 5108 18748 5160
rect 18788 5108 18840 5160
rect 21088 5219 21140 5228
rect 21088 5185 21097 5219
rect 21097 5185 21131 5219
rect 21131 5185 21140 5219
rect 21088 5176 21140 5185
rect 21272 5219 21324 5228
rect 21272 5185 21281 5219
rect 21281 5185 21315 5219
rect 21315 5185 21324 5219
rect 21272 5176 21324 5185
rect 22284 5176 22336 5228
rect 22468 5219 22520 5228
rect 22468 5185 22477 5219
rect 22477 5185 22511 5219
rect 22511 5185 22520 5219
rect 22468 5176 22520 5185
rect 22560 5219 22612 5228
rect 22560 5185 22569 5219
rect 22569 5185 22603 5219
rect 22603 5185 22612 5219
rect 22560 5176 22612 5185
rect 22468 5040 22520 5092
rect 1400 4972 1452 5024
rect 21272 4972 21324 5024
rect 23480 5176 23532 5228
rect 23664 5219 23716 5228
rect 23664 5185 23698 5219
rect 23698 5185 23716 5219
rect 23664 5176 23716 5185
rect 45652 5176 45704 5228
rect 46296 4972 46348 5024
rect 47676 5015 47728 5024
rect 47676 4981 47685 5015
rect 47685 4981 47719 5015
rect 47719 4981 47728 5015
rect 47676 4972 47728 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 22560 4768 22612 4820
rect 2504 4700 2556 4752
rect 1400 4675 1452 4684
rect 1400 4641 1409 4675
rect 1409 4641 1443 4675
rect 1443 4641 1452 4675
rect 1400 4632 1452 4641
rect 1584 4675 1636 4684
rect 1584 4641 1593 4675
rect 1593 4641 1627 4675
rect 1627 4641 1636 4675
rect 1584 4632 1636 4641
rect 2780 4675 2832 4684
rect 2780 4641 2789 4675
rect 2789 4641 2823 4675
rect 2823 4641 2832 4675
rect 2780 4632 2832 4641
rect 4620 4607 4672 4616
rect 4620 4573 4629 4607
rect 4629 4573 4663 4607
rect 4663 4573 4672 4607
rect 4620 4564 4672 4573
rect 20168 4700 20220 4752
rect 32220 4700 32272 4752
rect 27896 4632 27948 4684
rect 46296 4675 46348 4684
rect 20076 4564 20128 4616
rect 21824 4564 21876 4616
rect 23848 4564 23900 4616
rect 31208 4564 31260 4616
rect 46296 4641 46305 4675
rect 46305 4641 46339 4675
rect 46339 4641 46348 4675
rect 46296 4632 46348 4641
rect 47676 4632 47728 4684
rect 48136 4675 48188 4684
rect 48136 4641 48145 4675
rect 48145 4641 48179 4675
rect 48179 4641 48188 4675
rect 48136 4632 48188 4641
rect 14096 4496 14148 4548
rect 11704 4428 11756 4480
rect 12440 4471 12492 4480
rect 12440 4437 12449 4471
rect 12449 4437 12483 4471
rect 12483 4437 12492 4471
rect 12440 4428 12492 4437
rect 18144 4428 18196 4480
rect 40224 4428 40276 4480
rect 40500 4471 40552 4480
rect 40500 4437 40509 4471
rect 40509 4437 40543 4471
rect 40543 4437 40552 4471
rect 40500 4428 40552 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 19340 4224 19392 4276
rect 11704 4199 11756 4208
rect 11704 4165 11713 4199
rect 11713 4165 11747 4199
rect 11747 4165 11756 4199
rect 11704 4156 11756 4165
rect 4804 4131 4856 4140
rect 4804 4097 4813 4131
rect 4813 4097 4847 4131
rect 4847 4097 4856 4131
rect 4804 4088 4856 4097
rect 8116 4020 8168 4072
rect 9312 4063 9364 4072
rect 2596 3952 2648 4004
rect 8024 3952 8076 4004
rect 9312 4029 9321 4063
rect 9321 4029 9355 4063
rect 9355 4029 9364 4063
rect 9312 4020 9364 4029
rect 9404 4020 9456 4072
rect 10140 4020 10192 4072
rect 12532 4063 12584 4072
rect 12532 4029 12541 4063
rect 12541 4029 12575 4063
rect 12575 4029 12584 4063
rect 12532 4020 12584 4029
rect 18696 4088 18748 4140
rect 19432 4088 19484 4140
rect 19340 4020 19392 4072
rect 20904 4088 20956 4140
rect 20812 4020 20864 4072
rect 23940 4088 23992 4140
rect 28908 4088 28960 4140
rect 37280 4224 37332 4276
rect 37740 4224 37792 4276
rect 29460 4156 29512 4208
rect 29184 4088 29236 4140
rect 29828 4088 29880 4140
rect 30932 4131 30984 4140
rect 30932 4097 30941 4131
rect 30941 4097 30975 4131
rect 30975 4097 30984 4131
rect 30932 4088 30984 4097
rect 31760 4088 31812 4140
rect 36176 4131 36228 4140
rect 36176 4097 36185 4131
rect 36185 4097 36219 4131
rect 36219 4097 36228 4131
rect 36176 4088 36228 4097
rect 37832 4131 37884 4140
rect 37832 4097 37841 4131
rect 37841 4097 37875 4131
rect 37875 4097 37884 4131
rect 37832 4088 37884 4097
rect 35348 4020 35400 4072
rect 10692 3952 10744 4004
rect 10784 3952 10836 4004
rect 1400 3884 1452 3936
rect 3792 3884 3844 3936
rect 3976 3884 4028 3936
rect 4896 3927 4948 3936
rect 4896 3893 4905 3927
rect 4905 3893 4939 3927
rect 4939 3893 4948 3927
rect 4896 3884 4948 3893
rect 6460 3884 6512 3936
rect 10324 3884 10376 3936
rect 13268 3884 13320 3936
rect 14280 3884 14332 3936
rect 15108 3884 15160 3936
rect 17960 3884 18012 3936
rect 22560 3952 22612 4004
rect 30932 3952 30984 4004
rect 31116 3952 31168 4004
rect 19984 3884 20036 3936
rect 20260 3884 20312 3936
rect 20904 3927 20956 3936
rect 20904 3893 20913 3927
rect 20913 3893 20947 3927
rect 20947 3893 20956 3927
rect 20904 3884 20956 3893
rect 23572 3884 23624 3936
rect 25964 3884 26016 3936
rect 29736 3884 29788 3936
rect 31392 3884 31444 3936
rect 32404 3884 32456 3936
rect 32956 3927 33008 3936
rect 32956 3893 32965 3927
rect 32965 3893 32999 3927
rect 32999 3893 33008 3927
rect 32956 3884 33008 3893
rect 36452 3884 36504 3936
rect 38016 3884 38068 3936
rect 46756 4156 46808 4208
rect 38660 4063 38712 4072
rect 38660 4029 38669 4063
rect 38669 4029 38703 4063
rect 38703 4029 38712 4063
rect 38660 4020 38712 4029
rect 46388 4088 46440 4140
rect 46940 4088 46992 4140
rect 47492 4088 47544 4140
rect 47216 4020 47268 4072
rect 41604 3884 41656 3936
rect 42432 3884 42484 3936
rect 43996 3884 44048 3936
rect 44916 3927 44968 3936
rect 44916 3893 44925 3927
rect 44925 3893 44959 3927
rect 44959 3893 44968 3927
rect 44916 3884 44968 3893
rect 46480 3884 46532 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 3884 3680 3936 3732
rect 9312 3723 9364 3732
rect 3240 3612 3292 3664
rect 9312 3689 9321 3723
rect 9321 3689 9355 3723
rect 9355 3689 9364 3723
rect 9312 3680 9364 3689
rect 11612 3680 11664 3732
rect 13084 3680 13136 3732
rect 1400 3587 1452 3596
rect 1400 3553 1409 3587
rect 1409 3553 1443 3587
rect 1443 3553 1452 3587
rect 1400 3544 1452 3553
rect 1860 3587 1912 3596
rect 1860 3553 1869 3587
rect 1869 3553 1903 3587
rect 1903 3553 1912 3587
rect 1860 3544 1912 3553
rect 3792 3587 3844 3596
rect 3792 3553 3801 3587
rect 3801 3553 3835 3587
rect 3835 3553 3844 3587
rect 3792 3544 3844 3553
rect 3976 3587 4028 3596
rect 3976 3553 3985 3587
rect 3985 3553 4019 3587
rect 4019 3553 4028 3587
rect 3976 3544 4028 3553
rect 12164 3612 12216 3664
rect 12256 3612 12308 3664
rect 12440 3544 12492 3596
rect 12624 3612 12676 3664
rect 17868 3680 17920 3732
rect 21456 3680 21508 3732
rect 14096 3612 14148 3664
rect 26884 3612 26936 3664
rect 27528 3612 27580 3664
rect 31116 3612 31168 3664
rect 38660 3680 38712 3732
rect 43444 3680 43496 3732
rect 47032 3680 47084 3732
rect 48044 3612 48096 3664
rect 6092 3519 6144 3528
rect 6092 3485 6101 3519
rect 6101 3485 6135 3519
rect 6135 3485 6144 3519
rect 6092 3476 6144 3485
rect 6368 3476 6420 3528
rect 10784 3476 10836 3528
rect 15108 3587 15160 3596
rect 15108 3553 15117 3587
rect 15117 3553 15151 3587
rect 15151 3553 15160 3587
rect 15108 3544 15160 3553
rect 15476 3587 15528 3596
rect 15476 3553 15485 3587
rect 15485 3553 15519 3587
rect 15519 3553 15528 3587
rect 15476 3544 15528 3553
rect 20260 3587 20312 3596
rect 20260 3553 20269 3587
rect 20269 3553 20303 3587
rect 20303 3553 20312 3587
rect 20260 3544 20312 3553
rect 20628 3587 20680 3596
rect 20628 3553 20637 3587
rect 20637 3553 20671 3587
rect 20671 3553 20680 3587
rect 20628 3544 20680 3553
rect 25964 3587 26016 3596
rect 25964 3553 25973 3587
rect 25973 3553 26007 3587
rect 26007 3553 26016 3587
rect 25964 3544 26016 3553
rect 26424 3587 26476 3596
rect 26424 3553 26433 3587
rect 26433 3553 26467 3587
rect 26467 3553 26476 3587
rect 26424 3544 26476 3553
rect 14924 3519 14976 3528
rect 14924 3485 14933 3519
rect 14933 3485 14967 3519
rect 14967 3485 14976 3519
rect 14924 3476 14976 3485
rect 20076 3519 20128 3528
rect 20076 3485 20085 3519
rect 20085 3485 20119 3519
rect 20119 3485 20128 3519
rect 20076 3476 20128 3485
rect 23388 3476 23440 3528
rect 25780 3519 25832 3528
rect 25780 3485 25789 3519
rect 25789 3485 25823 3519
rect 25823 3485 25832 3519
rect 25780 3476 25832 3485
rect 2136 3408 2188 3460
rect 8944 3408 8996 3460
rect 18788 3408 18840 3460
rect 20812 3408 20864 3460
rect 25688 3408 25740 3460
rect 29000 3519 29052 3528
rect 29000 3485 29009 3519
rect 29009 3485 29043 3519
rect 29043 3485 29052 3519
rect 29000 3476 29052 3485
rect 29276 3476 29328 3528
rect 31576 3544 31628 3596
rect 36452 3587 36504 3596
rect 36452 3553 36461 3587
rect 36461 3553 36495 3587
rect 36495 3553 36504 3587
rect 36452 3544 36504 3553
rect 36728 3587 36780 3596
rect 36728 3553 36737 3587
rect 36737 3553 36771 3587
rect 36771 3553 36780 3587
rect 36728 3544 36780 3553
rect 37188 3544 37240 3596
rect 41604 3587 41656 3596
rect 31208 3519 31260 3528
rect 31208 3485 31217 3519
rect 31217 3485 31251 3519
rect 31251 3485 31260 3519
rect 31208 3476 31260 3485
rect 36268 3519 36320 3528
rect 36268 3485 36277 3519
rect 36277 3485 36311 3519
rect 36311 3485 36320 3519
rect 36268 3476 36320 3485
rect 41604 3553 41613 3587
rect 41613 3553 41647 3587
rect 41647 3553 41656 3587
rect 41604 3544 41656 3553
rect 41880 3587 41932 3596
rect 41880 3553 41889 3587
rect 41889 3553 41923 3587
rect 41923 3553 41932 3587
rect 41880 3544 41932 3553
rect 42064 3544 42116 3596
rect 46204 3544 46256 3596
rect 46480 3587 46532 3596
rect 46480 3553 46489 3587
rect 46489 3553 46523 3587
rect 46523 3553 46532 3587
rect 46480 3544 46532 3553
rect 43904 3519 43956 3528
rect 43904 3485 43913 3519
rect 43913 3485 43947 3519
rect 43947 3485 43956 3519
rect 43904 3476 43956 3485
rect 29644 3451 29696 3460
rect 29644 3417 29653 3451
rect 29653 3417 29687 3451
rect 29687 3417 29696 3451
rect 29644 3408 29696 3417
rect 29828 3408 29880 3460
rect 31392 3451 31444 3460
rect 1308 3340 1360 3392
rect 3332 3340 3384 3392
rect 6552 3340 6604 3392
rect 6920 3340 6972 3392
rect 12440 3340 12492 3392
rect 14648 3340 14700 3392
rect 25504 3340 25556 3392
rect 29460 3340 29512 3392
rect 29920 3340 29972 3392
rect 31392 3417 31401 3451
rect 31401 3417 31435 3451
rect 31435 3417 31444 3451
rect 31392 3408 31444 3417
rect 43444 3408 43496 3460
rect 46940 3408 46992 3460
rect 48320 3408 48372 3460
rect 40040 3340 40092 3392
rect 44180 3340 44232 3392
rect 45192 3340 45244 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 2136 3179 2188 3188
rect 2136 3145 2145 3179
rect 2145 3145 2179 3179
rect 2179 3145 2188 3179
rect 2136 3136 2188 3145
rect 2412 3136 2464 3188
rect 22560 3136 22612 3188
rect 22652 3136 22704 3188
rect 4896 3068 4948 3120
rect 6552 3111 6604 3120
rect 6552 3077 6561 3111
rect 6561 3077 6595 3111
rect 6595 3077 6604 3111
rect 6552 3068 6604 3077
rect 17868 3068 17920 3120
rect 18144 3111 18196 3120
rect 18144 3077 18153 3111
rect 18153 3077 18187 3111
rect 18187 3077 18196 3111
rect 18144 3068 18196 3077
rect 19984 3068 20036 3120
rect 1952 3000 2004 3052
rect 6368 3043 6420 3052
rect 6368 3009 6377 3043
rect 6377 3009 6411 3043
rect 6411 3009 6420 3043
rect 6368 3000 6420 3009
rect 8944 3043 8996 3052
rect 8944 3009 8953 3043
rect 8953 3009 8987 3043
rect 8987 3009 8996 3043
rect 8944 3000 8996 3009
rect 9680 3000 9732 3052
rect 12164 3000 12216 3052
rect 14188 3000 14240 3052
rect 14924 3000 14976 3052
rect 17960 3043 18012 3052
rect 17960 3009 17969 3043
rect 17969 3009 18003 3043
rect 18003 3009 18012 3043
rect 17960 3000 18012 3009
rect 20076 3000 20128 3052
rect 22560 3000 22612 3052
rect 4620 2932 4672 2984
rect 5172 2975 5224 2984
rect 5172 2941 5181 2975
rect 5181 2941 5215 2975
rect 5215 2941 5224 2975
rect 5172 2932 5224 2941
rect 6552 2932 6604 2984
rect 7748 2932 7800 2984
rect 12440 2975 12492 2984
rect 12440 2941 12449 2975
rect 12449 2941 12483 2975
rect 12483 2941 12492 2975
rect 12900 2975 12952 2984
rect 12440 2932 12492 2941
rect 12900 2941 12909 2975
rect 12909 2941 12943 2975
rect 12943 2941 12952 2975
rect 12900 2932 12952 2941
rect 18144 2932 18196 2984
rect 14648 2864 14700 2916
rect 23572 3111 23624 3120
rect 23572 3077 23581 3111
rect 23581 3077 23615 3111
rect 23615 3077 23624 3111
rect 23572 3068 23624 3077
rect 26148 3136 26200 3188
rect 28908 3136 28960 3188
rect 30840 3136 30892 3188
rect 36176 3136 36228 3188
rect 29920 3111 29972 3120
rect 23388 3043 23440 3052
rect 23388 3009 23397 3043
rect 23397 3009 23431 3043
rect 23431 3009 23440 3043
rect 23388 3000 23440 3009
rect 25780 3000 25832 3052
rect 23848 2975 23900 2984
rect 23848 2941 23857 2975
rect 23857 2941 23891 2975
rect 23891 2941 23900 2975
rect 23848 2932 23900 2941
rect 23204 2864 23256 2916
rect 29920 3077 29929 3111
rect 29929 3077 29963 3111
rect 29963 3077 29972 3111
rect 29920 3068 29972 3077
rect 32404 3111 32456 3120
rect 32404 3077 32413 3111
rect 32413 3077 32447 3111
rect 32447 3077 32456 3111
rect 32404 3068 32456 3077
rect 33048 3068 33100 3120
rect 40224 3111 40276 3120
rect 29736 3043 29788 3052
rect 29736 3009 29745 3043
rect 29745 3009 29779 3043
rect 29779 3009 29788 3043
rect 29736 3000 29788 3009
rect 36268 3000 36320 3052
rect 30288 2975 30340 2984
rect 30288 2941 30297 2975
rect 30297 2941 30331 2975
rect 30331 2941 30340 2975
rect 30288 2932 30340 2941
rect 32956 2932 33008 2984
rect 37740 2932 37792 2984
rect 30748 2864 30800 2916
rect 33508 2864 33560 2916
rect 10968 2796 11020 2848
rect 16580 2796 16632 2848
rect 22008 2796 22060 2848
rect 26884 2796 26936 2848
rect 33416 2796 33468 2848
rect 39580 2839 39632 2848
rect 39580 2805 39589 2839
rect 39589 2805 39623 2839
rect 39623 2805 39632 2839
rect 39580 2796 39632 2805
rect 40224 3077 40233 3111
rect 40233 3077 40267 3111
rect 40267 3077 40276 3111
rect 40224 3068 40276 3077
rect 40408 3136 40460 3188
rect 43904 3136 43956 3188
rect 46112 3136 46164 3188
rect 48044 3179 48096 3188
rect 48044 3145 48053 3179
rect 48053 3145 48087 3179
rect 48087 3145 48096 3179
rect 48044 3136 48096 3145
rect 44180 3111 44232 3120
rect 40500 2932 40552 2984
rect 41236 2975 41288 2984
rect 41236 2941 41245 2975
rect 41245 2941 41279 2975
rect 41279 2941 41288 2975
rect 41236 2932 41288 2941
rect 40408 2864 40460 2916
rect 42616 2796 42668 2848
rect 44180 3077 44189 3111
rect 44189 3077 44223 3111
rect 44223 3077 44232 3111
rect 44180 3068 44232 3077
rect 43168 3000 43220 3052
rect 43996 3043 44048 3052
rect 43996 3009 44005 3043
rect 44005 3009 44039 3043
rect 44039 3009 44048 3043
rect 43996 3000 44048 3009
rect 45744 3000 45796 3052
rect 49608 3000 49660 3052
rect 44456 2975 44508 2984
rect 44456 2941 44465 2975
rect 44465 2941 44499 2975
rect 44499 2941 44508 2975
rect 44456 2932 44508 2941
rect 43444 2907 43496 2916
rect 43444 2873 43453 2907
rect 43453 2873 43487 2907
rect 43487 2873 43496 2907
rect 43444 2864 43496 2873
rect 45652 2796 45704 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 3148 2592 3200 2644
rect 3700 2524 3752 2576
rect 4804 2567 4856 2576
rect 4804 2533 4813 2567
rect 4813 2533 4847 2567
rect 4847 2533 4856 2567
rect 4804 2524 4856 2533
rect 5816 2524 5868 2576
rect 6460 2499 6512 2508
rect 6460 2465 6469 2499
rect 6469 2465 6503 2499
rect 6503 2465 6512 2499
rect 6460 2456 6512 2465
rect 6920 2456 6972 2508
rect 7104 2456 7156 2508
rect 12164 2592 12216 2644
rect 22100 2592 22152 2644
rect 45836 2592 45888 2644
rect 12532 2456 12584 2508
rect 13544 2456 13596 2508
rect 1952 2388 2004 2440
rect 4528 2388 4580 2440
rect 1860 2363 1912 2372
rect 1860 2329 1869 2363
rect 1869 2329 1903 2363
rect 1903 2329 1912 2363
rect 1860 2320 1912 2329
rect 2228 2363 2280 2372
rect 2228 2329 2237 2363
rect 2237 2329 2271 2363
rect 2271 2329 2280 2363
rect 2228 2320 2280 2329
rect 8392 2320 8444 2372
rect 17408 2388 17460 2440
rect 14280 2363 14332 2372
rect 14280 2329 14289 2363
rect 14289 2329 14323 2363
rect 14323 2329 14332 2363
rect 14280 2320 14332 2329
rect 19984 2320 20036 2372
rect 20996 2524 21048 2576
rect 21272 2524 21324 2576
rect 20904 2456 20956 2508
rect 22008 2499 22060 2508
rect 22008 2465 22017 2499
rect 22017 2465 22051 2499
rect 22051 2465 22060 2499
rect 22008 2456 22060 2465
rect 23112 2524 23164 2576
rect 28080 2524 28132 2576
rect 32680 2524 32732 2576
rect 39948 2524 40000 2576
rect 24676 2456 24728 2508
rect 26148 2456 26200 2508
rect 28724 2456 28776 2508
rect 29000 2456 29052 2508
rect 29736 2499 29788 2508
rect 29736 2465 29745 2499
rect 29745 2465 29779 2499
rect 29779 2465 29788 2499
rect 29736 2456 29788 2465
rect 30932 2499 30984 2508
rect 30932 2465 30941 2499
rect 30941 2465 30975 2499
rect 30975 2465 30984 2499
rect 30932 2456 30984 2465
rect 32496 2456 32548 2508
rect 39580 2456 39632 2508
rect 40040 2499 40092 2508
rect 40040 2465 40049 2499
rect 40049 2465 40083 2499
rect 40083 2465 40092 2499
rect 40040 2456 40092 2465
rect 42432 2499 42484 2508
rect 42432 2465 42441 2499
rect 42441 2465 42475 2499
rect 42475 2465 42484 2499
rect 42432 2456 42484 2465
rect 42616 2499 42668 2508
rect 42616 2465 42625 2499
rect 42625 2465 42659 2499
rect 42659 2465 42668 2499
rect 42616 2456 42668 2465
rect 42708 2456 42760 2508
rect 44916 2456 44968 2508
rect 45192 2499 45244 2508
rect 45192 2465 45201 2499
rect 45201 2465 45235 2499
rect 45235 2465 45244 2499
rect 45192 2456 45244 2465
rect 45376 2456 45428 2508
rect 22928 2320 22980 2372
rect 25136 2320 25188 2372
rect 27068 2388 27120 2440
rect 28264 2388 28316 2440
rect 32864 2388 32916 2440
rect 15200 2252 15252 2304
rect 17684 2295 17736 2304
rect 17684 2261 17693 2295
rect 17693 2261 17727 2295
rect 17727 2261 17736 2295
rect 17684 2252 17736 2261
rect 24492 2252 24544 2304
rect 27712 2320 27764 2372
rect 28448 2320 28500 2372
rect 38660 2388 38712 2440
rect 38752 2431 38804 2440
rect 38752 2397 38761 2431
rect 38761 2397 38795 2431
rect 38795 2397 38804 2431
rect 38752 2388 38804 2397
rect 34152 2320 34204 2372
rect 34796 2320 34848 2372
rect 36084 2320 36136 2372
rect 47768 2363 47820 2372
rect 47768 2329 47777 2363
rect 47777 2329 47811 2363
rect 47811 2329 47820 2363
rect 47768 2320 47820 2329
rect 26148 2252 26200 2304
rect 47860 2295 47912 2304
rect 47860 2261 47869 2295
rect 47869 2261 47903 2295
rect 47903 2261 47912 2295
rect 47860 2252 47912 2261
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 24308 1980 24360 2032
rect 47860 1980 47912 2032
rect 22284 1912 22336 1964
rect 38752 1912 38804 1964
rect 17684 1844 17736 1896
rect 31668 1844 31720 1896
<< metal2 >>
rect 18 51200 74 52000
rect 662 51200 718 52000
rect 1306 51200 1362 52000
rect 1950 51354 2006 52000
rect 1950 51326 2176 51354
rect 1950 51200 2006 51326
rect 32 48278 60 51200
rect 676 49230 704 51200
rect 664 49224 716 49230
rect 664 49166 716 49172
rect 20 48272 72 48278
rect 20 48214 72 48220
rect 1320 48210 1348 51200
rect 1676 49088 1728 49094
rect 1676 49030 1728 49036
rect 1308 48204 1360 48210
rect 1308 48146 1360 48152
rect 1584 48068 1636 48074
rect 1584 48010 1636 48016
rect 1596 47802 1624 48010
rect 1584 47796 1636 47802
rect 1584 47738 1636 47744
rect 1398 47696 1454 47705
rect 1398 47631 1454 47640
rect 1412 46578 1440 47631
rect 1584 46980 1636 46986
rect 1584 46922 1636 46928
rect 1596 46714 1624 46922
rect 1584 46708 1636 46714
rect 1584 46650 1636 46656
rect 1400 46572 1452 46578
rect 1400 46514 1452 46520
rect 1584 46368 1636 46374
rect 1584 46310 1636 46316
rect 1492 45280 1544 45286
rect 1492 45222 1544 45228
rect 1400 42016 1452 42022
rect 1400 41958 1452 41964
rect 1412 41682 1440 41958
rect 1400 41676 1452 41682
rect 1400 41618 1452 41624
rect 1400 40928 1452 40934
rect 1400 40870 1452 40876
rect 1412 35170 1440 40870
rect 1504 35306 1532 45222
rect 1596 35494 1624 46310
rect 1584 35488 1636 35494
rect 1584 35430 1636 35436
rect 1504 35278 1624 35306
rect 1412 35142 1532 35170
rect 1400 35080 1452 35086
rect 1400 35022 1452 35028
rect 1412 34785 1440 35022
rect 1398 34776 1454 34785
rect 1398 34711 1454 34720
rect 1400 34400 1452 34406
rect 1400 34342 1452 34348
rect 1412 34066 1440 34342
rect 1400 34060 1452 34066
rect 1400 34002 1452 34008
rect 1400 31816 1452 31822
rect 1400 31758 1452 31764
rect 1412 31385 1440 31758
rect 1398 31376 1454 31385
rect 1398 31311 1454 31320
rect 1400 28960 1452 28966
rect 1400 28902 1452 28908
rect 1412 28626 1440 28902
rect 1400 28620 1452 28626
rect 1400 28562 1452 28568
rect 1400 27464 1452 27470
rect 1400 27406 1452 27412
rect 1308 26512 1360 26518
rect 1308 26454 1360 26460
rect 1320 25786 1348 26454
rect 1412 26450 1440 27406
rect 1400 26444 1452 26450
rect 1400 26386 1452 26392
rect 1398 25936 1454 25945
rect 1398 25871 1400 25880
rect 1452 25871 1454 25880
rect 1400 25842 1452 25848
rect 1320 25758 1440 25786
rect 1412 21078 1440 25758
rect 1504 23798 1532 35142
rect 1596 26518 1624 35278
rect 1584 26512 1636 26518
rect 1584 26454 1636 26460
rect 1584 26308 1636 26314
rect 1584 26250 1636 26256
rect 1596 26042 1624 26250
rect 1584 26036 1636 26042
rect 1584 25978 1636 25984
rect 1584 25696 1636 25702
rect 1584 25638 1636 25644
rect 1492 23792 1544 23798
rect 1492 23734 1544 23740
rect 1596 23322 1624 25638
rect 1584 23316 1636 23322
rect 1584 23258 1636 23264
rect 1400 21072 1452 21078
rect 1400 21014 1452 21020
rect 1584 18080 1636 18086
rect 1584 18022 1636 18028
rect 1596 17746 1624 18022
rect 1584 17740 1636 17746
rect 1584 17682 1636 17688
rect 1688 15638 1716 49030
rect 2148 47734 2176 51326
rect 2594 51200 2650 52000
rect 2870 51776 2926 51785
rect 2870 51711 2926 51720
rect 2884 48822 2912 51711
rect 3238 51200 3294 52000
rect 3882 51200 3938 52000
rect 4526 51354 4582 52000
rect 4526 51326 4660 51354
rect 4526 51200 4582 51326
rect 3252 49230 3280 51200
rect 3422 51096 3478 51105
rect 3422 51031 3478 51040
rect 3436 49774 3464 51031
rect 3424 49768 3476 49774
rect 3424 49710 3476 49716
rect 4214 49532 4522 49552
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49456 4522 49476
rect 3976 49292 4028 49298
rect 3976 49234 4028 49240
rect 4068 49292 4120 49298
rect 4068 49234 4120 49240
rect 3240 49224 3292 49230
rect 3240 49166 3292 49172
rect 3148 49088 3200 49094
rect 3148 49030 3200 49036
rect 2872 48816 2924 48822
rect 2872 48758 2924 48764
rect 3056 48680 3108 48686
rect 3056 48622 3108 48628
rect 3068 47802 3096 48622
rect 3056 47796 3108 47802
rect 3056 47738 3108 47744
rect 2136 47728 2188 47734
rect 2136 47670 2188 47676
rect 2504 47592 2556 47598
rect 2504 47534 2556 47540
rect 1952 47456 2004 47462
rect 1952 47398 2004 47404
rect 1860 47116 1912 47122
rect 1860 47058 1912 47064
rect 1872 47025 1900 47058
rect 1858 47016 1914 47025
rect 1858 46951 1914 46960
rect 1858 45656 1914 45665
rect 1858 45591 1914 45600
rect 1872 45558 1900 45591
rect 1860 45552 1912 45558
rect 1860 45494 1912 45500
rect 1858 44296 1914 44305
rect 1858 44231 1914 44240
rect 1872 43790 1900 44231
rect 1860 43784 1912 43790
rect 1860 43726 1912 43732
rect 1858 43616 1914 43625
rect 1858 43551 1914 43560
rect 1872 43382 1900 43551
rect 1860 43376 1912 43382
rect 1860 43318 1912 43324
rect 1860 41676 1912 41682
rect 1860 41618 1912 41624
rect 1872 41585 1900 41618
rect 1858 41576 1914 41585
rect 1858 41511 1914 41520
rect 1860 41132 1912 41138
rect 1860 41074 1912 41080
rect 1872 40905 1900 41074
rect 1858 40896 1914 40905
rect 1858 40831 1914 40840
rect 1860 40452 1912 40458
rect 1860 40394 1912 40400
rect 1872 40225 1900 40394
rect 1858 40216 1914 40225
rect 1858 40151 1914 40160
rect 1860 37868 1912 37874
rect 1860 37810 1912 37816
rect 1872 37505 1900 37810
rect 1858 37496 1914 37505
rect 1858 37431 1914 37440
rect 1860 37188 1912 37194
rect 1860 37130 1912 37136
rect 1872 36825 1900 37130
rect 1858 36816 1914 36825
rect 1858 36751 1914 36760
rect 1964 35894 1992 47398
rect 2136 46572 2188 46578
rect 2136 46514 2188 46520
rect 2044 44872 2096 44878
rect 2044 44814 2096 44820
rect 2056 44402 2084 44814
rect 2044 44396 2096 44402
rect 2044 44338 2096 44344
rect 2148 43246 2176 46514
rect 2228 44736 2280 44742
rect 2228 44678 2280 44684
rect 2240 44470 2268 44678
rect 2228 44464 2280 44470
rect 2228 44406 2280 44412
rect 2320 43716 2372 43722
rect 2320 43658 2372 43664
rect 2136 43240 2188 43246
rect 2136 43182 2188 43188
rect 2136 41132 2188 41138
rect 2136 41074 2188 41080
rect 2044 39840 2096 39846
rect 2044 39782 2096 39788
rect 2056 38962 2084 39782
rect 2044 38956 2096 38962
rect 2044 38898 2096 38904
rect 2044 36168 2096 36174
rect 2044 36110 2096 36116
rect 1872 35866 1992 35894
rect 1768 34536 1820 34542
rect 1768 34478 1820 34484
rect 1780 33522 1808 34478
rect 1768 33516 1820 33522
rect 1768 33458 1820 33464
rect 1768 30728 1820 30734
rect 1768 30670 1820 30676
rect 1780 30258 1808 30670
rect 1768 30252 1820 30258
rect 1768 30194 1820 30200
rect 1768 29640 1820 29646
rect 1768 29582 1820 29588
rect 1780 29170 1808 29582
rect 1768 29164 1820 29170
rect 1768 29106 1820 29112
rect 1768 27396 1820 27402
rect 1768 27338 1820 27344
rect 1780 26994 1808 27338
rect 1768 26988 1820 26994
rect 1768 26930 1820 26936
rect 1872 26234 1900 35866
rect 2056 35698 2084 36110
rect 2148 35894 2176 41074
rect 2228 39296 2280 39302
rect 2228 39238 2280 39244
rect 2240 39030 2268 39238
rect 2228 39024 2280 39030
rect 2228 38966 2280 38972
rect 2148 35866 2268 35894
rect 2044 35692 2096 35698
rect 2044 35634 2096 35640
rect 2044 34604 2096 34610
rect 2044 34546 2096 34552
rect 1952 33448 2004 33454
rect 1952 33390 2004 33396
rect 1964 33114 1992 33390
rect 1952 33108 2004 33114
rect 1952 33050 2004 33056
rect 2056 32994 2084 34546
rect 2136 34400 2188 34406
rect 2136 34342 2188 34348
rect 2148 34066 2176 34342
rect 2136 34060 2188 34066
rect 2136 34002 2188 34008
rect 2056 32966 2176 32994
rect 2044 32836 2096 32842
rect 2044 32778 2096 32784
rect 2056 32434 2084 32778
rect 2044 32428 2096 32434
rect 2044 32370 2096 32376
rect 1952 31816 2004 31822
rect 1952 31758 2004 31764
rect 1964 31346 1992 31758
rect 1952 31340 2004 31346
rect 1952 31282 2004 31288
rect 2148 31090 2176 32966
rect 2056 31062 2176 31090
rect 1952 29504 2004 29510
rect 1952 29446 2004 29452
rect 1964 29238 1992 29446
rect 1952 29232 2004 29238
rect 1952 29174 2004 29180
rect 2056 27470 2084 31062
rect 2136 30184 2188 30190
rect 2136 30126 2188 30132
rect 2148 29850 2176 30126
rect 2136 29844 2188 29850
rect 2136 29786 2188 29792
rect 2240 29730 2268 35866
rect 2332 31249 2360 43658
rect 2412 43104 2464 43110
rect 2412 43046 2464 43052
rect 2318 31240 2374 31249
rect 2318 31175 2374 31184
rect 2424 31090 2452 43046
rect 2148 29702 2268 29730
rect 2332 31062 2452 31090
rect 2044 27464 2096 27470
rect 2044 27406 2096 27412
rect 1952 27328 2004 27334
rect 1952 27270 2004 27276
rect 1964 27062 1992 27270
rect 1952 27056 2004 27062
rect 1952 26998 2004 27004
rect 1872 26206 1992 26234
rect 1768 25900 1820 25906
rect 1768 25842 1820 25848
rect 1780 22386 1808 25842
rect 1860 24132 1912 24138
rect 1860 24074 1912 24080
rect 1872 23905 1900 24074
rect 1858 23896 1914 23905
rect 1858 23831 1914 23840
rect 1964 23066 1992 26206
rect 2044 23520 2096 23526
rect 2044 23462 2096 23468
rect 2056 23186 2084 23462
rect 2044 23180 2096 23186
rect 2044 23122 2096 23128
rect 1964 23038 2084 23066
rect 1860 22636 1912 22642
rect 1860 22578 1912 22584
rect 1872 22545 1900 22578
rect 1858 22536 1914 22545
rect 1858 22471 1914 22480
rect 1780 22358 1900 22386
rect 1768 19848 1820 19854
rect 1768 19790 1820 19796
rect 1780 19378 1808 19790
rect 1768 19372 1820 19378
rect 1768 19314 1820 19320
rect 1872 19258 1900 22358
rect 1780 19230 1900 19258
rect 1952 19304 2004 19310
rect 1952 19246 2004 19252
rect 1676 15632 1728 15638
rect 1676 15574 1728 15580
rect 20 14000 72 14006
rect 20 13942 72 13948
rect 32 800 60 13942
rect 1676 13932 1728 13938
rect 1676 13874 1728 13880
rect 1584 13728 1636 13734
rect 1584 13670 1636 13676
rect 1596 13394 1624 13670
rect 1584 13388 1636 13394
rect 1584 13330 1636 13336
rect 1400 12776 1452 12782
rect 1400 12718 1452 12724
rect 1412 12345 1440 12718
rect 1398 12336 1454 12345
rect 1398 12271 1454 12280
rect 1400 10464 1452 10470
rect 1400 10406 1452 10412
rect 1412 10130 1440 10406
rect 1400 10124 1452 10130
rect 1400 10066 1452 10072
rect 664 9376 716 9382
rect 664 9318 716 9324
rect 676 800 704 9318
rect 1688 6914 1716 13874
rect 1780 11150 1808 19230
rect 1964 18970 1992 19246
rect 1952 18964 2004 18970
rect 1952 18906 2004 18912
rect 2056 18902 2084 23038
rect 2148 21434 2176 29702
rect 2332 29594 2360 31062
rect 2410 30968 2466 30977
rect 2410 30903 2466 30912
rect 2240 29566 2360 29594
rect 2240 21554 2268 29566
rect 2320 28484 2372 28490
rect 2320 28426 2372 28432
rect 2332 28218 2360 28426
rect 2320 28212 2372 28218
rect 2320 28154 2372 28160
rect 2320 27464 2372 27470
rect 2320 27406 2372 27412
rect 2332 21894 2360 27406
rect 2320 21888 2372 21894
rect 2320 21830 2372 21836
rect 2424 21622 2452 30903
rect 2516 22642 2544 47534
rect 3056 46504 3108 46510
rect 3056 46446 3108 46452
rect 2872 46368 2924 46374
rect 2872 46310 2924 46316
rect 2962 46336 3018 46345
rect 2884 46034 2912 46310
rect 2962 46271 3018 46280
rect 2976 46034 3004 46271
rect 2872 46028 2924 46034
rect 2872 45970 2924 45976
rect 2964 46028 3016 46034
rect 2964 45970 3016 45976
rect 2872 45892 2924 45898
rect 2872 45834 2924 45840
rect 2884 45490 2912 45834
rect 2872 45484 2924 45490
rect 2872 45426 2924 45432
rect 2778 44976 2834 44985
rect 2778 44911 2834 44920
rect 2792 44334 2820 44911
rect 2780 44328 2832 44334
rect 2780 44270 2832 44276
rect 2596 41540 2648 41546
rect 2596 41482 2648 41488
rect 2608 41274 2636 41482
rect 2596 41268 2648 41274
rect 2596 41210 2648 41216
rect 2778 39536 2834 39545
rect 2778 39471 2834 39480
rect 2792 38894 2820 39471
rect 2780 38888 2832 38894
rect 2780 38830 2832 38836
rect 2596 37732 2648 37738
rect 2596 37674 2648 37680
rect 2608 35894 2636 37674
rect 2778 36136 2834 36145
rect 2778 36071 2834 36080
rect 2608 35866 2728 35894
rect 2596 35488 2648 35494
rect 2596 35430 2648 35436
rect 2608 33318 2636 35430
rect 2596 33312 2648 33318
rect 2596 33254 2648 33260
rect 2596 33108 2648 33114
rect 2596 33050 2648 33056
rect 2608 32026 2636 33050
rect 2700 32502 2728 35866
rect 2792 35630 2820 36071
rect 2964 36032 3016 36038
rect 2964 35974 3016 35980
rect 2976 35766 3004 35974
rect 2964 35760 3016 35766
rect 2964 35702 3016 35708
rect 2780 35624 2832 35630
rect 2780 35566 2832 35572
rect 3068 34610 3096 46446
rect 3056 34604 3108 34610
rect 3056 34546 3108 34552
rect 2778 34096 2834 34105
rect 2778 34031 2780 34040
rect 2832 34031 2834 34040
rect 2780 34002 2832 34008
rect 2780 33448 2832 33454
rect 2778 33416 2780 33425
rect 2832 33416 2834 33425
rect 2778 33351 2834 33360
rect 2780 33312 2832 33318
rect 2780 33254 2832 33260
rect 2688 32496 2740 32502
rect 2688 32438 2740 32444
rect 2792 32314 2820 33254
rect 3054 32736 3110 32745
rect 3054 32671 3110 32680
rect 3068 32366 3096 32671
rect 2700 32286 2820 32314
rect 2964 32360 3016 32366
rect 2964 32302 3016 32308
rect 3056 32360 3108 32366
rect 3056 32302 3108 32308
rect 2596 32020 2648 32026
rect 2596 31962 2648 31968
rect 2700 29782 2728 32286
rect 2976 32026 3004 32302
rect 3054 32056 3110 32065
rect 2964 32020 3016 32026
rect 3054 31991 3110 32000
rect 2964 31962 3016 31968
rect 3068 31278 3096 31991
rect 2872 31272 2924 31278
rect 2872 31214 2924 31220
rect 3056 31272 3108 31278
rect 3056 31214 3108 31220
rect 2884 30938 2912 31214
rect 2872 30932 2924 30938
rect 2872 30874 2924 30880
rect 2780 30184 2832 30190
rect 2780 30126 2832 30132
rect 2792 30025 2820 30126
rect 2778 30016 2834 30025
rect 2778 29951 2834 29960
rect 2688 29776 2740 29782
rect 2688 29718 2740 29724
rect 2778 28656 2834 28665
rect 2778 28591 2780 28600
rect 2832 28591 2834 28600
rect 2780 28562 2832 28568
rect 2778 27296 2834 27305
rect 2778 27231 2834 27240
rect 2792 26926 2820 27231
rect 2780 26920 2832 26926
rect 2780 26862 2832 26868
rect 2778 26616 2834 26625
rect 2778 26551 2834 26560
rect 2792 26450 2820 26551
rect 2780 26444 2832 26450
rect 2780 26386 2832 26392
rect 2688 24132 2740 24138
rect 2688 24074 2740 24080
rect 2596 23044 2648 23050
rect 2596 22986 2648 22992
rect 2608 22778 2636 22986
rect 2596 22772 2648 22778
rect 2596 22714 2648 22720
rect 2504 22636 2556 22642
rect 2504 22578 2556 22584
rect 2412 21616 2464 21622
rect 2412 21558 2464 21564
rect 2228 21548 2280 21554
rect 2228 21490 2280 21496
rect 2148 21406 2360 21434
rect 2228 19304 2280 19310
rect 2228 19246 2280 19252
rect 2240 19145 2268 19246
rect 2226 19136 2282 19145
rect 2226 19071 2282 19080
rect 2044 18896 2096 18902
rect 2044 18838 2096 18844
rect 2136 18284 2188 18290
rect 2136 18226 2188 18232
rect 1860 17196 1912 17202
rect 1860 17138 1912 17144
rect 1872 17105 1900 17138
rect 1858 17096 1914 17105
rect 1858 17031 1914 17040
rect 2044 16584 2096 16590
rect 2044 16526 2096 16532
rect 2056 16114 2084 16526
rect 2044 16108 2096 16114
rect 2044 16050 2096 16056
rect 2148 13938 2176 18226
rect 2228 16448 2280 16454
rect 2228 16390 2280 16396
rect 2240 16182 2268 16390
rect 2228 16176 2280 16182
rect 2228 16118 2280 16124
rect 2136 13932 2188 13938
rect 2136 13874 2188 13880
rect 2332 11914 2360 21406
rect 2412 18760 2464 18766
rect 2412 18702 2464 18708
rect 2056 11886 2360 11914
rect 1768 11144 1820 11150
rect 1768 11086 1820 11092
rect 1860 11076 1912 11082
rect 1860 11018 1912 11024
rect 1952 11076 2004 11082
rect 1952 11018 2004 11024
rect 1872 10985 1900 11018
rect 1858 10976 1914 10985
rect 1858 10911 1914 10920
rect 1964 9518 1992 11018
rect 1952 9512 2004 9518
rect 1952 9454 2004 9460
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 1872 8265 1900 8434
rect 1858 8256 1914 8265
rect 2056 8242 2084 11886
rect 2424 11778 2452 18702
rect 2332 11750 2452 11778
rect 2136 10668 2188 10674
rect 2136 10610 2188 10616
rect 2148 8378 2176 10610
rect 2228 10464 2280 10470
rect 2228 10406 2280 10412
rect 2240 10130 2268 10406
rect 2228 10124 2280 10130
rect 2228 10066 2280 10072
rect 2148 8350 2268 8378
rect 2056 8214 2176 8242
rect 1858 8191 1914 8200
rect 1860 7812 1912 7818
rect 1860 7754 1912 7760
rect 1872 7585 1900 7754
rect 1858 7576 1914 7585
rect 1858 7511 1914 7520
rect 2044 7200 2096 7206
rect 2044 7142 2096 7148
rect 1688 6886 1992 6914
rect 1584 5568 1636 5574
rect 1584 5510 1636 5516
rect 1400 5024 1452 5030
rect 1400 4966 1452 4972
rect 1412 4690 1440 4966
rect 1596 4690 1624 5510
rect 1400 4684 1452 4690
rect 1400 4626 1452 4632
rect 1584 4684 1636 4690
rect 1584 4626 1636 4632
rect 1400 3936 1452 3942
rect 1400 3878 1452 3884
rect 1412 3602 1440 3878
rect 1400 3596 1452 3602
rect 1400 3538 1452 3544
rect 1860 3596 1912 3602
rect 1860 3538 1912 3544
rect 1872 3505 1900 3538
rect 1858 3496 1914 3505
rect 1858 3431 1914 3440
rect 1308 3392 1360 3398
rect 1308 3334 1360 3340
rect 1320 800 1348 3334
rect 1964 3058 1992 6886
rect 2056 6866 2084 7142
rect 2044 6860 2096 6866
rect 2044 6802 2096 6808
rect 2148 6322 2176 8214
rect 2240 6866 2268 8350
rect 2228 6860 2280 6866
rect 2228 6802 2280 6808
rect 2228 6724 2280 6730
rect 2228 6666 2280 6672
rect 2240 6458 2268 6666
rect 2228 6452 2280 6458
rect 2228 6394 2280 6400
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 2332 5710 2360 11750
rect 2412 6860 2464 6866
rect 2412 6802 2464 6808
rect 2320 5704 2372 5710
rect 2320 5646 2372 5652
rect 2136 3460 2188 3466
rect 2136 3402 2188 3408
rect 2148 3194 2176 3402
rect 2424 3194 2452 6802
rect 2516 4758 2544 22578
rect 2700 21690 2728 24074
rect 2778 23216 2834 23225
rect 2778 23151 2780 23160
rect 2832 23151 2834 23160
rect 2780 23122 2832 23128
rect 2688 21684 2740 21690
rect 2688 21626 2740 21632
rect 2872 18080 2924 18086
rect 2872 18022 2924 18028
rect 2884 17814 2912 18022
rect 2872 17808 2924 17814
rect 2778 17776 2834 17785
rect 2872 17750 2924 17756
rect 2778 17711 2780 17720
rect 2832 17711 2834 17720
rect 2780 17682 2832 17688
rect 2778 16416 2834 16425
rect 2778 16351 2834 16360
rect 2792 16046 2820 16351
rect 2780 16040 2832 16046
rect 2780 15982 2832 15988
rect 3160 14550 3188 49030
rect 3792 48680 3844 48686
rect 3792 48622 3844 48628
rect 3330 48376 3386 48385
rect 3330 48311 3386 48320
rect 3344 47734 3372 48311
rect 3332 47728 3384 47734
rect 3332 47670 3384 47676
rect 3804 47666 3832 48622
rect 3884 48612 3936 48618
rect 3884 48554 3936 48560
rect 3516 47660 3568 47666
rect 3516 47602 3568 47608
rect 3792 47660 3844 47666
rect 3792 47602 3844 47608
rect 3528 44742 3556 47602
rect 3896 47190 3924 48554
rect 3988 47258 4016 49234
rect 4080 49065 4108 49234
rect 4066 49056 4122 49065
rect 4066 48991 4122 49000
rect 4068 48680 4120 48686
rect 4068 48622 4120 48628
rect 3976 47252 4028 47258
rect 3976 47194 4028 47200
rect 3608 47184 3660 47190
rect 3608 47126 3660 47132
rect 3884 47184 3936 47190
rect 3884 47126 3936 47132
rect 3620 46578 3648 47126
rect 3608 46572 3660 46578
rect 3608 46514 3660 46520
rect 3516 44736 3568 44742
rect 3516 44678 3568 44684
rect 3422 38176 3478 38185
rect 3422 38111 3478 38120
rect 3332 29096 3384 29102
rect 3332 29038 3384 29044
rect 3148 14544 3200 14550
rect 3148 14486 3200 14492
rect 2872 13728 2924 13734
rect 2778 13696 2834 13705
rect 2872 13670 2924 13676
rect 2778 13631 2834 13640
rect 2792 13394 2820 13631
rect 2884 13462 2912 13670
rect 2872 13456 2924 13462
rect 2872 13398 2924 13404
rect 2780 13388 2832 13394
rect 2780 13330 2832 13336
rect 2964 10464 3016 10470
rect 2964 10406 3016 10412
rect 2778 10296 2834 10305
rect 2778 10231 2834 10240
rect 2792 10130 2820 10231
rect 2780 10124 2832 10130
rect 2780 10066 2832 10072
rect 2976 9654 3004 10406
rect 2964 9648 3016 9654
rect 2778 9616 2834 9625
rect 2964 9590 3016 9596
rect 2778 9551 2834 9560
rect 2792 9518 2820 9551
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 2778 6896 2834 6905
rect 2778 6831 2780 6840
rect 2832 6831 2834 6840
rect 2780 6802 2832 6808
rect 2964 5704 3016 5710
rect 2964 5646 3016 5652
rect 2778 5536 2834 5545
rect 2778 5471 2834 5480
rect 2792 5166 2820 5471
rect 2976 5370 3004 5646
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 2778 4856 2834 4865
rect 2778 4791 2834 4800
rect 2504 4752 2556 4758
rect 2504 4694 2556 4700
rect 2792 4690 2820 4791
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 2596 4004 2648 4010
rect 2596 3946 2648 3952
rect 2136 3188 2188 3194
rect 2136 3130 2188 3136
rect 2412 3188 2464 3194
rect 2412 3130 2464 3136
rect 1952 3052 2004 3058
rect 1952 2994 2004 3000
rect 1952 2440 2004 2446
rect 1952 2382 2004 2388
rect 2226 2408 2282 2417
rect 1860 2372 1912 2378
rect 1860 2314 1912 2320
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 1872 785 1900 2314
rect 1964 800 1992 2382
rect 2226 2343 2228 2352
rect 2280 2343 2282 2352
rect 2228 2314 2280 2320
rect 2608 800 2636 3946
rect 3240 3664 3292 3670
rect 3240 3606 3292 3612
rect 3148 2644 3200 2650
rect 3148 2586 3200 2592
rect 3160 2145 3188 2586
rect 3146 2136 3202 2145
rect 3146 2071 3202 2080
rect 3252 800 3280 3606
rect 3344 3398 3372 29038
rect 3436 21418 3464 38111
rect 3528 28082 3556 44678
rect 4080 30122 4108 48622
rect 4214 48444 4522 48464
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48368 4522 48388
rect 4436 48068 4488 48074
rect 4436 48010 4488 48016
rect 4448 47530 4476 48010
rect 4632 47666 4660 51326
rect 5170 51200 5226 52000
rect 5814 51200 5870 52000
rect 6458 51200 6514 52000
rect 7102 51200 7158 52000
rect 7746 51354 7802 52000
rect 8390 51354 8446 52000
rect 7746 51326 8248 51354
rect 7746 51200 7802 51326
rect 4710 50416 4766 50425
rect 4710 50351 4766 50360
rect 4724 48686 4752 50351
rect 4712 48680 4764 48686
rect 4712 48622 4764 48628
rect 5184 48210 5212 51200
rect 6472 49230 6500 51200
rect 6460 49224 6512 49230
rect 6460 49166 6512 49172
rect 5448 49156 5500 49162
rect 5448 49098 5500 49104
rect 6644 49156 6696 49162
rect 6644 49098 6696 49104
rect 5172 48204 5224 48210
rect 5172 48146 5224 48152
rect 5356 48136 5408 48142
rect 5356 48078 5408 48084
rect 4712 48000 4764 48006
rect 4712 47942 4764 47948
rect 4620 47660 4672 47666
rect 4620 47602 4672 47608
rect 4436 47524 4488 47530
rect 4436 47466 4488 47472
rect 4214 47356 4522 47376
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47280 4522 47300
rect 4724 46578 4752 47942
rect 4804 47456 4856 47462
rect 4804 47398 4856 47404
rect 4712 46572 4764 46578
rect 4712 46514 4764 46520
rect 4214 46268 4522 46288
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46192 4522 46212
rect 4214 45180 4522 45200
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45104 4522 45124
rect 4214 44092 4522 44112
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44016 4522 44036
rect 4214 43004 4522 43024
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42928 4522 42948
rect 4214 41916 4522 41936
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41840 4522 41860
rect 4214 40828 4522 40848
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40752 4522 40772
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4816 31482 4844 47398
rect 4896 47048 4948 47054
rect 4896 46990 4948 46996
rect 4908 46442 4936 46990
rect 4896 46436 4948 46442
rect 4896 46378 4948 46384
rect 4908 35894 4936 46378
rect 4908 35866 5028 35894
rect 4804 31476 4856 31482
rect 4804 31418 4856 31424
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4804 30252 4856 30258
rect 4804 30194 4856 30200
rect 4068 30116 4120 30122
rect 4068 30058 4120 30064
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4066 29336 4122 29345
rect 4066 29271 4122 29280
rect 4080 29170 4108 29271
rect 4068 29164 4120 29170
rect 4068 29106 4120 29112
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 3516 28076 3568 28082
rect 3516 28018 3568 28024
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 4816 22234 4844 30194
rect 4804 22228 4856 22234
rect 4804 22170 4856 22176
rect 3974 21856 4030 21865
rect 3974 21791 4030 21800
rect 3424 21412 3476 21418
rect 3424 21354 3476 21360
rect 3988 20874 4016 21791
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4066 21176 4122 21185
rect 4214 21168 4522 21188
rect 4066 21111 4122 21120
rect 3976 20868 4028 20874
rect 3976 20810 4028 20816
rect 4080 20806 4108 21111
rect 4068 20800 4120 20806
rect 4068 20742 4120 20748
rect 4896 20256 4948 20262
rect 4896 20198 4948 20204
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 4908 19922 4936 20198
rect 4896 19916 4948 19922
rect 4896 19858 4948 19864
rect 4066 19816 4122 19825
rect 4066 19751 4122 19760
rect 4080 19446 4108 19751
rect 4068 19440 4120 19446
rect 4068 19382 4120 19388
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 5000 18766 5028 35866
rect 5368 35222 5396 48078
rect 5460 47802 5488 49098
rect 6656 48754 6684 49098
rect 6920 49088 6972 49094
rect 6920 49030 6972 49036
rect 6644 48748 6696 48754
rect 6644 48690 6696 48696
rect 5540 48068 5592 48074
rect 5540 48010 5592 48016
rect 5448 47796 5500 47802
rect 5448 47738 5500 47744
rect 5448 47524 5500 47530
rect 5448 47466 5500 47472
rect 5460 42362 5488 47466
rect 5552 47258 5580 48010
rect 5540 47252 5592 47258
rect 5540 47194 5592 47200
rect 5448 42356 5500 42362
rect 5448 42298 5500 42304
rect 5540 39840 5592 39846
rect 5540 39782 5592 39788
rect 6092 39840 6144 39846
rect 6092 39782 6144 39788
rect 5552 39438 5580 39782
rect 5540 39432 5592 39438
rect 5540 39374 5592 39380
rect 5356 35216 5408 35222
rect 5356 35158 5408 35164
rect 5540 20800 5592 20806
rect 5540 20742 5592 20748
rect 5552 19922 5580 20742
rect 5540 19916 5592 19922
rect 5540 19858 5592 19864
rect 4988 18760 5040 18766
rect 4988 18702 5040 18708
rect 3976 18692 4028 18698
rect 3976 18634 4028 18640
rect 3700 17128 3752 17134
rect 3700 17070 3752 17076
rect 3424 9648 3476 9654
rect 3424 9590 3476 9596
rect 3436 8945 3464 9590
rect 3422 8936 3478 8945
rect 3422 8871 3478 8880
rect 3422 6216 3478 6225
rect 3422 6151 3478 6160
rect 3436 5914 3464 6151
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 3424 5364 3476 5370
rect 3424 5306 3476 5312
rect 3436 4185 3464 5306
rect 3422 4176 3478 4185
rect 3422 4111 3478 4120
rect 3332 3392 3384 3398
rect 3332 3334 3384 3340
rect 3712 2582 3740 17070
rect 3988 12850 4016 18634
rect 4066 18456 4122 18465
rect 4066 18391 4122 18400
rect 4080 18086 4108 18391
rect 4068 18080 4120 18086
rect 4068 18022 4120 18028
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 4068 13796 4120 13802
rect 4068 13738 4120 13744
rect 4080 13025 4108 13738
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4066 13016 4122 13025
rect 4066 12951 4122 12960
rect 3976 12844 4028 12850
rect 3976 12786 4028 12792
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 4804 5636 4856 5642
rect 4804 5578 4856 5584
rect 3884 5568 3936 5574
rect 3884 5510 3936 5516
rect 3896 5302 3924 5510
rect 3884 5296 3936 5302
rect 3884 5238 3936 5244
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 3804 3602 3832 3878
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3792 3596 3844 3602
rect 3792 3538 3844 3544
rect 3700 2576 3752 2582
rect 3700 2518 3752 2524
rect 3896 800 3924 3674
rect 3988 3602 4016 3878
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 3976 3596 4028 3602
rect 3976 3538 4028 3544
rect 4632 2990 4660 4558
rect 4816 4146 4844 5578
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 4908 3126 4936 3878
rect 6104 3534 6132 39782
rect 6736 25696 6788 25702
rect 6736 25638 6788 25644
rect 6748 25362 6776 25638
rect 6736 25356 6788 25362
rect 6736 25298 6788 25304
rect 6932 22982 6960 49030
rect 7116 48618 7144 51200
rect 7748 48680 7800 48686
rect 7748 48622 7800 48628
rect 7104 48612 7156 48618
rect 7104 48554 7156 48560
rect 7760 48278 7788 48622
rect 7748 48272 7800 48278
rect 7748 48214 7800 48220
rect 8220 48226 8248 51326
rect 8390 51326 8892 51354
rect 8390 51200 8446 51326
rect 8668 49292 8720 49298
rect 8668 49234 8720 49240
rect 8220 48198 8432 48226
rect 7104 48136 7156 48142
rect 7104 48078 7156 48084
rect 7116 25906 7144 48078
rect 7380 48000 7432 48006
rect 7380 47942 7432 47948
rect 7392 47666 7420 47942
rect 7472 47796 7524 47802
rect 7472 47738 7524 47744
rect 7380 47660 7432 47666
rect 7380 47602 7432 47608
rect 7484 47598 7512 47738
rect 7472 47592 7524 47598
rect 7472 47534 7524 47540
rect 7932 46368 7984 46374
rect 7932 46310 7984 46316
rect 7944 45490 7972 46310
rect 7932 45484 7984 45490
rect 7932 45426 7984 45432
rect 8404 45422 8432 48198
rect 8680 47802 8708 49234
rect 8668 47796 8720 47802
rect 8668 47738 8720 47744
rect 8116 45416 8168 45422
rect 8116 45358 8168 45364
rect 8392 45416 8444 45422
rect 8392 45358 8444 45364
rect 8128 45082 8156 45358
rect 8116 45076 8168 45082
rect 8116 45018 8168 45024
rect 8864 31754 8892 51326
rect 9034 51200 9090 52000
rect 9678 51200 9734 52000
rect 10322 51200 10378 52000
rect 10966 51354 11022 52000
rect 10428 51326 11022 51354
rect 9220 49768 9272 49774
rect 9220 49710 9272 49716
rect 8944 49088 8996 49094
rect 8944 49030 8996 49036
rect 8956 48754 8984 49030
rect 8944 48748 8996 48754
rect 8944 48690 8996 48696
rect 9128 48680 9180 48686
rect 9128 48622 9180 48628
rect 9140 48346 9168 48622
rect 9128 48340 9180 48346
rect 9128 48282 9180 48288
rect 8944 48136 8996 48142
rect 8944 48078 8996 48084
rect 9128 48136 9180 48142
rect 9128 48078 9180 48084
rect 8956 47666 8984 48078
rect 8944 47660 8996 47666
rect 8944 47602 8996 47608
rect 9036 47592 9088 47598
rect 9036 47534 9088 47540
rect 9048 47258 9076 47534
rect 9036 47252 9088 47258
rect 9036 47194 9088 47200
rect 9140 47122 9168 48078
rect 9232 47598 9260 49710
rect 9692 48686 9720 51200
rect 9864 49224 9916 49230
rect 9864 49166 9916 49172
rect 9680 48680 9732 48686
rect 9680 48622 9732 48628
rect 9876 48210 9904 49166
rect 10336 48210 10364 51200
rect 9864 48204 9916 48210
rect 9864 48146 9916 48152
rect 10324 48204 10376 48210
rect 10324 48146 10376 48152
rect 9956 48068 10008 48074
rect 9956 48010 10008 48016
rect 9968 47802 9996 48010
rect 9956 47796 10008 47802
rect 9956 47738 10008 47744
rect 9220 47592 9272 47598
rect 9220 47534 9272 47540
rect 9128 47116 9180 47122
rect 9128 47058 9180 47064
rect 9140 45554 9168 47058
rect 9404 47048 9456 47054
rect 9404 46990 9456 46996
rect 9048 45526 9168 45554
rect 8944 44872 8996 44878
rect 8944 44814 8996 44820
rect 8956 43926 8984 44814
rect 8944 43920 8996 43926
rect 8944 43862 8996 43868
rect 9048 32978 9076 45526
rect 9036 32972 9088 32978
rect 9036 32914 9088 32920
rect 8864 31726 9076 31754
rect 8484 31272 8536 31278
rect 8484 31214 8536 31220
rect 8496 30190 8524 31214
rect 7748 30184 7800 30190
rect 7748 30126 7800 30132
rect 8484 30184 8536 30190
rect 8484 30126 8536 30132
rect 7760 29102 7788 30126
rect 8944 29504 8996 29510
rect 8944 29446 8996 29452
rect 8956 29238 8984 29446
rect 8944 29232 8996 29238
rect 8944 29174 8996 29180
rect 7748 29096 7800 29102
rect 7748 29038 7800 29044
rect 7288 27872 7340 27878
rect 7288 27814 7340 27820
rect 7300 27402 7328 27814
rect 7760 27470 7788 29038
rect 8852 29028 8904 29034
rect 8852 28970 8904 28976
rect 8300 28756 8352 28762
rect 8300 28698 8352 28704
rect 8312 28218 8340 28698
rect 8864 28694 8892 28970
rect 8852 28688 8904 28694
rect 8852 28630 8904 28636
rect 8300 28212 8352 28218
rect 8352 28172 8432 28200
rect 8300 28154 8352 28160
rect 8300 28076 8352 28082
rect 8300 28018 8352 28024
rect 7748 27464 7800 27470
rect 7748 27406 7800 27412
rect 7288 27396 7340 27402
rect 7288 27338 7340 27344
rect 7760 26382 7788 27406
rect 8312 26858 8340 28018
rect 8404 27062 8432 28172
rect 8760 27872 8812 27878
rect 8760 27814 8812 27820
rect 8772 27130 8800 27814
rect 9048 27538 9076 31726
rect 9128 29640 9180 29646
rect 9128 29582 9180 29588
rect 9140 28762 9168 29582
rect 9128 28756 9180 28762
rect 9128 28698 9180 28704
rect 9312 28008 9364 28014
rect 9312 27950 9364 27956
rect 9036 27532 9088 27538
rect 9036 27474 9088 27480
rect 9324 27334 9352 27950
rect 9312 27328 9364 27334
rect 9312 27270 9364 27276
rect 8760 27124 8812 27130
rect 8760 27066 8812 27072
rect 8392 27056 8444 27062
rect 8392 26998 8444 27004
rect 8300 26852 8352 26858
rect 8300 26794 8352 26800
rect 7748 26376 7800 26382
rect 7748 26318 7800 26324
rect 7104 25900 7156 25906
rect 7104 25842 7156 25848
rect 7116 25498 7144 25842
rect 7104 25492 7156 25498
rect 7104 25434 7156 25440
rect 7760 24818 7788 26318
rect 9220 26308 9272 26314
rect 9220 26250 9272 26256
rect 9232 26042 9260 26250
rect 9220 26036 9272 26042
rect 9220 25978 9272 25984
rect 8116 25356 8168 25362
rect 8116 25298 8168 25304
rect 7748 24812 7800 24818
rect 7748 24754 7800 24760
rect 6920 22976 6972 22982
rect 6920 22918 6972 22924
rect 7840 22092 7892 22098
rect 7840 22034 7892 22040
rect 7852 21978 7880 22034
rect 7116 21950 7880 21978
rect 8024 22024 8076 22030
rect 8024 21966 8076 21972
rect 7116 21622 7144 21950
rect 7196 21888 7248 21894
rect 7196 21830 7248 21836
rect 7288 21888 7340 21894
rect 7288 21830 7340 21836
rect 7208 21622 7236 21830
rect 7104 21616 7156 21622
rect 7104 21558 7156 21564
rect 7196 21616 7248 21622
rect 7196 21558 7248 21564
rect 7300 21554 7328 21830
rect 7288 21548 7340 21554
rect 7288 21490 7340 21496
rect 7472 21480 7524 21486
rect 7472 21422 7524 21428
rect 7484 21146 7512 21422
rect 7472 21140 7524 21146
rect 7472 21082 7524 21088
rect 6828 20936 6880 20942
rect 6828 20878 6880 20884
rect 6840 18290 6868 20878
rect 7932 20596 7984 20602
rect 7932 20538 7984 20544
rect 6828 18284 6880 18290
rect 6828 18226 6880 18232
rect 7472 18284 7524 18290
rect 7472 18226 7524 18232
rect 6828 18080 6880 18086
rect 6828 18022 6880 18028
rect 6920 18080 6972 18086
rect 6920 18022 6972 18028
rect 6840 17746 6868 18022
rect 6828 17740 6880 17746
rect 6828 17682 6880 17688
rect 6932 17610 6960 18022
rect 7484 17814 7512 18226
rect 7472 17808 7524 17814
rect 7472 17750 7524 17756
rect 6920 17604 6972 17610
rect 6920 17546 6972 17552
rect 7944 15094 7972 20538
rect 8036 19922 8064 21966
rect 8024 19916 8076 19922
rect 8024 19858 8076 19864
rect 8036 19378 8064 19858
rect 8024 19372 8076 19378
rect 8024 19314 8076 19320
rect 8036 18358 8064 19314
rect 8024 18352 8076 18358
rect 8024 18294 8076 18300
rect 8128 17218 8156 25298
rect 8944 25152 8996 25158
rect 8944 25094 8996 25100
rect 8956 24818 8984 25094
rect 8944 24812 8996 24818
rect 8944 24754 8996 24760
rect 9128 24608 9180 24614
rect 9128 24550 9180 24556
rect 8852 24200 8904 24206
rect 8852 24142 8904 24148
rect 8864 23866 8892 24142
rect 9140 24138 9168 24550
rect 9324 24342 9352 27270
rect 9416 24954 9444 46990
rect 10428 45554 10456 51326
rect 10966 51200 11022 51326
rect 11610 51200 11666 52000
rect 12254 51354 12310 52000
rect 12898 51354 12954 52000
rect 12254 51326 12388 51354
rect 12254 51200 12310 51326
rect 11624 49230 11652 51200
rect 11612 49224 11664 49230
rect 11612 49166 11664 49172
rect 12164 49156 12216 49162
rect 12164 49098 12216 49104
rect 11520 48680 11572 48686
rect 11520 48622 11572 48628
rect 11704 48680 11756 48686
rect 11704 48622 11756 48628
rect 11532 47666 11560 48622
rect 11716 48346 11744 48622
rect 11704 48340 11756 48346
rect 11704 48282 11756 48288
rect 11980 48136 12032 48142
rect 11980 48078 12032 48084
rect 11520 47660 11572 47666
rect 11520 47602 11572 47608
rect 11992 47598 12020 48078
rect 11980 47592 12032 47598
rect 11980 47534 12032 47540
rect 9876 45526 10456 45554
rect 9876 33862 9904 45526
rect 11992 35894 12020 47534
rect 12176 35894 12204 49098
rect 12360 48668 12388 51326
rect 12728 51326 12954 51354
rect 12728 49298 12756 51326
rect 12898 51200 12954 51326
rect 13542 51354 13598 52000
rect 14186 51354 14242 52000
rect 13542 51326 13768 51354
rect 13542 51200 13598 51326
rect 13740 49314 13768 51326
rect 14016 51326 14242 51354
rect 13740 49298 13860 49314
rect 12716 49292 12768 49298
rect 13740 49292 13872 49298
rect 13740 49286 13820 49292
rect 12716 49234 12768 49240
rect 13820 49234 13872 49240
rect 12992 49224 13044 49230
rect 12992 49166 13044 49172
rect 12440 48680 12492 48686
rect 12360 48640 12440 48668
rect 12440 48622 12492 48628
rect 11992 35866 12112 35894
rect 12176 35866 12388 35894
rect 11704 35692 11756 35698
rect 11704 35634 11756 35640
rect 11716 35154 11744 35634
rect 11704 35148 11756 35154
rect 11704 35090 11756 35096
rect 11888 33924 11940 33930
rect 11888 33866 11940 33872
rect 9864 33856 9916 33862
rect 9864 33798 9916 33804
rect 11900 33658 11928 33866
rect 11888 33652 11940 33658
rect 11888 33594 11940 33600
rect 11704 33516 11756 33522
rect 11704 33458 11756 33464
rect 11716 33318 11744 33458
rect 11704 33312 11756 33318
rect 11704 33254 11756 33260
rect 11520 31680 11572 31686
rect 11520 31622 11572 31628
rect 11532 31414 11560 31622
rect 11520 31408 11572 31414
rect 11520 31350 11572 31356
rect 10324 31340 10376 31346
rect 10324 31282 10376 31288
rect 10140 31136 10192 31142
rect 10140 31078 10192 31084
rect 9680 30660 9732 30666
rect 9680 30602 9732 30608
rect 10048 30660 10100 30666
rect 10152 30648 10180 31078
rect 10336 30938 10364 31282
rect 10324 30932 10376 30938
rect 10324 30874 10376 30880
rect 10416 30728 10468 30734
rect 10416 30670 10468 30676
rect 10784 30728 10836 30734
rect 11152 30728 11204 30734
rect 10784 30670 10836 30676
rect 10980 30676 11152 30682
rect 10980 30670 11204 30676
rect 10100 30620 10180 30648
rect 10048 30602 10100 30608
rect 9692 30326 9720 30602
rect 9680 30320 9732 30326
rect 9680 30262 9732 30268
rect 9864 29232 9916 29238
rect 9864 29174 9916 29180
rect 9680 29096 9732 29102
rect 9680 29038 9732 29044
rect 9692 27962 9720 29038
rect 9772 28960 9824 28966
rect 9772 28902 9824 28908
rect 9784 28626 9812 28902
rect 9772 28620 9824 28626
rect 9772 28562 9824 28568
rect 9784 28082 9812 28562
rect 9876 28082 9904 29174
rect 9956 28416 10008 28422
rect 9956 28358 10008 28364
rect 9772 28076 9824 28082
rect 9772 28018 9824 28024
rect 9864 28076 9916 28082
rect 9864 28018 9916 28024
rect 9692 27934 9812 27962
rect 9680 27872 9732 27878
rect 9680 27814 9732 27820
rect 9692 26926 9720 27814
rect 9680 26920 9732 26926
rect 9680 26862 9732 26868
rect 9680 26784 9732 26790
rect 9680 26726 9732 26732
rect 9692 25906 9720 26726
rect 9680 25900 9732 25906
rect 9680 25842 9732 25848
rect 9404 24948 9456 24954
rect 9404 24890 9456 24896
rect 9312 24336 9364 24342
rect 9312 24278 9364 24284
rect 9128 24132 9180 24138
rect 9128 24074 9180 24080
rect 8852 23860 8904 23866
rect 8852 23802 8904 23808
rect 9220 23724 9272 23730
rect 9324 23712 9352 24278
rect 9404 24064 9456 24070
rect 9404 24006 9456 24012
rect 9416 23730 9444 24006
rect 9272 23684 9352 23712
rect 9220 23666 9272 23672
rect 9324 23526 9352 23684
rect 9404 23724 9456 23730
rect 9404 23666 9456 23672
rect 9312 23520 9364 23526
rect 9312 23462 9364 23468
rect 9416 22094 9444 23666
rect 9496 22636 9548 22642
rect 9496 22578 9548 22584
rect 9508 22166 9536 22578
rect 9784 22438 9812 27934
rect 9876 27674 9904 28018
rect 9864 27668 9916 27674
rect 9864 27610 9916 27616
rect 9876 26994 9904 27610
rect 9968 27470 9996 28358
rect 9956 27464 10008 27470
rect 9956 27406 10008 27412
rect 9864 26988 9916 26994
rect 9864 26930 9916 26936
rect 9956 22568 10008 22574
rect 9956 22510 10008 22516
rect 9772 22432 9824 22438
rect 9772 22374 9824 22380
rect 9496 22160 9548 22166
rect 9496 22102 9548 22108
rect 9324 22066 9444 22094
rect 8760 20392 8812 20398
rect 8760 20334 8812 20340
rect 8944 20392 8996 20398
rect 8944 20334 8996 20340
rect 8772 19514 8800 20334
rect 8956 20058 8984 20334
rect 8944 20052 8996 20058
rect 8944 19994 8996 20000
rect 9220 19712 9272 19718
rect 9220 19654 9272 19660
rect 8760 19508 8812 19514
rect 8760 19450 8812 19456
rect 9232 19446 9260 19654
rect 9220 19440 9272 19446
rect 9220 19382 9272 19388
rect 9324 18766 9352 22066
rect 9404 19848 9456 19854
rect 9508 19836 9536 22102
rect 9968 22030 9996 22510
rect 9956 22024 10008 22030
rect 9956 21966 10008 21972
rect 9956 21888 10008 21894
rect 9956 21830 10008 21836
rect 9968 21554 9996 21830
rect 9956 21548 10008 21554
rect 9956 21490 10008 21496
rect 9456 19808 9536 19836
rect 9588 19848 9640 19854
rect 9404 19790 9456 19796
rect 9588 19790 9640 19796
rect 9680 19848 9732 19854
rect 9680 19790 9732 19796
rect 9600 18834 9628 19790
rect 9692 19514 9720 19790
rect 9680 19508 9732 19514
rect 9680 19450 9732 19456
rect 9772 19372 9824 19378
rect 9772 19314 9824 19320
rect 9784 19258 9812 19314
rect 9784 19230 9996 19258
rect 9588 18828 9640 18834
rect 9588 18770 9640 18776
rect 9312 18760 9364 18766
rect 9312 18702 9364 18708
rect 9496 18760 9548 18766
rect 9496 18702 9548 18708
rect 9036 18624 9088 18630
rect 9036 18566 9088 18572
rect 9048 18290 9076 18566
rect 9508 18426 9536 18702
rect 9496 18420 9548 18426
rect 9496 18362 9548 18368
rect 9036 18284 9088 18290
rect 9036 18226 9088 18232
rect 9600 18154 9628 18770
rect 9864 18284 9916 18290
rect 9864 18226 9916 18232
rect 9588 18148 9640 18154
rect 9588 18090 9640 18096
rect 8208 18080 8260 18086
rect 8208 18022 8260 18028
rect 9404 18080 9456 18086
rect 9404 18022 9456 18028
rect 8036 17190 8156 17218
rect 7932 15088 7984 15094
rect 7932 15030 7984 15036
rect 7944 13326 7972 15030
rect 7932 13320 7984 13326
rect 7932 13262 7984 13268
rect 8036 4010 8064 17190
rect 8220 17082 8248 18022
rect 9416 17610 9444 18022
rect 9404 17604 9456 17610
rect 9404 17546 9456 17552
rect 9588 17536 9640 17542
rect 9588 17478 9640 17484
rect 9600 17202 9628 17478
rect 9876 17270 9904 18226
rect 9968 17882 9996 19230
rect 9956 17876 10008 17882
rect 9956 17818 10008 17824
rect 9864 17264 9916 17270
rect 9864 17206 9916 17212
rect 9588 17196 9640 17202
rect 9588 17138 9640 17144
rect 8128 17054 8248 17082
rect 8128 13938 8156 17054
rect 9600 15570 9628 17138
rect 9680 16108 9732 16114
rect 9680 16050 9732 16056
rect 9588 15564 9640 15570
rect 9588 15506 9640 15512
rect 9404 15428 9456 15434
rect 9404 15370 9456 15376
rect 9416 15162 9444 15370
rect 9404 15156 9456 15162
rect 9404 15098 9456 15104
rect 9692 15026 9720 16050
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 9692 14482 9720 14962
rect 9680 14476 9732 14482
rect 9680 14418 9732 14424
rect 8116 13932 8168 13938
rect 8116 13874 8168 13880
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 8312 13530 8340 13806
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 8116 13320 8168 13326
rect 8116 13262 8168 13268
rect 8128 4078 8156 13262
rect 10060 12434 10088 30602
rect 10232 30252 10284 30258
rect 10232 30194 10284 30200
rect 10244 29850 10272 30194
rect 10232 29844 10284 29850
rect 10232 29786 10284 29792
rect 10428 29510 10456 30670
rect 10796 30258 10824 30670
rect 10980 30654 11192 30670
rect 10876 30592 10928 30598
rect 10876 30534 10928 30540
rect 10600 30252 10652 30258
rect 10600 30194 10652 30200
rect 10784 30252 10836 30258
rect 10784 30194 10836 30200
rect 10612 30054 10640 30194
rect 10600 30048 10652 30054
rect 10600 29990 10652 29996
rect 10692 30048 10744 30054
rect 10692 29990 10744 29996
rect 10508 29844 10560 29850
rect 10508 29786 10560 29792
rect 10520 29646 10548 29786
rect 10508 29640 10560 29646
rect 10508 29582 10560 29588
rect 10232 29504 10284 29510
rect 10232 29446 10284 29452
rect 10416 29504 10468 29510
rect 10416 29446 10468 29452
rect 10244 29306 10272 29446
rect 10232 29300 10284 29306
rect 10232 29242 10284 29248
rect 10244 28558 10272 29242
rect 10520 28966 10548 29582
rect 10508 28960 10560 28966
rect 10508 28902 10560 28908
rect 10232 28552 10284 28558
rect 10232 28494 10284 28500
rect 10140 26920 10192 26926
rect 10140 26862 10192 26868
rect 10152 26518 10180 26862
rect 10140 26512 10192 26518
rect 10140 26454 10192 26460
rect 10244 25378 10272 28494
rect 10612 28200 10640 29990
rect 10704 29646 10732 29990
rect 10796 29714 10824 30194
rect 10784 29708 10836 29714
rect 10784 29650 10836 29656
rect 10888 29646 10916 30534
rect 10692 29640 10744 29646
rect 10692 29582 10744 29588
rect 10876 29640 10928 29646
rect 10876 29582 10928 29588
rect 10980 28490 11008 30654
rect 11532 29170 11560 31350
rect 11716 29578 11744 33254
rect 11888 31340 11940 31346
rect 11888 31282 11940 31288
rect 11900 30938 11928 31282
rect 11888 30932 11940 30938
rect 11888 30874 11940 30880
rect 11704 29572 11756 29578
rect 11704 29514 11756 29520
rect 11520 29164 11572 29170
rect 11520 29106 11572 29112
rect 11612 29164 11664 29170
rect 11612 29106 11664 29112
rect 11624 28762 11652 29106
rect 11612 28756 11664 28762
rect 11612 28698 11664 28704
rect 11520 28552 11572 28558
rect 11520 28494 11572 28500
rect 10968 28484 11020 28490
rect 10968 28426 11020 28432
rect 10612 28172 10824 28200
rect 10416 27396 10468 27402
rect 10416 27338 10468 27344
rect 10324 27056 10376 27062
rect 10324 26998 10376 27004
rect 10336 26042 10364 26998
rect 10428 26994 10456 27338
rect 10692 27328 10744 27334
rect 10692 27270 10744 27276
rect 10416 26988 10468 26994
rect 10416 26930 10468 26936
rect 10704 26858 10732 27270
rect 10692 26852 10744 26858
rect 10692 26794 10744 26800
rect 10796 26738 10824 28172
rect 10980 27606 11008 28426
rect 11532 28218 11560 28494
rect 11980 28416 12032 28422
rect 11980 28358 12032 28364
rect 11520 28212 11572 28218
rect 11520 28154 11572 28160
rect 11888 28144 11940 28150
rect 11888 28086 11940 28092
rect 10968 27600 11020 27606
rect 10968 27542 11020 27548
rect 10876 27464 10928 27470
rect 10876 27406 10928 27412
rect 10704 26710 10824 26738
rect 10324 26036 10376 26042
rect 10324 25978 10376 25984
rect 10324 25696 10376 25702
rect 10324 25638 10376 25644
rect 10508 25696 10560 25702
rect 10508 25638 10560 25644
rect 10336 25498 10364 25638
rect 10324 25492 10376 25498
rect 10324 25434 10376 25440
rect 10244 25350 10364 25378
rect 10336 24614 10364 25350
rect 10520 25294 10548 25638
rect 10508 25288 10560 25294
rect 10508 25230 10560 25236
rect 10600 24744 10652 24750
rect 10600 24686 10652 24692
rect 10232 24608 10284 24614
rect 10232 24550 10284 24556
rect 10324 24608 10376 24614
rect 10324 24550 10376 24556
rect 10244 24274 10272 24550
rect 10232 24268 10284 24274
rect 10232 24210 10284 24216
rect 10508 24268 10560 24274
rect 10508 24210 10560 24216
rect 10140 24200 10192 24206
rect 10140 24142 10192 24148
rect 10324 24200 10376 24206
rect 10324 24142 10376 24148
rect 10152 23526 10180 24142
rect 10336 23610 10364 24142
rect 10416 23724 10468 23730
rect 10416 23666 10468 23672
rect 10244 23582 10364 23610
rect 10140 23520 10192 23526
rect 10140 23462 10192 23468
rect 10140 21956 10192 21962
rect 10140 21898 10192 21904
rect 10152 18358 10180 21898
rect 10244 21554 10272 23582
rect 10428 23526 10456 23666
rect 10520 23662 10548 24210
rect 10612 23730 10640 24686
rect 10600 23724 10652 23730
rect 10600 23666 10652 23672
rect 10508 23656 10560 23662
rect 10508 23598 10560 23604
rect 10324 23520 10376 23526
rect 10324 23462 10376 23468
rect 10416 23520 10468 23526
rect 10416 23462 10468 23468
rect 10336 23186 10364 23462
rect 10324 23180 10376 23186
rect 10324 23122 10376 23128
rect 10428 22574 10456 23462
rect 10612 22778 10640 23666
rect 10600 22772 10652 22778
rect 10600 22714 10652 22720
rect 10416 22568 10468 22574
rect 10416 22510 10468 22516
rect 10416 22432 10468 22438
rect 10416 22374 10468 22380
rect 10232 21548 10284 21554
rect 10232 21490 10284 21496
rect 10428 20398 10456 22374
rect 10508 20460 10560 20466
rect 10508 20402 10560 20408
rect 10416 20392 10468 20398
rect 10416 20334 10468 20340
rect 10232 19848 10284 19854
rect 10232 19790 10284 19796
rect 10416 19848 10468 19854
rect 10520 19802 10548 20402
rect 10468 19796 10548 19802
rect 10416 19790 10548 19796
rect 10244 18766 10272 19790
rect 10428 19774 10548 19790
rect 10520 19378 10548 19774
rect 10508 19372 10560 19378
rect 10508 19314 10560 19320
rect 10232 18760 10284 18766
rect 10232 18702 10284 18708
rect 10140 18352 10192 18358
rect 10140 18294 10192 18300
rect 10244 18290 10272 18702
rect 10520 18290 10548 19314
rect 10232 18284 10284 18290
rect 10232 18226 10284 18232
rect 10508 18284 10560 18290
rect 10508 18226 10560 18232
rect 10140 16516 10192 16522
rect 10140 16458 10192 16464
rect 10152 16250 10180 16458
rect 10140 16244 10192 16250
rect 10140 16186 10192 16192
rect 10244 15366 10272 18226
rect 10520 17202 10548 18226
rect 10508 17196 10560 17202
rect 10508 17138 10560 17144
rect 10232 15360 10284 15366
rect 10232 15302 10284 15308
rect 10060 12406 10272 12434
rect 10244 6914 10272 12406
rect 10152 6886 10272 6914
rect 10152 4078 10180 6886
rect 8116 4072 8168 4078
rect 8116 4014 8168 4020
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 9404 4072 9456 4078
rect 9404 4014 9456 4020
rect 10140 4072 10192 4078
rect 10140 4014 10192 4020
rect 8024 4004 8076 4010
rect 8024 3946 8076 3952
rect 6460 3936 6512 3942
rect 6460 3878 6512 3884
rect 6092 3528 6144 3534
rect 6092 3470 6144 3476
rect 6368 3528 6420 3534
rect 6368 3470 6420 3476
rect 4896 3120 4948 3126
rect 4896 3062 4948 3068
rect 6380 3058 6408 3470
rect 6368 3052 6420 3058
rect 6368 2994 6420 3000
rect 4620 2984 4672 2990
rect 4620 2926 4672 2932
rect 5172 2984 5224 2990
rect 5172 2926 5224 2932
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 4804 2576 4856 2582
rect 4802 2544 4804 2553
rect 4856 2544 4858 2553
rect 4802 2479 4858 2488
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 4540 800 4568 2382
rect 5184 800 5212 2926
rect 5816 2576 5868 2582
rect 5816 2518 5868 2524
rect 5828 800 5856 2518
rect 6472 2514 6500 3878
rect 9324 3738 9352 4014
rect 9312 3732 9364 3738
rect 9312 3674 9364 3680
rect 8944 3460 8996 3466
rect 8944 3402 8996 3408
rect 6552 3392 6604 3398
rect 6552 3334 6604 3340
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 6564 3126 6592 3334
rect 6552 3120 6604 3126
rect 6552 3062 6604 3068
rect 6552 2984 6604 2990
rect 6552 2926 6604 2932
rect 6460 2508 6512 2514
rect 6460 2450 6512 2456
rect 6564 2394 6592 2926
rect 6932 2514 6960 3334
rect 8956 3058 8984 3402
rect 8944 3052 8996 3058
rect 8944 2994 8996 3000
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 7104 2508 7156 2514
rect 7104 2450 7156 2456
rect 6472 2366 6592 2394
rect 6472 800 6500 2366
rect 7116 800 7144 2450
rect 7760 800 7788 2926
rect 8392 2372 8444 2378
rect 8392 2314 8444 2320
rect 8404 800 8432 2314
rect 9048 870 9168 898
rect 9048 800 9076 870
rect 1858 776 1914 785
rect 1858 711 1914 720
rect 1950 0 2006 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9140 762 9168 870
rect 9416 762 9444 4014
rect 10704 4010 10732 26710
rect 10888 26518 10916 27406
rect 10980 27402 11008 27542
rect 10968 27396 11020 27402
rect 10968 27338 11020 27344
rect 11900 27130 11928 28086
rect 11992 27878 12020 28358
rect 11980 27872 12032 27878
rect 11980 27814 12032 27820
rect 11888 27124 11940 27130
rect 11888 27066 11940 27072
rect 11980 27056 12032 27062
rect 11980 26998 12032 27004
rect 11428 26580 11480 26586
rect 11428 26522 11480 26528
rect 10784 26512 10836 26518
rect 10784 26454 10836 26460
rect 10876 26512 10928 26518
rect 10876 26454 10928 26460
rect 10796 24818 10824 26454
rect 10888 25906 10916 26454
rect 10968 26240 11020 26246
rect 10968 26182 11020 26188
rect 10876 25900 10928 25906
rect 10876 25842 10928 25848
rect 10980 25294 11008 26182
rect 11440 25294 11468 26522
rect 11796 26308 11848 26314
rect 11796 26250 11848 26256
rect 11704 25764 11756 25770
rect 11704 25706 11756 25712
rect 10968 25288 11020 25294
rect 10968 25230 11020 25236
rect 11428 25288 11480 25294
rect 11428 25230 11480 25236
rect 10784 24812 10836 24818
rect 10784 24754 10836 24760
rect 10796 23730 10824 24754
rect 10980 24290 11008 25230
rect 11716 25158 11744 25706
rect 11808 25294 11836 26250
rect 11992 25974 12020 26998
rect 11980 25968 12032 25974
rect 11980 25910 12032 25916
rect 11992 25498 12020 25910
rect 11980 25492 12032 25498
rect 11980 25434 12032 25440
rect 11796 25288 11848 25294
rect 11796 25230 11848 25236
rect 11704 25152 11756 25158
rect 11704 25094 11756 25100
rect 11796 24676 11848 24682
rect 11796 24618 11848 24624
rect 11152 24336 11204 24342
rect 10980 24284 11152 24290
rect 10980 24278 11204 24284
rect 10980 24274 11192 24278
rect 11808 24274 11836 24618
rect 11888 24608 11940 24614
rect 11888 24550 11940 24556
rect 10968 24268 11192 24274
rect 11020 24262 11192 24268
rect 11244 24268 11296 24274
rect 10968 24210 11020 24216
rect 11244 24210 11296 24216
rect 11796 24268 11848 24274
rect 11796 24210 11848 24216
rect 10876 24200 10928 24206
rect 10876 24142 10928 24148
rect 10888 23730 10916 24142
rect 10968 24132 11020 24138
rect 11256 24120 11284 24210
rect 11428 24132 11480 24138
rect 11256 24092 11428 24120
rect 10968 24074 11020 24080
rect 11428 24074 11480 24080
rect 10784 23724 10836 23730
rect 10784 23666 10836 23672
rect 10876 23724 10928 23730
rect 10876 23666 10928 23672
rect 10796 23118 10824 23666
rect 10980 23662 11008 24074
rect 11704 24064 11756 24070
rect 11702 24032 11704 24041
rect 11756 24032 11758 24041
rect 11702 23967 11758 23976
rect 11704 23724 11756 23730
rect 11704 23666 11756 23672
rect 10968 23656 11020 23662
rect 10968 23598 11020 23604
rect 11716 23254 11744 23666
rect 11704 23248 11756 23254
rect 11704 23190 11756 23196
rect 10784 23112 10836 23118
rect 10784 23054 10836 23060
rect 10782 22672 10838 22681
rect 10782 22607 10784 22616
rect 10836 22607 10838 22616
rect 10784 22578 10836 22584
rect 10968 22568 11020 22574
rect 10968 22510 11020 22516
rect 10980 21962 11008 22510
rect 10968 21956 11020 21962
rect 10968 21898 11020 21904
rect 11612 21412 11664 21418
rect 11612 21354 11664 21360
rect 11624 21078 11652 21354
rect 11612 21072 11664 21078
rect 11612 21014 11664 21020
rect 11612 20868 11664 20874
rect 11612 20810 11664 20816
rect 11520 19780 11572 19786
rect 11520 19722 11572 19728
rect 10968 19712 11020 19718
rect 10968 19654 11020 19660
rect 10980 19417 11008 19654
rect 11532 19514 11560 19722
rect 11520 19508 11572 19514
rect 11520 19450 11572 19456
rect 10966 19408 11022 19417
rect 10966 19343 11022 19352
rect 11336 18624 11388 18630
rect 11336 18566 11388 18572
rect 11348 17610 11376 18566
rect 11336 17604 11388 17610
rect 11336 17546 11388 17552
rect 11520 17536 11572 17542
rect 11520 17478 11572 17484
rect 11532 15570 11560 17478
rect 11624 16590 11652 20810
rect 11704 20460 11756 20466
rect 11704 20402 11756 20408
rect 11716 20058 11744 20402
rect 11704 20052 11756 20058
rect 11704 19994 11756 20000
rect 11808 19378 11836 24210
rect 11900 24206 11928 24550
rect 11888 24200 11940 24206
rect 11888 24142 11940 24148
rect 11888 24064 11940 24070
rect 11888 24006 11940 24012
rect 11900 23186 11928 24006
rect 11888 23180 11940 23186
rect 11888 23122 11940 23128
rect 11980 20256 12032 20262
rect 11980 20198 12032 20204
rect 11992 19378 12020 20198
rect 11796 19372 11848 19378
rect 11796 19314 11848 19320
rect 11980 19372 12032 19378
rect 11980 19314 12032 19320
rect 11888 18760 11940 18766
rect 11888 18702 11940 18708
rect 11900 18426 11928 18702
rect 11888 18420 11940 18426
rect 11888 18362 11940 18368
rect 11704 18284 11756 18290
rect 11704 18226 11756 18232
rect 11716 17542 11744 18226
rect 11704 17536 11756 17542
rect 11704 17478 11756 17484
rect 12084 16726 12112 35866
rect 12164 32224 12216 32230
rect 12164 32166 12216 32172
rect 12176 31822 12204 32166
rect 12164 31816 12216 31822
rect 12164 31758 12216 31764
rect 12256 31748 12308 31754
rect 12256 31690 12308 31696
rect 12268 31414 12296 31690
rect 12256 31408 12308 31414
rect 12256 31350 12308 31356
rect 12164 30864 12216 30870
rect 12162 30832 12164 30841
rect 12216 30832 12218 30841
rect 12162 30767 12218 30776
rect 12268 30326 12296 31350
rect 12256 30320 12308 30326
rect 12256 30262 12308 30268
rect 12256 29572 12308 29578
rect 12256 29514 12308 29520
rect 12268 28558 12296 29514
rect 12256 28552 12308 28558
rect 12256 28494 12308 28500
rect 12268 28218 12296 28494
rect 12256 28212 12308 28218
rect 12256 28154 12308 28160
rect 12164 28008 12216 28014
rect 12164 27950 12216 27956
rect 12176 26382 12204 27950
rect 12164 26376 12216 26382
rect 12164 26318 12216 26324
rect 12256 26240 12308 26246
rect 12256 26182 12308 26188
rect 12268 26042 12296 26182
rect 12256 26036 12308 26042
rect 12256 25978 12308 25984
rect 12164 21480 12216 21486
rect 12164 21422 12216 21428
rect 12176 21146 12204 21422
rect 12256 21344 12308 21350
rect 12256 21286 12308 21292
rect 12268 21146 12296 21286
rect 12164 21140 12216 21146
rect 12164 21082 12216 21088
rect 12256 21140 12308 21146
rect 12256 21082 12308 21088
rect 12360 20942 12388 35866
rect 13004 34746 13032 49166
rect 14016 48754 14044 51326
rect 14186 51200 14242 51326
rect 14830 51354 14886 52000
rect 14830 51326 14964 51354
rect 14830 51200 14886 51326
rect 14372 49224 14424 49230
rect 14372 49166 14424 49172
rect 14384 48822 14412 49166
rect 14372 48816 14424 48822
rect 14372 48758 14424 48764
rect 14004 48748 14056 48754
rect 14004 48690 14056 48696
rect 14936 48210 14964 51326
rect 15474 51200 15530 52000
rect 16118 51200 16174 52000
rect 16762 51200 16818 52000
rect 17406 51200 17462 52000
rect 18050 51200 18106 52000
rect 18694 51200 18750 52000
rect 19338 51200 19394 52000
rect 19982 51200 20038 52000
rect 20626 51200 20682 52000
rect 21270 51200 21326 52000
rect 21914 51200 21970 52000
rect 22558 51200 22614 52000
rect 23202 51200 23258 52000
rect 23846 51200 23902 52000
rect 24490 51354 24546 52000
rect 24490 51326 24808 51354
rect 24490 51200 24546 51326
rect 14924 48204 14976 48210
rect 14924 48146 14976 48152
rect 14464 48136 14516 48142
rect 14464 48078 14516 48084
rect 14372 48068 14424 48074
rect 14372 48010 14424 48016
rect 14384 47258 14412 48010
rect 14476 47666 14504 48078
rect 14464 47660 14516 47666
rect 14464 47602 14516 47608
rect 14372 47252 14424 47258
rect 14372 47194 14424 47200
rect 14280 47048 14332 47054
rect 14280 46990 14332 46996
rect 14292 46510 14320 46990
rect 15488 46986 15516 51200
rect 16132 48754 16160 51200
rect 16580 49224 16632 49230
rect 16580 49166 16632 49172
rect 16672 49224 16724 49230
rect 16672 49166 16724 49172
rect 16120 48748 16172 48754
rect 16120 48690 16172 48696
rect 16592 48210 16620 49166
rect 16684 48754 16712 49166
rect 16776 48770 16804 51200
rect 16672 48748 16724 48754
rect 16776 48742 16988 48770
rect 16672 48690 16724 48696
rect 16960 48686 16988 48742
rect 16856 48680 16908 48686
rect 16856 48622 16908 48628
rect 16948 48680 17000 48686
rect 16948 48622 17000 48628
rect 16580 48204 16632 48210
rect 16580 48146 16632 48152
rect 16868 47802 16896 48622
rect 17132 48272 17184 48278
rect 17132 48214 17184 48220
rect 16856 47796 16908 47802
rect 16856 47738 16908 47744
rect 16672 47660 16724 47666
rect 16672 47602 16724 47608
rect 16684 47258 16712 47602
rect 17144 47598 17172 48214
rect 17420 48210 17448 51200
rect 18064 49298 18092 51200
rect 18052 49292 18104 49298
rect 18052 49234 18104 49240
rect 19352 49230 19380 51200
rect 19996 49230 20024 51200
rect 20444 49292 20496 49298
rect 20444 49234 20496 49240
rect 19340 49224 19392 49230
rect 19340 49166 19392 49172
rect 19984 49224 20036 49230
rect 19984 49166 20036 49172
rect 20168 49088 20220 49094
rect 20168 49030 20220 49036
rect 20352 49088 20404 49094
rect 20352 49030 20404 49036
rect 19574 48988 19882 49008
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48912 19882 48932
rect 20180 48890 20208 49030
rect 20168 48884 20220 48890
rect 20168 48826 20220 48832
rect 18604 48612 18656 48618
rect 18604 48554 18656 48560
rect 17408 48204 17460 48210
rect 17408 48146 17460 48152
rect 17408 48068 17460 48074
rect 17408 48010 17460 48016
rect 17420 47802 17448 48010
rect 17408 47796 17460 47802
rect 17408 47738 17460 47744
rect 17316 47660 17368 47666
rect 17316 47602 17368 47608
rect 17132 47592 17184 47598
rect 17132 47534 17184 47540
rect 17224 47524 17276 47530
rect 17224 47466 17276 47472
rect 16672 47252 16724 47258
rect 16672 47194 16724 47200
rect 15476 46980 15528 46986
rect 15476 46922 15528 46928
rect 16580 46980 16632 46986
rect 16580 46922 16632 46928
rect 14280 46504 14332 46510
rect 14280 46446 14332 46452
rect 15108 44940 15160 44946
rect 15108 44882 15160 44888
rect 15120 43858 15148 44882
rect 15108 43852 15160 43858
rect 15108 43794 15160 43800
rect 15752 42016 15804 42022
rect 15752 41958 15804 41964
rect 15764 41682 15792 41958
rect 16592 41682 16620 46922
rect 15752 41676 15804 41682
rect 15752 41618 15804 41624
rect 16580 41676 16632 41682
rect 16580 41618 16632 41624
rect 15568 41608 15620 41614
rect 15568 41550 15620 41556
rect 15200 41200 15252 41206
rect 15200 41142 15252 41148
rect 15016 41132 15068 41138
rect 15016 41074 15068 41080
rect 12992 34740 13044 34746
rect 12992 34682 13044 34688
rect 14464 34536 14516 34542
rect 14464 34478 14516 34484
rect 14476 33658 14504 34478
rect 14464 33652 14516 33658
rect 14464 33594 14516 33600
rect 14096 32428 14148 32434
rect 14096 32370 14148 32376
rect 14108 32026 14136 32370
rect 14096 32020 14148 32026
rect 14096 31962 14148 31968
rect 13176 31884 13228 31890
rect 13176 31826 13228 31832
rect 12624 31680 12676 31686
rect 12624 31622 12676 31628
rect 12440 30728 12492 30734
rect 12440 30670 12492 30676
rect 12452 30598 12480 30670
rect 12636 30666 12664 31622
rect 13188 31482 13216 31826
rect 14556 31816 14608 31822
rect 14556 31758 14608 31764
rect 13176 31476 13228 31482
rect 13176 31418 13228 31424
rect 14096 31476 14148 31482
rect 14096 31418 14148 31424
rect 13360 31340 13412 31346
rect 13360 31282 13412 31288
rect 13280 30870 13308 30901
rect 13268 30864 13320 30870
rect 13266 30832 13268 30841
rect 13320 30832 13322 30841
rect 13372 30802 13400 31282
rect 13266 30767 13322 30776
rect 13360 30796 13412 30802
rect 13280 30734 13308 30767
rect 13360 30738 13412 30744
rect 14108 30734 14136 31418
rect 14372 31408 14424 31414
rect 14372 31350 14424 31356
rect 13268 30728 13320 30734
rect 13268 30670 13320 30676
rect 14096 30728 14148 30734
rect 14096 30670 14148 30676
rect 12624 30660 12676 30666
rect 12624 30602 12676 30608
rect 12440 30592 12492 30598
rect 12440 30534 12492 30540
rect 12452 30122 12480 30534
rect 12440 30116 12492 30122
rect 12440 30058 12492 30064
rect 13728 29776 13780 29782
rect 13728 29718 13780 29724
rect 12440 29708 12492 29714
rect 12440 29650 12492 29656
rect 12452 28422 12480 29650
rect 13636 29504 13688 29510
rect 13636 29446 13688 29452
rect 13648 29170 13676 29446
rect 13740 29306 13768 29718
rect 14384 29646 14412 31350
rect 14568 31210 14596 31758
rect 14556 31204 14608 31210
rect 14556 31146 14608 31152
rect 14372 29640 14424 29646
rect 14372 29582 14424 29588
rect 14568 29510 14596 31146
rect 14372 29504 14424 29510
rect 14372 29446 14424 29452
rect 14556 29504 14608 29510
rect 14556 29446 14608 29452
rect 13728 29300 13780 29306
rect 13728 29242 13780 29248
rect 14384 29170 14412 29446
rect 12900 29164 12952 29170
rect 12900 29106 12952 29112
rect 13636 29164 13688 29170
rect 13636 29106 13688 29112
rect 14372 29164 14424 29170
rect 14372 29106 14424 29112
rect 12532 28960 12584 28966
rect 12532 28902 12584 28908
rect 12544 28558 12572 28902
rect 12532 28552 12584 28558
rect 12532 28494 12584 28500
rect 12440 28416 12492 28422
rect 12440 28358 12492 28364
rect 12544 27946 12572 28494
rect 12716 28484 12768 28490
rect 12716 28426 12768 28432
rect 12728 28082 12756 28426
rect 12716 28076 12768 28082
rect 12716 28018 12768 28024
rect 12532 27940 12584 27946
rect 12532 27882 12584 27888
rect 12544 27614 12572 27882
rect 12716 27668 12768 27674
rect 12544 27586 12664 27614
rect 12716 27610 12768 27616
rect 12532 27532 12584 27538
rect 12532 27474 12584 27480
rect 12544 26382 12572 27474
rect 12636 27402 12664 27586
rect 12624 27396 12676 27402
rect 12624 27338 12676 27344
rect 12532 26376 12584 26382
rect 12532 26318 12584 26324
rect 12532 26240 12584 26246
rect 12532 26182 12584 26188
rect 12440 25968 12492 25974
rect 12440 25910 12492 25916
rect 12452 25838 12480 25910
rect 12440 25832 12492 25838
rect 12440 25774 12492 25780
rect 12544 25770 12572 26182
rect 12728 26042 12756 27610
rect 12912 27606 12940 29106
rect 13360 28960 13412 28966
rect 13360 28902 13412 28908
rect 13372 28626 13400 28902
rect 13360 28620 13412 28626
rect 13360 28562 13412 28568
rect 14004 28620 14056 28626
rect 14004 28562 14056 28568
rect 12992 28484 13044 28490
rect 12992 28426 13044 28432
rect 13004 28218 13032 28426
rect 12992 28212 13044 28218
rect 12992 28154 13044 28160
rect 12992 28076 13044 28082
rect 12992 28018 13044 28024
rect 12900 27600 12952 27606
rect 12900 27542 12952 27548
rect 12808 27328 12860 27334
rect 12808 27270 12860 27276
rect 12820 27130 12848 27270
rect 12808 27124 12860 27130
rect 12808 27066 12860 27072
rect 13004 27062 13032 28018
rect 12992 27056 13044 27062
rect 12992 26998 13044 27004
rect 13372 26858 13400 28562
rect 14016 28082 14044 28562
rect 14280 28552 14332 28558
rect 14280 28494 14332 28500
rect 14096 28144 14148 28150
rect 14096 28086 14148 28092
rect 14004 28076 14056 28082
rect 14004 28018 14056 28024
rect 14108 26976 14136 28086
rect 14292 27606 14320 28494
rect 14384 28218 14412 29106
rect 14372 28212 14424 28218
rect 14372 28154 14424 28160
rect 14280 27600 14332 27606
rect 14280 27542 14332 27548
rect 14188 26988 14240 26994
rect 14108 26948 14188 26976
rect 14188 26930 14240 26936
rect 13360 26852 13412 26858
rect 13360 26794 13412 26800
rect 13372 26382 13400 26794
rect 14292 26382 14320 27542
rect 14372 26988 14424 26994
rect 14372 26930 14424 26936
rect 14384 26586 14412 26930
rect 14464 26784 14516 26790
rect 14464 26726 14516 26732
rect 14372 26580 14424 26586
rect 14372 26522 14424 26528
rect 14476 26382 14504 26726
rect 13360 26376 13412 26382
rect 13360 26318 13412 26324
rect 14280 26376 14332 26382
rect 14280 26318 14332 26324
rect 14464 26376 14516 26382
rect 14464 26318 14516 26324
rect 13176 26308 13228 26314
rect 13176 26250 13228 26256
rect 12716 26036 12768 26042
rect 12716 25978 12768 25984
rect 12808 25900 12860 25906
rect 12808 25842 12860 25848
rect 12532 25764 12584 25770
rect 12532 25706 12584 25712
rect 12624 25696 12676 25702
rect 12624 25638 12676 25644
rect 12636 23730 12664 25638
rect 12820 25226 12848 25842
rect 13188 25702 13216 26250
rect 13176 25696 13228 25702
rect 13176 25638 13228 25644
rect 12900 25492 12952 25498
rect 12900 25434 12952 25440
rect 12912 25294 12940 25434
rect 12900 25288 12952 25294
rect 12900 25230 12952 25236
rect 12808 25220 12860 25226
rect 12808 25162 12860 25168
rect 12900 25152 12952 25158
rect 12900 25094 12952 25100
rect 12912 24410 12940 25094
rect 12900 24404 12952 24410
rect 12900 24346 12952 24352
rect 12900 24200 12952 24206
rect 12900 24142 12952 24148
rect 12912 23866 12940 24142
rect 12900 23860 12952 23866
rect 12900 23802 12952 23808
rect 12624 23724 12676 23730
rect 12624 23666 12676 23672
rect 12440 23520 12492 23526
rect 12440 23462 12492 23468
rect 12452 23050 12480 23462
rect 12992 23112 13044 23118
rect 12992 23054 13044 23060
rect 13084 23112 13136 23118
rect 13084 23054 13136 23060
rect 12440 23044 12492 23050
rect 12440 22986 12492 22992
rect 12808 21004 12860 21010
rect 12808 20946 12860 20952
rect 12348 20936 12400 20942
rect 12348 20878 12400 20884
rect 12820 20262 12848 20946
rect 12900 20800 12952 20806
rect 12900 20742 12952 20748
rect 12912 20534 12940 20742
rect 12900 20528 12952 20534
rect 12900 20470 12952 20476
rect 13004 20466 13032 23054
rect 13096 22710 13124 23054
rect 13084 22704 13136 22710
rect 13084 22646 13136 22652
rect 13084 21480 13136 21486
rect 13084 21422 13136 21428
rect 12992 20460 13044 20466
rect 12992 20402 13044 20408
rect 12808 20256 12860 20262
rect 12808 20198 12860 20204
rect 12530 19408 12586 19417
rect 12164 19372 12216 19378
rect 12530 19343 12586 19352
rect 12164 19314 12216 19320
rect 12176 18766 12204 19314
rect 12256 19304 12308 19310
rect 12256 19246 12308 19252
rect 12164 18760 12216 18766
rect 12164 18702 12216 18708
rect 12268 18698 12296 19246
rect 12256 18692 12308 18698
rect 12256 18634 12308 18640
rect 12440 17672 12492 17678
rect 12440 17614 12492 17620
rect 12072 16720 12124 16726
rect 12072 16662 12124 16668
rect 11612 16584 11664 16590
rect 11612 16526 11664 16532
rect 12452 16182 12480 17614
rect 12440 16176 12492 16182
rect 12440 16118 12492 16124
rect 10968 15564 11020 15570
rect 10968 15506 11020 15512
rect 11520 15564 11572 15570
rect 11520 15506 11572 15512
rect 10980 5370 11008 15506
rect 11704 15428 11756 15434
rect 11704 15370 11756 15376
rect 11716 15162 11744 15370
rect 11704 15156 11756 15162
rect 11704 15098 11756 15104
rect 12544 14482 12572 19343
rect 12820 18834 12848 20198
rect 13004 19854 13032 20402
rect 12992 19848 13044 19854
rect 12992 19790 13044 19796
rect 12808 18828 12860 18834
rect 12808 18770 12860 18776
rect 12900 18624 12952 18630
rect 12900 18566 12952 18572
rect 12912 18358 12940 18566
rect 12900 18352 12952 18358
rect 12900 18294 12952 18300
rect 13004 18290 13032 19790
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 13004 17678 13032 18226
rect 12992 17672 13044 17678
rect 12992 17614 13044 17620
rect 13004 17202 13032 17614
rect 12992 17196 13044 17202
rect 12992 17138 13044 17144
rect 12532 14476 12584 14482
rect 12532 14418 12584 14424
rect 12624 14272 12676 14278
rect 12624 14214 12676 14220
rect 12636 14006 12664 14214
rect 12624 14000 12676 14006
rect 12624 13942 12676 13948
rect 12440 12708 12492 12714
rect 12440 12650 12492 12656
rect 12452 9654 12480 12650
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 10968 5364 11020 5370
rect 10968 5306 11020 5312
rect 11704 4480 11756 4486
rect 11704 4422 11756 4428
rect 12440 4480 12492 4486
rect 12440 4422 12492 4428
rect 11716 4214 11744 4422
rect 11704 4208 11756 4214
rect 11704 4150 11756 4156
rect 10692 4004 10744 4010
rect 10692 3946 10744 3952
rect 10784 4004 10836 4010
rect 10784 3946 10836 3952
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 9692 800 9720 2994
rect 10336 800 10364 3878
rect 10796 3534 10824 3946
rect 11612 3732 11664 3738
rect 11612 3674 11664 3680
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 10968 2848 11020 2854
rect 10968 2790 11020 2796
rect 10980 800 11008 2790
rect 11624 800 11652 3674
rect 12164 3664 12216 3670
rect 12164 3606 12216 3612
rect 12256 3664 12308 3670
rect 12256 3606 12308 3612
rect 12176 3369 12204 3606
rect 12162 3360 12218 3369
rect 12162 3295 12218 3304
rect 12164 3052 12216 3058
rect 12164 2994 12216 3000
rect 12176 2650 12204 2994
rect 12164 2644 12216 2650
rect 12164 2586 12216 2592
rect 12268 800 12296 3606
rect 12452 3602 12480 4422
rect 12532 4072 12584 4078
rect 12532 4014 12584 4020
rect 12440 3596 12492 3602
rect 12440 3538 12492 3544
rect 12440 3392 12492 3398
rect 12440 3334 12492 3340
rect 12452 2990 12480 3334
rect 12440 2984 12492 2990
rect 12440 2926 12492 2932
rect 12544 2514 12572 4014
rect 13096 3738 13124 21422
rect 13188 14006 13216 25638
rect 13372 25294 13400 26318
rect 13728 26036 13780 26042
rect 13728 25978 13780 25984
rect 13360 25288 13412 25294
rect 13360 25230 13412 25236
rect 13740 25226 13768 25978
rect 14096 25900 14148 25906
rect 14096 25842 14148 25848
rect 14108 25294 14136 25842
rect 14568 25702 14596 29446
rect 14648 28484 14700 28490
rect 14648 28426 14700 28432
rect 14740 28484 14792 28490
rect 14740 28426 14792 28432
rect 14660 28218 14688 28426
rect 14648 28212 14700 28218
rect 14648 28154 14700 28160
rect 14752 27402 14780 28426
rect 14740 27396 14792 27402
rect 14740 27338 14792 27344
rect 14280 25696 14332 25702
rect 14280 25638 14332 25644
rect 14556 25696 14608 25702
rect 14556 25638 14608 25644
rect 14292 25294 14320 25638
rect 14096 25288 14148 25294
rect 14096 25230 14148 25236
rect 14280 25288 14332 25294
rect 14280 25230 14332 25236
rect 13728 25220 13780 25226
rect 13728 25162 13780 25168
rect 13820 25152 13872 25158
rect 13820 25094 13872 25100
rect 13832 24274 13860 25094
rect 14108 24970 14136 25230
rect 14108 24942 14320 24970
rect 14188 24812 14240 24818
rect 14188 24754 14240 24760
rect 14096 24608 14148 24614
rect 14096 24550 14148 24556
rect 13820 24268 13872 24274
rect 13820 24210 13872 24216
rect 14108 24206 14136 24550
rect 14200 24274 14228 24754
rect 14188 24268 14240 24274
rect 14188 24210 14240 24216
rect 13912 24200 13964 24206
rect 13912 24142 13964 24148
rect 14096 24200 14148 24206
rect 14096 24142 14148 24148
rect 13820 23860 13872 23866
rect 13820 23802 13872 23808
rect 13268 23180 13320 23186
rect 13268 23122 13320 23128
rect 13280 22710 13308 23122
rect 13832 22778 13860 23802
rect 13820 22772 13872 22778
rect 13820 22714 13872 22720
rect 13268 22704 13320 22710
rect 13268 22646 13320 22652
rect 13728 22568 13780 22574
rect 13726 22536 13728 22545
rect 13780 22536 13782 22545
rect 13726 22471 13782 22480
rect 13832 22438 13860 22714
rect 13924 22438 13952 24142
rect 14096 23724 14148 23730
rect 14096 23666 14148 23672
rect 14108 22710 14136 23666
rect 14096 22704 14148 22710
rect 14096 22646 14148 22652
rect 13820 22432 13872 22438
rect 13820 22374 13872 22380
rect 13912 22432 13964 22438
rect 13912 22374 13964 22380
rect 14096 22024 14148 22030
rect 14096 21966 14148 21972
rect 13820 21548 13872 21554
rect 13820 21490 13872 21496
rect 13452 21072 13504 21078
rect 13452 21014 13504 21020
rect 13544 21072 13596 21078
rect 13544 21014 13596 21020
rect 13464 20806 13492 21014
rect 13556 20942 13584 21014
rect 13544 20936 13596 20942
rect 13544 20878 13596 20884
rect 13452 20800 13504 20806
rect 13452 20742 13504 20748
rect 13544 19372 13596 19378
rect 13544 19314 13596 19320
rect 13556 19174 13584 19314
rect 13832 19310 13860 21490
rect 14108 21350 14136 21966
rect 14200 21554 14228 24210
rect 14292 23798 14320 24942
rect 14280 23792 14332 23798
rect 14280 23734 14332 23740
rect 14648 23792 14700 23798
rect 14648 23734 14700 23740
rect 14292 23118 14320 23734
rect 14372 23520 14424 23526
rect 14372 23462 14424 23468
rect 14280 23112 14332 23118
rect 14280 23054 14332 23060
rect 14280 22772 14332 22778
rect 14280 22714 14332 22720
rect 14292 22506 14320 22714
rect 14384 22710 14412 23462
rect 14464 22976 14516 22982
rect 14464 22918 14516 22924
rect 14476 22778 14504 22918
rect 14464 22772 14516 22778
rect 14464 22714 14516 22720
rect 14372 22704 14424 22710
rect 14372 22646 14424 22652
rect 14464 22636 14516 22642
rect 14464 22578 14516 22584
rect 14280 22500 14332 22506
rect 14280 22442 14332 22448
rect 14476 21962 14504 22578
rect 14556 22092 14608 22098
rect 14556 22034 14608 22040
rect 14464 21956 14516 21962
rect 14464 21898 14516 21904
rect 14568 21842 14596 22034
rect 14476 21814 14596 21842
rect 14476 21554 14504 21814
rect 14556 21684 14608 21690
rect 14556 21626 14608 21632
rect 14188 21548 14240 21554
rect 14188 21490 14240 21496
rect 14464 21548 14516 21554
rect 14464 21490 14516 21496
rect 14096 21344 14148 21350
rect 14096 21286 14148 21292
rect 14096 20868 14148 20874
rect 14096 20810 14148 20816
rect 14372 20868 14424 20874
rect 14476 20856 14504 21490
rect 14424 20828 14504 20856
rect 14372 20810 14424 20816
rect 14108 19514 14136 20810
rect 14476 20262 14504 20828
rect 14568 20806 14596 21626
rect 14660 21486 14688 23734
rect 14752 23118 14780 27338
rect 14832 25832 14884 25838
rect 14832 25774 14884 25780
rect 14844 24886 14872 25774
rect 14832 24880 14884 24886
rect 14832 24822 14884 24828
rect 14844 24206 14872 24822
rect 15028 24818 15056 41074
rect 15212 35086 15240 41142
rect 15580 40916 15608 41550
rect 15660 40928 15712 40934
rect 15580 40888 15660 40916
rect 15660 40870 15712 40876
rect 16684 36174 16712 47194
rect 17236 46986 17264 47466
rect 17328 47190 17356 47602
rect 17316 47184 17368 47190
rect 17316 47126 17368 47132
rect 17224 46980 17276 46986
rect 17224 46922 17276 46928
rect 17132 40384 17184 40390
rect 17132 40326 17184 40332
rect 17144 39522 17172 40326
rect 17224 39840 17276 39846
rect 17224 39782 17276 39788
rect 17236 39642 17264 39782
rect 17224 39636 17276 39642
rect 17224 39578 17276 39584
rect 17144 39494 17264 39522
rect 16672 36168 16724 36174
rect 16672 36110 16724 36116
rect 15844 35488 15896 35494
rect 15844 35430 15896 35436
rect 15856 35222 15884 35430
rect 15844 35216 15896 35222
rect 15844 35158 15896 35164
rect 15200 35080 15252 35086
rect 15200 35022 15252 35028
rect 15212 34610 15240 35022
rect 15856 34678 15884 35158
rect 15844 34672 15896 34678
rect 15844 34614 15896 34620
rect 15200 34604 15252 34610
rect 15200 34546 15252 34552
rect 15212 34066 15240 34546
rect 15200 34060 15252 34066
rect 15200 34002 15252 34008
rect 15212 32502 15240 34002
rect 15856 33538 15884 34614
rect 16580 34536 16632 34542
rect 16580 34478 16632 34484
rect 16592 33862 16620 34478
rect 16672 33924 16724 33930
rect 16672 33866 16724 33872
rect 16580 33856 16632 33862
rect 16580 33798 16632 33804
rect 15764 33522 15884 33538
rect 16028 33584 16080 33590
rect 16028 33526 16080 33532
rect 15752 33516 15884 33522
rect 15804 33510 15884 33516
rect 15752 33458 15804 33464
rect 15292 33380 15344 33386
rect 15292 33322 15344 33328
rect 15200 32496 15252 32502
rect 15200 32438 15252 32444
rect 15200 32224 15252 32230
rect 15200 32166 15252 32172
rect 15212 31890 15240 32166
rect 15304 31958 15332 33322
rect 15384 32428 15436 32434
rect 15384 32370 15436 32376
rect 15292 31952 15344 31958
rect 15292 31894 15344 31900
rect 15200 31884 15252 31890
rect 15200 31826 15252 31832
rect 15304 31414 15332 31894
rect 15396 31482 15424 32370
rect 15568 32360 15620 32366
rect 15568 32302 15620 32308
rect 15476 32224 15528 32230
rect 15476 32166 15528 32172
rect 15384 31476 15436 31482
rect 15384 31418 15436 31424
rect 15292 31408 15344 31414
rect 15292 31350 15344 31356
rect 15396 31278 15424 31418
rect 15384 31272 15436 31278
rect 15384 31214 15436 31220
rect 15488 31142 15516 32166
rect 15580 31686 15608 32302
rect 15764 31754 15792 33458
rect 15936 33448 15988 33454
rect 15936 33390 15988 33396
rect 15948 32910 15976 33390
rect 16040 33046 16068 33526
rect 16592 33522 16620 33798
rect 16580 33516 16632 33522
rect 16580 33458 16632 33464
rect 16684 33386 16712 33866
rect 16764 33652 16816 33658
rect 16764 33594 16816 33600
rect 16672 33380 16724 33386
rect 16672 33322 16724 33328
rect 16028 33040 16080 33046
rect 16028 32982 16080 32988
rect 15936 32904 15988 32910
rect 15936 32846 15988 32852
rect 15948 32570 15976 32846
rect 15936 32564 15988 32570
rect 15936 32506 15988 32512
rect 15672 31726 15792 31754
rect 15844 31748 15896 31754
rect 15568 31680 15620 31686
rect 15568 31622 15620 31628
rect 15580 31346 15608 31622
rect 15568 31340 15620 31346
rect 15568 31282 15620 31288
rect 15476 31136 15528 31142
rect 15476 31078 15528 31084
rect 15476 30728 15528 30734
rect 15396 30676 15476 30682
rect 15396 30670 15528 30676
rect 15396 30654 15516 30670
rect 15396 29646 15424 30654
rect 15384 29640 15436 29646
rect 15384 29582 15436 29588
rect 15292 26308 15344 26314
rect 15292 26250 15344 26256
rect 15304 26042 15332 26250
rect 15292 26036 15344 26042
rect 15292 25978 15344 25984
rect 15016 24812 15068 24818
rect 15016 24754 15068 24760
rect 15304 24206 15332 25978
rect 14832 24200 14884 24206
rect 14832 24142 14884 24148
rect 15292 24200 15344 24206
rect 15292 24142 15344 24148
rect 14924 24132 14976 24138
rect 14924 24074 14976 24080
rect 14832 24064 14884 24070
rect 14832 24006 14884 24012
rect 14844 23866 14872 24006
rect 14832 23860 14884 23866
rect 14832 23802 14884 23808
rect 14936 23798 14964 24074
rect 14924 23792 14976 23798
rect 14924 23734 14976 23740
rect 15304 23730 15332 24142
rect 15292 23724 15344 23730
rect 15292 23666 15344 23672
rect 14740 23112 14792 23118
rect 14740 23054 14792 23060
rect 14922 22536 14978 22545
rect 14832 22500 14884 22506
rect 14922 22471 14924 22480
rect 14832 22442 14884 22448
rect 14976 22471 14978 22480
rect 14924 22442 14976 22448
rect 14844 21690 14872 22442
rect 15292 22160 15344 22166
rect 15292 22102 15344 22108
rect 14832 21684 14884 21690
rect 14832 21626 14884 21632
rect 15304 21486 15332 22102
rect 15396 22094 15424 29582
rect 15476 29232 15528 29238
rect 15474 29200 15476 29209
rect 15528 29200 15530 29209
rect 15474 29135 15530 29144
rect 15672 28966 15700 31726
rect 15844 31690 15896 31696
rect 15752 31340 15804 31346
rect 15752 31282 15804 31288
rect 15764 30954 15792 31282
rect 15856 31210 15884 31690
rect 15936 31476 15988 31482
rect 15936 31418 15988 31424
rect 15948 31210 15976 31418
rect 15844 31204 15896 31210
rect 15844 31146 15896 31152
rect 15936 31204 15988 31210
rect 15936 31146 15988 31152
rect 15764 30926 15884 30954
rect 15752 29164 15804 29170
rect 15752 29106 15804 29112
rect 15660 28960 15712 28966
rect 15660 28902 15712 28908
rect 15660 28756 15712 28762
rect 15660 28698 15712 28704
rect 15476 26920 15528 26926
rect 15528 26868 15608 26874
rect 15476 26862 15608 26868
rect 15488 26846 15608 26862
rect 15580 26246 15608 26846
rect 15568 26240 15620 26246
rect 15568 26182 15620 26188
rect 15580 25906 15608 26182
rect 15568 25900 15620 25906
rect 15568 25842 15620 25848
rect 15672 25838 15700 28698
rect 15764 28558 15792 29106
rect 15752 28552 15804 28558
rect 15752 28494 15804 28500
rect 15752 25900 15804 25906
rect 15856 25888 15884 30926
rect 15936 30660 15988 30666
rect 15936 30602 15988 30608
rect 15948 30394 15976 30602
rect 15936 30388 15988 30394
rect 15936 30330 15988 30336
rect 16040 30258 16068 32982
rect 16776 32570 16804 33594
rect 16764 32564 16816 32570
rect 16764 32506 16816 32512
rect 16856 32428 16908 32434
rect 16856 32370 16908 32376
rect 16868 31482 16896 32370
rect 17132 31816 17184 31822
rect 17132 31758 17184 31764
rect 16856 31476 16908 31482
rect 16856 31418 16908 31424
rect 16212 31408 16264 31414
rect 16212 31350 16264 31356
rect 16120 31340 16172 31346
rect 16120 31282 16172 31288
rect 16132 30938 16160 31282
rect 16120 30932 16172 30938
rect 16120 30874 16172 30880
rect 16028 30252 16080 30258
rect 16028 30194 16080 30200
rect 16028 29640 16080 29646
rect 16028 29582 16080 29588
rect 16040 29102 16068 29582
rect 16028 29096 16080 29102
rect 16028 29038 16080 29044
rect 16028 28960 16080 28966
rect 16028 28902 16080 28908
rect 15804 25860 15884 25888
rect 15752 25842 15804 25848
rect 15660 25832 15712 25838
rect 15660 25774 15712 25780
rect 15764 24750 15792 25842
rect 15752 24744 15804 24750
rect 15752 24686 15804 24692
rect 15568 24064 15620 24070
rect 15568 24006 15620 24012
rect 15580 23798 15608 24006
rect 15568 23792 15620 23798
rect 15568 23734 15620 23740
rect 15936 23520 15988 23526
rect 15936 23462 15988 23468
rect 15660 23180 15712 23186
rect 15660 23122 15712 23128
rect 15396 22066 15608 22094
rect 15384 21548 15436 21554
rect 15384 21490 15436 21496
rect 14648 21480 14700 21486
rect 14648 21422 14700 21428
rect 15292 21480 15344 21486
rect 15292 21422 15344 21428
rect 14556 20800 14608 20806
rect 14556 20742 14608 20748
rect 14464 20256 14516 20262
rect 14464 20198 14516 20204
rect 14372 19780 14424 19786
rect 14372 19722 14424 19728
rect 14384 19514 14412 19722
rect 14096 19508 14148 19514
rect 14096 19450 14148 19456
rect 14372 19508 14424 19514
rect 14372 19450 14424 19456
rect 13820 19304 13872 19310
rect 13820 19246 13872 19252
rect 13544 19168 13596 19174
rect 13544 19110 13596 19116
rect 13556 18766 13584 19110
rect 13832 18766 13860 19246
rect 13544 18760 13596 18766
rect 13544 18702 13596 18708
rect 13820 18760 13872 18766
rect 13820 18702 13872 18708
rect 14108 18698 14136 19450
rect 14188 19440 14240 19446
rect 14188 19382 14240 19388
rect 14096 18692 14148 18698
rect 14096 18634 14148 18640
rect 13728 16584 13780 16590
rect 13728 16526 13780 16532
rect 13740 16250 13768 16526
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 14200 16046 14228 19382
rect 14372 19372 14424 19378
rect 14372 19314 14424 19320
rect 14384 18426 14412 19314
rect 14372 18420 14424 18426
rect 14372 18362 14424 18368
rect 14476 18306 14504 20198
rect 14556 19780 14608 19786
rect 14660 19768 14688 21422
rect 15200 19984 15252 19990
rect 15200 19926 15252 19932
rect 14608 19740 14688 19768
rect 14556 19722 14608 19728
rect 14568 19446 14596 19722
rect 15108 19712 15160 19718
rect 15108 19654 15160 19660
rect 14556 19440 14608 19446
rect 14556 19382 14608 19388
rect 15120 19378 15148 19654
rect 15108 19372 15160 19378
rect 15108 19314 15160 19320
rect 14740 18760 14792 18766
rect 14740 18702 14792 18708
rect 14292 18278 14504 18306
rect 14188 16040 14240 16046
rect 14188 15982 14240 15988
rect 14292 15502 14320 18278
rect 14648 17196 14700 17202
rect 14648 17138 14700 17144
rect 14660 16794 14688 17138
rect 14648 16788 14700 16794
rect 14648 16730 14700 16736
rect 14752 16658 14780 18702
rect 15212 17762 15240 19926
rect 15304 19310 15332 21422
rect 15396 21350 15424 21490
rect 15384 21344 15436 21350
rect 15384 21286 15436 21292
rect 15476 20256 15528 20262
rect 15476 20198 15528 20204
rect 15488 19786 15516 20198
rect 15476 19780 15528 19786
rect 15476 19722 15528 19728
rect 15292 19304 15344 19310
rect 15292 19246 15344 19252
rect 15384 19304 15436 19310
rect 15384 19246 15436 19252
rect 15212 17734 15332 17762
rect 15200 17604 15252 17610
rect 15200 17546 15252 17552
rect 15108 17536 15160 17542
rect 15108 17478 15160 17484
rect 14832 16720 14884 16726
rect 14832 16662 14884 16668
rect 14740 16652 14792 16658
rect 14740 16594 14792 16600
rect 14844 16114 14872 16662
rect 15120 16590 15148 17478
rect 15108 16584 15160 16590
rect 15108 16526 15160 16532
rect 15212 16454 15240 17546
rect 15200 16448 15252 16454
rect 15200 16390 15252 16396
rect 14464 16108 14516 16114
rect 14464 16050 14516 16056
rect 14832 16108 14884 16114
rect 14832 16050 14884 16056
rect 14280 15496 14332 15502
rect 14476 15480 14504 16050
rect 15212 15706 15240 16390
rect 15200 15700 15252 15706
rect 15200 15642 15252 15648
rect 14648 15496 14700 15502
rect 14280 15438 14332 15444
rect 14464 15474 14516 15480
rect 13268 15428 13320 15434
rect 14648 15438 14700 15444
rect 14464 15416 14516 15422
rect 13268 15370 13320 15376
rect 13176 14000 13228 14006
rect 13176 13942 13228 13948
rect 13280 3942 13308 15370
rect 14096 15360 14148 15366
rect 14096 15302 14148 15308
rect 13728 15156 13780 15162
rect 13728 15098 13780 15104
rect 13740 14822 13768 15098
rect 14108 15026 14136 15302
rect 14660 15162 14688 15438
rect 14648 15156 14700 15162
rect 14648 15098 14700 15104
rect 14280 15088 14332 15094
rect 14280 15030 14332 15036
rect 14096 15020 14148 15026
rect 14096 14962 14148 14968
rect 13728 14816 13780 14822
rect 13728 14758 13780 14764
rect 13740 14074 13768 14758
rect 14096 14272 14148 14278
rect 14096 14214 14148 14220
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 14108 12850 14136 14214
rect 14292 13394 14320 15030
rect 15212 14958 15240 15642
rect 15304 15502 15332 17734
rect 15396 16590 15424 19246
rect 15580 17762 15608 22066
rect 15672 21690 15700 23122
rect 15948 22710 15976 23462
rect 15936 22704 15988 22710
rect 15936 22646 15988 22652
rect 16040 22438 16068 28902
rect 16028 22432 16080 22438
rect 16028 22374 16080 22380
rect 15660 21684 15712 21690
rect 15660 21626 15712 21632
rect 15750 20632 15806 20641
rect 15750 20567 15806 20576
rect 15764 20466 15792 20567
rect 15752 20460 15804 20466
rect 15752 20402 15804 20408
rect 15936 20460 15988 20466
rect 15936 20402 15988 20408
rect 15948 20058 15976 20402
rect 15936 20052 15988 20058
rect 15936 19994 15988 20000
rect 16224 19922 16252 31350
rect 17144 30326 17172 31758
rect 17132 30320 17184 30326
rect 17132 30262 17184 30268
rect 16304 30252 16356 30258
rect 16304 30194 16356 30200
rect 16316 29714 16344 30194
rect 16304 29708 16356 29714
rect 16304 29650 16356 29656
rect 16764 29504 16816 29510
rect 16764 29446 16816 29452
rect 16580 29232 16632 29238
rect 16580 29174 16632 29180
rect 16592 28218 16620 29174
rect 16580 28212 16632 28218
rect 16580 28154 16632 28160
rect 16776 28150 16804 29446
rect 16946 29200 17002 29209
rect 16946 29135 16948 29144
rect 17000 29135 17002 29144
rect 16948 29106 17000 29112
rect 16764 28144 16816 28150
rect 16764 28086 16816 28092
rect 16776 27470 16804 28086
rect 17144 27606 17172 30262
rect 17236 29714 17264 39494
rect 18616 38962 18644 48554
rect 20260 48544 20312 48550
rect 20260 48486 20312 48492
rect 20272 48210 20300 48486
rect 20260 48204 20312 48210
rect 20260 48146 20312 48152
rect 20168 48068 20220 48074
rect 20168 48010 20220 48016
rect 19574 47900 19882 47920
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47824 19882 47844
rect 20180 47802 20208 48010
rect 20168 47796 20220 47802
rect 20168 47738 20220 47744
rect 20076 47660 20128 47666
rect 20076 47602 20128 47608
rect 19574 46812 19882 46832
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46736 19882 46756
rect 19340 46504 19392 46510
rect 19340 46446 19392 46452
rect 19708 46504 19760 46510
rect 19708 46446 19760 46452
rect 18604 38956 18656 38962
rect 18604 38898 18656 38904
rect 18604 38344 18656 38350
rect 18604 38286 18656 38292
rect 17408 36916 17460 36922
rect 17408 36858 17460 36864
rect 17420 32026 17448 36858
rect 18616 36786 18644 38286
rect 18696 38276 18748 38282
rect 18696 38218 18748 38224
rect 18708 38010 18736 38218
rect 18696 38004 18748 38010
rect 18696 37946 18748 37952
rect 18880 37868 18932 37874
rect 18880 37810 18932 37816
rect 18604 36780 18656 36786
rect 18604 36722 18656 36728
rect 18604 35624 18656 35630
rect 18604 35566 18656 35572
rect 17776 35284 17828 35290
rect 17776 35226 17828 35232
rect 17684 34604 17736 34610
rect 17684 34546 17736 34552
rect 17500 34400 17552 34406
rect 17500 34342 17552 34348
rect 17512 33930 17540 34342
rect 17696 34202 17724 34546
rect 17788 34474 17816 35226
rect 18616 35086 18644 35566
rect 18604 35080 18656 35086
rect 18604 35022 18656 35028
rect 18696 34944 18748 34950
rect 18696 34886 18748 34892
rect 18708 34746 18736 34886
rect 18892 34762 18920 37810
rect 19248 37120 19300 37126
rect 19248 37062 19300 37068
rect 19260 36854 19288 37062
rect 19248 36848 19300 36854
rect 19248 36790 19300 36796
rect 19156 36100 19208 36106
rect 19156 36042 19208 36048
rect 19168 35578 19196 36042
rect 19248 36032 19300 36038
rect 19248 35974 19300 35980
rect 19260 35766 19288 35974
rect 19248 35760 19300 35766
rect 19248 35702 19300 35708
rect 19168 35550 19288 35578
rect 19156 35080 19208 35086
rect 19156 35022 19208 35028
rect 18696 34740 18748 34746
rect 18892 34734 19012 34762
rect 18696 34682 18748 34688
rect 17776 34468 17828 34474
rect 17776 34410 17828 34416
rect 17684 34196 17736 34202
rect 17684 34138 17736 34144
rect 17500 33924 17552 33930
rect 17500 33866 17552 33872
rect 17512 33454 17540 33866
rect 17500 33448 17552 33454
rect 17500 33390 17552 33396
rect 17408 32020 17460 32026
rect 17408 31962 17460 31968
rect 17420 30666 17448 31962
rect 17408 30660 17460 30666
rect 17408 30602 17460 30608
rect 17592 30592 17644 30598
rect 17592 30534 17644 30540
rect 17224 29708 17276 29714
rect 17224 29650 17276 29656
rect 17316 28960 17368 28966
rect 17316 28902 17368 28908
rect 17132 27600 17184 27606
rect 17132 27542 17184 27548
rect 16764 27464 16816 27470
rect 16764 27406 16816 27412
rect 16672 26784 16724 26790
rect 16672 26726 16724 26732
rect 16684 26382 16712 26726
rect 16672 26376 16724 26382
rect 16672 26318 16724 26324
rect 16776 25906 16804 27406
rect 17040 27328 17092 27334
rect 17040 27270 17092 27276
rect 17052 26994 17080 27270
rect 17020 26988 17080 26994
rect 17072 26948 17080 26988
rect 17020 26930 17072 26936
rect 17144 26586 17172 27542
rect 17328 26994 17356 28902
rect 17604 27538 17632 30534
rect 17592 27532 17644 27538
rect 17592 27474 17644 27480
rect 17604 26994 17632 27474
rect 17316 26988 17368 26994
rect 17316 26930 17368 26936
rect 17592 26988 17644 26994
rect 17592 26930 17644 26936
rect 17224 26852 17276 26858
rect 17224 26794 17276 26800
rect 17132 26580 17184 26586
rect 17132 26522 17184 26528
rect 16764 25900 16816 25906
rect 16764 25842 16816 25848
rect 17144 25838 17172 26522
rect 17236 26042 17264 26794
rect 17224 26036 17276 26042
rect 17224 25978 17276 25984
rect 17132 25832 17184 25838
rect 17132 25774 17184 25780
rect 17040 25492 17092 25498
rect 17040 25434 17092 25440
rect 17052 25158 17080 25434
rect 17040 25152 17092 25158
rect 17040 25094 17092 25100
rect 17316 24200 17368 24206
rect 17316 24142 17368 24148
rect 16672 24132 16724 24138
rect 16672 24074 16724 24080
rect 16578 24032 16634 24041
rect 16578 23967 16634 23976
rect 16592 23186 16620 23967
rect 16684 23866 16712 24074
rect 16672 23860 16724 23866
rect 16672 23802 16724 23808
rect 17132 23724 17184 23730
rect 17132 23666 17184 23672
rect 17144 23254 17172 23666
rect 17328 23594 17356 24142
rect 17408 24064 17460 24070
rect 17406 24032 17408 24041
rect 17460 24032 17462 24041
rect 17406 23967 17462 23976
rect 17316 23588 17368 23594
rect 17316 23530 17368 23536
rect 17132 23248 17184 23254
rect 17132 23190 17184 23196
rect 16580 23180 16632 23186
rect 16580 23122 16632 23128
rect 17224 23180 17276 23186
rect 17224 23122 17276 23128
rect 16856 23112 16908 23118
rect 16856 23054 16908 23060
rect 16580 23044 16632 23050
rect 16580 22986 16632 22992
rect 16592 22094 16620 22986
rect 16592 22066 16712 22094
rect 16684 22030 16712 22066
rect 16672 22024 16724 22030
rect 16672 21966 16724 21972
rect 16488 21548 16540 21554
rect 16488 21490 16540 21496
rect 16212 19916 16264 19922
rect 16212 19858 16264 19864
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 15752 18624 15804 18630
rect 15752 18566 15804 18572
rect 15488 17734 15608 17762
rect 15764 17746 15792 18566
rect 15948 18426 15976 19790
rect 16500 19378 16528 21490
rect 16764 21344 16816 21350
rect 16764 21286 16816 21292
rect 16672 21072 16724 21078
rect 16672 21014 16724 21020
rect 16684 20505 16712 21014
rect 16776 20874 16804 21286
rect 16868 21010 16896 23054
rect 17236 22778 17264 23122
rect 17328 23118 17356 23530
rect 17316 23112 17368 23118
rect 17316 23054 17368 23060
rect 17224 22772 17276 22778
rect 17224 22714 17276 22720
rect 17224 22092 17276 22098
rect 17224 22034 17276 22040
rect 17236 21622 17264 22034
rect 17592 21956 17644 21962
rect 17592 21898 17644 21904
rect 17224 21616 17276 21622
rect 17224 21558 17276 21564
rect 17408 21616 17460 21622
rect 17408 21558 17460 21564
rect 16856 21004 16908 21010
rect 16856 20946 16908 20952
rect 17420 20942 17448 21558
rect 17604 20942 17632 21898
rect 17408 20936 17460 20942
rect 17408 20878 17460 20884
rect 17592 20936 17644 20942
rect 17592 20878 17644 20884
rect 16764 20868 16816 20874
rect 16764 20810 16816 20816
rect 17500 20868 17552 20874
rect 17500 20810 17552 20816
rect 17512 20602 17540 20810
rect 17132 20596 17184 20602
rect 17132 20538 17184 20544
rect 17500 20596 17552 20602
rect 17500 20538 17552 20544
rect 16670 20496 16726 20505
rect 16670 20431 16726 20440
rect 16684 20058 16712 20431
rect 16672 20052 16724 20058
rect 16672 19994 16724 20000
rect 17144 19990 17172 20538
rect 17316 20460 17368 20466
rect 17316 20402 17368 20408
rect 17224 20256 17276 20262
rect 17224 20198 17276 20204
rect 17132 19984 17184 19990
rect 17132 19926 17184 19932
rect 16856 19780 16908 19786
rect 16856 19722 16908 19728
rect 16948 19780 17000 19786
rect 16948 19722 17000 19728
rect 16868 19514 16896 19722
rect 16856 19508 16908 19514
rect 16856 19450 16908 19456
rect 16960 19446 16988 19722
rect 16948 19440 17000 19446
rect 16948 19382 17000 19388
rect 16488 19372 16540 19378
rect 16488 19314 16540 19320
rect 16120 19236 16172 19242
rect 16120 19178 16172 19184
rect 16132 18766 16160 19178
rect 16120 18760 16172 18766
rect 16120 18702 16172 18708
rect 15936 18420 15988 18426
rect 15936 18362 15988 18368
rect 15752 17740 15804 17746
rect 15384 16584 15436 16590
rect 15384 16526 15436 16532
rect 15292 15496 15344 15502
rect 15292 15438 15344 15444
rect 15200 14952 15252 14958
rect 15200 14894 15252 14900
rect 14924 14408 14976 14414
rect 14924 14350 14976 14356
rect 14936 13938 14964 14350
rect 15200 14340 15252 14346
rect 15200 14282 15252 14288
rect 14924 13932 14976 13938
rect 14924 13874 14976 13880
rect 15212 13870 15240 14282
rect 15200 13864 15252 13870
rect 15200 13806 15252 13812
rect 15016 13728 15068 13734
rect 15016 13670 15068 13676
rect 14280 13388 14332 13394
rect 14280 13330 14332 13336
rect 15028 13258 15056 13670
rect 15212 13326 15240 13806
rect 15200 13320 15252 13326
rect 15200 13262 15252 13268
rect 15016 13252 15068 13258
rect 15016 13194 15068 13200
rect 15304 12918 15332 15438
rect 15488 13938 15516 17734
rect 15752 17682 15804 17688
rect 15568 17672 15620 17678
rect 15568 17614 15620 17620
rect 15580 17066 15608 17614
rect 15568 17060 15620 17066
rect 15568 17002 15620 17008
rect 16396 16652 16448 16658
rect 16396 16594 16448 16600
rect 16408 16522 16436 16594
rect 16396 16516 16448 16522
rect 16396 16458 16448 16464
rect 15660 16448 15712 16454
rect 15660 16390 15712 16396
rect 15672 16182 15700 16390
rect 15660 16176 15712 16182
rect 15660 16118 15712 16124
rect 16408 16114 16436 16458
rect 16396 16108 16448 16114
rect 16396 16050 16448 16056
rect 16408 15570 16436 16050
rect 16396 15564 16448 15570
rect 16396 15506 16448 15512
rect 16500 15502 16528 19314
rect 16856 18692 16908 18698
rect 16856 18634 16908 18640
rect 16868 18426 16896 18634
rect 17236 18426 17264 20198
rect 17328 19174 17356 20402
rect 17500 19780 17552 19786
rect 17500 19722 17552 19728
rect 17512 19378 17540 19722
rect 17500 19372 17552 19378
rect 17500 19314 17552 19320
rect 17316 19168 17368 19174
rect 17316 19110 17368 19116
rect 17500 19168 17552 19174
rect 17500 19110 17552 19116
rect 16856 18420 16908 18426
rect 16856 18362 16908 18368
rect 17224 18420 17276 18426
rect 17224 18362 17276 18368
rect 17512 18290 17540 19110
rect 17040 18284 17092 18290
rect 17040 18226 17092 18232
rect 17500 18284 17552 18290
rect 17500 18226 17552 18232
rect 16856 17196 16908 17202
rect 16856 17138 16908 17144
rect 16672 17128 16724 17134
rect 16672 17070 16724 17076
rect 16488 15496 16540 15502
rect 16488 15438 16540 15444
rect 16684 15026 16712 17070
rect 16868 16794 16896 17138
rect 16856 16788 16908 16794
rect 16856 16730 16908 16736
rect 17052 16574 17080 18226
rect 17316 16584 17368 16590
rect 17052 16546 17172 16574
rect 16948 15360 17000 15366
rect 16948 15302 17000 15308
rect 16960 15094 16988 15302
rect 16948 15088 17000 15094
rect 16948 15030 17000 15036
rect 16672 15020 16724 15026
rect 16672 14962 16724 14968
rect 16684 14074 16712 14962
rect 16672 14068 16724 14074
rect 16672 14010 16724 14016
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 15488 13546 15516 13874
rect 15488 13530 15608 13546
rect 15488 13524 15620 13530
rect 15488 13518 15568 13524
rect 15568 13466 15620 13472
rect 15292 12912 15344 12918
rect 15292 12854 15344 12860
rect 16684 12850 16712 14010
rect 14096 12844 14148 12850
rect 14096 12786 14148 12792
rect 16672 12844 16724 12850
rect 16672 12786 16724 12792
rect 14280 12776 14332 12782
rect 14280 12718 14332 12724
rect 14292 12442 14320 12718
rect 14280 12436 14332 12442
rect 14280 12378 14332 12384
rect 16684 11694 16712 12786
rect 16672 11688 16724 11694
rect 16672 11630 16724 11636
rect 17040 11688 17092 11694
rect 17040 11630 17092 11636
rect 17052 10130 17080 11630
rect 17144 11150 17172 16546
rect 17316 16526 17368 16532
rect 17328 16250 17356 16526
rect 17316 16244 17368 16250
rect 17316 16186 17368 16192
rect 17316 16108 17368 16114
rect 17316 16050 17368 16056
rect 17328 15706 17356 16050
rect 17316 15700 17368 15706
rect 17316 15642 17368 15648
rect 17328 15434 17356 15642
rect 17316 15428 17368 15434
rect 17316 15370 17368 15376
rect 17500 15428 17552 15434
rect 17500 15370 17552 15376
rect 17224 15360 17276 15366
rect 17224 15302 17276 15308
rect 17236 13258 17264 15302
rect 17512 15162 17540 15370
rect 17500 15156 17552 15162
rect 17500 15098 17552 15104
rect 17512 13938 17540 15098
rect 17500 13932 17552 13938
rect 17500 13874 17552 13880
rect 17224 13252 17276 13258
rect 17224 13194 17276 13200
rect 17236 11762 17264 13194
rect 17224 11756 17276 11762
rect 17224 11698 17276 11704
rect 17132 11144 17184 11150
rect 17132 11086 17184 11092
rect 17040 10124 17092 10130
rect 17040 10066 17092 10072
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 15200 6112 15252 6118
rect 15200 6054 15252 6060
rect 14096 4548 14148 4554
rect 14096 4490 14148 4496
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 13084 3732 13136 3738
rect 13084 3674 13136 3680
rect 14108 3670 14136 4490
rect 14280 3936 14332 3942
rect 14280 3878 14332 3884
rect 15108 3936 15160 3942
rect 15108 3878 15160 3884
rect 12624 3664 12676 3670
rect 12624 3606 12676 3612
rect 14096 3664 14148 3670
rect 14096 3606 14148 3612
rect 12636 3369 12664 3606
rect 12622 3360 12678 3369
rect 12622 3295 12678 3304
rect 14188 3052 14240 3058
rect 14188 2994 14240 3000
rect 12900 2984 12952 2990
rect 12900 2926 12952 2932
rect 12532 2508 12584 2514
rect 12532 2450 12584 2456
rect 12912 800 12940 2926
rect 13544 2508 13596 2514
rect 13544 2450 13596 2456
rect 13556 800 13584 2450
rect 14200 800 14228 2994
rect 14292 2378 14320 3878
rect 15120 3602 15148 3878
rect 15108 3596 15160 3602
rect 15108 3538 15160 3544
rect 14924 3528 14976 3534
rect 14924 3470 14976 3476
rect 14648 3392 14700 3398
rect 14648 3334 14700 3340
rect 14660 2922 14688 3334
rect 14936 3058 14964 3470
rect 14924 3052 14976 3058
rect 14924 2994 14976 3000
rect 14648 2916 14700 2922
rect 14648 2858 14700 2864
rect 14280 2372 14332 2378
rect 14280 2314 14332 2320
rect 15212 2310 15240 6054
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 15200 2304 15252 2310
rect 15200 2246 15252 2252
rect 15488 800 15516 3538
rect 16592 2854 16620 9318
rect 17696 8362 17724 34138
rect 18144 34128 18196 34134
rect 18144 34070 18196 34076
rect 17868 33856 17920 33862
rect 17868 33798 17920 33804
rect 17880 33522 17908 33798
rect 17868 33516 17920 33522
rect 17868 33458 17920 33464
rect 18052 33448 18104 33454
rect 18052 33390 18104 33396
rect 18064 32366 18092 33390
rect 18052 32360 18104 32366
rect 18052 32302 18104 32308
rect 18064 31822 18092 32302
rect 18052 31816 18104 31822
rect 18052 31758 18104 31764
rect 18064 31346 18092 31758
rect 18052 31340 18104 31346
rect 18052 31282 18104 31288
rect 17776 30252 17828 30258
rect 17776 30194 17828 30200
rect 17788 30122 17816 30194
rect 17776 30116 17828 30122
rect 17776 30058 17828 30064
rect 17776 29640 17828 29646
rect 17776 29582 17828 29588
rect 17788 28694 17816 29582
rect 18156 29306 18184 34070
rect 18328 32904 18380 32910
rect 18328 32846 18380 32852
rect 18512 32904 18564 32910
rect 18512 32846 18564 32852
rect 18340 31929 18368 32846
rect 18524 32570 18552 32846
rect 18512 32564 18564 32570
rect 18512 32506 18564 32512
rect 18696 32360 18748 32366
rect 18696 32302 18748 32308
rect 18708 32026 18736 32302
rect 18788 32224 18840 32230
rect 18788 32166 18840 32172
rect 18880 32224 18932 32230
rect 18880 32166 18932 32172
rect 18696 32020 18748 32026
rect 18696 31962 18748 31968
rect 18326 31920 18382 31929
rect 18326 31855 18382 31864
rect 18800 31822 18828 32166
rect 18788 31816 18840 31822
rect 18788 31758 18840 31764
rect 18892 31754 18920 32166
rect 18880 31748 18932 31754
rect 18880 31690 18932 31696
rect 18892 31482 18920 31690
rect 18880 31476 18932 31482
rect 18880 31418 18932 31424
rect 18420 31136 18472 31142
rect 18420 31078 18472 31084
rect 18432 30326 18460 31078
rect 18420 30320 18472 30326
rect 18420 30262 18472 30268
rect 18604 30116 18656 30122
rect 18604 30058 18656 30064
rect 18616 29646 18644 30058
rect 18604 29640 18656 29646
rect 18604 29582 18656 29588
rect 18328 29504 18380 29510
rect 18328 29446 18380 29452
rect 18144 29300 18196 29306
rect 18144 29242 18196 29248
rect 18052 28960 18104 28966
rect 18052 28902 18104 28908
rect 17776 28688 17828 28694
rect 17776 28630 17828 28636
rect 17788 27334 17816 28630
rect 18064 28558 18092 28902
rect 18052 28552 18104 28558
rect 18052 28494 18104 28500
rect 18156 28150 18184 29242
rect 18340 28626 18368 29446
rect 18604 29164 18656 29170
rect 18604 29106 18656 29112
rect 18616 28762 18644 29106
rect 18604 28756 18656 28762
rect 18604 28698 18656 28704
rect 18328 28620 18380 28626
rect 18328 28562 18380 28568
rect 18144 28144 18196 28150
rect 18144 28086 18196 28092
rect 17868 27464 17920 27470
rect 17868 27406 17920 27412
rect 17776 27328 17828 27334
rect 17776 27270 17828 27276
rect 17788 27062 17816 27270
rect 17776 27056 17828 27062
rect 17776 26998 17828 27004
rect 17788 25226 17816 26998
rect 17880 26926 17908 27406
rect 18236 27328 18288 27334
rect 18236 27270 18288 27276
rect 18248 26994 18276 27270
rect 18236 26988 18288 26994
rect 18236 26930 18288 26936
rect 18512 26988 18564 26994
rect 18512 26930 18564 26936
rect 17868 26920 17920 26926
rect 17868 26862 17920 26868
rect 18524 26858 18552 26930
rect 18512 26852 18564 26858
rect 18512 26794 18564 26800
rect 18236 26784 18288 26790
rect 18236 26726 18288 26732
rect 18328 26784 18380 26790
rect 18328 26726 18380 26732
rect 17960 26308 18012 26314
rect 17960 26250 18012 26256
rect 17972 25362 18000 26250
rect 18052 26240 18104 26246
rect 18052 26182 18104 26188
rect 18064 25906 18092 26182
rect 18248 25906 18276 26726
rect 18052 25900 18104 25906
rect 18052 25842 18104 25848
rect 18236 25900 18288 25906
rect 18236 25842 18288 25848
rect 17960 25356 18012 25362
rect 17960 25298 18012 25304
rect 18340 25294 18368 26726
rect 18788 26240 18840 26246
rect 18788 26182 18840 26188
rect 18328 25288 18380 25294
rect 18328 25230 18380 25236
rect 17776 25220 17828 25226
rect 17776 25162 17828 25168
rect 18696 24200 18748 24206
rect 18696 24142 18748 24148
rect 18236 24132 18288 24138
rect 18236 24074 18288 24080
rect 18052 24064 18104 24070
rect 18052 24006 18104 24012
rect 18064 23798 18092 24006
rect 18248 23866 18276 24074
rect 18236 23860 18288 23866
rect 18236 23802 18288 23808
rect 18052 23792 18104 23798
rect 18052 23734 18104 23740
rect 18144 23724 18196 23730
rect 18144 23666 18196 23672
rect 17868 23656 17920 23662
rect 17868 23598 17920 23604
rect 17880 23118 17908 23598
rect 17868 23112 17920 23118
rect 17868 23054 17920 23060
rect 17960 22976 18012 22982
rect 17960 22918 18012 22924
rect 18052 22976 18104 22982
rect 18052 22918 18104 22924
rect 17972 22778 18000 22918
rect 17960 22772 18012 22778
rect 17960 22714 18012 22720
rect 18064 22658 18092 22918
rect 17972 22630 18092 22658
rect 17972 22506 18000 22630
rect 18156 22506 18184 23666
rect 18248 22642 18276 23802
rect 18708 23798 18736 24142
rect 18696 23792 18748 23798
rect 18696 23734 18748 23740
rect 18418 22672 18474 22681
rect 18236 22636 18288 22642
rect 18236 22578 18288 22584
rect 18328 22636 18380 22642
rect 18418 22607 18474 22616
rect 18328 22578 18380 22584
rect 17960 22500 18012 22506
rect 17960 22442 18012 22448
rect 18144 22500 18196 22506
rect 18144 22442 18196 22448
rect 17972 22030 18000 22442
rect 17960 22024 18012 22030
rect 17960 21966 18012 21972
rect 17776 20800 17828 20806
rect 17776 20742 17828 20748
rect 17788 19786 17816 20742
rect 17958 20632 18014 20641
rect 17868 20596 17920 20602
rect 17958 20567 17960 20576
rect 17868 20538 17920 20544
rect 18012 20567 18014 20576
rect 17960 20538 18012 20544
rect 17880 20262 17908 20538
rect 18156 20505 18184 22442
rect 18248 22114 18276 22578
rect 18340 22234 18368 22578
rect 18432 22506 18460 22607
rect 18420 22500 18472 22506
rect 18420 22442 18472 22448
rect 18328 22228 18380 22234
rect 18328 22170 18380 22176
rect 18512 22160 18564 22166
rect 18248 22108 18512 22114
rect 18248 22102 18564 22108
rect 18248 22086 18552 22102
rect 18236 21344 18288 21350
rect 18236 21286 18288 21292
rect 18248 20788 18276 21286
rect 18328 20800 18380 20806
rect 18248 20760 18328 20788
rect 18142 20496 18198 20505
rect 18142 20431 18144 20440
rect 18196 20431 18198 20440
rect 18144 20402 18196 20408
rect 18052 20392 18104 20398
rect 18052 20334 18104 20340
rect 17868 20256 17920 20262
rect 17868 20198 17920 20204
rect 18064 20058 18092 20334
rect 18052 20052 18104 20058
rect 18052 19994 18104 20000
rect 17776 19780 17828 19786
rect 17776 19722 17828 19728
rect 18144 19372 18196 19378
rect 18144 19314 18196 19320
rect 18156 18154 18184 19314
rect 18144 18148 18196 18154
rect 18144 18090 18196 18096
rect 17868 17876 17920 17882
rect 17868 17818 17920 17824
rect 17880 16590 17908 17818
rect 18156 17814 18184 18090
rect 18144 17808 18196 17814
rect 18144 17750 18196 17756
rect 17960 17604 18012 17610
rect 17960 17546 18012 17552
rect 17972 16794 18000 17546
rect 17960 16788 18012 16794
rect 17960 16730 18012 16736
rect 17868 16584 17920 16590
rect 17868 16526 17920 16532
rect 17880 16250 17908 16526
rect 17868 16244 17920 16250
rect 17868 16186 17920 16192
rect 17868 16108 17920 16114
rect 17868 16050 17920 16056
rect 17880 15978 17908 16050
rect 17868 15972 17920 15978
rect 17868 15914 17920 15920
rect 17880 15434 17908 15914
rect 17868 15428 17920 15434
rect 17868 15370 17920 15376
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 17972 14482 18000 14962
rect 17960 14476 18012 14482
rect 17960 14418 18012 14424
rect 17868 13184 17920 13190
rect 17868 13126 17920 13132
rect 17880 12918 17908 13126
rect 17868 12912 17920 12918
rect 17868 12854 17920 12860
rect 18052 12640 18104 12646
rect 18052 12582 18104 12588
rect 18064 12306 18092 12582
rect 18052 12300 18104 12306
rect 18052 12242 18104 12248
rect 17868 12164 17920 12170
rect 17868 12106 17920 12112
rect 17776 9512 17828 9518
rect 17776 9454 17828 9460
rect 17788 9178 17816 9454
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 17684 8356 17736 8362
rect 17684 8298 17736 8304
rect 17684 7744 17736 7750
rect 17684 7686 17736 7692
rect 17696 7410 17724 7686
rect 17684 7404 17736 7410
rect 17684 7346 17736 7352
rect 17880 3738 17908 12106
rect 18248 12102 18276 20760
rect 18328 20742 18380 20748
rect 18604 19780 18656 19786
rect 18604 19722 18656 19728
rect 18328 16992 18380 16998
rect 18328 16934 18380 16940
rect 18340 16182 18368 16934
rect 18512 16788 18564 16794
rect 18512 16730 18564 16736
rect 18328 16176 18380 16182
rect 18328 16118 18380 16124
rect 18420 16108 18472 16114
rect 18420 16050 18472 16056
rect 18328 13320 18380 13326
rect 18328 13262 18380 13268
rect 18340 12442 18368 13262
rect 18328 12436 18380 12442
rect 18328 12378 18380 12384
rect 18236 12096 18288 12102
rect 18236 12038 18288 12044
rect 17960 11348 18012 11354
rect 17960 11290 18012 11296
rect 17972 8974 18000 11290
rect 18248 11150 18276 12038
rect 18432 11642 18460 16050
rect 18524 14414 18552 16730
rect 18616 15026 18644 19722
rect 18604 15020 18656 15026
rect 18604 14962 18656 14968
rect 18604 14816 18656 14822
rect 18604 14758 18656 14764
rect 18512 14408 18564 14414
rect 18512 14350 18564 14356
rect 18616 13870 18644 14758
rect 18696 14340 18748 14346
rect 18696 14282 18748 14288
rect 18708 14006 18736 14282
rect 18696 14000 18748 14006
rect 18696 13942 18748 13948
rect 18604 13864 18656 13870
rect 18604 13806 18656 13812
rect 18604 13388 18656 13394
rect 18604 13330 18656 13336
rect 18512 13320 18564 13326
rect 18512 13262 18564 13268
rect 18340 11614 18460 11642
rect 18236 11144 18288 11150
rect 18236 11086 18288 11092
rect 18340 10554 18368 11614
rect 18420 11552 18472 11558
rect 18420 11494 18472 11500
rect 18156 10526 18368 10554
rect 17960 8968 18012 8974
rect 17960 8910 18012 8916
rect 17972 6798 18000 8910
rect 18052 7880 18104 7886
rect 18052 7822 18104 7828
rect 18064 7546 18092 7822
rect 18052 7540 18104 7546
rect 18052 7482 18104 7488
rect 18156 7154 18184 10526
rect 18432 10470 18460 11494
rect 18524 11014 18552 13262
rect 18616 11286 18644 13330
rect 18708 12918 18736 13942
rect 18696 12912 18748 12918
rect 18696 12854 18748 12860
rect 18800 12434 18828 26182
rect 18708 12406 18828 12434
rect 18880 12436 18932 12442
rect 18604 11280 18656 11286
rect 18604 11222 18656 11228
rect 18512 11008 18564 11014
rect 18512 10950 18564 10956
rect 18616 10538 18644 11222
rect 18604 10532 18656 10538
rect 18604 10474 18656 10480
rect 18328 10464 18380 10470
rect 18328 10406 18380 10412
rect 18420 10464 18472 10470
rect 18420 10406 18472 10412
rect 18340 10062 18368 10406
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 18420 9920 18472 9926
rect 18420 9862 18472 9868
rect 18432 9654 18460 9862
rect 18420 9648 18472 9654
rect 18420 9590 18472 9596
rect 18236 9512 18288 9518
rect 18236 9454 18288 9460
rect 18248 9382 18276 9454
rect 18236 9376 18288 9382
rect 18236 9318 18288 9324
rect 18420 8560 18472 8566
rect 18472 8520 18552 8548
rect 18420 8502 18472 8508
rect 18328 8424 18380 8430
rect 18326 8392 18328 8401
rect 18380 8392 18382 8401
rect 18326 8327 18382 8336
rect 18524 8378 18552 8520
rect 18616 8378 18644 10474
rect 18524 8350 18644 8378
rect 18524 8294 18552 8350
rect 18432 8266 18552 8294
rect 18432 7864 18460 8266
rect 18420 7858 18472 7864
rect 18420 7800 18472 7806
rect 18236 7540 18288 7546
rect 18236 7482 18288 7488
rect 18064 7126 18184 7154
rect 17960 6792 18012 6798
rect 17960 6734 18012 6740
rect 17960 3936 18012 3942
rect 17960 3878 18012 3884
rect 17868 3732 17920 3738
rect 17868 3674 17920 3680
rect 17868 3120 17920 3126
rect 17868 3062 17920 3068
rect 17880 2938 17908 3062
rect 17972 3058 18000 3878
rect 17960 3052 18012 3058
rect 17960 2994 18012 3000
rect 18064 2938 18092 7126
rect 18248 7018 18276 7482
rect 18156 6990 18276 7018
rect 18156 6322 18184 6990
rect 18328 6656 18380 6662
rect 18328 6598 18380 6604
rect 18340 6390 18368 6598
rect 18328 6384 18380 6390
rect 18328 6326 18380 6332
rect 18144 6316 18196 6322
rect 18144 6258 18196 6264
rect 18708 5166 18736 12406
rect 18880 12378 18932 12384
rect 18892 11354 18920 12378
rect 18880 11348 18932 11354
rect 18880 11290 18932 11296
rect 18880 11008 18932 11014
rect 18880 10950 18932 10956
rect 18788 10668 18840 10674
rect 18788 10610 18840 10616
rect 18800 10266 18828 10610
rect 18788 10260 18840 10266
rect 18788 10202 18840 10208
rect 18892 8498 18920 10950
rect 18788 8492 18840 8498
rect 18788 8434 18840 8440
rect 18880 8492 18932 8498
rect 18880 8434 18932 8440
rect 18800 8362 18828 8434
rect 18788 8356 18840 8362
rect 18788 8298 18840 8304
rect 18984 8090 19012 34734
rect 19064 34740 19116 34746
rect 19064 34682 19116 34688
rect 19076 32910 19104 34682
rect 19168 32994 19196 35022
rect 19260 34678 19288 35550
rect 19248 34672 19300 34678
rect 19248 34614 19300 34620
rect 19168 32978 19288 32994
rect 19168 32972 19300 32978
rect 19168 32966 19248 32972
rect 19248 32914 19300 32920
rect 19064 32904 19116 32910
rect 19064 32846 19116 32852
rect 19156 32768 19208 32774
rect 19156 32710 19208 32716
rect 19168 32434 19196 32710
rect 19156 32428 19208 32434
rect 19156 32370 19208 32376
rect 19154 31920 19210 31929
rect 19260 31890 19288 32914
rect 19154 31855 19210 31864
rect 19248 31884 19300 31890
rect 19168 23050 19196 31855
rect 19248 31826 19300 31832
rect 19352 30682 19380 46446
rect 19720 46170 19748 46446
rect 19708 46164 19760 46170
rect 19708 46106 19760 46112
rect 20088 45966 20116 47602
rect 20076 45960 20128 45966
rect 20076 45902 20128 45908
rect 19574 45724 19882 45744
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45648 19882 45668
rect 19574 44636 19882 44656
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44560 19882 44580
rect 19574 43548 19882 43568
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43472 19882 43492
rect 20088 42634 20116 45902
rect 20168 43784 20220 43790
rect 20168 43726 20220 43732
rect 20180 43314 20208 43726
rect 20168 43308 20220 43314
rect 20168 43250 20220 43256
rect 20180 42702 20208 43250
rect 20168 42696 20220 42702
rect 20168 42638 20220 42644
rect 20076 42628 20128 42634
rect 20076 42570 20128 42576
rect 19574 42460 19882 42480
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42384 19882 42404
rect 19574 41372 19882 41392
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41296 19882 41316
rect 19574 40284 19882 40304
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40208 19882 40228
rect 19984 39364 20036 39370
rect 19984 39306 20036 39312
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 19996 39098 20024 39306
rect 19984 39092 20036 39098
rect 19984 39034 20036 39040
rect 19984 38208 20036 38214
rect 19984 38150 20036 38156
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 19996 37942 20024 38150
rect 19800 37936 19852 37942
rect 19800 37878 19852 37884
rect 19984 37936 20036 37942
rect 19984 37878 20036 37884
rect 19616 37732 19668 37738
rect 19616 37674 19668 37680
rect 19628 37398 19656 37674
rect 19616 37392 19668 37398
rect 19616 37334 19668 37340
rect 19812 37262 19840 37878
rect 19432 37256 19484 37262
rect 19432 37198 19484 37204
rect 19800 37256 19852 37262
rect 19800 37198 19852 37204
rect 19444 35698 19472 37198
rect 19984 37188 20036 37194
rect 19984 37130 20036 37136
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19432 35692 19484 35698
rect 19432 35634 19484 35640
rect 19996 35086 20024 37130
rect 19984 35080 20036 35086
rect 19984 35022 20036 35028
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 19432 34604 19484 34610
rect 19432 34546 19484 34552
rect 19444 33522 19472 34546
rect 19996 34134 20024 35022
rect 19984 34128 20036 34134
rect 19984 34070 20036 34076
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 19432 33516 19484 33522
rect 19432 33458 19484 33464
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 19432 32428 19484 32434
rect 19432 32370 19484 32376
rect 19892 32428 19944 32434
rect 19892 32370 19944 32376
rect 19444 31686 19472 32370
rect 19904 32230 19932 32370
rect 19892 32224 19944 32230
rect 19892 32166 19944 32172
rect 20088 31754 20116 42570
rect 19996 31726 20116 31754
rect 19432 31680 19484 31686
rect 19432 31622 19484 31628
rect 19260 30654 19380 30682
rect 19444 30666 19472 31622
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19524 30864 19576 30870
rect 19524 30806 19576 30812
rect 19432 30660 19484 30666
rect 19260 30138 19288 30654
rect 19536 30648 19564 30806
rect 19432 30602 19484 30608
rect 19516 30620 19564 30648
rect 19340 30592 19392 30598
rect 19516 30546 19544 30620
rect 19340 30534 19392 30540
rect 19352 30326 19380 30534
rect 19444 30518 19544 30546
rect 19340 30320 19392 30326
rect 19340 30262 19392 30268
rect 19260 30110 19380 30138
rect 19352 29578 19380 30110
rect 19340 29572 19392 29578
rect 19340 29514 19392 29520
rect 19352 29306 19380 29514
rect 19340 29300 19392 29306
rect 19340 29242 19392 29248
rect 19444 27520 19472 30518
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 19444 27492 19564 27520
rect 19536 27402 19564 27492
rect 19432 27396 19484 27402
rect 19432 27338 19484 27344
rect 19524 27396 19576 27402
rect 19524 27338 19576 27344
rect 19444 26042 19472 27338
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19432 26036 19484 26042
rect 19432 25978 19484 25984
rect 19444 25362 19472 25978
rect 19996 25838 20024 31726
rect 20076 31204 20128 31210
rect 20076 31146 20128 31152
rect 20088 30598 20116 31146
rect 20076 30592 20128 30598
rect 20076 30534 20128 30540
rect 20076 30048 20128 30054
rect 20076 29990 20128 29996
rect 20088 29510 20116 29990
rect 20076 29504 20128 29510
rect 20076 29446 20128 29452
rect 20088 29238 20116 29446
rect 20076 29232 20128 29238
rect 20076 29174 20128 29180
rect 20088 28558 20116 29174
rect 20076 28552 20128 28558
rect 20076 28494 20128 28500
rect 20088 26382 20116 28494
rect 20180 27470 20208 42638
rect 20364 41414 20392 49030
rect 20272 41386 20392 41414
rect 20272 27946 20300 41386
rect 20352 39840 20404 39846
rect 20352 39782 20404 39788
rect 20364 38962 20392 39782
rect 20352 38956 20404 38962
rect 20352 38898 20404 38904
rect 20352 37868 20404 37874
rect 20352 37810 20404 37816
rect 20364 36854 20392 37810
rect 20352 36848 20404 36854
rect 20352 36790 20404 36796
rect 20456 36242 20484 49234
rect 20640 48210 20668 51200
rect 21272 49768 21324 49774
rect 21272 49710 21324 49716
rect 20812 48612 20864 48618
rect 20812 48554 20864 48560
rect 20628 48204 20680 48210
rect 20628 48146 20680 48152
rect 20536 43376 20588 43382
rect 20536 43318 20588 43324
rect 20548 40066 20576 43318
rect 20628 41608 20680 41614
rect 20680 41556 20760 41562
rect 20628 41550 20760 41556
rect 20640 41534 20760 41550
rect 20548 40038 20668 40066
rect 20536 39976 20588 39982
rect 20536 39918 20588 39924
rect 20548 37874 20576 39918
rect 20640 38978 20668 40038
rect 20732 39438 20760 41534
rect 20824 41138 20852 48554
rect 21284 46646 21312 49710
rect 21928 48142 21956 51200
rect 22572 49298 22600 51200
rect 22560 49292 22612 49298
rect 22560 49234 22612 49240
rect 22008 49224 22060 49230
rect 22008 49166 22060 49172
rect 22020 48754 22048 49166
rect 22192 49156 22244 49162
rect 22192 49098 22244 49104
rect 22008 48748 22060 48754
rect 22008 48690 22060 48696
rect 21916 48136 21968 48142
rect 21916 48078 21968 48084
rect 21640 48000 21692 48006
rect 21640 47942 21692 47948
rect 21272 46640 21324 46646
rect 21272 46582 21324 46588
rect 21364 42696 21416 42702
rect 21364 42638 21416 42644
rect 21376 41614 21404 42638
rect 21456 42152 21508 42158
rect 21456 42094 21508 42100
rect 21364 41608 21416 41614
rect 21364 41550 21416 41556
rect 20904 41540 20956 41546
rect 20904 41482 20956 41488
rect 20812 41132 20864 41138
rect 20812 41074 20864 41080
rect 20916 41002 20944 41482
rect 21180 41132 21232 41138
rect 21180 41074 21232 41080
rect 20904 40996 20956 41002
rect 20904 40938 20956 40944
rect 20720 39432 20772 39438
rect 20720 39374 20772 39380
rect 20640 38950 20760 38978
rect 20628 38888 20680 38894
rect 20628 38830 20680 38836
rect 20536 37868 20588 37874
rect 20536 37810 20588 37816
rect 20640 37754 20668 38830
rect 20548 37738 20668 37754
rect 20536 37732 20668 37738
rect 20588 37726 20668 37732
rect 20536 37674 20588 37680
rect 20548 36378 20576 37674
rect 20732 37618 20760 38950
rect 21192 37670 21220 41074
rect 21468 41070 21496 42094
rect 21652 41414 21680 47942
rect 22204 47802 22232 49098
rect 22928 48816 22980 48822
rect 22928 48758 22980 48764
rect 22192 47796 22244 47802
rect 22192 47738 22244 47744
rect 22008 47592 22060 47598
rect 21928 47552 22008 47580
rect 21732 47048 21784 47054
rect 21732 46990 21784 46996
rect 21744 46730 21772 46990
rect 21928 46918 21956 47552
rect 22008 47534 22060 47540
rect 22008 46980 22060 46986
rect 22940 46934 22968 48758
rect 23216 48618 23244 51200
rect 23860 49366 23888 51200
rect 23848 49360 23900 49366
rect 23848 49302 23900 49308
rect 24780 49298 24808 51326
rect 25134 51200 25190 52000
rect 25778 51200 25834 52000
rect 26422 51200 26478 52000
rect 27066 51354 27122 52000
rect 27066 51326 27568 51354
rect 27066 51200 27122 51326
rect 24768 49292 24820 49298
rect 24768 49234 24820 49240
rect 24400 49224 24452 49230
rect 24400 49166 24452 49172
rect 23480 49088 23532 49094
rect 23480 49030 23532 49036
rect 23204 48612 23256 48618
rect 23204 48554 23256 48560
rect 22008 46922 22060 46928
rect 21916 46912 21968 46918
rect 21916 46854 21968 46860
rect 22020 46730 22048 46922
rect 21744 46702 22048 46730
rect 22848 46906 22968 46934
rect 21744 42226 21772 46702
rect 22376 44940 22428 44946
rect 22376 44882 22428 44888
rect 22008 43308 22060 43314
rect 22060 43268 22140 43296
rect 22008 43250 22060 43256
rect 21824 42628 21876 42634
rect 21824 42570 21876 42576
rect 21836 42362 21864 42570
rect 22112 42362 22140 43268
rect 22284 43104 22336 43110
rect 22284 43046 22336 43052
rect 21824 42356 21876 42362
rect 21824 42298 21876 42304
rect 22100 42356 22152 42362
rect 22100 42298 22152 42304
rect 21732 42220 21784 42226
rect 21732 42162 21784 42168
rect 22008 41472 22060 41478
rect 22008 41414 22060 41420
rect 21652 41386 21772 41414
rect 21456 41064 21508 41070
rect 21456 41006 21508 41012
rect 21272 40112 21324 40118
rect 21272 40054 21324 40060
rect 21284 39574 21312 40054
rect 21272 39568 21324 39574
rect 21272 39510 21324 39516
rect 21284 38758 21312 39510
rect 21272 38752 21324 38758
rect 21272 38694 21324 38700
rect 21364 38276 21416 38282
rect 21364 38218 21416 38224
rect 21376 37874 21404 38218
rect 21364 37868 21416 37874
rect 21364 37810 21416 37816
rect 20640 37590 20760 37618
rect 21180 37664 21232 37670
rect 21180 37606 21232 37612
rect 20536 36372 20588 36378
rect 20536 36314 20588 36320
rect 20444 36236 20496 36242
rect 20444 36178 20496 36184
rect 20444 35692 20496 35698
rect 20444 35634 20496 35640
rect 20456 34610 20484 35634
rect 20640 35034 20668 37590
rect 20812 37120 20864 37126
rect 20812 37062 20864 37068
rect 20824 36718 20852 37062
rect 20812 36712 20864 36718
rect 20812 36654 20864 36660
rect 20812 36100 20864 36106
rect 20812 36042 20864 36048
rect 20824 35834 20852 36042
rect 20812 35828 20864 35834
rect 20812 35770 20864 35776
rect 20812 35488 20864 35494
rect 20812 35430 20864 35436
rect 20824 35290 20852 35430
rect 20812 35284 20864 35290
rect 20812 35226 20864 35232
rect 20548 35006 20668 35034
rect 20444 34604 20496 34610
rect 20444 34546 20496 34552
rect 20548 33318 20576 35006
rect 20628 34944 20680 34950
rect 20628 34886 20680 34892
rect 20640 34678 20668 34886
rect 20628 34672 20680 34678
rect 20628 34614 20680 34620
rect 20904 33924 20956 33930
rect 20904 33866 20956 33872
rect 20536 33312 20588 33318
rect 20536 33254 20588 33260
rect 20628 32768 20680 32774
rect 20628 32710 20680 32716
rect 20640 32502 20668 32710
rect 20628 32496 20680 32502
rect 20628 32438 20680 32444
rect 20916 32230 20944 33866
rect 20904 32224 20956 32230
rect 20904 32166 20956 32172
rect 20812 31340 20864 31346
rect 20812 31282 20864 31288
rect 20352 31272 20404 31278
rect 20352 31214 20404 31220
rect 20364 30734 20392 31214
rect 20352 30728 20404 30734
rect 20352 30670 20404 30676
rect 20824 30666 20852 31282
rect 20916 31142 20944 32166
rect 21088 31340 21140 31346
rect 21088 31282 21140 31288
rect 20904 31136 20956 31142
rect 20904 31078 20956 31084
rect 21100 30938 21128 31282
rect 21088 30932 21140 30938
rect 21088 30874 21140 30880
rect 20536 30660 20588 30666
rect 20536 30602 20588 30608
rect 20720 30660 20772 30666
rect 20720 30602 20772 30608
rect 20812 30660 20864 30666
rect 20812 30602 20864 30608
rect 20548 30122 20576 30602
rect 20536 30116 20588 30122
rect 20536 30058 20588 30064
rect 20628 30048 20680 30054
rect 20628 29990 20680 29996
rect 20352 29844 20404 29850
rect 20352 29786 20404 29792
rect 20364 29170 20392 29786
rect 20352 29164 20404 29170
rect 20352 29106 20404 29112
rect 20352 28960 20404 28966
rect 20352 28902 20404 28908
rect 20364 28490 20392 28902
rect 20352 28484 20404 28490
rect 20352 28426 20404 28432
rect 20260 27940 20312 27946
rect 20260 27882 20312 27888
rect 20168 27464 20220 27470
rect 20168 27406 20220 27412
rect 20180 26994 20208 27406
rect 20536 27056 20588 27062
rect 20536 26998 20588 27004
rect 20168 26988 20220 26994
rect 20168 26930 20220 26936
rect 20076 26376 20128 26382
rect 20076 26318 20128 26324
rect 20180 26042 20208 26930
rect 20260 26852 20312 26858
rect 20260 26794 20312 26800
rect 20168 26036 20220 26042
rect 20168 25978 20220 25984
rect 19984 25832 20036 25838
rect 19984 25774 20036 25780
rect 20168 25764 20220 25770
rect 20168 25706 20220 25712
rect 19432 25356 19484 25362
rect 19432 25298 19484 25304
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19984 24200 20036 24206
rect 19984 24142 20036 24148
rect 19432 24132 19484 24138
rect 19432 24074 19484 24080
rect 19444 23254 19472 24074
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 19524 23520 19576 23526
rect 19524 23462 19576 23468
rect 19432 23248 19484 23254
rect 19432 23190 19484 23196
rect 19536 23066 19564 23462
rect 19444 23050 19564 23066
rect 19156 23044 19208 23050
rect 19156 22986 19208 22992
rect 19340 23044 19392 23050
rect 19340 22986 19392 22992
rect 19432 23044 19564 23050
rect 19484 23038 19564 23044
rect 19432 22986 19484 22992
rect 19352 21962 19380 22986
rect 19444 22506 19472 22986
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19892 22636 19944 22642
rect 19892 22578 19944 22584
rect 19904 22545 19932 22578
rect 19890 22536 19946 22545
rect 19432 22500 19484 22506
rect 19890 22471 19946 22480
rect 19432 22442 19484 22448
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 19340 21956 19392 21962
rect 19340 21898 19392 21904
rect 19352 21690 19380 21898
rect 19340 21684 19392 21690
rect 19340 21626 19392 21632
rect 19444 20618 19472 21966
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19260 20590 19472 20618
rect 19260 20466 19288 20590
rect 19340 20528 19392 20534
rect 19340 20470 19392 20476
rect 19248 20460 19300 20466
rect 19248 20402 19300 20408
rect 19352 19854 19380 20470
rect 19616 20460 19668 20466
rect 19616 20402 19668 20408
rect 19432 20392 19484 20398
rect 19432 20334 19484 20340
rect 19340 19848 19392 19854
rect 19340 19790 19392 19796
rect 19156 19712 19208 19718
rect 19156 19654 19208 19660
rect 19064 16448 19116 16454
rect 19064 16390 19116 16396
rect 19076 16250 19104 16390
rect 19064 16244 19116 16250
rect 19064 16186 19116 16192
rect 19168 14498 19196 19654
rect 19352 19446 19380 19790
rect 19340 19440 19392 19446
rect 19340 19382 19392 19388
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 19352 18630 19380 19246
rect 19444 19174 19472 20334
rect 19628 20058 19656 20402
rect 19616 20052 19668 20058
rect 19616 19994 19668 20000
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19798 19408 19854 19417
rect 19798 19343 19854 19352
rect 19812 19174 19840 19343
rect 19432 19168 19484 19174
rect 19432 19110 19484 19116
rect 19800 19168 19852 19174
rect 19800 19110 19852 19116
rect 19812 18766 19840 19110
rect 19996 18902 20024 24142
rect 20076 22568 20128 22574
rect 20076 22510 20128 22516
rect 20088 22166 20116 22510
rect 20076 22160 20128 22166
rect 20076 22102 20128 22108
rect 20180 21554 20208 25706
rect 20272 24206 20300 26794
rect 20548 26518 20576 26998
rect 20536 26512 20588 26518
rect 20536 26454 20588 26460
rect 20444 25832 20496 25838
rect 20444 25774 20496 25780
rect 20352 25696 20404 25702
rect 20352 25638 20404 25644
rect 20364 25362 20392 25638
rect 20352 25356 20404 25362
rect 20352 25298 20404 25304
rect 20260 24200 20312 24206
rect 20260 24142 20312 24148
rect 20352 24132 20404 24138
rect 20352 24074 20404 24080
rect 20260 23860 20312 23866
rect 20260 23802 20312 23808
rect 20168 21548 20220 21554
rect 20168 21490 20220 21496
rect 20180 20942 20208 21490
rect 20168 20936 20220 20942
rect 20168 20878 20220 20884
rect 19984 18896 20036 18902
rect 19984 18838 20036 18844
rect 19800 18760 19852 18766
rect 19852 18720 20024 18748
rect 19800 18702 19852 18708
rect 19340 18624 19392 18630
rect 19340 18566 19392 18572
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19996 18290 20024 18720
rect 20168 18624 20220 18630
rect 20168 18566 20220 18572
rect 20180 18290 20208 18566
rect 19984 18284 20036 18290
rect 19984 18226 20036 18232
rect 20168 18284 20220 18290
rect 20168 18226 20220 18232
rect 20168 18080 20220 18086
rect 20168 18022 20220 18028
rect 19340 17672 19392 17678
rect 19340 17614 19392 17620
rect 19248 16652 19300 16658
rect 19352 16640 19380 17614
rect 20076 17604 20128 17610
rect 20076 17546 20128 17552
rect 19432 17536 19484 17542
rect 19432 17478 19484 17484
rect 19984 17536 20036 17542
rect 19984 17478 20036 17484
rect 19444 16794 19472 17478
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19890 17232 19946 17241
rect 19890 17167 19946 17176
rect 19904 17134 19932 17167
rect 19892 17128 19944 17134
rect 19892 17070 19944 17076
rect 19432 16788 19484 16794
rect 19432 16730 19484 16736
rect 19300 16612 19472 16640
rect 19248 16594 19300 16600
rect 19340 16516 19392 16522
rect 19340 16458 19392 16464
rect 19352 14618 19380 16458
rect 19444 15026 19472 16612
rect 19904 16522 19932 17070
rect 19892 16516 19944 16522
rect 19892 16458 19944 16464
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19996 16182 20024 17478
rect 20088 17066 20116 17546
rect 20076 17060 20128 17066
rect 20076 17002 20128 17008
rect 20076 16516 20128 16522
rect 20076 16458 20128 16464
rect 20088 16250 20116 16458
rect 20076 16244 20128 16250
rect 20076 16186 20128 16192
rect 19984 16176 20036 16182
rect 19984 16118 20036 16124
rect 19524 16108 19576 16114
rect 19524 16050 19576 16056
rect 19536 15502 19564 16050
rect 20076 16040 20128 16046
rect 20076 15982 20128 15988
rect 19524 15496 19576 15502
rect 19524 15438 19576 15444
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19432 15020 19484 15026
rect 19432 14962 19484 14968
rect 19892 15020 19944 15026
rect 19892 14962 19944 14968
rect 19984 15020 20036 15026
rect 19984 14962 20036 14968
rect 19340 14612 19392 14618
rect 19340 14554 19392 14560
rect 19168 14470 19380 14498
rect 19904 14482 19932 14962
rect 19996 14550 20024 14962
rect 19984 14544 20036 14550
rect 19984 14486 20036 14492
rect 19352 13138 19380 14470
rect 19892 14476 19944 14482
rect 19892 14418 19944 14424
rect 19904 14362 19932 14418
rect 19904 14334 20024 14362
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 19260 13110 19380 13138
rect 19156 12776 19208 12782
rect 19156 12718 19208 12724
rect 19168 12170 19196 12718
rect 19260 12646 19288 13110
rect 19340 12980 19392 12986
rect 19340 12922 19392 12928
rect 19248 12640 19300 12646
rect 19248 12582 19300 12588
rect 19156 12164 19208 12170
rect 19156 12106 19208 12112
rect 19168 11234 19196 12106
rect 19248 11756 19300 11762
rect 19248 11698 19300 11704
rect 19260 11354 19288 11698
rect 19248 11348 19300 11354
rect 19248 11290 19300 11296
rect 19168 11206 19288 11234
rect 19064 10668 19116 10674
rect 19064 10610 19116 10616
rect 19076 10470 19104 10610
rect 19064 10464 19116 10470
rect 19064 10406 19116 10412
rect 18972 8084 19024 8090
rect 18972 8026 19024 8032
rect 19076 7818 19104 10406
rect 19260 9994 19288 11206
rect 19352 10674 19380 12922
rect 19444 12434 19472 13806
rect 19708 13728 19760 13734
rect 19708 13670 19760 13676
rect 19720 13326 19748 13670
rect 19708 13320 19760 13326
rect 19708 13262 19760 13268
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 19996 12986 20024 14334
rect 20088 13734 20116 15982
rect 20076 13728 20128 13734
rect 20076 13670 20128 13676
rect 19984 12980 20036 12986
rect 19984 12922 20036 12928
rect 20076 12640 20128 12646
rect 20180 12617 20208 18022
rect 20272 13297 20300 23802
rect 20364 21962 20392 24074
rect 20352 21956 20404 21962
rect 20352 21898 20404 21904
rect 20364 21690 20392 21898
rect 20352 21684 20404 21690
rect 20352 21626 20404 21632
rect 20352 21344 20404 21350
rect 20352 21286 20404 21292
rect 20364 20534 20392 21286
rect 20352 20528 20404 20534
rect 20352 20470 20404 20476
rect 20352 18760 20404 18766
rect 20352 18702 20404 18708
rect 20364 17202 20392 18702
rect 20352 17196 20404 17202
rect 20352 17138 20404 17144
rect 20364 16114 20392 17138
rect 20352 16108 20404 16114
rect 20352 16050 20404 16056
rect 20364 15706 20392 16050
rect 20352 15700 20404 15706
rect 20352 15642 20404 15648
rect 20364 14414 20392 15642
rect 20352 14408 20404 14414
rect 20352 14350 20404 14356
rect 20258 13288 20314 13297
rect 20258 13223 20314 13232
rect 20260 13184 20312 13190
rect 20260 13126 20312 13132
rect 20076 12582 20128 12588
rect 20166 12608 20222 12617
rect 19444 12406 19564 12434
rect 19536 12170 19564 12406
rect 20088 12322 20116 12582
rect 20166 12543 20222 12552
rect 20088 12294 20208 12322
rect 20272 12306 20300 13126
rect 20350 12608 20406 12617
rect 20350 12543 20406 12552
rect 20076 12232 20128 12238
rect 20076 12174 20128 12180
rect 19524 12164 19576 12170
rect 19524 12106 19576 12112
rect 19984 12096 20036 12102
rect 19984 12038 20036 12044
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19892 11756 19944 11762
rect 19892 11698 19944 11704
rect 19430 11112 19486 11121
rect 19430 11047 19432 11056
rect 19484 11047 19486 11056
rect 19432 11018 19484 11024
rect 19904 10996 19932 11698
rect 19996 11218 20024 12038
rect 20088 11898 20116 12174
rect 20076 11892 20128 11898
rect 20076 11834 20128 11840
rect 19984 11212 20036 11218
rect 19984 11154 20036 11160
rect 20076 11212 20128 11218
rect 20076 11154 20128 11160
rect 19904 10968 20024 10996
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19340 10668 19392 10674
rect 19340 10610 19392 10616
rect 19352 10130 19380 10610
rect 19430 10432 19486 10441
rect 19430 10367 19486 10376
rect 19340 10124 19392 10130
rect 19340 10066 19392 10072
rect 19248 9988 19300 9994
rect 19248 9930 19300 9936
rect 19260 7886 19288 9930
rect 19352 8498 19380 10066
rect 19340 8492 19392 8498
rect 19340 8434 19392 8440
rect 19248 7880 19300 7886
rect 19248 7822 19300 7828
rect 18788 7812 18840 7818
rect 18788 7754 18840 7760
rect 19064 7812 19116 7818
rect 19064 7754 19116 7760
rect 18800 7274 18828 7754
rect 19352 7478 19380 8434
rect 19444 7546 19472 10367
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19616 8288 19668 8294
rect 19616 8230 19668 8236
rect 19628 8090 19656 8230
rect 19616 8084 19668 8090
rect 19616 8026 19668 8032
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19432 7540 19484 7546
rect 19432 7482 19484 7488
rect 19340 7472 19392 7478
rect 19340 7414 19392 7420
rect 18788 7268 18840 7274
rect 18788 7210 18840 7216
rect 19352 6866 19380 7414
rect 19340 6860 19392 6866
rect 19340 6802 19392 6808
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19432 6180 19484 6186
rect 19432 6122 19484 6128
rect 19340 5568 19392 5574
rect 19340 5510 19392 5516
rect 19352 5302 19380 5510
rect 19340 5296 19392 5302
rect 19340 5238 19392 5244
rect 18696 5160 18748 5166
rect 18696 5102 18748 5108
rect 18788 5160 18840 5166
rect 18788 5102 18840 5108
rect 18144 4480 18196 4486
rect 18144 4422 18196 4428
rect 18156 3126 18184 4422
rect 18696 4140 18748 4146
rect 18696 4082 18748 4088
rect 18144 3120 18196 3126
rect 18144 3062 18196 3068
rect 17880 2910 18092 2938
rect 18144 2984 18196 2990
rect 18144 2926 18196 2932
rect 16580 2848 16632 2854
rect 16580 2790 16632 2796
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 17420 800 17448 2382
rect 17684 2304 17736 2310
rect 17684 2246 17736 2252
rect 17696 1902 17724 2246
rect 17684 1896 17736 1902
rect 17684 1838 17736 1844
rect 18156 1578 18184 2926
rect 18064 1550 18184 1578
rect 18064 800 18092 1550
rect 18708 800 18736 4082
rect 18800 3466 18828 5102
rect 19340 4276 19392 4282
rect 19340 4218 19392 4224
rect 19352 4078 19380 4218
rect 19444 4146 19472 6122
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 19432 4140 19484 4146
rect 19432 4082 19484 4088
rect 19340 4072 19392 4078
rect 19340 4014 19392 4020
rect 19996 3942 20024 10968
rect 20088 5710 20116 11154
rect 20180 11150 20208 12294
rect 20260 12300 20312 12306
rect 20260 12242 20312 12248
rect 20260 12164 20312 12170
rect 20260 12106 20312 12112
rect 20168 11144 20220 11150
rect 20168 11086 20220 11092
rect 20272 10826 20300 12106
rect 20180 10798 20300 10826
rect 20076 5704 20128 5710
rect 20076 5646 20128 5652
rect 20088 4622 20116 5646
rect 20180 4758 20208 10798
rect 20364 7954 20392 12543
rect 20456 11218 20484 25774
rect 20548 18086 20576 26454
rect 20640 25226 20668 29990
rect 20732 29646 20760 30602
rect 20904 29844 20956 29850
rect 20904 29786 20956 29792
rect 20916 29646 20944 29786
rect 20720 29640 20772 29646
rect 20720 29582 20772 29588
rect 20904 29640 20956 29646
rect 20904 29582 20956 29588
rect 20812 29504 20864 29510
rect 20812 29446 20864 29452
rect 20824 29170 20852 29446
rect 20812 29164 20864 29170
rect 20812 29106 20864 29112
rect 20916 28762 20944 29582
rect 20996 29164 21048 29170
rect 20996 29106 21048 29112
rect 20904 28756 20956 28762
rect 20904 28698 20956 28704
rect 21008 28150 21036 29106
rect 21192 29034 21220 37606
rect 21376 37194 21404 37810
rect 21364 37188 21416 37194
rect 21364 37130 21416 37136
rect 21272 34400 21324 34406
rect 21272 34342 21324 34348
rect 21284 34066 21312 34342
rect 21272 34060 21324 34066
rect 21272 34002 21324 34008
rect 21270 31784 21326 31793
rect 21270 31719 21326 31728
rect 21284 31686 21312 31719
rect 21272 31680 21324 31686
rect 21272 31622 21324 31628
rect 21284 31346 21312 31622
rect 21272 31340 21324 31346
rect 21272 31282 21324 31288
rect 21272 30660 21324 30666
rect 21272 30602 21324 30608
rect 21180 29028 21232 29034
rect 21180 28970 21232 28976
rect 20996 28144 21048 28150
rect 20996 28086 21048 28092
rect 20812 27396 20864 27402
rect 20812 27338 20864 27344
rect 20628 25220 20680 25226
rect 20628 25162 20680 25168
rect 20628 24676 20680 24682
rect 20628 24618 20680 24624
rect 20640 24138 20668 24618
rect 20628 24132 20680 24138
rect 20628 24074 20680 24080
rect 20640 22982 20668 24074
rect 20824 23866 20852 27338
rect 21180 24064 21232 24070
rect 21180 24006 21232 24012
rect 20812 23860 20864 23866
rect 20812 23802 20864 23808
rect 21192 23662 21220 24006
rect 21284 23882 21312 30602
rect 21376 30258 21404 37130
rect 21468 36122 21496 41006
rect 21548 37392 21600 37398
rect 21548 37334 21600 37340
rect 21560 37126 21588 37334
rect 21548 37120 21600 37126
rect 21548 37062 21600 37068
rect 21560 36310 21588 37062
rect 21548 36304 21600 36310
rect 21548 36246 21600 36252
rect 21468 36094 21588 36122
rect 21456 35692 21508 35698
rect 21456 35634 21508 35640
rect 21468 35154 21496 35634
rect 21560 35494 21588 36094
rect 21640 36100 21692 36106
rect 21640 36042 21692 36048
rect 21548 35488 21600 35494
rect 21548 35430 21600 35436
rect 21456 35148 21508 35154
rect 21456 35090 21508 35096
rect 21652 35086 21680 36042
rect 21640 35080 21692 35086
rect 21640 35022 21692 35028
rect 21744 33998 21772 41386
rect 22020 41138 22048 41414
rect 22008 41132 22060 41138
rect 22008 41074 22060 41080
rect 22112 40934 22140 42298
rect 22296 42226 22324 43046
rect 22284 42220 22336 42226
rect 22284 42162 22336 42168
rect 22100 40928 22152 40934
rect 22100 40870 22152 40876
rect 22008 40044 22060 40050
rect 22008 39986 22060 39992
rect 21824 39432 21876 39438
rect 21824 39374 21876 39380
rect 21836 38894 21864 39374
rect 21916 38956 21968 38962
rect 22020 38944 22048 39986
rect 22192 39296 22244 39302
rect 22192 39238 22244 39244
rect 21968 38916 22048 38944
rect 21916 38898 21968 38904
rect 21824 38888 21876 38894
rect 21824 38830 21876 38836
rect 21836 38350 21864 38830
rect 21824 38344 21876 38350
rect 21824 38286 21876 38292
rect 21916 38344 21968 38350
rect 21916 38286 21968 38292
rect 21836 37262 21864 38286
rect 21928 37466 21956 38286
rect 22020 38010 22048 38916
rect 22100 38956 22152 38962
rect 22100 38898 22152 38904
rect 22112 38554 22140 38898
rect 22100 38548 22152 38554
rect 22100 38490 22152 38496
rect 22204 38350 22232 39238
rect 22192 38344 22244 38350
rect 22192 38286 22244 38292
rect 22008 38004 22060 38010
rect 22008 37946 22060 37952
rect 21916 37460 21968 37466
rect 21916 37402 21968 37408
rect 21824 37256 21876 37262
rect 21824 37198 21876 37204
rect 21836 36718 21864 37198
rect 21824 36712 21876 36718
rect 21824 36654 21876 36660
rect 21836 34542 21864 36654
rect 21916 36032 21968 36038
rect 21916 35974 21968 35980
rect 21824 34536 21876 34542
rect 21824 34478 21876 34484
rect 21732 33992 21784 33998
rect 21732 33934 21784 33940
rect 21548 32496 21600 32502
rect 21732 32496 21784 32502
rect 21600 32444 21732 32450
rect 21548 32438 21784 32444
rect 21560 32422 21772 32438
rect 21836 31890 21864 34478
rect 21928 34134 21956 35974
rect 22008 35488 22060 35494
rect 22008 35430 22060 35436
rect 21916 34128 21968 34134
rect 21916 34070 21968 34076
rect 21916 32428 21968 32434
rect 21916 32370 21968 32376
rect 21824 31884 21876 31890
rect 21824 31826 21876 31832
rect 21928 31822 21956 32370
rect 21916 31816 21968 31822
rect 21916 31758 21968 31764
rect 21456 31680 21508 31686
rect 21456 31622 21508 31628
rect 21468 31210 21496 31622
rect 21548 31476 21600 31482
rect 21548 31418 21600 31424
rect 21456 31204 21508 31210
rect 21456 31146 21508 31152
rect 21468 30870 21496 31146
rect 21456 30864 21508 30870
rect 21456 30806 21508 30812
rect 21364 30252 21416 30258
rect 21364 30194 21416 30200
rect 21468 28966 21496 30806
rect 21560 30666 21588 31418
rect 21824 31136 21876 31142
rect 21824 31078 21876 31084
rect 21548 30660 21600 30666
rect 21548 30602 21600 30608
rect 21456 28960 21508 28966
rect 21456 28902 21508 28908
rect 21836 28626 21864 31078
rect 22020 30054 22048 35430
rect 22284 34740 22336 34746
rect 22284 34682 22336 34688
rect 22100 34604 22152 34610
rect 22100 34546 22152 34552
rect 22112 34202 22140 34546
rect 22100 34196 22152 34202
rect 22100 34138 22152 34144
rect 22192 34196 22244 34202
rect 22192 34138 22244 34144
rect 22008 30048 22060 30054
rect 22008 29990 22060 29996
rect 22008 29708 22060 29714
rect 22008 29650 22060 29656
rect 22020 29170 22048 29650
rect 22204 29232 22232 34138
rect 22296 34066 22324 34682
rect 22284 34060 22336 34066
rect 22284 34002 22336 34008
rect 22296 33590 22324 34002
rect 22284 33584 22336 33590
rect 22284 33526 22336 33532
rect 22388 32298 22416 44882
rect 22744 43308 22796 43314
rect 22744 43250 22796 43256
rect 22756 42566 22784 43250
rect 22744 42560 22796 42566
rect 22744 42502 22796 42508
rect 22756 42090 22784 42502
rect 22744 42084 22796 42090
rect 22744 42026 22796 42032
rect 22744 41540 22796 41546
rect 22744 41482 22796 41488
rect 22756 41274 22784 41482
rect 22744 41268 22796 41274
rect 22744 41210 22796 41216
rect 22848 41138 22876 46906
rect 23388 42628 23440 42634
rect 23388 42570 23440 42576
rect 23400 42362 23428 42570
rect 23388 42356 23440 42362
rect 23388 42298 23440 42304
rect 23204 41472 23256 41478
rect 23204 41414 23256 41420
rect 22836 41132 22888 41138
rect 22836 41074 22888 41080
rect 23017 41135 23069 41141
rect 23069 41092 23152 41120
rect 23017 41077 23069 41083
rect 23124 40934 23152 41092
rect 23216 41070 23244 41414
rect 23296 41132 23348 41138
rect 23296 41074 23348 41080
rect 23204 41064 23256 41070
rect 23204 41006 23256 41012
rect 23308 41002 23336 41074
rect 23296 40996 23348 41002
rect 23296 40938 23348 40944
rect 22468 40928 22520 40934
rect 22468 40870 22520 40876
rect 23112 40928 23164 40934
rect 23112 40870 23164 40876
rect 22480 39438 22508 40870
rect 22468 39432 22520 39438
rect 22468 39374 22520 39380
rect 22480 38554 22508 39374
rect 22468 38548 22520 38554
rect 22468 38490 22520 38496
rect 23020 38480 23072 38486
rect 23020 38422 23072 38428
rect 23032 38282 23060 38422
rect 23020 38276 23072 38282
rect 23020 38218 23072 38224
rect 23032 37754 23060 38218
rect 22848 37726 23060 37754
rect 22652 37188 22704 37194
rect 22652 37130 22704 37136
rect 22664 36854 22692 37130
rect 22652 36848 22704 36854
rect 22652 36790 22704 36796
rect 22468 36780 22520 36786
rect 22468 36722 22520 36728
rect 22480 36378 22508 36722
rect 22468 36372 22520 36378
rect 22468 36314 22520 36320
rect 22744 36372 22796 36378
rect 22744 36314 22796 36320
rect 22756 36174 22784 36314
rect 22744 36168 22796 36174
rect 22744 36110 22796 36116
rect 22848 35562 22876 37726
rect 22928 37120 22980 37126
rect 22928 37062 22980 37068
rect 22940 36174 22968 37062
rect 23020 36304 23072 36310
rect 23020 36246 23072 36252
rect 22928 36168 22980 36174
rect 22928 36110 22980 36116
rect 23032 36106 23060 36246
rect 23020 36100 23072 36106
rect 23020 36042 23072 36048
rect 23124 35894 23152 40870
rect 23308 40730 23336 40938
rect 23296 40724 23348 40730
rect 23296 40666 23348 40672
rect 23388 40452 23440 40458
rect 23388 40394 23440 40400
rect 23204 40044 23256 40050
rect 23204 39986 23256 39992
rect 23216 39642 23244 39986
rect 23296 39976 23348 39982
rect 23296 39918 23348 39924
rect 23308 39642 23336 39918
rect 23204 39636 23256 39642
rect 23204 39578 23256 39584
rect 23296 39636 23348 39642
rect 23296 39578 23348 39584
rect 23400 38962 23428 40394
rect 23492 39438 23520 49030
rect 23664 48680 23716 48686
rect 23664 48622 23716 48628
rect 23676 48278 23704 48622
rect 23664 48272 23716 48278
rect 23664 48214 23716 48220
rect 23848 48136 23900 48142
rect 23848 48078 23900 48084
rect 23756 45484 23808 45490
rect 23756 45426 23808 45432
rect 23768 44810 23796 45426
rect 23756 44804 23808 44810
rect 23756 44746 23808 44752
rect 23768 44402 23796 44746
rect 23756 44396 23808 44402
rect 23756 44338 23808 44344
rect 23768 43790 23796 44338
rect 23860 44334 23888 48078
rect 24216 47660 24268 47666
rect 24216 47602 24268 47608
rect 24124 45416 24176 45422
rect 24124 45358 24176 45364
rect 23848 44328 23900 44334
rect 23848 44270 23900 44276
rect 23756 43784 23808 43790
rect 23756 43726 23808 43732
rect 23572 43716 23624 43722
rect 23572 43658 23624 43664
rect 23480 39432 23532 39438
rect 23480 39374 23532 39380
rect 23480 39296 23532 39302
rect 23480 39238 23532 39244
rect 23388 38956 23440 38962
rect 23388 38898 23440 38904
rect 23296 37188 23348 37194
rect 23296 37130 23348 37136
rect 23308 36582 23336 37130
rect 23204 36576 23256 36582
rect 23204 36518 23256 36524
rect 23296 36576 23348 36582
rect 23296 36518 23348 36524
rect 23216 36310 23244 36518
rect 23296 36372 23348 36378
rect 23296 36314 23348 36320
rect 23204 36304 23256 36310
rect 23204 36246 23256 36252
rect 23032 35866 23152 35894
rect 22836 35556 22888 35562
rect 22836 35498 22888 35504
rect 22560 35080 22612 35086
rect 22560 35022 22612 35028
rect 22572 33998 22600 35022
rect 22652 35012 22704 35018
rect 22652 34954 22704 34960
rect 22560 33992 22612 33998
rect 22560 33934 22612 33940
rect 22572 32434 22600 33934
rect 22664 33862 22692 34954
rect 23032 34202 23060 35866
rect 23204 34944 23256 34950
rect 23204 34886 23256 34892
rect 23216 34746 23244 34886
rect 23204 34740 23256 34746
rect 23204 34682 23256 34688
rect 23112 34400 23164 34406
rect 23112 34342 23164 34348
rect 23020 34196 23072 34202
rect 23020 34138 23072 34144
rect 23124 33998 23152 34342
rect 23112 33992 23164 33998
rect 23112 33934 23164 33940
rect 22652 33856 22704 33862
rect 22652 33798 22704 33804
rect 23124 33658 23152 33934
rect 23112 33652 23164 33658
rect 23112 33594 23164 33600
rect 23112 33516 23164 33522
rect 23112 33458 23164 33464
rect 22652 32564 22704 32570
rect 22652 32506 22704 32512
rect 23020 32564 23072 32570
rect 23020 32506 23072 32512
rect 22560 32428 22612 32434
rect 22560 32370 22612 32376
rect 22468 32360 22520 32366
rect 22468 32302 22520 32308
rect 22376 32292 22428 32298
rect 22376 32234 22428 32240
rect 22480 31686 22508 32302
rect 22560 31810 22612 31816
rect 22560 31752 22612 31758
rect 22376 31680 22428 31686
rect 22376 31622 22428 31628
rect 22468 31680 22520 31686
rect 22468 31622 22520 31628
rect 22201 29173 22232 29232
rect 22008 29164 22060 29170
rect 22008 29106 22060 29112
rect 22189 29167 22241 29173
rect 22189 29109 22241 29115
rect 22284 29164 22336 29170
rect 22100 29028 22152 29034
rect 22100 28970 22152 28976
rect 21824 28620 21876 28626
rect 21824 28562 21876 28568
rect 21836 27538 21864 28562
rect 22112 28558 22140 28970
rect 22100 28552 22152 28558
rect 22100 28494 22152 28500
rect 22204 28082 22232 29109
rect 22284 29106 22336 29112
rect 22296 28218 22324 29106
rect 22284 28212 22336 28218
rect 22284 28154 22336 28160
rect 22192 28076 22244 28082
rect 22192 28018 22244 28024
rect 22284 28076 22336 28082
rect 22284 28018 22336 28024
rect 22100 27872 22152 27878
rect 22100 27814 22152 27820
rect 21824 27532 21876 27538
rect 21824 27474 21876 27480
rect 22112 27402 22140 27814
rect 22100 27396 22152 27402
rect 22100 27338 22152 27344
rect 22296 27130 22324 28018
rect 22284 27124 22336 27130
rect 22284 27066 22336 27072
rect 22284 26240 22336 26246
rect 22388 26234 22416 31622
rect 22572 30938 22600 31752
rect 22560 30932 22612 30938
rect 22560 30874 22612 30880
rect 22664 30734 22692 32506
rect 23032 32434 23060 32506
rect 23020 32428 23072 32434
rect 23020 32370 23072 32376
rect 22836 32360 22888 32366
rect 22836 32302 22888 32308
rect 22744 31816 22796 31822
rect 22742 31784 22744 31793
rect 22796 31784 22798 31793
rect 22848 31754 22876 32302
rect 22928 31952 22980 31958
rect 22928 31894 22980 31900
rect 22742 31719 22798 31728
rect 22836 31748 22888 31754
rect 22756 31686 22784 31719
rect 22836 31690 22888 31696
rect 22744 31680 22796 31686
rect 22744 31622 22796 31628
rect 22756 30734 22784 31622
rect 22940 31346 22968 31894
rect 22928 31340 22980 31346
rect 22928 31282 22980 31288
rect 23124 30802 23152 33458
rect 23202 32600 23258 32609
rect 23202 32535 23258 32544
rect 23216 32434 23244 32535
rect 23204 32428 23256 32434
rect 23204 32370 23256 32376
rect 23112 30796 23164 30802
rect 23112 30738 23164 30744
rect 22652 30728 22704 30734
rect 22652 30670 22704 30676
rect 22744 30728 22796 30734
rect 22744 30670 22796 30676
rect 23124 30326 23152 30738
rect 23112 30320 23164 30326
rect 23112 30262 23164 30268
rect 23124 29714 23152 30262
rect 23112 29708 23164 29714
rect 23112 29650 23164 29656
rect 22928 29504 22980 29510
rect 22928 29446 22980 29452
rect 22940 29170 22968 29446
rect 22560 29164 22612 29170
rect 22560 29106 22612 29112
rect 22928 29164 22980 29170
rect 22928 29106 22980 29112
rect 22572 28150 22600 29106
rect 22560 28144 22612 28150
rect 22560 28086 22612 28092
rect 22940 28082 22968 29106
rect 22928 28076 22980 28082
rect 22928 28018 22980 28024
rect 22836 28008 22888 28014
rect 22836 27950 22888 27956
rect 22388 26206 22600 26234
rect 22284 26182 22336 26188
rect 21824 26036 21876 26042
rect 21824 25978 21876 25984
rect 21548 25356 21600 25362
rect 21548 25298 21600 25304
rect 21284 23854 21404 23882
rect 21272 23724 21324 23730
rect 21272 23666 21324 23672
rect 21180 23656 21232 23662
rect 21180 23598 21232 23604
rect 20904 23588 20956 23594
rect 20904 23530 20956 23536
rect 20720 23520 20772 23526
rect 20720 23462 20772 23468
rect 20732 23050 20760 23462
rect 20720 23044 20772 23050
rect 20720 22986 20772 22992
rect 20812 23044 20864 23050
rect 20812 22986 20864 22992
rect 20628 22976 20680 22982
rect 20628 22918 20680 22924
rect 20824 22794 20852 22986
rect 20732 22766 20852 22794
rect 20732 22710 20760 22766
rect 20720 22704 20772 22710
rect 20720 22646 20772 22652
rect 20916 22506 20944 23530
rect 21284 22794 21312 23666
rect 21008 22766 21312 22794
rect 20904 22500 20956 22506
rect 20904 22442 20956 22448
rect 20812 22432 20864 22438
rect 20810 22400 20812 22409
rect 20864 22400 20866 22409
rect 20810 22335 20866 22344
rect 21008 22094 21036 22766
rect 21284 22642 21312 22766
rect 21088 22636 21140 22642
rect 21088 22578 21140 22584
rect 21272 22636 21324 22642
rect 21272 22578 21324 22584
rect 21100 22234 21128 22578
rect 21088 22228 21140 22234
rect 21088 22170 21140 22176
rect 21376 22094 21404 23854
rect 20916 22066 21036 22094
rect 21192 22066 21404 22094
rect 20628 22024 20680 22030
rect 20628 21966 20680 21972
rect 20640 21842 20668 21966
rect 20640 21814 20760 21842
rect 20628 21684 20680 21690
rect 20628 21626 20680 21632
rect 20640 21146 20668 21626
rect 20732 21350 20760 21814
rect 20812 21480 20864 21486
rect 20812 21422 20864 21428
rect 20720 21344 20772 21350
rect 20720 21286 20772 21292
rect 20628 21140 20680 21146
rect 20628 21082 20680 21088
rect 20732 21026 20760 21286
rect 20824 21146 20852 21422
rect 20812 21140 20864 21146
rect 20812 21082 20864 21088
rect 20640 20998 20760 21026
rect 20640 18986 20668 20998
rect 20812 19712 20864 19718
rect 20812 19654 20864 19660
rect 20824 19446 20852 19654
rect 20812 19440 20864 19446
rect 20812 19382 20864 19388
rect 20640 18958 20760 18986
rect 20824 18970 20852 19382
rect 20628 18896 20680 18902
rect 20628 18838 20680 18844
rect 20536 18080 20588 18086
rect 20536 18022 20588 18028
rect 20640 17082 20668 18838
rect 20548 17054 20668 17082
rect 20548 11898 20576 17054
rect 20732 16946 20760 18958
rect 20812 18964 20864 18970
rect 20812 18906 20864 18912
rect 20812 18624 20864 18630
rect 20812 18566 20864 18572
rect 20824 17610 20852 18566
rect 20812 17604 20864 17610
rect 20812 17546 20864 17552
rect 20824 17270 20852 17546
rect 20812 17264 20864 17270
rect 20812 17206 20864 17212
rect 20812 17060 20864 17066
rect 20812 17002 20864 17008
rect 20640 16918 20760 16946
rect 20640 13938 20668 16918
rect 20824 16794 20852 17002
rect 20812 16788 20864 16794
rect 20812 16730 20864 16736
rect 20916 16250 20944 22066
rect 20996 22024 21048 22030
rect 20996 21966 21048 21972
rect 21008 20942 21036 21966
rect 20996 20936 21048 20942
rect 20996 20878 21048 20884
rect 21008 20806 21036 20878
rect 20996 20800 21048 20806
rect 20996 20742 21048 20748
rect 21088 20256 21140 20262
rect 21088 20198 21140 20204
rect 21100 19786 21128 20198
rect 21088 19780 21140 19786
rect 21088 19722 21140 19728
rect 20996 19712 21048 19718
rect 20996 19654 21048 19660
rect 21008 19514 21036 19654
rect 20996 19508 21048 19514
rect 20996 19450 21048 19456
rect 21100 19378 21128 19722
rect 21088 19372 21140 19378
rect 21088 19314 21140 19320
rect 20996 18760 21048 18766
rect 20996 18702 21048 18708
rect 21008 17241 21036 18702
rect 21088 18692 21140 18698
rect 21088 18634 21140 18640
rect 21100 18086 21128 18634
rect 21088 18080 21140 18086
rect 21088 18022 21140 18028
rect 20994 17232 21050 17241
rect 20994 17167 21050 17176
rect 20904 16244 20956 16250
rect 20904 16186 20956 16192
rect 20720 16108 20772 16114
rect 20720 16050 20772 16056
rect 20732 15570 20760 16050
rect 20720 15564 20772 15570
rect 20720 15506 20772 15512
rect 20904 15474 20956 15480
rect 20956 15422 21036 15450
rect 20904 15416 20956 15422
rect 20904 15360 20956 15366
rect 20904 15302 20956 15308
rect 20916 14414 20944 15302
rect 21008 14958 21036 15422
rect 20996 14952 21048 14958
rect 20996 14894 21048 14900
rect 20904 14408 20956 14414
rect 20904 14350 20956 14356
rect 21008 14278 21036 14894
rect 20996 14272 21048 14278
rect 20996 14214 21048 14220
rect 21008 14074 21036 14214
rect 20996 14068 21048 14074
rect 20996 14010 21048 14016
rect 20628 13932 20680 13938
rect 20628 13874 20680 13880
rect 20536 11892 20588 11898
rect 20536 11834 20588 11840
rect 20640 11778 20668 13874
rect 20720 13320 20772 13326
rect 20720 13262 20772 13268
rect 20732 12442 20760 13262
rect 20996 12912 21048 12918
rect 20996 12854 21048 12860
rect 20720 12436 20772 12442
rect 20720 12378 20772 12384
rect 20548 11762 20668 11778
rect 20536 11756 20668 11762
rect 20588 11750 20668 11756
rect 20536 11698 20588 11704
rect 20444 11212 20496 11218
rect 20444 11154 20496 11160
rect 20444 11008 20496 11014
rect 20444 10950 20496 10956
rect 20456 10742 20484 10950
rect 20444 10736 20496 10742
rect 20444 10678 20496 10684
rect 20548 10554 20576 11698
rect 20732 11694 20760 12378
rect 21008 11762 21036 12854
rect 20996 11756 21048 11762
rect 20996 11698 21048 11704
rect 20628 11688 20680 11694
rect 20628 11630 20680 11636
rect 20720 11688 20772 11694
rect 20720 11630 20772 11636
rect 20640 10810 20668 11630
rect 20904 11552 20956 11558
rect 20904 11494 20956 11500
rect 20916 11150 20944 11494
rect 20904 11144 20956 11150
rect 20904 11086 20956 11092
rect 20628 10804 20680 10810
rect 20628 10746 20680 10752
rect 20456 10526 20576 10554
rect 20640 10538 20668 10746
rect 20628 10532 20680 10538
rect 20456 10062 20484 10526
rect 20628 10474 20680 10480
rect 20444 10056 20496 10062
rect 20444 9998 20496 10004
rect 21086 8392 21142 8401
rect 20720 8356 20772 8362
rect 21086 8327 21142 8336
rect 20720 8298 20772 8304
rect 20732 8090 20760 8298
rect 20720 8084 20772 8090
rect 20720 8026 20772 8032
rect 20352 7948 20404 7954
rect 20352 7890 20404 7896
rect 20732 7886 20760 8026
rect 20720 7880 20772 7886
rect 20720 7822 20772 7828
rect 20996 7812 21048 7818
rect 20996 7754 21048 7760
rect 20260 7744 20312 7750
rect 20260 7686 20312 7692
rect 20272 7478 20300 7686
rect 21008 7546 21036 7754
rect 21100 7750 21128 8327
rect 21088 7744 21140 7750
rect 21088 7686 21140 7692
rect 20996 7540 21048 7546
rect 20996 7482 21048 7488
rect 20260 7472 20312 7478
rect 20312 7432 20392 7460
rect 20260 7414 20312 7420
rect 20260 6860 20312 6866
rect 20260 6802 20312 6808
rect 20272 5778 20300 6802
rect 20364 6662 20392 7432
rect 20904 7404 20956 7410
rect 20904 7346 20956 7352
rect 20916 7002 20944 7346
rect 21088 7200 21140 7206
rect 21088 7142 21140 7148
rect 20904 6996 20956 7002
rect 20904 6938 20956 6944
rect 20628 6724 20680 6730
rect 20628 6666 20680 6672
rect 20352 6656 20404 6662
rect 20352 6598 20404 6604
rect 20536 6112 20588 6118
rect 20536 6054 20588 6060
rect 20260 5772 20312 5778
rect 20260 5714 20312 5720
rect 20548 5710 20576 6054
rect 20536 5704 20588 5710
rect 20536 5646 20588 5652
rect 20640 5370 20668 6666
rect 20628 5364 20680 5370
rect 20628 5306 20680 5312
rect 20168 4752 20220 4758
rect 20168 4694 20220 4700
rect 20076 4616 20128 4622
rect 20076 4558 20128 4564
rect 20916 4146 20944 6938
rect 21100 5234 21128 7142
rect 21088 5228 21140 5234
rect 21088 5170 21140 5176
rect 20904 4140 20956 4146
rect 20904 4082 20956 4088
rect 20812 4072 20864 4078
rect 20812 4014 20864 4020
rect 19984 3936 20036 3942
rect 19984 3878 20036 3884
rect 20260 3936 20312 3942
rect 20260 3878 20312 3884
rect 18788 3460 18840 3466
rect 18788 3402 18840 3408
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 19996 3126 20024 3878
rect 20272 3602 20300 3878
rect 20260 3596 20312 3602
rect 20260 3538 20312 3544
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 20076 3528 20128 3534
rect 20076 3470 20128 3476
rect 19984 3120 20036 3126
rect 19984 3062 20036 3068
rect 20088 3058 20116 3470
rect 20076 3052 20128 3058
rect 20076 2994 20128 3000
rect 19984 2372 20036 2378
rect 19984 2314 20036 2320
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 19996 800 20024 2314
rect 20640 800 20668 3538
rect 20824 3466 20852 4014
rect 20904 3936 20956 3942
rect 20904 3878 20956 3884
rect 20812 3460 20864 3466
rect 20812 3402 20864 3408
rect 20916 2514 20944 3878
rect 21192 2774 21220 22066
rect 21272 21548 21324 21554
rect 21272 21490 21324 21496
rect 21284 21146 21312 21490
rect 21272 21140 21324 21146
rect 21272 21082 21324 21088
rect 21284 20942 21312 21082
rect 21272 20936 21324 20942
rect 21272 20878 21324 20884
rect 21284 18630 21312 20878
rect 21364 20800 21416 20806
rect 21364 20742 21416 20748
rect 21272 18624 21324 18630
rect 21272 18566 21324 18572
rect 21272 18080 21324 18086
rect 21270 18048 21272 18057
rect 21324 18048 21326 18057
rect 21270 17983 21326 17992
rect 21272 16244 21324 16250
rect 21272 16186 21324 16192
rect 21284 6322 21312 16186
rect 21376 14006 21404 20742
rect 21454 19816 21510 19825
rect 21454 19751 21510 19760
rect 21468 16046 21496 19751
rect 21560 18737 21588 25298
rect 21836 25226 21864 25978
rect 22296 25974 22324 26182
rect 22284 25968 22336 25974
rect 22284 25910 22336 25916
rect 22468 25900 22520 25906
rect 22468 25842 22520 25848
rect 22480 25362 22508 25842
rect 22468 25356 22520 25362
rect 22468 25298 22520 25304
rect 21824 25220 21876 25226
rect 21824 25162 21876 25168
rect 21640 25152 21692 25158
rect 21640 25094 21692 25100
rect 21652 19854 21680 25094
rect 22100 24880 22152 24886
rect 22020 24828 22100 24834
rect 22020 24822 22152 24828
rect 22020 24806 22140 24822
rect 21824 24744 21876 24750
rect 21824 24686 21876 24692
rect 21836 23730 21864 24686
rect 21824 23724 21876 23730
rect 21824 23666 21876 23672
rect 21732 20460 21784 20466
rect 21732 20402 21784 20408
rect 21916 20460 21968 20466
rect 21916 20402 21968 20408
rect 21744 19990 21772 20402
rect 21732 19984 21784 19990
rect 21732 19926 21784 19932
rect 21640 19848 21692 19854
rect 21640 19790 21692 19796
rect 21732 19848 21784 19854
rect 21732 19790 21784 19796
rect 21744 19446 21772 19790
rect 21824 19780 21876 19786
rect 21824 19722 21876 19728
rect 21732 19440 21784 19446
rect 21732 19382 21784 19388
rect 21836 19378 21864 19722
rect 21928 19514 21956 20402
rect 22020 20330 22048 24806
rect 22100 24132 22152 24138
rect 22100 24074 22152 24080
rect 22008 20324 22060 20330
rect 22008 20266 22060 20272
rect 22008 19984 22060 19990
rect 22008 19926 22060 19932
rect 21916 19508 21968 19514
rect 21916 19450 21968 19456
rect 22020 19378 22048 19926
rect 21824 19372 21876 19378
rect 21824 19314 21876 19320
rect 22008 19372 22060 19378
rect 22008 19314 22060 19320
rect 22020 19174 22048 19314
rect 22008 19168 22060 19174
rect 22008 19110 22060 19116
rect 21732 18964 21784 18970
rect 21732 18906 21784 18912
rect 21744 18766 21772 18906
rect 21732 18760 21784 18766
rect 21546 18728 21602 18737
rect 21732 18702 21784 18708
rect 21546 18663 21602 18672
rect 21640 18624 21692 18630
rect 21640 18566 21692 18572
rect 21652 18358 21680 18566
rect 21640 18352 21692 18358
rect 21640 18294 21692 18300
rect 21730 18320 21786 18329
rect 21730 18255 21786 18264
rect 21744 17542 21772 18255
rect 21732 17536 21784 17542
rect 21732 17478 21784 17484
rect 21744 17270 21772 17478
rect 21732 17264 21784 17270
rect 21732 17206 21784 17212
rect 21456 16040 21508 16046
rect 21456 15982 21508 15988
rect 21916 15496 21968 15502
rect 21916 15438 21968 15444
rect 21548 15428 21600 15434
rect 21548 15370 21600 15376
rect 21824 15428 21876 15434
rect 21824 15370 21876 15376
rect 21560 15162 21588 15370
rect 21548 15156 21600 15162
rect 21548 15098 21600 15104
rect 21836 14890 21864 15370
rect 21928 15026 21956 15438
rect 22008 15360 22060 15366
rect 22008 15302 22060 15308
rect 21916 15020 21968 15026
rect 21916 14962 21968 14968
rect 21824 14884 21876 14890
rect 21824 14826 21876 14832
rect 21928 14074 21956 14962
rect 22020 14346 22048 15302
rect 22008 14340 22060 14346
rect 22008 14282 22060 14288
rect 21916 14068 21968 14074
rect 21916 14010 21968 14016
rect 21364 14000 21416 14006
rect 21364 13942 21416 13948
rect 21376 12918 21404 13942
rect 21364 12912 21416 12918
rect 21364 12854 21416 12860
rect 21916 12164 21968 12170
rect 21916 12106 21968 12112
rect 21928 11898 21956 12106
rect 21916 11892 21968 11898
rect 21916 11834 21968 11840
rect 21456 11076 21508 11082
rect 21456 11018 21508 11024
rect 21272 6316 21324 6322
rect 21272 6258 21324 6264
rect 21284 5234 21312 6258
rect 21272 5228 21324 5234
rect 21272 5170 21324 5176
rect 21284 5030 21312 5170
rect 21272 5024 21324 5030
rect 21272 4966 21324 4972
rect 21468 3738 21496 11018
rect 22008 10532 22060 10538
rect 22008 10474 22060 10480
rect 21824 10464 21876 10470
rect 21824 10406 21876 10412
rect 21836 10062 21864 10406
rect 22020 10062 22048 10474
rect 21824 10056 21876 10062
rect 21824 9998 21876 10004
rect 22008 10056 22060 10062
rect 22008 9998 22060 10004
rect 21640 7744 21692 7750
rect 21640 7686 21692 7692
rect 21652 6474 21680 7686
rect 21652 6446 21956 6474
rect 21652 5846 21680 6446
rect 21928 6322 21956 6446
rect 21824 6316 21876 6322
rect 21824 6258 21876 6264
rect 21916 6316 21968 6322
rect 21916 6258 21968 6264
rect 21640 5840 21692 5846
rect 21640 5782 21692 5788
rect 21836 4622 21864 6258
rect 21824 4616 21876 4622
rect 21824 4558 21876 4564
rect 21456 3732 21508 3738
rect 21456 3674 21508 3680
rect 22008 2848 22060 2854
rect 22008 2790 22060 2796
rect 21008 2746 21220 2774
rect 21008 2582 21036 2746
rect 20996 2576 21048 2582
rect 20996 2518 21048 2524
rect 21272 2576 21324 2582
rect 21272 2518 21324 2524
rect 20904 2508 20956 2514
rect 20904 2450 20956 2456
rect 21284 800 21312 2518
rect 22020 2514 22048 2790
rect 22112 2650 22140 24074
rect 22376 23112 22428 23118
rect 22376 23054 22428 23060
rect 22190 21992 22246 22001
rect 22190 21927 22192 21936
rect 22244 21927 22246 21936
rect 22284 21956 22336 21962
rect 22192 21898 22244 21904
rect 22284 21898 22336 21904
rect 22296 21622 22324 21898
rect 22388 21622 22416 23054
rect 22572 22094 22600 26206
rect 22744 24404 22796 24410
rect 22744 24346 22796 24352
rect 22572 22066 22692 22094
rect 22284 21616 22336 21622
rect 22284 21558 22336 21564
rect 22376 21616 22428 21622
rect 22428 21576 22508 21604
rect 22376 21558 22428 21564
rect 22376 21480 22428 21486
rect 22374 21448 22376 21457
rect 22428 21448 22430 21457
rect 22374 21383 22430 21392
rect 22374 21176 22430 21185
rect 22374 21111 22376 21120
rect 22428 21111 22430 21120
rect 22376 21082 22428 21088
rect 22376 21004 22428 21010
rect 22376 20946 22428 20952
rect 22388 20262 22416 20946
rect 22192 20256 22244 20262
rect 22192 20198 22244 20204
rect 22376 20256 22428 20262
rect 22376 20198 22428 20204
rect 22204 19446 22232 20198
rect 22284 19712 22336 19718
rect 22284 19654 22336 19660
rect 22192 19440 22244 19446
rect 22192 19382 22244 19388
rect 22192 19236 22244 19242
rect 22192 19178 22244 19184
rect 22204 18358 22232 19178
rect 22192 18352 22244 18358
rect 22192 18294 22244 18300
rect 22296 16114 22324 19654
rect 22388 18834 22416 20198
rect 22480 19417 22508 21576
rect 22560 21548 22612 21554
rect 22560 21490 22612 21496
rect 22572 21146 22600 21490
rect 22560 21140 22612 21146
rect 22560 21082 22612 21088
rect 22560 20868 22612 20874
rect 22560 20810 22612 20816
rect 22572 20330 22600 20810
rect 22560 20324 22612 20330
rect 22560 20266 22612 20272
rect 22466 19408 22522 19417
rect 22466 19343 22468 19352
rect 22520 19343 22522 19352
rect 22468 19314 22520 19320
rect 22376 18828 22428 18834
rect 22376 18770 22428 18776
rect 22480 16658 22508 19314
rect 22560 18760 22612 18766
rect 22560 18702 22612 18708
rect 22572 18426 22600 18702
rect 22560 18420 22612 18426
rect 22560 18362 22612 18368
rect 22468 16652 22520 16658
rect 22468 16594 22520 16600
rect 22284 16108 22336 16114
rect 22284 16050 22336 16056
rect 22296 15026 22324 16050
rect 22192 15020 22244 15026
rect 22192 14962 22244 14968
rect 22284 15020 22336 15026
rect 22284 14962 22336 14968
rect 22204 14550 22232 14962
rect 22468 14884 22520 14890
rect 22468 14826 22520 14832
rect 22192 14544 22244 14550
rect 22192 14486 22244 14492
rect 22192 11688 22244 11694
rect 22192 11630 22244 11636
rect 22204 11150 22232 11630
rect 22192 11144 22244 11150
rect 22192 11086 22244 11092
rect 22204 7342 22232 11086
rect 22376 11076 22428 11082
rect 22376 11018 22428 11024
rect 22284 11008 22336 11014
rect 22284 10950 22336 10956
rect 22296 10674 22324 10950
rect 22284 10668 22336 10674
rect 22284 10610 22336 10616
rect 22284 10532 22336 10538
rect 22284 10474 22336 10480
rect 22296 9994 22324 10474
rect 22388 10266 22416 11018
rect 22480 10674 22508 14826
rect 22468 10668 22520 10674
rect 22468 10610 22520 10616
rect 22376 10260 22428 10266
rect 22376 10202 22428 10208
rect 22284 9988 22336 9994
rect 22284 9930 22336 9936
rect 22192 7336 22244 7342
rect 22192 7278 22244 7284
rect 22204 6730 22232 7278
rect 22192 6724 22244 6730
rect 22192 6666 22244 6672
rect 22204 6254 22232 6666
rect 22296 6390 22324 9930
rect 22284 6384 22336 6390
rect 22284 6326 22336 6332
rect 22468 6384 22520 6390
rect 22468 6326 22520 6332
rect 22192 6248 22244 6254
rect 22192 6190 22244 6196
rect 22192 5636 22244 5642
rect 22192 5578 22244 5584
rect 22204 5370 22232 5578
rect 22192 5364 22244 5370
rect 22192 5306 22244 5312
rect 22480 5234 22508 6326
rect 22284 5228 22336 5234
rect 22284 5170 22336 5176
rect 22468 5228 22520 5234
rect 22468 5170 22520 5176
rect 22560 5228 22612 5234
rect 22560 5170 22612 5176
rect 22100 2644 22152 2650
rect 22100 2586 22152 2592
rect 22008 2508 22060 2514
rect 22008 2450 22060 2456
rect 22296 1970 22324 5170
rect 22480 5098 22508 5170
rect 22468 5092 22520 5098
rect 22468 5034 22520 5040
rect 22572 4826 22600 5170
rect 22560 4820 22612 4826
rect 22560 4762 22612 4768
rect 22560 4004 22612 4010
rect 22560 3946 22612 3952
rect 22572 3194 22600 3946
rect 22664 3194 22692 22066
rect 22756 14414 22784 24346
rect 22848 17252 22876 27950
rect 22940 27402 22968 28018
rect 22928 27396 22980 27402
rect 22928 27338 22980 27344
rect 23308 22094 23336 36314
rect 23400 33454 23428 38898
rect 23492 38758 23520 39238
rect 23480 38752 23532 38758
rect 23480 38694 23532 38700
rect 23492 38418 23520 38694
rect 23480 38412 23532 38418
rect 23480 38354 23532 38360
rect 23480 35080 23532 35086
rect 23480 35022 23532 35028
rect 23388 33448 23440 33454
rect 23388 33390 23440 33396
rect 23388 32836 23440 32842
rect 23388 32778 23440 32784
rect 23400 24410 23428 32778
rect 23492 32473 23520 35022
rect 23478 32464 23534 32473
rect 23478 32399 23534 32408
rect 23478 32056 23534 32065
rect 23478 31991 23534 32000
rect 23492 31822 23520 31991
rect 23480 31816 23532 31822
rect 23480 31758 23532 31764
rect 23584 30818 23612 43658
rect 24032 42696 24084 42702
rect 24032 42638 24084 42644
rect 23848 42288 23900 42294
rect 23848 42230 23900 42236
rect 23664 42152 23716 42158
rect 23664 42094 23716 42100
rect 23676 41546 23704 42094
rect 23860 41818 23888 42230
rect 24044 42226 24072 42638
rect 23940 42220 23992 42226
rect 23940 42162 23992 42168
rect 24032 42220 24084 42226
rect 24032 42162 24084 42168
rect 23848 41812 23900 41818
rect 23848 41754 23900 41760
rect 23664 41540 23716 41546
rect 23664 41482 23716 41488
rect 23952 41478 23980 42162
rect 24044 41750 24072 42162
rect 24032 41744 24084 41750
rect 24032 41686 24084 41692
rect 24032 41608 24084 41614
rect 24032 41550 24084 41556
rect 23848 41472 23900 41478
rect 23848 41414 23900 41420
rect 23940 41472 23992 41478
rect 23940 41414 23992 41420
rect 23860 41138 23888 41414
rect 23664 41132 23716 41138
rect 23664 41074 23716 41080
rect 23848 41132 23900 41138
rect 23848 41074 23900 41080
rect 23676 40390 23704 41074
rect 23664 40384 23716 40390
rect 23664 40326 23716 40332
rect 23676 39953 23704 40326
rect 23860 40118 23888 41074
rect 23848 40112 23900 40118
rect 23848 40054 23900 40060
rect 23662 39944 23718 39953
rect 23662 39879 23718 39888
rect 23846 39944 23902 39953
rect 23846 39879 23902 39888
rect 23664 39296 23716 39302
rect 23664 39238 23716 39244
rect 23676 38282 23704 39238
rect 23756 38888 23808 38894
rect 23756 38830 23808 38836
rect 23664 38276 23716 38282
rect 23664 38218 23716 38224
rect 23768 36530 23796 38830
rect 23676 36502 23796 36530
rect 23676 30938 23704 36502
rect 23860 35086 23888 39879
rect 23952 39438 23980 41414
rect 23940 39432 23992 39438
rect 23940 39374 23992 39380
rect 23952 38486 23980 39374
rect 23940 38480 23992 38486
rect 23940 38422 23992 38428
rect 23940 37800 23992 37806
rect 23940 37742 23992 37748
rect 23952 37262 23980 37742
rect 23940 37256 23992 37262
rect 23940 37198 23992 37204
rect 23940 36848 23992 36854
rect 23940 36790 23992 36796
rect 23848 35080 23900 35086
rect 23848 35022 23900 35028
rect 23952 34610 23980 36790
rect 23940 34604 23992 34610
rect 23940 34546 23992 34552
rect 23940 33992 23992 33998
rect 23940 33934 23992 33940
rect 23756 33108 23808 33114
rect 23756 33050 23808 33056
rect 23768 32502 23796 33050
rect 23848 32836 23900 32842
rect 23848 32778 23900 32784
rect 23860 32570 23888 32778
rect 23848 32564 23900 32570
rect 23848 32506 23900 32512
rect 23756 32496 23808 32502
rect 23952 32450 23980 33934
rect 23756 32438 23808 32444
rect 23860 32422 23980 32450
rect 23756 32224 23808 32230
rect 23756 32166 23808 32172
rect 23768 31822 23796 32166
rect 23756 31816 23808 31822
rect 23756 31758 23808 31764
rect 23664 30932 23716 30938
rect 23664 30874 23716 30880
rect 23584 30790 23796 30818
rect 23664 30728 23716 30734
rect 23664 30670 23716 30676
rect 23572 30592 23624 30598
rect 23572 30534 23624 30540
rect 23480 29640 23532 29646
rect 23478 29608 23480 29617
rect 23532 29608 23534 29617
rect 23478 29543 23534 29552
rect 23480 28416 23532 28422
rect 23480 28358 23532 28364
rect 23492 28082 23520 28358
rect 23480 28076 23532 28082
rect 23480 28018 23532 28024
rect 23492 27538 23520 28018
rect 23480 27532 23532 27538
rect 23480 27474 23532 27480
rect 23480 27328 23532 27334
rect 23480 27270 23532 27276
rect 23492 26926 23520 27270
rect 23480 26920 23532 26926
rect 23480 26862 23532 26868
rect 23480 25900 23532 25906
rect 23480 25842 23532 25848
rect 23388 24404 23440 24410
rect 23388 24346 23440 24352
rect 23492 23798 23520 25842
rect 23480 23792 23532 23798
rect 23480 23734 23532 23740
rect 23492 23186 23520 23734
rect 23584 23594 23612 30534
rect 23676 26738 23704 30670
rect 23768 26874 23796 30790
rect 23860 26994 23888 32422
rect 23940 32020 23992 32026
rect 23940 31962 23992 31968
rect 23952 31414 23980 31962
rect 23940 31408 23992 31414
rect 23940 31350 23992 31356
rect 23940 27124 23992 27130
rect 23940 27066 23992 27072
rect 23848 26988 23900 26994
rect 23848 26930 23900 26936
rect 23768 26846 23888 26874
rect 23676 26710 23796 26738
rect 23572 23588 23624 23594
rect 23572 23530 23624 23536
rect 23480 23180 23532 23186
rect 23480 23122 23532 23128
rect 23664 22976 23716 22982
rect 23664 22918 23716 22924
rect 23216 22066 23336 22094
rect 23112 21616 23164 21622
rect 23112 21558 23164 21564
rect 23018 21448 23074 21457
rect 23018 21383 23074 21392
rect 23032 21350 23060 21383
rect 22928 21344 22980 21350
rect 22928 21286 22980 21292
rect 23020 21344 23072 21350
rect 23020 21286 23072 21292
rect 22940 20942 22968 21286
rect 22928 20936 22980 20942
rect 22928 20878 22980 20884
rect 23032 20534 23060 21286
rect 23124 21185 23152 21558
rect 23110 21176 23166 21185
rect 23110 21111 23166 21120
rect 23020 20528 23072 20534
rect 23020 20470 23072 20476
rect 23112 20528 23164 20534
rect 23112 20470 23164 20476
rect 22928 20256 22980 20262
rect 22928 20198 22980 20204
rect 22940 19825 22968 20198
rect 22926 19816 22982 19825
rect 22926 19751 22982 19760
rect 22928 19372 22980 19378
rect 22928 19314 22980 19320
rect 22940 18970 22968 19314
rect 23124 19174 23152 20470
rect 23112 19168 23164 19174
rect 23112 19110 23164 19116
rect 22928 18964 22980 18970
rect 22928 18906 22980 18912
rect 22928 18624 22980 18630
rect 22926 18592 22928 18601
rect 22980 18592 22982 18601
rect 22926 18527 22982 18536
rect 22848 17224 22968 17252
rect 22744 14408 22796 14414
rect 22744 14350 22796 14356
rect 22836 14272 22888 14278
rect 22836 14214 22888 14220
rect 22848 14006 22876 14214
rect 22836 14000 22888 14006
rect 22836 13942 22888 13948
rect 22836 7812 22888 7818
rect 22836 7754 22888 7760
rect 22848 6186 22876 7754
rect 22836 6180 22888 6186
rect 22836 6122 22888 6128
rect 22560 3188 22612 3194
rect 22560 3130 22612 3136
rect 22652 3188 22704 3194
rect 22652 3130 22704 3136
rect 22560 3052 22612 3058
rect 22560 2994 22612 3000
rect 22284 1964 22336 1970
rect 22284 1906 22336 1912
rect 22572 800 22600 2994
rect 22940 2378 22968 17224
rect 23020 17196 23072 17202
rect 23020 17138 23072 17144
rect 23032 17105 23060 17138
rect 23018 17096 23074 17105
rect 23018 17031 23074 17040
rect 23124 16454 23152 19110
rect 23112 16448 23164 16454
rect 23112 16390 23164 16396
rect 23020 14612 23072 14618
rect 23020 14554 23072 14560
rect 23032 14074 23060 14554
rect 23020 14068 23072 14074
rect 23020 14010 23072 14016
rect 23020 13320 23072 13326
rect 23020 13262 23072 13268
rect 23032 10674 23060 13262
rect 23216 12434 23244 22066
rect 23676 22001 23704 22918
rect 23768 22094 23796 26710
rect 23860 25362 23888 26846
rect 23952 26246 23980 27066
rect 23940 26240 23992 26246
rect 23940 26182 23992 26188
rect 23848 25356 23900 25362
rect 23848 25298 23900 25304
rect 23940 23112 23992 23118
rect 23940 23054 23992 23060
rect 23952 22778 23980 23054
rect 23940 22772 23992 22778
rect 23940 22714 23992 22720
rect 24044 22094 24072 41550
rect 24136 41414 24164 45358
rect 24228 42242 24256 47602
rect 24308 47456 24360 47462
rect 24308 47398 24360 47404
rect 24320 47258 24348 47398
rect 24412 47258 24440 49166
rect 24584 49156 24636 49162
rect 24584 49098 24636 49104
rect 24596 47802 24624 49098
rect 25792 48822 25820 51200
rect 26436 48822 26464 51200
rect 27540 49586 27568 51326
rect 27710 51200 27766 52000
rect 28354 51200 28410 52000
rect 28998 51200 29054 52000
rect 29642 51200 29698 52000
rect 30930 51200 30986 52000
rect 31574 51200 31630 52000
rect 32218 51200 32274 52000
rect 32862 51200 32918 52000
rect 33506 51354 33562 52000
rect 34150 51354 34206 52000
rect 33506 51326 33824 51354
rect 33506 51200 33562 51326
rect 27540 49558 27660 49586
rect 27632 49298 27660 49558
rect 27620 49292 27672 49298
rect 27620 49234 27672 49240
rect 26976 49224 27028 49230
rect 26976 49166 27028 49172
rect 26792 48884 26844 48890
rect 26792 48826 26844 48832
rect 25780 48816 25832 48822
rect 25780 48758 25832 48764
rect 26424 48816 26476 48822
rect 26424 48758 26476 48764
rect 25412 48544 25464 48550
rect 25412 48486 25464 48492
rect 25504 48544 25556 48550
rect 25504 48486 25556 48492
rect 25320 48272 25372 48278
rect 25320 48214 25372 48220
rect 24952 48068 25004 48074
rect 24952 48010 25004 48016
rect 24584 47796 24636 47802
rect 24584 47738 24636 47744
rect 24768 47796 24820 47802
rect 24768 47738 24820 47744
rect 24308 47252 24360 47258
rect 24308 47194 24360 47200
rect 24400 47252 24452 47258
rect 24400 47194 24452 47200
rect 24780 47122 24808 47738
rect 24964 47734 24992 48010
rect 25228 48000 25280 48006
rect 25228 47942 25280 47948
rect 24952 47728 25004 47734
rect 24952 47670 25004 47676
rect 24860 47252 24912 47258
rect 24860 47194 24912 47200
rect 24768 47116 24820 47122
rect 24768 47058 24820 47064
rect 24872 47054 24900 47194
rect 24860 47048 24912 47054
rect 24860 46990 24912 46996
rect 24768 44328 24820 44334
rect 24768 44270 24820 44276
rect 24676 43308 24728 43314
rect 24676 43250 24728 43256
rect 24584 43240 24636 43246
rect 24584 43182 24636 43188
rect 24228 42214 24348 42242
rect 24136 41386 24256 41414
rect 24228 41274 24256 41386
rect 24216 41268 24268 41274
rect 24216 41210 24268 41216
rect 24216 34604 24268 34610
rect 24216 34546 24268 34552
rect 24228 34202 24256 34546
rect 24216 34196 24268 34202
rect 24216 34138 24268 34144
rect 24320 34082 24348 42214
rect 24596 41546 24624 43182
rect 24688 42294 24716 43250
rect 24676 42288 24728 42294
rect 24676 42230 24728 42236
rect 24780 42140 24808 44270
rect 24964 43722 24992 47670
rect 25240 47666 25268 47942
rect 25228 47660 25280 47666
rect 25228 47602 25280 47608
rect 25136 47592 25188 47598
rect 25136 47534 25188 47540
rect 24952 43716 25004 43722
rect 24952 43658 25004 43664
rect 24860 43308 24912 43314
rect 24860 43250 24912 43256
rect 25044 43308 25096 43314
rect 25044 43250 25096 43256
rect 24872 42634 24900 43250
rect 24952 43104 25004 43110
rect 24952 43046 25004 43052
rect 24964 42702 24992 43046
rect 24952 42696 25004 42702
rect 24952 42638 25004 42644
rect 24860 42628 24912 42634
rect 24860 42570 24912 42576
rect 24688 42112 24808 42140
rect 24584 41540 24636 41546
rect 24584 41482 24636 41488
rect 24492 40112 24544 40118
rect 24492 40054 24544 40060
rect 24400 39908 24452 39914
rect 24400 39850 24452 39856
rect 24412 39370 24440 39850
rect 24400 39364 24452 39370
rect 24400 39306 24452 39312
rect 24400 37120 24452 37126
rect 24400 37062 24452 37068
rect 24412 36922 24440 37062
rect 24400 36916 24452 36922
rect 24400 36858 24452 36864
rect 24504 36802 24532 40054
rect 24584 39296 24636 39302
rect 24584 39238 24636 39244
rect 24596 38758 24624 39238
rect 24688 38894 24716 42112
rect 24952 42016 25004 42022
rect 24952 41958 25004 41964
rect 24768 41744 24820 41750
rect 24768 41686 24820 41692
rect 24780 39846 24808 41686
rect 24964 41614 24992 41958
rect 25056 41614 25084 43250
rect 24952 41608 25004 41614
rect 24952 41550 25004 41556
rect 25044 41608 25096 41614
rect 25044 41550 25096 41556
rect 24860 40044 24912 40050
rect 24860 39986 24912 39992
rect 24768 39840 24820 39846
rect 24768 39782 24820 39788
rect 24780 39438 24808 39782
rect 24768 39432 24820 39438
rect 24768 39374 24820 39380
rect 24780 38962 24808 39374
rect 24872 39370 24900 39986
rect 25148 39574 25176 47534
rect 25240 47054 25268 47602
rect 25228 47048 25280 47054
rect 25228 46990 25280 46996
rect 25240 46646 25268 46990
rect 25228 46640 25280 46646
rect 25228 46582 25280 46588
rect 25240 45966 25268 46582
rect 25228 45960 25280 45966
rect 25228 45902 25280 45908
rect 25228 41200 25280 41206
rect 25228 41142 25280 41148
rect 25240 40934 25268 41142
rect 25228 40928 25280 40934
rect 25228 40870 25280 40876
rect 25136 39568 25188 39574
rect 25136 39510 25188 39516
rect 24860 39364 24912 39370
rect 24860 39306 24912 39312
rect 24952 39364 25004 39370
rect 24952 39306 25004 39312
rect 24768 38956 24820 38962
rect 24768 38898 24820 38904
rect 24676 38888 24728 38894
rect 24676 38830 24728 38836
rect 24584 38752 24636 38758
rect 24584 38694 24636 38700
rect 24596 37942 24624 38694
rect 24676 38344 24728 38350
rect 24676 38286 24728 38292
rect 24688 37942 24716 38286
rect 24584 37936 24636 37942
rect 24584 37878 24636 37884
rect 24676 37936 24728 37942
rect 24676 37878 24728 37884
rect 24780 37262 24808 38898
rect 24768 37256 24820 37262
rect 24768 37198 24820 37204
rect 24584 37188 24636 37194
rect 24584 37130 24636 37136
rect 24596 36922 24624 37130
rect 24584 36916 24636 36922
rect 24584 36858 24636 36864
rect 24780 36854 24808 37198
rect 24860 37120 24912 37126
rect 24860 37062 24912 37068
rect 24768 36848 24820 36854
rect 24400 36780 24452 36786
rect 24504 36774 24624 36802
rect 24768 36790 24820 36796
rect 24400 36722 24452 36728
rect 24412 36378 24440 36722
rect 24400 36372 24452 36378
rect 24400 36314 24452 36320
rect 24228 34054 24348 34082
rect 24124 33040 24176 33046
rect 24124 32982 24176 32988
rect 24136 32570 24164 32982
rect 24124 32564 24176 32570
rect 24124 32506 24176 32512
rect 24122 32464 24178 32473
rect 24122 32399 24178 32408
rect 24136 27062 24164 32399
rect 24228 27130 24256 34054
rect 24492 33584 24544 33590
rect 24492 33526 24544 33532
rect 24308 33312 24360 33318
rect 24308 33254 24360 33260
rect 24320 32434 24348 33254
rect 24504 32434 24532 33526
rect 24308 32428 24360 32434
rect 24308 32370 24360 32376
rect 24492 32428 24544 32434
rect 24492 32370 24544 32376
rect 24308 32292 24360 32298
rect 24308 32234 24360 32240
rect 24216 27124 24268 27130
rect 24216 27066 24268 27072
rect 24124 27056 24176 27062
rect 24124 26998 24176 27004
rect 24216 26988 24268 26994
rect 24216 26930 24268 26936
rect 24124 23656 24176 23662
rect 24124 23598 24176 23604
rect 24136 22778 24164 23598
rect 24124 22772 24176 22778
rect 24124 22714 24176 22720
rect 23768 22066 23980 22094
rect 24044 22066 24164 22094
rect 23478 21992 23534 22001
rect 23478 21927 23534 21936
rect 23662 21992 23718 22001
rect 23662 21927 23718 21936
rect 23386 17504 23442 17513
rect 23386 17439 23442 17448
rect 23400 17338 23428 17439
rect 23492 17354 23520 21927
rect 23664 21344 23716 21350
rect 23664 21286 23716 21292
rect 23676 21146 23704 21286
rect 23664 21140 23716 21146
rect 23664 21082 23716 21088
rect 23572 19168 23624 19174
rect 23572 19110 23624 19116
rect 23584 18340 23612 19110
rect 23676 18630 23704 21082
rect 23848 20460 23900 20466
rect 23848 20402 23900 20408
rect 23756 20392 23808 20398
rect 23756 20334 23808 20340
rect 23664 18624 23716 18630
rect 23664 18566 23716 18572
rect 23584 18312 23704 18340
rect 23676 18222 23704 18312
rect 23664 18216 23716 18222
rect 23664 18158 23716 18164
rect 23388 17332 23440 17338
rect 23492 17326 23612 17354
rect 23676 17338 23704 18158
rect 23388 17274 23440 17280
rect 23480 17264 23532 17270
rect 23480 17206 23532 17212
rect 23388 17196 23440 17202
rect 23388 17138 23440 17144
rect 23400 16833 23428 17138
rect 23386 16824 23442 16833
rect 23386 16759 23442 16768
rect 23492 14550 23520 17206
rect 23480 14544 23532 14550
rect 23480 14486 23532 14492
rect 23388 14408 23440 14414
rect 23388 14350 23440 14356
rect 23400 13938 23428 14350
rect 23388 13932 23440 13938
rect 23388 13874 23440 13880
rect 23584 13530 23612 17326
rect 23664 17332 23716 17338
rect 23664 17274 23716 17280
rect 23664 16448 23716 16454
rect 23664 16390 23716 16396
rect 23676 16130 23704 16390
rect 23768 16250 23796 20334
rect 23860 19786 23888 20402
rect 23952 19938 23980 22066
rect 24032 20392 24084 20398
rect 24032 20334 24084 20340
rect 24044 20058 24072 20334
rect 24032 20052 24084 20058
rect 24032 19994 24084 20000
rect 23952 19910 24072 19938
rect 23848 19780 23900 19786
rect 23848 19722 23900 19728
rect 23940 19712 23992 19718
rect 23940 19654 23992 19660
rect 23952 18698 23980 19654
rect 24044 18873 24072 19910
rect 24030 18864 24086 18873
rect 24030 18799 24086 18808
rect 24032 18760 24084 18766
rect 24032 18702 24084 18708
rect 23940 18692 23992 18698
rect 23940 18634 23992 18640
rect 23848 18624 23900 18630
rect 23848 18566 23900 18572
rect 23860 18154 23888 18566
rect 23952 18290 23980 18634
rect 23940 18284 23992 18290
rect 23940 18226 23992 18232
rect 23848 18148 23900 18154
rect 23848 18090 23900 18096
rect 23860 17218 23888 18090
rect 23952 17338 23980 18226
rect 24044 18154 24072 18702
rect 24032 18148 24084 18154
rect 24032 18090 24084 18096
rect 23940 17332 23992 17338
rect 23940 17274 23992 17280
rect 23860 17190 23980 17218
rect 23848 16992 23900 16998
rect 23848 16934 23900 16940
rect 23860 16590 23888 16934
rect 23848 16584 23900 16590
rect 23848 16526 23900 16532
rect 23952 16522 23980 17190
rect 24044 16969 24072 18090
rect 24136 17542 24164 22066
rect 24228 18465 24256 26930
rect 24214 18456 24270 18465
rect 24214 18391 24270 18400
rect 24216 18284 24268 18290
rect 24216 18226 24268 18232
rect 24124 17536 24176 17542
rect 24124 17478 24176 17484
rect 24124 17332 24176 17338
rect 24124 17274 24176 17280
rect 24030 16960 24086 16969
rect 24030 16895 24086 16904
rect 23940 16516 23992 16522
rect 23940 16458 23992 16464
rect 23756 16244 23808 16250
rect 23756 16186 23808 16192
rect 23676 16102 23888 16130
rect 23664 15496 23716 15502
rect 23664 15438 23716 15444
rect 23572 13524 23624 13530
rect 23572 13466 23624 13472
rect 23584 12986 23612 13466
rect 23572 12980 23624 12986
rect 23572 12922 23624 12928
rect 23572 12844 23624 12850
rect 23572 12786 23624 12792
rect 23584 12753 23612 12786
rect 23570 12744 23626 12753
rect 23570 12679 23626 12688
rect 23480 12640 23532 12646
rect 23480 12582 23532 12588
rect 23124 12406 23244 12434
rect 23020 10668 23072 10674
rect 23020 10610 23072 10616
rect 23124 2582 23152 12406
rect 23492 12238 23520 12582
rect 23676 12238 23704 15438
rect 23756 13184 23808 13190
rect 23756 13126 23808 13132
rect 23768 12918 23796 13126
rect 23756 12912 23808 12918
rect 23756 12854 23808 12860
rect 23768 12782 23796 12854
rect 23756 12776 23808 12782
rect 23756 12718 23808 12724
rect 23480 12232 23532 12238
rect 23480 12174 23532 12180
rect 23664 12232 23716 12238
rect 23664 12174 23716 12180
rect 23492 11914 23520 12174
rect 23492 11886 23612 11914
rect 23480 11824 23532 11830
rect 23480 11766 23532 11772
rect 23492 11150 23520 11766
rect 23480 11144 23532 11150
rect 23480 11086 23532 11092
rect 23480 10736 23532 10742
rect 23480 10678 23532 10684
rect 23388 10464 23440 10470
rect 23388 10406 23440 10412
rect 23296 9920 23348 9926
rect 23296 9862 23348 9868
rect 23204 9580 23256 9586
rect 23204 9522 23256 9528
rect 23216 9178 23244 9522
rect 23308 9518 23336 9862
rect 23296 9512 23348 9518
rect 23296 9454 23348 9460
rect 23204 9172 23256 9178
rect 23204 9114 23256 9120
rect 23308 8974 23336 9454
rect 23296 8968 23348 8974
rect 23296 8910 23348 8916
rect 23204 6656 23256 6662
rect 23204 6598 23256 6604
rect 23216 6322 23244 6598
rect 23400 6322 23428 10406
rect 23492 7410 23520 10678
rect 23584 9466 23612 11886
rect 23664 11008 23716 11014
rect 23664 10950 23716 10956
rect 23676 10470 23704 10950
rect 23664 10464 23716 10470
rect 23664 10406 23716 10412
rect 23676 10130 23704 10406
rect 23664 10124 23716 10130
rect 23664 10066 23716 10072
rect 23768 9654 23796 12718
rect 23860 11286 23888 16102
rect 24136 15570 24164 17274
rect 24228 16998 24256 18226
rect 24216 16992 24268 16998
rect 24216 16934 24268 16940
rect 24214 16824 24270 16833
rect 24214 16759 24216 16768
rect 24268 16759 24270 16768
rect 24216 16730 24268 16736
rect 24216 16516 24268 16522
rect 24216 16458 24268 16464
rect 24124 15564 24176 15570
rect 24124 15506 24176 15512
rect 23940 13388 23992 13394
rect 23940 13330 23992 13336
rect 23952 12782 23980 13330
rect 23940 12776 23992 12782
rect 23992 12736 24164 12764
rect 23940 12718 23992 12724
rect 23938 12336 23994 12345
rect 23938 12271 23994 12280
rect 23848 11280 23900 11286
rect 23848 11222 23900 11228
rect 23860 11150 23888 11222
rect 23848 11144 23900 11150
rect 23848 11086 23900 11092
rect 23848 11008 23900 11014
rect 23848 10950 23900 10956
rect 23860 10674 23888 10950
rect 23848 10668 23900 10674
rect 23848 10610 23900 10616
rect 23848 9988 23900 9994
rect 23848 9930 23900 9936
rect 23756 9648 23808 9654
rect 23756 9590 23808 9596
rect 23584 9438 23796 9466
rect 23572 9036 23624 9042
rect 23572 8978 23624 8984
rect 23584 8906 23612 8978
rect 23768 8906 23796 9438
rect 23572 8900 23624 8906
rect 23756 8900 23808 8906
rect 23624 8860 23704 8888
rect 23572 8842 23624 8848
rect 23676 8498 23704 8860
rect 23756 8842 23808 8848
rect 23768 8634 23796 8842
rect 23756 8628 23808 8634
rect 23756 8570 23808 8576
rect 23664 8492 23716 8498
rect 23664 8434 23716 8440
rect 23676 7750 23704 8434
rect 23664 7744 23716 7750
rect 23664 7686 23716 7692
rect 23480 7404 23532 7410
rect 23480 7346 23532 7352
rect 23204 6316 23256 6322
rect 23204 6258 23256 6264
rect 23388 6316 23440 6322
rect 23388 6258 23440 6264
rect 23492 5710 23520 7346
rect 23664 6112 23716 6118
rect 23664 6054 23716 6060
rect 23480 5704 23532 5710
rect 23480 5646 23532 5652
rect 23492 5234 23520 5646
rect 23676 5234 23704 6054
rect 23860 5574 23888 9930
rect 23848 5568 23900 5574
rect 23848 5510 23900 5516
rect 23480 5228 23532 5234
rect 23480 5170 23532 5176
rect 23664 5228 23716 5234
rect 23664 5170 23716 5176
rect 23860 4622 23888 5510
rect 23848 4616 23900 4622
rect 23848 4558 23900 4564
rect 23952 4146 23980 12271
rect 24030 11112 24086 11121
rect 24030 11047 24032 11056
rect 24084 11047 24086 11056
rect 24032 11018 24084 11024
rect 24044 9994 24072 11018
rect 24136 10130 24164 12736
rect 24228 11286 24256 16458
rect 24216 11280 24268 11286
rect 24216 11222 24268 11228
rect 24124 10124 24176 10130
rect 24124 10066 24176 10072
rect 24032 9988 24084 9994
rect 24032 9930 24084 9936
rect 24136 7954 24164 10066
rect 24228 8566 24256 11222
rect 24216 8560 24268 8566
rect 24216 8502 24268 8508
rect 24124 7948 24176 7954
rect 24124 7890 24176 7896
rect 24136 7206 24164 7890
rect 24124 7200 24176 7206
rect 24124 7142 24176 7148
rect 23940 4140 23992 4146
rect 23940 4082 23992 4088
rect 23572 3936 23624 3942
rect 23572 3878 23624 3884
rect 23388 3528 23440 3534
rect 23388 3470 23440 3476
rect 23400 3058 23428 3470
rect 23584 3126 23612 3878
rect 23572 3120 23624 3126
rect 23572 3062 23624 3068
rect 23388 3052 23440 3058
rect 23388 2994 23440 3000
rect 23848 2984 23900 2990
rect 23848 2926 23900 2932
rect 23204 2916 23256 2922
rect 23204 2858 23256 2864
rect 23112 2576 23164 2582
rect 23112 2518 23164 2524
rect 22928 2372 22980 2378
rect 22928 2314 22980 2320
rect 23216 800 23244 2858
rect 23860 800 23888 2926
rect 24320 2038 24348 32234
rect 24596 29510 24624 36774
rect 24872 36174 24900 37062
rect 24676 36168 24728 36174
rect 24676 36110 24728 36116
rect 24860 36168 24912 36174
rect 24860 36110 24912 36116
rect 24400 29504 24452 29510
rect 24400 29446 24452 29452
rect 24584 29504 24636 29510
rect 24584 29446 24636 29452
rect 24412 29238 24440 29446
rect 24400 29232 24452 29238
rect 24400 29174 24452 29180
rect 24492 29096 24544 29102
rect 24492 29038 24544 29044
rect 24504 28626 24532 29038
rect 24492 28620 24544 28626
rect 24492 28562 24544 28568
rect 24400 28076 24452 28082
rect 24400 28018 24452 28024
rect 24412 24682 24440 28018
rect 24504 27470 24532 28562
rect 24584 28484 24636 28490
rect 24584 28426 24636 28432
rect 24596 28218 24624 28426
rect 24584 28212 24636 28218
rect 24584 28154 24636 28160
rect 24492 27464 24544 27470
rect 24492 27406 24544 27412
rect 24504 26450 24532 27406
rect 24688 26874 24716 36110
rect 24964 36106 24992 39306
rect 24952 36100 25004 36106
rect 24952 36042 25004 36048
rect 24768 34128 24820 34134
rect 24768 34070 24820 34076
rect 24780 32774 24808 34070
rect 25044 33992 25096 33998
rect 25044 33934 25096 33940
rect 25056 33590 25084 33934
rect 25044 33584 25096 33590
rect 25044 33526 25096 33532
rect 24768 32768 24820 32774
rect 24768 32710 24820 32716
rect 25044 31204 25096 31210
rect 25044 31146 25096 31152
rect 25056 30666 25084 31146
rect 25044 30660 25096 30666
rect 25044 30602 25096 30608
rect 24952 29708 25004 29714
rect 24952 29650 25004 29656
rect 24860 29640 24912 29646
rect 24860 29582 24912 29588
rect 24768 29504 24820 29510
rect 24768 29446 24820 29452
rect 24780 26994 24808 29446
rect 24872 29306 24900 29582
rect 24860 29300 24912 29306
rect 24860 29242 24912 29248
rect 24964 29186 24992 29650
rect 25136 29640 25188 29646
rect 25134 29608 25136 29617
rect 25188 29608 25190 29617
rect 25134 29543 25190 29552
rect 25044 29504 25096 29510
rect 25044 29446 25096 29452
rect 24872 29158 24992 29186
rect 24872 28966 24900 29158
rect 24860 28960 24912 28966
rect 24860 28902 24912 28908
rect 24872 28082 24900 28902
rect 24860 28076 24912 28082
rect 24860 28018 24912 28024
rect 24952 28076 25004 28082
rect 24952 28018 25004 28024
rect 24964 27674 24992 28018
rect 24952 27668 25004 27674
rect 24952 27610 25004 27616
rect 25056 27130 25084 29446
rect 25148 28082 25176 29543
rect 25136 28076 25188 28082
rect 25136 28018 25188 28024
rect 25044 27124 25096 27130
rect 25044 27066 25096 27072
rect 24768 26988 24820 26994
rect 24768 26930 24820 26936
rect 24596 26846 24716 26874
rect 24492 26444 24544 26450
rect 24492 26386 24544 26392
rect 24504 25974 24532 26386
rect 24492 25968 24544 25974
rect 24492 25910 24544 25916
rect 24492 25220 24544 25226
rect 24492 25162 24544 25168
rect 24400 24676 24452 24682
rect 24400 24618 24452 24624
rect 24504 24562 24532 25162
rect 24412 24534 24532 24562
rect 24412 22642 24440 24534
rect 24492 23724 24544 23730
rect 24492 23666 24544 23672
rect 24504 23594 24532 23666
rect 24492 23588 24544 23594
rect 24492 23530 24544 23536
rect 24400 22636 24452 22642
rect 24400 22578 24452 22584
rect 24412 17338 24440 22578
rect 24596 22094 24624 26846
rect 24676 26784 24728 26790
rect 24676 26726 24728 26732
rect 25044 26784 25096 26790
rect 25044 26726 25096 26732
rect 24688 26382 24716 26726
rect 24676 26376 24728 26382
rect 24676 26318 24728 26324
rect 24860 25696 24912 25702
rect 24860 25638 24912 25644
rect 24872 25294 24900 25638
rect 24860 25288 24912 25294
rect 24860 25230 24912 25236
rect 24768 24200 24820 24206
rect 24768 24142 24820 24148
rect 24780 23526 24808 24142
rect 24860 24064 24912 24070
rect 24860 24006 24912 24012
rect 24872 23798 24900 24006
rect 24860 23792 24912 23798
rect 24860 23734 24912 23740
rect 25056 23730 25084 26726
rect 25044 23724 25096 23730
rect 25044 23666 25096 23672
rect 24768 23520 24820 23526
rect 24768 23462 24820 23468
rect 24780 22710 24808 23462
rect 24952 23044 25004 23050
rect 24952 22986 25004 22992
rect 24768 22704 24820 22710
rect 24768 22646 24820 22652
rect 24768 22568 24820 22574
rect 24768 22510 24820 22516
rect 24596 22066 24716 22094
rect 24584 19168 24636 19174
rect 24584 19110 24636 19116
rect 24596 18698 24624 19110
rect 24584 18692 24636 18698
rect 24584 18634 24636 18640
rect 24596 18086 24624 18634
rect 24584 18080 24636 18086
rect 24584 18022 24636 18028
rect 24596 17746 24624 18022
rect 24584 17740 24636 17746
rect 24584 17682 24636 17688
rect 24492 17604 24544 17610
rect 24492 17546 24544 17552
rect 24504 17338 24532 17546
rect 24584 17536 24636 17542
rect 24584 17478 24636 17484
rect 24400 17332 24452 17338
rect 24400 17274 24452 17280
rect 24492 17332 24544 17338
rect 24492 17274 24544 17280
rect 24398 17096 24454 17105
rect 24398 17031 24454 17040
rect 24412 16794 24440 17031
rect 24504 16833 24532 17274
rect 24490 16824 24546 16833
rect 24400 16788 24452 16794
rect 24490 16759 24546 16768
rect 24400 16730 24452 16736
rect 24398 16552 24454 16561
rect 24398 16487 24400 16496
rect 24452 16487 24454 16496
rect 24492 16516 24544 16522
rect 24400 16458 24452 16464
rect 24492 16458 24544 16464
rect 24504 16425 24532 16458
rect 24490 16416 24546 16425
rect 24490 16351 24546 16360
rect 24492 16040 24544 16046
rect 24492 15982 24544 15988
rect 24504 15434 24532 15982
rect 24492 15428 24544 15434
rect 24492 15370 24544 15376
rect 24400 15360 24452 15366
rect 24400 15302 24452 15308
rect 24412 13938 24440 15302
rect 24400 13932 24452 13938
rect 24400 13874 24452 13880
rect 24492 12844 24544 12850
rect 24492 12786 24544 12792
rect 24504 12442 24532 12786
rect 24492 12436 24544 12442
rect 24492 12378 24544 12384
rect 24400 11144 24452 11150
rect 24400 11086 24452 11092
rect 24412 9654 24440 11086
rect 24492 10464 24544 10470
rect 24492 10406 24544 10412
rect 24400 9648 24452 9654
rect 24400 9590 24452 9596
rect 24504 9586 24532 10406
rect 24596 9994 24624 17478
rect 24584 9988 24636 9994
rect 24584 9930 24636 9936
rect 24492 9580 24544 9586
rect 24492 9522 24544 9528
rect 24584 9580 24636 9586
rect 24584 9522 24636 9528
rect 24400 9512 24452 9518
rect 24400 9454 24452 9460
rect 24412 9382 24440 9454
rect 24400 9376 24452 9382
rect 24400 9318 24452 9324
rect 24492 9376 24544 9382
rect 24492 9318 24544 9324
rect 24400 9172 24452 9178
rect 24400 9114 24452 9120
rect 24412 8498 24440 9114
rect 24504 9042 24532 9318
rect 24492 9036 24544 9042
rect 24492 8978 24544 8984
rect 24400 8492 24452 8498
rect 24400 8434 24452 8440
rect 24400 8288 24452 8294
rect 24400 8230 24452 8236
rect 24412 7886 24440 8230
rect 24596 8022 24624 9522
rect 24584 8016 24636 8022
rect 24584 7958 24636 7964
rect 24400 7880 24452 7886
rect 24400 7822 24452 7828
rect 24492 7880 24544 7886
rect 24492 7822 24544 7828
rect 24504 6934 24532 7822
rect 24596 7546 24624 7958
rect 24584 7540 24636 7546
rect 24584 7482 24636 7488
rect 24492 6928 24544 6934
rect 24492 6870 24544 6876
rect 24688 2514 24716 22066
rect 24780 19514 24808 22510
rect 24964 22506 24992 22986
rect 24952 22500 25004 22506
rect 24952 22442 25004 22448
rect 24860 22024 24912 22030
rect 24860 21966 24912 21972
rect 24872 21622 24900 21966
rect 24860 21616 24912 21622
rect 24860 21558 24912 21564
rect 24952 21548 25004 21554
rect 24952 21490 25004 21496
rect 24964 20398 24992 21490
rect 25056 20942 25084 23666
rect 25228 22772 25280 22778
rect 25228 22714 25280 22720
rect 25240 22642 25268 22714
rect 25228 22636 25280 22642
rect 25228 22578 25280 22584
rect 25136 22568 25188 22574
rect 25136 22510 25188 22516
rect 25148 22030 25176 22510
rect 25228 22500 25280 22506
rect 25228 22442 25280 22448
rect 25240 22409 25268 22442
rect 25226 22400 25282 22409
rect 25226 22335 25282 22344
rect 25332 22094 25360 48214
rect 25424 48210 25452 48486
rect 25412 48204 25464 48210
rect 25412 48146 25464 48152
rect 25412 47524 25464 47530
rect 25412 47466 25464 47472
rect 25424 46034 25452 47466
rect 25412 46028 25464 46034
rect 25412 45970 25464 45976
rect 25240 22066 25360 22094
rect 25136 22024 25188 22030
rect 25136 21966 25188 21972
rect 25044 20936 25096 20942
rect 25044 20878 25096 20884
rect 25148 20534 25176 21966
rect 25240 21690 25268 22066
rect 25320 21956 25372 21962
rect 25320 21898 25372 21904
rect 25332 21865 25360 21898
rect 25318 21856 25374 21865
rect 25318 21791 25374 21800
rect 25228 21684 25280 21690
rect 25228 21626 25280 21632
rect 25136 20528 25188 20534
rect 25136 20470 25188 20476
rect 24952 20392 25004 20398
rect 24952 20334 25004 20340
rect 24768 19508 24820 19514
rect 24768 19450 24820 19456
rect 24780 16114 24808 19450
rect 25044 19372 25096 19378
rect 25044 19314 25096 19320
rect 25056 18834 25084 19314
rect 25044 18828 25096 18834
rect 25044 18770 25096 18776
rect 24952 18624 25004 18630
rect 24950 18592 24952 18601
rect 25004 18592 25006 18601
rect 25056 18578 25084 18770
rect 25056 18550 25176 18578
rect 24950 18527 25006 18536
rect 24858 18184 24914 18193
rect 24858 18119 24914 18128
rect 24872 17678 24900 18119
rect 24860 17672 24912 17678
rect 24964 17649 24992 18527
rect 25044 18284 25096 18290
rect 25044 18226 25096 18232
rect 25056 17678 25084 18226
rect 25044 17672 25096 17678
rect 24860 17614 24912 17620
rect 24950 17640 25006 17649
rect 25044 17614 25096 17620
rect 24950 17575 25006 17584
rect 24860 17536 24912 17542
rect 24964 17524 24992 17575
rect 24964 17496 25084 17524
rect 24860 17478 24912 17484
rect 24872 16946 24900 17478
rect 24872 16918 24992 16946
rect 24858 16824 24914 16833
rect 24858 16759 24914 16768
rect 24872 16590 24900 16759
rect 24860 16584 24912 16590
rect 24860 16526 24912 16532
rect 24964 16182 24992 16918
rect 24952 16176 25004 16182
rect 24952 16118 25004 16124
rect 24768 16108 24820 16114
rect 24768 16050 24820 16056
rect 24860 15972 24912 15978
rect 24860 15914 24912 15920
rect 24768 15904 24820 15910
rect 24768 15846 24820 15852
rect 24780 15502 24808 15846
rect 24768 15496 24820 15502
rect 24872 15484 24900 15914
rect 24964 15706 24992 16118
rect 25056 15910 25084 17496
rect 25148 17134 25176 18550
rect 25320 18284 25372 18290
rect 25320 18226 25372 18232
rect 25228 17876 25280 17882
rect 25228 17818 25280 17824
rect 25240 17542 25268 17818
rect 25228 17536 25280 17542
rect 25228 17478 25280 17484
rect 25136 17128 25188 17134
rect 25136 17070 25188 17076
rect 25228 17060 25280 17066
rect 25228 17002 25280 17008
rect 25240 16726 25268 17002
rect 25228 16720 25280 16726
rect 25228 16662 25280 16668
rect 25044 15904 25096 15910
rect 25044 15846 25096 15852
rect 24952 15700 25004 15706
rect 24952 15642 25004 15648
rect 24952 15496 25004 15502
rect 24872 15456 24952 15484
rect 24768 15438 24820 15444
rect 24952 15438 25004 15444
rect 24768 14544 24820 14550
rect 24768 14486 24820 14492
rect 24780 13870 24808 14486
rect 24768 13864 24820 13870
rect 24768 13806 24820 13812
rect 24780 11830 24808 13806
rect 24768 11824 24820 11830
rect 24768 11766 24820 11772
rect 24860 10668 24912 10674
rect 24860 10610 24912 10616
rect 24768 9920 24820 9926
rect 24768 9862 24820 9868
rect 24780 9654 24808 9862
rect 24872 9722 24900 10610
rect 24964 10606 24992 15438
rect 25136 14816 25188 14822
rect 25136 14758 25188 14764
rect 25148 14278 25176 14758
rect 25136 14272 25188 14278
rect 25136 14214 25188 14220
rect 25228 13728 25280 13734
rect 25228 13670 25280 13676
rect 25240 13326 25268 13670
rect 25228 13320 25280 13326
rect 25228 13262 25280 13268
rect 25136 13252 25188 13258
rect 25136 13194 25188 13200
rect 25044 13184 25096 13190
rect 25044 13126 25096 13132
rect 24952 10600 25004 10606
rect 24952 10542 25004 10548
rect 25056 10452 25084 13126
rect 25148 12850 25176 13194
rect 25136 12844 25188 12850
rect 25136 12786 25188 12792
rect 25134 12744 25190 12753
rect 25134 12679 25136 12688
rect 25188 12679 25190 12688
rect 25136 12650 25188 12656
rect 25136 11348 25188 11354
rect 25136 11290 25188 11296
rect 24964 10424 25084 10452
rect 24964 10130 24992 10424
rect 24952 10124 25004 10130
rect 24952 10066 25004 10072
rect 25148 9926 25176 11290
rect 25228 11144 25280 11150
rect 25228 11086 25280 11092
rect 25240 10742 25268 11086
rect 25228 10736 25280 10742
rect 25228 10678 25280 10684
rect 25240 10266 25268 10678
rect 25228 10260 25280 10266
rect 25228 10202 25280 10208
rect 25136 9920 25188 9926
rect 25136 9862 25188 9868
rect 24860 9716 24912 9722
rect 24860 9658 24912 9664
rect 24768 9648 24820 9654
rect 24768 9590 24820 9596
rect 24780 9110 24808 9590
rect 24860 9580 24912 9586
rect 24860 9522 24912 9528
rect 24768 9104 24820 9110
rect 24768 9046 24820 9052
rect 24872 8956 24900 9522
rect 25148 9518 25176 9862
rect 25136 9512 25188 9518
rect 25136 9454 25188 9460
rect 24780 8928 24900 8956
rect 24780 8634 24808 8928
rect 24768 8628 24820 8634
rect 24768 8570 24820 8576
rect 25332 7818 25360 18226
rect 25424 10282 25452 45970
rect 25516 24070 25544 48486
rect 26700 47592 26752 47598
rect 26700 47534 26752 47540
rect 26712 47258 26740 47534
rect 26148 47252 26200 47258
rect 26148 47194 26200 47200
rect 26700 47252 26752 47258
rect 26700 47194 26752 47200
rect 26160 45490 26188 47194
rect 26148 45484 26200 45490
rect 26148 45426 26200 45432
rect 25596 44736 25648 44742
rect 25596 44678 25648 44684
rect 25608 31754 25636 44678
rect 25688 42696 25740 42702
rect 25688 42638 25740 42644
rect 25700 42362 25728 42638
rect 26148 42560 26200 42566
rect 26148 42502 26200 42508
rect 26516 42560 26568 42566
rect 26516 42502 26568 42508
rect 25688 42356 25740 42362
rect 25688 42298 25740 42304
rect 25964 42016 26016 42022
rect 25964 41958 26016 41964
rect 25976 41682 26004 41958
rect 26160 41818 26188 42502
rect 26148 41812 26200 41818
rect 26148 41754 26200 41760
rect 25964 41676 26016 41682
rect 25964 41618 26016 41624
rect 26528 41614 26556 42502
rect 26516 41608 26568 41614
rect 26516 41550 26568 41556
rect 26516 41472 26568 41478
rect 26516 41414 26568 41420
rect 25780 40044 25832 40050
rect 25780 39986 25832 39992
rect 26056 40044 26108 40050
rect 26056 39986 26108 39992
rect 25688 38956 25740 38962
rect 25688 38898 25740 38904
rect 25700 38554 25728 38898
rect 25688 38548 25740 38554
rect 25688 38490 25740 38496
rect 25792 38486 25820 39986
rect 25964 39840 26016 39846
rect 25964 39782 26016 39788
rect 25976 39438 26004 39782
rect 25964 39432 26016 39438
rect 25964 39374 26016 39380
rect 26068 39098 26096 39986
rect 26424 39432 26476 39438
rect 26424 39374 26476 39380
rect 26436 39098 26464 39374
rect 26056 39092 26108 39098
rect 26056 39034 26108 39040
rect 26424 39092 26476 39098
rect 26424 39034 26476 39040
rect 25872 38956 25924 38962
rect 25872 38898 25924 38904
rect 25780 38480 25832 38486
rect 25780 38422 25832 38428
rect 25792 38010 25820 38422
rect 25780 38004 25832 38010
rect 25780 37946 25832 37952
rect 25884 37890 25912 38898
rect 26068 38214 26096 39034
rect 26056 38208 26108 38214
rect 26056 38150 26108 38156
rect 25792 37862 25912 37890
rect 26240 37936 26292 37942
rect 26240 37878 26292 37884
rect 25792 37194 25820 37862
rect 25780 37188 25832 37194
rect 25780 37130 25832 37136
rect 26056 37188 26108 37194
rect 26056 37130 26108 37136
rect 26068 36378 26096 37130
rect 26252 37074 26280 37878
rect 26424 37868 26476 37874
rect 26424 37810 26476 37816
rect 26332 37664 26384 37670
rect 26332 37606 26384 37612
rect 26344 37194 26372 37606
rect 26332 37188 26384 37194
rect 26332 37130 26384 37136
rect 26252 37046 26372 37074
rect 26056 36372 26108 36378
rect 26056 36314 26108 36320
rect 26240 36100 26292 36106
rect 26240 36042 26292 36048
rect 26252 35630 26280 36042
rect 26240 35624 26292 35630
rect 26240 35566 26292 35572
rect 26240 35080 26292 35086
rect 26240 35022 26292 35028
rect 26252 34610 26280 35022
rect 26344 35018 26372 37046
rect 26436 35766 26464 37810
rect 26424 35760 26476 35766
rect 26424 35702 26476 35708
rect 26332 35012 26384 35018
rect 26332 34954 26384 34960
rect 26240 34604 26292 34610
rect 26240 34546 26292 34552
rect 25688 34400 25740 34406
rect 25688 34342 25740 34348
rect 25700 34134 25728 34342
rect 25688 34128 25740 34134
rect 25688 34070 25740 34076
rect 25700 33862 25728 34070
rect 25688 33856 25740 33862
rect 25688 33798 25740 33804
rect 26436 33590 26464 35702
rect 26528 34678 26556 41414
rect 26700 37256 26752 37262
rect 26700 37198 26752 37204
rect 26712 36922 26740 37198
rect 26700 36916 26752 36922
rect 26700 36858 26752 36864
rect 26608 36032 26660 36038
rect 26608 35974 26660 35980
rect 26620 35766 26648 35974
rect 26608 35760 26660 35766
rect 26608 35702 26660 35708
rect 26712 35698 26740 36858
rect 26700 35692 26752 35698
rect 26700 35634 26752 35640
rect 26516 34672 26568 34678
rect 26516 34614 26568 34620
rect 26424 33584 26476 33590
rect 26424 33526 26476 33532
rect 25780 33516 25832 33522
rect 25780 33458 25832 33464
rect 25792 32774 25820 33458
rect 25780 32768 25832 32774
rect 25780 32710 25832 32716
rect 25686 32600 25742 32609
rect 25686 32535 25742 32544
rect 25700 32026 25728 32535
rect 25792 32502 25820 32710
rect 25780 32496 25832 32502
rect 25780 32438 25832 32444
rect 26436 32434 26464 33526
rect 26424 32428 26476 32434
rect 26424 32370 26476 32376
rect 25780 32292 25832 32298
rect 25780 32234 25832 32240
rect 25792 32065 25820 32234
rect 26148 32224 26200 32230
rect 26148 32166 26200 32172
rect 25778 32056 25834 32065
rect 25688 32020 25740 32026
rect 25778 31991 25834 32000
rect 25688 31962 25740 31968
rect 25608 31726 25728 31754
rect 25596 30048 25648 30054
rect 25596 29990 25648 29996
rect 25608 29646 25636 29990
rect 25596 29640 25648 29646
rect 25596 29582 25648 29588
rect 25594 27024 25650 27033
rect 25594 26959 25596 26968
rect 25648 26959 25650 26968
rect 25596 26930 25648 26936
rect 25608 26790 25636 26930
rect 25596 26784 25648 26790
rect 25596 26726 25648 26732
rect 25504 24064 25556 24070
rect 25504 24006 25556 24012
rect 25504 23792 25556 23798
rect 25504 23734 25556 23740
rect 25516 23662 25544 23734
rect 25596 23724 25648 23730
rect 25596 23666 25648 23672
rect 25504 23656 25556 23662
rect 25504 23598 25556 23604
rect 25516 22642 25544 23598
rect 25608 23322 25636 23666
rect 25596 23316 25648 23322
rect 25596 23258 25648 23264
rect 25504 22636 25556 22642
rect 25504 22578 25556 22584
rect 25502 22128 25558 22137
rect 25502 22063 25558 22072
rect 25516 22030 25544 22063
rect 25504 22024 25556 22030
rect 25504 21966 25556 21972
rect 25596 18080 25648 18086
rect 25596 18022 25648 18028
rect 25608 17882 25636 18022
rect 25596 17876 25648 17882
rect 25596 17818 25648 17824
rect 25504 17672 25556 17678
rect 25504 17614 25556 17620
rect 25516 17202 25544 17614
rect 25608 17241 25636 17818
rect 25594 17232 25650 17241
rect 25504 17196 25556 17202
rect 25594 17167 25596 17176
rect 25504 17138 25556 17144
rect 25648 17167 25650 17176
rect 25596 17138 25648 17144
rect 25516 16454 25544 17138
rect 25608 17107 25636 17138
rect 25504 16448 25556 16454
rect 25504 16390 25556 16396
rect 25504 15156 25556 15162
rect 25504 15098 25556 15104
rect 25516 14074 25544 15098
rect 25504 14068 25556 14074
rect 25504 14010 25556 14016
rect 25504 11552 25556 11558
rect 25504 11494 25556 11500
rect 25516 11150 25544 11494
rect 25504 11144 25556 11150
rect 25504 11086 25556 11092
rect 25504 10668 25556 10674
rect 25504 10610 25556 10616
rect 25516 10452 25544 10610
rect 25516 10424 25636 10452
rect 25424 10254 25544 10282
rect 25412 10192 25464 10198
rect 25412 10134 25464 10140
rect 25424 9654 25452 10134
rect 25412 9648 25464 9654
rect 25412 9590 25464 9596
rect 25412 9512 25464 9518
rect 25412 9454 25464 9460
rect 25424 8974 25452 9454
rect 25412 8968 25464 8974
rect 25412 8910 25464 8916
rect 25320 7812 25372 7818
rect 25320 7754 25372 7760
rect 25136 7744 25188 7750
rect 25136 7686 25188 7692
rect 25148 7478 25176 7686
rect 25136 7472 25188 7478
rect 25136 7414 25188 7420
rect 24768 6724 24820 6730
rect 24768 6666 24820 6672
rect 24780 5370 24808 6666
rect 24768 5364 24820 5370
rect 24768 5306 24820 5312
rect 25516 3398 25544 10254
rect 25608 10198 25636 10424
rect 25596 10192 25648 10198
rect 25596 10134 25648 10140
rect 25700 3466 25728 31726
rect 26160 31346 26188 32166
rect 26240 31680 26292 31686
rect 26240 31622 26292 31628
rect 26252 31346 26280 31622
rect 26148 31340 26200 31346
rect 26148 31282 26200 31288
rect 26240 31340 26292 31346
rect 26240 31282 26292 31288
rect 25780 31136 25832 31142
rect 25780 31078 25832 31084
rect 25792 30666 25820 31078
rect 25780 30660 25832 30666
rect 25780 30602 25832 30608
rect 26056 28416 26108 28422
rect 26056 28358 26108 28364
rect 25780 27940 25832 27946
rect 25780 27882 25832 27888
rect 25792 22982 25820 27882
rect 26068 27606 26096 28358
rect 26056 27600 26108 27606
rect 26056 27542 26108 27548
rect 26068 27402 26096 27542
rect 26056 27396 26108 27402
rect 26056 27338 26108 27344
rect 26528 26994 26556 34614
rect 26056 26988 26108 26994
rect 26056 26930 26108 26936
rect 26516 26988 26568 26994
rect 26516 26930 26568 26936
rect 26068 26586 26096 26930
rect 26056 26580 26108 26586
rect 26056 26522 26108 26528
rect 26804 26330 26832 48826
rect 26884 47660 26936 47666
rect 26884 47602 26936 47608
rect 26896 43790 26924 47602
rect 26988 46578 27016 49166
rect 27160 49156 27212 49162
rect 27160 49098 27212 49104
rect 27172 47666 27200 49098
rect 27620 48612 27672 48618
rect 27620 48554 27672 48560
rect 27160 47660 27212 47666
rect 27160 47602 27212 47608
rect 27528 47592 27580 47598
rect 27528 47534 27580 47540
rect 27540 47054 27568 47534
rect 27528 47048 27580 47054
rect 27528 46990 27580 46996
rect 26976 46572 27028 46578
rect 26976 46514 27028 46520
rect 26884 43784 26936 43790
rect 26884 43726 26936 43732
rect 27160 43308 27212 43314
rect 27160 43250 27212 43256
rect 27436 43308 27488 43314
rect 27436 43250 27488 43256
rect 26976 43104 27028 43110
rect 26976 43046 27028 43052
rect 26988 42702 27016 43046
rect 26884 42696 26936 42702
rect 26884 42638 26936 42644
rect 26976 42696 27028 42702
rect 26976 42638 27028 42644
rect 26896 41206 26924 42638
rect 27172 41478 27200 43250
rect 27448 41818 27476 43250
rect 27528 42696 27580 42702
rect 27528 42638 27580 42644
rect 27436 41812 27488 41818
rect 27436 41754 27488 41760
rect 27448 41698 27476 41754
rect 27356 41670 27476 41698
rect 27160 41472 27212 41478
rect 27160 41414 27212 41420
rect 26884 41200 26936 41206
rect 26884 41142 26936 41148
rect 27356 40730 27384 41670
rect 27540 41546 27568 42638
rect 27528 41540 27580 41546
rect 27528 41482 27580 41488
rect 27540 41414 27568 41482
rect 27448 41386 27568 41414
rect 27448 41002 27476 41386
rect 27436 40996 27488 41002
rect 27436 40938 27488 40944
rect 27344 40724 27396 40730
rect 27344 40666 27396 40672
rect 26976 40112 27028 40118
rect 26976 40054 27028 40060
rect 26988 39098 27016 40054
rect 27252 39500 27304 39506
rect 27252 39442 27304 39448
rect 27160 39364 27212 39370
rect 27160 39306 27212 39312
rect 26976 39092 27028 39098
rect 26976 39034 27028 39040
rect 27172 38486 27200 39306
rect 27160 38480 27212 38486
rect 27160 38422 27212 38428
rect 26976 37188 27028 37194
rect 26976 37130 27028 37136
rect 26988 36854 27016 37130
rect 26976 36848 27028 36854
rect 26976 36790 27028 36796
rect 27068 36848 27120 36854
rect 27068 36790 27120 36796
rect 26884 36712 26936 36718
rect 26884 36654 26936 36660
rect 26896 35630 26924 36654
rect 27080 36174 27108 36790
rect 27264 36242 27292 39442
rect 27436 39296 27488 39302
rect 27436 39238 27488 39244
rect 27448 38962 27476 39238
rect 27436 38956 27488 38962
rect 27436 38898 27488 38904
rect 27448 38010 27476 38898
rect 27436 38004 27488 38010
rect 27436 37946 27488 37952
rect 27344 37868 27396 37874
rect 27344 37810 27396 37816
rect 27356 37262 27384 37810
rect 27528 37800 27580 37806
rect 27528 37742 27580 37748
rect 27344 37256 27396 37262
rect 27344 37198 27396 37204
rect 27436 37120 27488 37126
rect 27436 37062 27488 37068
rect 27448 36786 27476 37062
rect 27436 36780 27488 36786
rect 27436 36722 27488 36728
rect 27540 36242 27568 37742
rect 27632 36530 27660 48554
rect 27724 48210 27752 51200
rect 27712 48204 27764 48210
rect 27712 48146 27764 48152
rect 28080 48136 28132 48142
rect 28080 48078 28132 48084
rect 28092 47666 28120 48078
rect 28172 48068 28224 48074
rect 28172 48010 28224 48016
rect 28080 47660 28132 47666
rect 28080 47602 28132 47608
rect 28184 47546 28212 48010
rect 28092 47518 28212 47546
rect 28368 47530 28396 51200
rect 29012 48822 29040 51200
rect 29000 48816 29052 48822
rect 29000 48758 29052 48764
rect 29656 48686 29684 51200
rect 30944 49298 30972 51200
rect 30564 49292 30616 49298
rect 30564 49234 30616 49240
rect 30932 49292 30984 49298
rect 30932 49234 30984 49240
rect 29920 49156 29972 49162
rect 29920 49098 29972 49104
rect 29368 48680 29420 48686
rect 29368 48622 29420 48628
rect 29644 48680 29696 48686
rect 29644 48622 29696 48628
rect 29276 48612 29328 48618
rect 29276 48554 29328 48560
rect 28448 48544 28500 48550
rect 28448 48486 28500 48492
rect 28356 47524 28408 47530
rect 28092 46374 28120 47518
rect 28356 47466 28408 47472
rect 28264 47048 28316 47054
rect 28264 46990 28316 46996
rect 28080 46368 28132 46374
rect 28080 46310 28132 46316
rect 27988 42696 28040 42702
rect 27988 42638 28040 42644
rect 27896 42628 27948 42634
rect 27896 42570 27948 42576
rect 27804 42560 27856 42566
rect 27804 42502 27856 42508
rect 27816 42226 27844 42502
rect 27804 42220 27856 42226
rect 27804 42162 27856 42168
rect 27712 42084 27764 42090
rect 27712 42026 27764 42032
rect 27724 41682 27752 42026
rect 27908 41818 27936 42570
rect 28000 42226 28028 42638
rect 27988 42220 28040 42226
rect 27988 42162 28040 42168
rect 27896 41812 27948 41818
rect 27896 41754 27948 41760
rect 27712 41676 27764 41682
rect 27712 41618 27764 41624
rect 27724 41414 27752 41618
rect 28092 41414 28120 46310
rect 27724 41386 27844 41414
rect 27816 38554 27844 41386
rect 27908 41386 28120 41414
rect 27804 38548 27856 38554
rect 27804 38490 27856 38496
rect 27632 36502 27844 36530
rect 27252 36236 27304 36242
rect 27252 36178 27304 36184
rect 27528 36236 27580 36242
rect 27528 36178 27580 36184
rect 27068 36168 27120 36174
rect 27068 36110 27120 36116
rect 26884 35624 26936 35630
rect 26884 35566 26936 35572
rect 27540 35290 27568 36178
rect 27528 35284 27580 35290
rect 27528 35226 27580 35232
rect 26976 35012 27028 35018
rect 26976 34954 27028 34960
rect 26884 34060 26936 34066
rect 26884 34002 26936 34008
rect 26896 33386 26924 34002
rect 26884 33380 26936 33386
rect 26884 33322 26936 33328
rect 26896 33153 26924 33322
rect 26882 33144 26938 33153
rect 26882 33079 26938 33088
rect 26896 32366 26924 33079
rect 26884 32360 26936 32366
rect 26884 32302 26936 32308
rect 26884 32224 26936 32230
rect 26884 32166 26936 32172
rect 26896 31822 26924 32166
rect 26884 31816 26936 31822
rect 26884 31758 26936 31764
rect 26988 31278 27016 34954
rect 27712 33992 27764 33998
rect 27712 33934 27764 33940
rect 27436 33924 27488 33930
rect 27436 33866 27488 33872
rect 27160 33856 27212 33862
rect 27160 33798 27212 33804
rect 27172 32910 27200 33798
rect 27448 33658 27476 33866
rect 27436 33652 27488 33658
rect 27436 33594 27488 33600
rect 27724 33590 27752 33934
rect 27712 33584 27764 33590
rect 27712 33526 27764 33532
rect 27068 32904 27120 32910
rect 27068 32846 27120 32852
rect 27160 32904 27212 32910
rect 27160 32846 27212 32852
rect 27620 32904 27672 32910
rect 27620 32846 27672 32852
rect 26976 31272 27028 31278
rect 26976 31214 27028 31220
rect 27080 30734 27108 32846
rect 27632 32570 27660 32846
rect 27620 32564 27672 32570
rect 27620 32506 27672 32512
rect 27724 32434 27752 33526
rect 27344 32428 27396 32434
rect 27344 32370 27396 32376
rect 27712 32428 27764 32434
rect 27712 32370 27764 32376
rect 27252 31272 27304 31278
rect 27252 31214 27304 31220
rect 27068 30728 27120 30734
rect 27068 30670 27120 30676
rect 27160 30592 27212 30598
rect 27160 30534 27212 30540
rect 27172 26450 27200 30534
rect 27264 29714 27292 31214
rect 27356 31210 27384 32370
rect 27620 32224 27672 32230
rect 27620 32166 27672 32172
rect 27528 31748 27580 31754
rect 27528 31690 27580 31696
rect 27436 31680 27488 31686
rect 27436 31622 27488 31628
rect 27344 31204 27396 31210
rect 27344 31146 27396 31152
rect 27448 30598 27476 31622
rect 27540 31278 27568 31690
rect 27528 31272 27580 31278
rect 27528 31214 27580 31220
rect 27540 30870 27568 31214
rect 27528 30864 27580 30870
rect 27528 30806 27580 30812
rect 27528 30728 27580 30734
rect 27528 30670 27580 30676
rect 27436 30592 27488 30598
rect 27436 30534 27488 30540
rect 27540 30394 27568 30670
rect 27528 30388 27580 30394
rect 27528 30330 27580 30336
rect 27344 30252 27396 30258
rect 27344 30194 27396 30200
rect 27252 29708 27304 29714
rect 27252 29650 27304 29656
rect 27356 29170 27384 30194
rect 27540 30190 27568 30330
rect 27632 30258 27660 32166
rect 27724 31346 27752 32370
rect 27712 31340 27764 31346
rect 27712 31282 27764 31288
rect 27620 30252 27672 30258
rect 27620 30194 27672 30200
rect 27528 30184 27580 30190
rect 27528 30126 27580 30132
rect 27344 29164 27396 29170
rect 27344 29106 27396 29112
rect 27160 26444 27212 26450
rect 27160 26386 27212 26392
rect 26804 26302 27292 26330
rect 26240 26240 26292 26246
rect 26240 26182 26292 26188
rect 25872 26036 25924 26042
rect 25872 25978 25924 25984
rect 25884 25906 25912 25978
rect 25872 25900 25924 25906
rect 25872 25842 25924 25848
rect 26056 25900 26108 25906
rect 26056 25842 26108 25848
rect 26068 25498 26096 25842
rect 26252 25838 26280 26182
rect 26884 25900 26936 25906
rect 26884 25842 26936 25848
rect 26240 25832 26292 25838
rect 26240 25774 26292 25780
rect 26056 25492 26108 25498
rect 26056 25434 26108 25440
rect 25872 25356 25924 25362
rect 25872 25298 25924 25304
rect 25884 24818 25912 25298
rect 26896 25294 26924 25842
rect 26884 25288 26936 25294
rect 26884 25230 26936 25236
rect 26896 24818 26924 25230
rect 27160 25152 27212 25158
rect 27160 25094 27212 25100
rect 25872 24812 25924 24818
rect 25872 24754 25924 24760
rect 26884 24812 26936 24818
rect 26884 24754 26936 24760
rect 25884 23526 25912 24754
rect 26240 24744 26292 24750
rect 26068 24704 26240 24732
rect 26068 24614 26096 24704
rect 26240 24686 26292 24692
rect 26332 24676 26384 24682
rect 26332 24618 26384 24624
rect 26056 24608 26108 24614
rect 26056 24550 26108 24556
rect 26068 24154 26096 24550
rect 26344 24342 26372 24618
rect 26332 24336 26384 24342
rect 26332 24278 26384 24284
rect 26148 24200 26200 24206
rect 25976 24148 26148 24154
rect 25976 24142 26200 24148
rect 25976 24126 26188 24142
rect 27068 24132 27120 24138
rect 25872 23520 25924 23526
rect 25872 23462 25924 23468
rect 25872 23316 25924 23322
rect 25872 23258 25924 23264
rect 25780 22976 25832 22982
rect 25780 22918 25832 22924
rect 25884 22642 25912 23258
rect 25872 22636 25924 22642
rect 25872 22578 25924 22584
rect 25976 22094 26004 24126
rect 27068 24074 27120 24080
rect 26056 24064 26108 24070
rect 26056 24006 26108 24012
rect 26792 24064 26844 24070
rect 26792 24006 26844 24012
rect 25884 22066 26004 22094
rect 26068 22094 26096 24006
rect 26804 23118 26832 24006
rect 27080 23322 27108 24074
rect 27068 23316 27120 23322
rect 27068 23258 27120 23264
rect 26792 23112 26844 23118
rect 26792 23054 26844 23060
rect 27068 23112 27120 23118
rect 27068 23054 27120 23060
rect 26700 22772 26752 22778
rect 26700 22714 26752 22720
rect 26148 22704 26200 22710
rect 26148 22646 26200 22652
rect 26160 22438 26188 22646
rect 26148 22432 26200 22438
rect 26148 22374 26200 22380
rect 26712 22166 26740 22714
rect 26700 22160 26752 22166
rect 26700 22102 26752 22108
rect 26332 22094 26384 22098
rect 26068 22066 26280 22094
rect 25780 21140 25832 21146
rect 25780 21082 25832 21088
rect 25792 20942 25820 21082
rect 25780 20936 25832 20942
rect 25780 20878 25832 20884
rect 25884 18290 25912 22066
rect 26068 21690 26096 22066
rect 26252 22030 26280 22066
rect 26332 22092 26648 22094
rect 26384 22066 26648 22092
rect 26332 22034 26384 22040
rect 26240 22024 26292 22030
rect 26424 22024 26476 22030
rect 26240 21966 26292 21972
rect 26344 21972 26424 21978
rect 26344 21966 26476 21972
rect 26344 21950 26464 21966
rect 26240 21888 26292 21894
rect 26240 21830 26292 21836
rect 26252 21690 26280 21830
rect 26056 21684 26108 21690
rect 26056 21626 26108 21632
rect 26240 21684 26292 21690
rect 26240 21626 26292 21632
rect 26054 21584 26110 21593
rect 26054 21519 26056 21528
rect 26108 21519 26110 21528
rect 26148 21548 26200 21554
rect 26056 21490 26108 21496
rect 26148 21490 26200 21496
rect 26160 20942 26188 21490
rect 26344 21486 26372 21950
rect 26424 21888 26476 21894
rect 26424 21830 26476 21836
rect 26516 21888 26568 21894
rect 26516 21830 26568 21836
rect 26436 21622 26464 21830
rect 26424 21616 26476 21622
rect 26528 21593 26556 21830
rect 26620 21729 26648 22066
rect 26606 21720 26662 21729
rect 26606 21655 26662 21664
rect 26424 21558 26476 21564
rect 26514 21584 26570 21593
rect 26514 21519 26570 21528
rect 26332 21480 26384 21486
rect 26332 21422 26384 21428
rect 26424 21480 26476 21486
rect 26424 21422 26476 21428
rect 26698 21448 26754 21457
rect 26148 20936 26200 20942
rect 26148 20878 26200 20884
rect 26240 20868 26292 20874
rect 26436 20856 26464 21422
rect 26698 21383 26754 21392
rect 26712 21078 26740 21383
rect 26700 21072 26752 21078
rect 26700 21014 26752 21020
rect 26292 20828 26464 20856
rect 26240 20810 26292 20816
rect 26240 19848 26292 19854
rect 26240 19790 26292 19796
rect 26252 19310 26280 19790
rect 26240 19304 26292 19310
rect 26240 19246 26292 19252
rect 26804 18766 26832 23054
rect 26882 22536 26938 22545
rect 26882 22471 26938 22480
rect 26896 22166 26924 22471
rect 26884 22160 26936 22166
rect 26884 22102 26936 22108
rect 26884 21616 26936 21622
rect 26884 21558 26936 21564
rect 26896 21010 26924 21558
rect 26976 21412 27028 21418
rect 26976 21354 27028 21360
rect 26988 21321 27016 21354
rect 26974 21312 27030 21321
rect 26974 21247 27030 21256
rect 26884 21004 26936 21010
rect 26884 20946 26936 20952
rect 26976 19712 27028 19718
rect 26976 19654 27028 19660
rect 26988 19446 27016 19654
rect 26976 19440 27028 19446
rect 26976 19382 27028 19388
rect 26988 18766 27016 19382
rect 27080 19310 27108 23054
rect 27172 19446 27200 25094
rect 27264 22094 27292 26302
rect 27356 25242 27384 29106
rect 27436 28416 27488 28422
rect 27436 28358 27488 28364
rect 27448 27033 27476 28358
rect 27540 28014 27568 30126
rect 27620 29232 27672 29238
rect 27620 29174 27672 29180
rect 27632 28558 27660 29174
rect 27620 28552 27672 28558
rect 27620 28494 27672 28500
rect 27620 28076 27672 28082
rect 27620 28018 27672 28024
rect 27528 28008 27580 28014
rect 27528 27950 27580 27956
rect 27632 27606 27660 28018
rect 27620 27600 27672 27606
rect 27620 27542 27672 27548
rect 27712 27600 27764 27606
rect 27712 27542 27764 27548
rect 27724 27130 27752 27542
rect 27712 27124 27764 27130
rect 27712 27066 27764 27072
rect 27434 27024 27490 27033
rect 27434 26959 27490 26968
rect 27712 25764 27764 25770
rect 27712 25706 27764 25712
rect 27620 25696 27672 25702
rect 27620 25638 27672 25644
rect 27632 25498 27660 25638
rect 27724 25498 27752 25706
rect 27620 25492 27672 25498
rect 27620 25434 27672 25440
rect 27712 25492 27764 25498
rect 27712 25434 27764 25440
rect 27356 25214 27476 25242
rect 27344 25152 27396 25158
rect 27344 25094 27396 25100
rect 27356 24818 27384 25094
rect 27344 24812 27396 24818
rect 27344 24754 27396 24760
rect 27448 23118 27476 25214
rect 27712 24880 27764 24886
rect 27712 24822 27764 24828
rect 27528 24064 27580 24070
rect 27528 24006 27580 24012
rect 27540 23730 27568 24006
rect 27724 23746 27752 24822
rect 27816 24750 27844 36502
rect 27908 27962 27936 41386
rect 27988 39432 28040 39438
rect 27988 39374 28040 39380
rect 28000 38894 28028 39374
rect 28080 39364 28132 39370
rect 28080 39306 28132 39312
rect 28092 39098 28120 39306
rect 28080 39092 28132 39098
rect 28080 39034 28132 39040
rect 27988 38888 28040 38894
rect 27988 38830 28040 38836
rect 28080 37868 28132 37874
rect 28080 37810 28132 37816
rect 27988 37188 28040 37194
rect 27988 37130 28040 37136
rect 28000 36854 28028 37130
rect 28092 37126 28120 37810
rect 28080 37120 28132 37126
rect 28080 37062 28132 37068
rect 27988 36848 28040 36854
rect 27988 36790 28040 36796
rect 28172 36848 28224 36854
rect 28172 36790 28224 36796
rect 28184 36378 28212 36790
rect 28080 36372 28132 36378
rect 28080 36314 28132 36320
rect 28172 36372 28224 36378
rect 28172 36314 28224 36320
rect 28092 36258 28120 36314
rect 27988 36236 28040 36242
rect 28092 36230 28212 36258
rect 27988 36178 28040 36184
rect 28000 35834 28028 36178
rect 28184 36106 28212 36230
rect 28172 36100 28224 36106
rect 28172 36042 28224 36048
rect 27988 35828 28040 35834
rect 27988 35770 28040 35776
rect 28184 35630 28212 36042
rect 28172 35624 28224 35630
rect 28172 35566 28224 35572
rect 28184 35154 28212 35566
rect 28172 35148 28224 35154
rect 28172 35090 28224 35096
rect 28172 34536 28224 34542
rect 28172 34478 28224 34484
rect 28184 33998 28212 34478
rect 28172 33992 28224 33998
rect 28172 33934 28224 33940
rect 27988 33516 28040 33522
rect 27988 33458 28040 33464
rect 28172 33516 28224 33522
rect 28172 33458 28224 33464
rect 28000 32774 28028 33458
rect 28080 33448 28132 33454
rect 28080 33390 28132 33396
rect 27988 32768 28040 32774
rect 27988 32710 28040 32716
rect 28092 32570 28120 33390
rect 28080 32564 28132 32570
rect 28080 32506 28132 32512
rect 28184 32450 28212 33458
rect 28000 32422 28212 32450
rect 28000 31754 28028 32422
rect 28172 32224 28224 32230
rect 28172 32166 28224 32172
rect 28000 31726 28120 31754
rect 28092 29238 28120 31726
rect 28184 31226 28212 32166
rect 28276 31346 28304 46990
rect 28356 36168 28408 36174
rect 28356 36110 28408 36116
rect 28368 35834 28396 36110
rect 28356 35828 28408 35834
rect 28356 35770 28408 35776
rect 28368 33658 28396 35770
rect 28356 33652 28408 33658
rect 28356 33594 28408 33600
rect 28356 32360 28408 32366
rect 28356 32302 28408 32308
rect 28264 31340 28316 31346
rect 28264 31282 28316 31288
rect 28184 31198 28304 31226
rect 28172 31136 28224 31142
rect 28172 31078 28224 31084
rect 28184 30734 28212 31078
rect 28172 30728 28224 30734
rect 28172 30670 28224 30676
rect 28172 29640 28224 29646
rect 28172 29582 28224 29588
rect 28080 29232 28132 29238
rect 28080 29174 28132 29180
rect 27988 29164 28040 29170
rect 27988 29106 28040 29112
rect 28000 28762 28028 29106
rect 28092 28966 28120 29174
rect 28184 29034 28212 29582
rect 28172 29028 28224 29034
rect 28172 28970 28224 28976
rect 28080 28960 28132 28966
rect 28080 28902 28132 28908
rect 27988 28756 28040 28762
rect 27988 28698 28040 28704
rect 27908 27934 28212 27962
rect 27896 27872 27948 27878
rect 27896 27814 27948 27820
rect 27908 25838 27936 27814
rect 27988 27464 28040 27470
rect 27988 27406 28040 27412
rect 28000 27033 28028 27406
rect 27986 27024 28042 27033
rect 27986 26959 27988 26968
rect 28040 26959 28042 26968
rect 27988 26930 28040 26936
rect 27988 26784 28040 26790
rect 27988 26726 28040 26732
rect 28000 25906 28028 26726
rect 27988 25900 28040 25906
rect 27988 25842 28040 25848
rect 27896 25832 27948 25838
rect 27896 25774 27948 25780
rect 27908 24750 27936 25774
rect 27804 24744 27856 24750
rect 27804 24686 27856 24692
rect 27896 24744 27948 24750
rect 27896 24686 27948 24692
rect 27804 24608 27856 24614
rect 27804 24550 27856 24556
rect 27816 23866 27844 24550
rect 27908 24206 27936 24686
rect 28080 24608 28132 24614
rect 28080 24550 28132 24556
rect 27896 24200 27948 24206
rect 27896 24142 27948 24148
rect 27804 23860 27856 23866
rect 27804 23802 27856 23808
rect 27896 23860 27948 23866
rect 27896 23802 27948 23808
rect 27908 23746 27936 23802
rect 27528 23724 27580 23730
rect 27724 23718 27936 23746
rect 27528 23666 27580 23672
rect 27712 23588 27764 23594
rect 27712 23530 27764 23536
rect 27436 23112 27488 23118
rect 27436 23054 27488 23060
rect 27264 22066 27568 22094
rect 27252 21888 27304 21894
rect 27252 21830 27304 21836
rect 27264 21554 27292 21830
rect 27342 21584 27398 21593
rect 27252 21548 27304 21554
rect 27342 21519 27398 21528
rect 27252 21490 27304 21496
rect 27264 20874 27292 21490
rect 27356 21486 27384 21519
rect 27344 21480 27396 21486
rect 27344 21422 27396 21428
rect 27344 21344 27396 21350
rect 27344 21286 27396 21292
rect 27356 21162 27384 21286
rect 27356 21146 27476 21162
rect 27540 21146 27568 22066
rect 27620 21480 27672 21486
rect 27620 21422 27672 21428
rect 27356 21140 27488 21146
rect 27356 21134 27436 21140
rect 27436 21082 27488 21088
rect 27528 21140 27580 21146
rect 27528 21082 27580 21088
rect 27448 20913 27476 21082
rect 27632 21010 27660 21422
rect 27620 21004 27672 21010
rect 27620 20946 27672 20952
rect 27434 20904 27490 20913
rect 27252 20868 27304 20874
rect 27434 20839 27490 20848
rect 27252 20810 27304 20816
rect 27724 19922 27752 23530
rect 27908 23050 27936 23718
rect 28092 23118 28120 24550
rect 28080 23112 28132 23118
rect 28080 23054 28132 23060
rect 27896 23044 27948 23050
rect 27896 22986 27948 22992
rect 27804 22024 27856 22030
rect 27804 21966 27856 21972
rect 27816 20942 27844 21966
rect 27804 20936 27856 20942
rect 27804 20878 27856 20884
rect 27908 20890 27936 22986
rect 28184 22094 28212 27934
rect 28276 26042 28304 31198
rect 28368 30938 28396 32302
rect 28356 30932 28408 30938
rect 28356 30874 28408 30880
rect 28356 29572 28408 29578
rect 28356 29514 28408 29520
rect 28368 29306 28396 29514
rect 28356 29300 28408 29306
rect 28356 29242 28408 29248
rect 28356 29028 28408 29034
rect 28356 28970 28408 28976
rect 28368 27538 28396 28970
rect 28356 27532 28408 27538
rect 28356 27474 28408 27480
rect 28264 26036 28316 26042
rect 28264 25978 28316 25984
rect 28276 24886 28304 25978
rect 28356 25288 28408 25294
rect 28354 25256 28356 25265
rect 28408 25256 28410 25265
rect 28354 25191 28410 25200
rect 28264 24880 28316 24886
rect 28264 24822 28316 24828
rect 28276 23594 28304 24822
rect 28264 23588 28316 23594
rect 28264 23530 28316 23536
rect 28092 22066 28212 22094
rect 27908 20862 28028 20890
rect 27896 20800 27948 20806
rect 27896 20742 27948 20748
rect 27908 20534 27936 20742
rect 27896 20528 27948 20534
rect 27896 20470 27948 20476
rect 27804 20256 27856 20262
rect 27804 20198 27856 20204
rect 27712 19916 27764 19922
rect 27712 19858 27764 19864
rect 27344 19848 27396 19854
rect 27344 19790 27396 19796
rect 27160 19440 27212 19446
rect 27160 19382 27212 19388
rect 27068 19304 27120 19310
rect 27068 19246 27120 19252
rect 26332 18760 26384 18766
rect 26792 18760 26844 18766
rect 26332 18702 26384 18708
rect 26422 18728 26478 18737
rect 26056 18420 26108 18426
rect 26056 18362 26108 18368
rect 26240 18420 26292 18426
rect 26240 18362 26292 18368
rect 26068 18329 26096 18362
rect 26054 18320 26110 18329
rect 25872 18284 25924 18290
rect 26054 18255 26110 18264
rect 25872 18226 25924 18232
rect 26148 18216 26200 18222
rect 26146 18184 26148 18193
rect 26200 18184 26202 18193
rect 25780 18148 25832 18154
rect 26146 18119 26202 18128
rect 25780 18090 25832 18096
rect 25792 17728 25820 18090
rect 26252 17882 26280 18362
rect 26344 18222 26372 18702
rect 26792 18702 26844 18708
rect 26976 18760 27028 18766
rect 26976 18702 27028 18708
rect 26422 18663 26478 18672
rect 26332 18216 26384 18222
rect 26332 18158 26384 18164
rect 26436 17882 26464 18663
rect 26700 18216 26752 18222
rect 26700 18158 26752 18164
rect 26240 17876 26292 17882
rect 26240 17818 26292 17824
rect 26424 17876 26476 17882
rect 26424 17818 26476 17824
rect 26712 17814 26740 18158
rect 26332 17808 26384 17814
rect 26332 17750 26384 17756
rect 26700 17808 26752 17814
rect 26700 17750 26752 17756
rect 25872 17740 25924 17746
rect 25792 17700 25872 17728
rect 25792 17066 25820 17700
rect 25872 17682 25924 17688
rect 26240 17672 26292 17678
rect 26238 17640 26240 17649
rect 26292 17640 26294 17649
rect 26238 17575 26294 17584
rect 25872 17332 25924 17338
rect 25872 17274 25924 17280
rect 25780 17060 25832 17066
rect 25780 17002 25832 17008
rect 25884 16425 25912 17274
rect 26344 16998 26372 17750
rect 26804 17678 26832 18702
rect 27252 18284 27304 18290
rect 27252 18226 27304 18232
rect 26424 17672 26476 17678
rect 26424 17614 26476 17620
rect 26792 17672 26844 17678
rect 26792 17614 26844 17620
rect 27068 17672 27120 17678
rect 27068 17614 27120 17620
rect 26436 17202 26464 17614
rect 26884 17604 26936 17610
rect 26884 17546 26936 17552
rect 26976 17604 27028 17610
rect 26976 17546 27028 17552
rect 26424 17196 26476 17202
rect 26424 17138 26476 17144
rect 26332 16992 26384 16998
rect 26332 16934 26384 16940
rect 26896 16590 26924 17546
rect 26988 17513 27016 17546
rect 26974 17504 27030 17513
rect 26974 17439 27030 17448
rect 27080 17241 27108 17614
rect 27264 17338 27292 18226
rect 27356 17814 27384 19790
rect 27816 19718 27844 20198
rect 27804 19712 27856 19718
rect 27804 19654 27856 19660
rect 27620 19236 27672 19242
rect 27620 19178 27672 19184
rect 27528 18760 27580 18766
rect 27448 18720 27528 18748
rect 27448 18630 27476 18720
rect 27528 18702 27580 18708
rect 27436 18624 27488 18630
rect 27436 18566 27488 18572
rect 27448 18086 27476 18566
rect 27436 18080 27488 18086
rect 27436 18022 27488 18028
rect 27526 18048 27582 18057
rect 27344 17808 27396 17814
rect 27344 17750 27396 17756
rect 27252 17332 27304 17338
rect 27252 17274 27304 17280
rect 27066 17232 27122 17241
rect 26976 17196 27028 17202
rect 27066 17167 27068 17176
rect 26976 17138 27028 17144
rect 27120 17167 27122 17176
rect 27068 17138 27120 17144
rect 26884 16584 26936 16590
rect 26884 16526 26936 16532
rect 26148 16448 26200 16454
rect 25870 16416 25926 16425
rect 26148 16390 26200 16396
rect 25870 16351 25926 16360
rect 26160 15638 26188 16390
rect 26700 16244 26752 16250
rect 26700 16186 26752 16192
rect 26148 15632 26200 15638
rect 26148 15574 26200 15580
rect 26056 15020 26108 15026
rect 26160 15008 26188 15574
rect 26516 15496 26568 15502
rect 26516 15438 26568 15444
rect 26528 15366 26556 15438
rect 26424 15360 26476 15366
rect 26424 15302 26476 15308
rect 26516 15360 26568 15366
rect 26516 15302 26568 15308
rect 26240 15156 26292 15162
rect 26240 15098 26292 15104
rect 26108 14980 26188 15008
rect 26056 14962 26108 14968
rect 26252 14958 26280 15098
rect 26436 15026 26464 15302
rect 26424 15020 26476 15026
rect 26424 14962 26476 14968
rect 26608 15020 26660 15026
rect 26608 14962 26660 14968
rect 26240 14952 26292 14958
rect 26240 14894 26292 14900
rect 26332 14952 26384 14958
rect 26332 14894 26384 14900
rect 26516 14952 26568 14958
rect 26516 14894 26568 14900
rect 26148 14340 26200 14346
rect 26148 14282 26200 14288
rect 26160 14074 26188 14282
rect 26148 14068 26200 14074
rect 26148 14010 26200 14016
rect 26344 13530 26372 14894
rect 26528 14550 26556 14894
rect 26516 14544 26568 14550
rect 26516 14486 26568 14492
rect 26528 13938 26556 14486
rect 26620 14278 26648 14962
rect 26608 14272 26660 14278
rect 26608 14214 26660 14220
rect 26516 13932 26568 13938
rect 26516 13874 26568 13880
rect 26332 13524 26384 13530
rect 26332 13466 26384 13472
rect 26620 13326 26648 14214
rect 26608 13320 26660 13326
rect 26608 13262 26660 13268
rect 26332 12776 26384 12782
rect 26332 12718 26384 12724
rect 26344 12434 26372 12718
rect 26712 12442 26740 16186
rect 26884 15496 26936 15502
rect 26988 15484 27016 17138
rect 27080 16590 27108 17138
rect 27068 16584 27120 16590
rect 27068 16526 27120 16532
rect 27158 16552 27214 16561
rect 27158 16487 27214 16496
rect 27172 16454 27200 16487
rect 27160 16448 27212 16454
rect 27160 16390 27212 16396
rect 27252 16108 27304 16114
rect 27252 16050 27304 16056
rect 26936 15456 27016 15484
rect 27068 15496 27120 15502
rect 26884 15438 26936 15444
rect 27068 15438 27120 15444
rect 26792 14816 26844 14822
rect 26790 14784 26792 14793
rect 26844 14784 26846 14793
rect 26790 14719 26846 14728
rect 26896 13870 26924 15438
rect 27080 15094 27108 15438
rect 27264 15366 27292 16050
rect 27344 15904 27396 15910
rect 27344 15846 27396 15852
rect 27356 15706 27384 15846
rect 27344 15700 27396 15706
rect 27344 15642 27396 15648
rect 27252 15360 27304 15366
rect 27252 15302 27304 15308
rect 27160 15156 27212 15162
rect 27160 15098 27212 15104
rect 27068 15088 27120 15094
rect 27068 15030 27120 15036
rect 26976 14816 27028 14822
rect 26976 14758 27028 14764
rect 26988 14346 27016 14758
rect 26976 14340 27028 14346
rect 26976 14282 27028 14288
rect 26884 13864 26936 13870
rect 26884 13806 26936 13812
rect 26884 13320 26936 13326
rect 26884 13262 26936 13268
rect 26792 12912 26844 12918
rect 26792 12854 26844 12860
rect 26804 12646 26832 12854
rect 26792 12640 26844 12646
rect 26792 12582 26844 12588
rect 26160 12406 26372 12434
rect 26700 12436 26752 12442
rect 25964 11756 26016 11762
rect 25964 11698 26016 11704
rect 25976 11354 26004 11698
rect 25964 11348 26016 11354
rect 25964 11290 26016 11296
rect 25872 10668 25924 10674
rect 25872 10610 25924 10616
rect 25884 8838 25912 10610
rect 25872 8832 25924 8838
rect 25872 8774 25924 8780
rect 26056 8424 26108 8430
rect 26056 8366 26108 8372
rect 26068 7410 26096 8366
rect 26160 7750 26188 12406
rect 26700 12378 26752 12384
rect 26896 12306 26924 13262
rect 26884 12300 26936 12306
rect 26884 12242 26936 12248
rect 26700 12232 26752 12238
rect 26700 12174 26752 12180
rect 26424 11688 26476 11694
rect 26424 11630 26476 11636
rect 26332 11008 26384 11014
rect 26332 10950 26384 10956
rect 26344 10826 26372 10950
rect 26252 10810 26372 10826
rect 26436 10810 26464 11630
rect 26240 10804 26372 10810
rect 26292 10798 26372 10804
rect 26240 10746 26292 10752
rect 26240 10668 26292 10674
rect 26240 10610 26292 10616
rect 26252 10130 26280 10610
rect 26240 10124 26292 10130
rect 26240 10066 26292 10072
rect 26148 7744 26200 7750
rect 26148 7686 26200 7692
rect 26056 7404 26108 7410
rect 26056 7346 26108 7352
rect 26240 7404 26292 7410
rect 26240 7346 26292 7352
rect 26148 7336 26200 7342
rect 26148 7278 26200 7284
rect 26160 7206 26188 7278
rect 26148 7200 26200 7206
rect 26148 7142 26200 7148
rect 26252 6798 26280 7346
rect 26344 6866 26372 10798
rect 26424 10804 26476 10810
rect 26424 10746 26476 10752
rect 26712 10742 26740 12174
rect 26884 12164 26936 12170
rect 26884 12106 26936 12112
rect 26896 11626 26924 12106
rect 26884 11620 26936 11626
rect 26884 11562 26936 11568
rect 26988 11082 27016 14282
rect 27068 14272 27120 14278
rect 27068 14214 27120 14220
rect 27080 14074 27108 14214
rect 27068 14068 27120 14074
rect 27068 14010 27120 14016
rect 27172 13530 27200 15098
rect 27264 14249 27292 15302
rect 27250 14240 27306 14249
rect 27250 14175 27306 14184
rect 27160 13524 27212 13530
rect 27160 13466 27212 13472
rect 27252 12980 27304 12986
rect 27252 12922 27304 12928
rect 27264 12646 27292 12922
rect 27252 12640 27304 12646
rect 27252 12582 27304 12588
rect 27160 11552 27212 11558
rect 27160 11494 27212 11500
rect 26976 11076 27028 11082
rect 26976 11018 27028 11024
rect 27172 10810 27200 11494
rect 27264 11014 27292 12582
rect 27448 12434 27476 18022
rect 27526 17983 27582 17992
rect 27540 17202 27568 17983
rect 27528 17196 27580 17202
rect 27528 17138 27580 17144
rect 27632 16590 27660 19178
rect 27896 18692 27948 18698
rect 27896 18634 27948 18640
rect 27710 18320 27766 18329
rect 27710 18255 27766 18264
rect 27724 18222 27752 18255
rect 27712 18216 27764 18222
rect 27764 18176 27844 18204
rect 27712 18158 27764 18164
rect 27816 17746 27844 18176
rect 27712 17740 27764 17746
rect 27712 17682 27764 17688
rect 27804 17740 27856 17746
rect 27804 17682 27856 17688
rect 27724 17338 27752 17682
rect 27712 17332 27764 17338
rect 27712 17274 27764 17280
rect 27620 16584 27672 16590
rect 27620 16526 27672 16532
rect 27528 15564 27580 15570
rect 27528 15506 27580 15512
rect 27540 15162 27568 15506
rect 27528 15156 27580 15162
rect 27528 15098 27580 15104
rect 27540 13938 27568 15098
rect 27632 14822 27660 16526
rect 27908 15994 27936 18634
rect 28000 18086 28028 20862
rect 27988 18080 28040 18086
rect 27988 18022 28040 18028
rect 27988 17536 28040 17542
rect 27988 17478 28040 17484
rect 28000 17338 28028 17478
rect 27988 17332 28040 17338
rect 27988 17274 28040 17280
rect 28000 17066 28028 17274
rect 27988 17060 28040 17066
rect 27988 17002 28040 17008
rect 27986 16688 28042 16697
rect 27986 16623 27988 16632
rect 28040 16623 28042 16632
rect 27988 16594 28040 16600
rect 27724 15966 27936 15994
rect 27620 14816 27672 14822
rect 27620 14758 27672 14764
rect 27620 14408 27672 14414
rect 27620 14350 27672 14356
rect 27528 13932 27580 13938
rect 27528 13874 27580 13880
rect 27632 13818 27660 14350
rect 27540 13790 27660 13818
rect 27540 13734 27568 13790
rect 27528 13728 27580 13734
rect 27528 13670 27580 13676
rect 27620 13524 27672 13530
rect 27620 13466 27672 13472
rect 27448 12406 27568 12434
rect 27540 12238 27568 12406
rect 27528 12232 27580 12238
rect 27528 12174 27580 12180
rect 27540 11762 27568 12174
rect 27528 11756 27580 11762
rect 27528 11698 27580 11704
rect 27540 11218 27568 11698
rect 27632 11558 27660 13466
rect 27724 13394 27752 15966
rect 27896 15904 27948 15910
rect 27896 15846 27948 15852
rect 27804 15428 27856 15434
rect 27804 15370 27856 15376
rect 27816 15337 27844 15370
rect 27802 15328 27858 15337
rect 27802 15263 27858 15272
rect 27804 15156 27856 15162
rect 27804 15098 27856 15104
rect 27816 15026 27844 15098
rect 27804 15020 27856 15026
rect 27804 14962 27856 14968
rect 27908 14414 27936 15846
rect 27988 15700 28040 15706
rect 27988 15642 28040 15648
rect 28000 14414 28028 15642
rect 27896 14408 27948 14414
rect 27896 14350 27948 14356
rect 27988 14408 28040 14414
rect 27988 14350 28040 14356
rect 27804 14272 27856 14278
rect 27896 14272 27948 14278
rect 27804 14214 27856 14220
rect 27894 14240 27896 14249
rect 27948 14240 27950 14249
rect 27816 13938 27844 14214
rect 27894 14175 27950 14184
rect 27896 14068 27948 14074
rect 27896 14010 27948 14016
rect 27804 13932 27856 13938
rect 27804 13874 27856 13880
rect 27908 13462 27936 14010
rect 28000 13870 28028 14350
rect 27988 13864 28040 13870
rect 27988 13806 28040 13812
rect 27896 13456 27948 13462
rect 27896 13398 27948 13404
rect 27712 13388 27764 13394
rect 27712 13330 27764 13336
rect 27724 12850 27752 13330
rect 27712 12844 27764 12850
rect 27712 12786 27764 12792
rect 27724 12170 27752 12786
rect 27988 12640 28040 12646
rect 27988 12582 28040 12588
rect 27712 12164 27764 12170
rect 27712 12106 27764 12112
rect 27620 11552 27672 11558
rect 27620 11494 27672 11500
rect 27896 11552 27948 11558
rect 27896 11494 27948 11500
rect 27528 11212 27580 11218
rect 27528 11154 27580 11160
rect 27908 11082 27936 11494
rect 28000 11150 28028 12582
rect 27988 11144 28040 11150
rect 27988 11086 28040 11092
rect 27528 11076 27580 11082
rect 27528 11018 27580 11024
rect 27896 11076 27948 11082
rect 27896 11018 27948 11024
rect 27252 11008 27304 11014
rect 27252 10950 27304 10956
rect 27160 10804 27212 10810
rect 27160 10746 27212 10752
rect 26700 10736 26752 10742
rect 26700 10678 26752 10684
rect 26976 10668 27028 10674
rect 26976 10610 27028 10616
rect 26792 10600 26844 10606
rect 26792 10542 26844 10548
rect 26804 9994 26832 10542
rect 26988 9994 27016 10610
rect 27172 10062 27200 10746
rect 27436 10192 27488 10198
rect 27436 10134 27488 10140
rect 27160 10056 27212 10062
rect 27160 9998 27212 10004
rect 26792 9988 26844 9994
rect 26792 9930 26844 9936
rect 26976 9988 27028 9994
rect 26976 9930 27028 9936
rect 26804 9382 26832 9930
rect 27160 9580 27212 9586
rect 27160 9522 27212 9528
rect 26792 9376 26844 9382
rect 26792 9318 26844 9324
rect 26976 9376 27028 9382
rect 26976 9318 27028 9324
rect 26988 8974 27016 9318
rect 26976 8968 27028 8974
rect 26976 8910 27028 8916
rect 27172 8566 27200 9522
rect 27448 8634 27476 10134
rect 27436 8628 27488 8634
rect 27436 8570 27488 8576
rect 27160 8560 27212 8566
rect 27160 8502 27212 8508
rect 27068 7268 27120 7274
rect 27068 7210 27120 7216
rect 26332 6860 26384 6866
rect 26332 6802 26384 6808
rect 27080 6798 27108 7210
rect 27172 6798 27200 8502
rect 27540 8090 27568 11018
rect 27712 11008 27764 11014
rect 27712 10950 27764 10956
rect 27724 10266 27752 10950
rect 28000 10674 28028 11086
rect 27988 10668 28040 10674
rect 27988 10610 28040 10616
rect 27804 10464 27856 10470
rect 27804 10406 27856 10412
rect 27896 10464 27948 10470
rect 27896 10406 27948 10412
rect 27712 10260 27764 10266
rect 27712 10202 27764 10208
rect 27816 10062 27844 10406
rect 27804 10056 27856 10062
rect 27804 9998 27856 10004
rect 27620 9988 27672 9994
rect 27620 9930 27672 9936
rect 27712 9988 27764 9994
rect 27712 9930 27764 9936
rect 27632 8430 27660 9930
rect 27724 8974 27752 9930
rect 27908 9926 27936 10406
rect 28092 10146 28120 22066
rect 28264 21956 28316 21962
rect 28264 21898 28316 21904
rect 28172 21548 28224 21554
rect 28172 21490 28224 21496
rect 28184 21185 28212 21490
rect 28276 21350 28304 21898
rect 28460 21622 28488 48486
rect 28540 47592 28592 47598
rect 28540 47534 28592 47540
rect 28552 47054 28580 47534
rect 28540 47048 28592 47054
rect 28540 46990 28592 46996
rect 28816 43444 28868 43450
rect 28816 43386 28868 43392
rect 28828 42702 28856 43386
rect 29092 42764 29144 42770
rect 29092 42706 29144 42712
rect 28816 42696 28868 42702
rect 28816 42638 28868 42644
rect 28828 42294 28856 42638
rect 28816 42288 28868 42294
rect 28816 42230 28868 42236
rect 28828 40662 28856 42230
rect 29104 42022 29132 42706
rect 29182 42392 29238 42401
rect 29182 42327 29184 42336
rect 29236 42327 29238 42336
rect 29184 42298 29236 42304
rect 29092 42016 29144 42022
rect 29092 41958 29144 41964
rect 29000 41540 29052 41546
rect 29000 41482 29052 41488
rect 29012 41274 29040 41482
rect 29104 41478 29132 41958
rect 29092 41472 29144 41478
rect 29092 41414 29144 41420
rect 29000 41268 29052 41274
rect 29000 41210 29052 41216
rect 29104 41138 29132 41414
rect 29184 41268 29236 41274
rect 29184 41210 29236 41216
rect 29092 41132 29144 41138
rect 29092 41074 29144 41080
rect 28816 40656 28868 40662
rect 28816 40598 28868 40604
rect 28828 39370 28856 40598
rect 29196 40526 29224 41210
rect 29184 40520 29236 40526
rect 29184 40462 29236 40468
rect 28816 39364 28868 39370
rect 28816 39306 28868 39312
rect 29092 39092 29144 39098
rect 29092 39034 29144 39040
rect 28908 38888 28960 38894
rect 28908 38830 28960 38836
rect 28816 38344 28868 38350
rect 28816 38286 28868 38292
rect 28828 38010 28856 38286
rect 28816 38004 28868 38010
rect 28816 37946 28868 37952
rect 28540 37120 28592 37126
rect 28592 37068 28672 37074
rect 28540 37062 28672 37068
rect 28552 37046 28672 37062
rect 28540 34604 28592 34610
rect 28540 34546 28592 34552
rect 28552 33114 28580 34546
rect 28540 33108 28592 33114
rect 28540 33050 28592 33056
rect 28540 32564 28592 32570
rect 28540 32506 28592 32512
rect 28552 31890 28580 32506
rect 28540 31884 28592 31890
rect 28540 31826 28592 31832
rect 28644 31482 28672 37046
rect 28816 36780 28868 36786
rect 28816 36722 28868 36728
rect 28828 36582 28856 36722
rect 28816 36576 28868 36582
rect 28816 36518 28868 36524
rect 28920 36530 28948 38830
rect 29000 38344 29052 38350
rect 29000 38286 29052 38292
rect 29012 37466 29040 38286
rect 29104 37942 29132 39034
rect 29288 38944 29316 48554
rect 29380 48278 29408 48622
rect 29932 48346 29960 49098
rect 29920 48340 29972 48346
rect 29920 48282 29972 48288
rect 29368 48272 29420 48278
rect 29368 48214 29420 48220
rect 30104 48136 30156 48142
rect 29550 48104 29606 48113
rect 30104 48078 30156 48084
rect 29550 48039 29606 48048
rect 29564 47598 29592 48039
rect 30116 47734 30144 48078
rect 30104 47728 30156 47734
rect 30104 47670 30156 47676
rect 29552 47592 29604 47598
rect 29552 47534 29604 47540
rect 30116 44946 30144 47670
rect 30576 47666 30604 49234
rect 31944 49224 31996 49230
rect 31944 49166 31996 49172
rect 31956 48210 31984 49166
rect 32128 49088 32180 49094
rect 32128 49030 32180 49036
rect 32140 48754 32168 49030
rect 32128 48748 32180 48754
rect 32128 48690 32180 48696
rect 32232 48210 32260 51200
rect 32876 48686 32904 51200
rect 32312 48680 32364 48686
rect 32312 48622 32364 48628
rect 32864 48680 32916 48686
rect 32864 48622 32916 48628
rect 32324 48278 32352 48622
rect 33796 48550 33824 51326
rect 34072 51326 34206 51354
rect 33784 48544 33836 48550
rect 33784 48486 33836 48492
rect 32312 48272 32364 48278
rect 32312 48214 32364 48220
rect 31944 48204 31996 48210
rect 31944 48146 31996 48152
rect 32220 48204 32272 48210
rect 32220 48146 32272 48152
rect 30748 48136 30800 48142
rect 30748 48078 30800 48084
rect 33784 48136 33836 48142
rect 33784 48078 33836 48084
rect 30760 47802 30788 48078
rect 32220 48068 32272 48074
rect 32220 48010 32272 48016
rect 32128 48000 32180 48006
rect 32128 47942 32180 47948
rect 30748 47796 30800 47802
rect 30748 47738 30800 47744
rect 30564 47660 30616 47666
rect 30564 47602 30616 47608
rect 30104 44940 30156 44946
rect 30104 44882 30156 44888
rect 29368 42696 29420 42702
rect 29368 42638 29420 42644
rect 29552 42696 29604 42702
rect 29552 42638 29604 42644
rect 29380 42362 29408 42638
rect 29368 42356 29420 42362
rect 29368 42298 29420 42304
rect 29564 41682 29592 42638
rect 30196 42560 30248 42566
rect 30196 42502 30248 42508
rect 29644 42356 29696 42362
rect 29644 42298 29696 42304
rect 29920 42356 29972 42362
rect 29920 42298 29972 42304
rect 29552 41676 29604 41682
rect 29552 41618 29604 41624
rect 29564 41070 29592 41618
rect 29552 41064 29604 41070
rect 29552 41006 29604 41012
rect 29656 39098 29684 42298
rect 29932 42226 29960 42298
rect 29920 42220 29972 42226
rect 29920 42162 29972 42168
rect 30208 42158 30236 42502
rect 30196 42152 30248 42158
rect 30196 42094 30248 42100
rect 30208 41414 30236 42094
rect 30288 42016 30340 42022
rect 30288 41958 30340 41964
rect 30300 41818 30328 41958
rect 30288 41812 30340 41818
rect 30288 41754 30340 41760
rect 30760 41414 30788 47738
rect 32140 47666 32168 47942
rect 32232 47802 32260 48010
rect 32220 47796 32272 47802
rect 32220 47738 32272 47744
rect 33796 47666 33824 48078
rect 31852 47660 31904 47666
rect 31852 47602 31904 47608
rect 32128 47660 32180 47666
rect 32128 47602 32180 47608
rect 33140 47660 33192 47666
rect 33140 47602 33192 47608
rect 33784 47660 33836 47666
rect 33784 47602 33836 47608
rect 30838 42392 30894 42401
rect 30838 42327 30840 42336
rect 30892 42327 30894 42336
rect 30840 42298 30892 42304
rect 30932 41472 30984 41478
rect 30932 41414 30984 41420
rect 31864 41414 31892 47602
rect 33152 47122 33180 47602
rect 33140 47116 33192 47122
rect 33140 47058 33192 47064
rect 33692 47116 33744 47122
rect 33692 47058 33744 47064
rect 33324 41472 33376 41478
rect 33324 41414 33376 41420
rect 30208 41386 30328 41414
rect 30300 41154 30328 41386
rect 30208 41126 30328 41154
rect 30668 41386 30788 41414
rect 29828 40452 29880 40458
rect 29828 40394 29880 40400
rect 29840 40186 29868 40394
rect 29828 40180 29880 40186
rect 29828 40122 29880 40128
rect 29828 40044 29880 40050
rect 29828 39986 29880 39992
rect 29644 39092 29696 39098
rect 29644 39034 29696 39040
rect 29196 38916 29316 38944
rect 29092 37936 29144 37942
rect 29092 37878 29144 37884
rect 29000 37460 29052 37466
rect 29000 37402 29052 37408
rect 29012 37194 29040 37402
rect 29092 37324 29144 37330
rect 29092 37266 29144 37272
rect 29000 37188 29052 37194
rect 29000 37130 29052 37136
rect 28920 36502 28994 36530
rect 28966 36394 28994 36502
rect 29104 36394 29132 37266
rect 29196 36666 29224 38916
rect 29840 38894 29868 39986
rect 30208 39914 30236 41126
rect 30288 41064 30340 41070
rect 30288 41006 30340 41012
rect 30196 39908 30248 39914
rect 30196 39850 30248 39856
rect 30300 39506 30328 41006
rect 30288 39500 30340 39506
rect 30288 39442 30340 39448
rect 29828 38888 29880 38894
rect 29828 38830 29880 38836
rect 29276 38820 29328 38826
rect 29276 38762 29328 38768
rect 29288 38418 29316 38762
rect 29276 38412 29328 38418
rect 29276 38354 29328 38360
rect 29288 37398 29316 38354
rect 29736 37868 29788 37874
rect 29736 37810 29788 37816
rect 29276 37392 29328 37398
rect 29276 37334 29328 37340
rect 29748 37194 29776 37810
rect 29840 37806 29868 38830
rect 30300 38350 30328 39442
rect 30380 39364 30432 39370
rect 30380 39306 30432 39312
rect 30392 39098 30420 39306
rect 30380 39092 30432 39098
rect 30380 39034 30432 39040
rect 30380 38956 30432 38962
rect 30380 38898 30432 38904
rect 30288 38344 30340 38350
rect 30288 38286 30340 38292
rect 30300 37874 30328 38286
rect 30392 38214 30420 38898
rect 30380 38208 30432 38214
rect 30380 38150 30432 38156
rect 30288 37868 30340 37874
rect 30288 37810 30340 37816
rect 29828 37800 29880 37806
rect 29828 37742 29880 37748
rect 29840 37330 29868 37742
rect 29828 37324 29880 37330
rect 29828 37266 29880 37272
rect 29736 37188 29788 37194
rect 29736 37130 29788 37136
rect 29368 37120 29420 37126
rect 29368 37062 29420 37068
rect 29380 36786 29408 37062
rect 29368 36780 29420 36786
rect 29368 36722 29420 36728
rect 29552 36780 29604 36786
rect 29552 36722 29604 36728
rect 29196 36638 29408 36666
rect 28966 36366 29132 36394
rect 28908 35556 28960 35562
rect 28908 35498 28960 35504
rect 28724 35012 28776 35018
rect 28724 34954 28776 34960
rect 28736 32434 28764 34954
rect 28920 34542 28948 35498
rect 29380 35222 29408 36638
rect 29564 36310 29592 36722
rect 29552 36304 29604 36310
rect 29552 36246 29604 36252
rect 29748 35698 29776 37130
rect 30104 36780 30156 36786
rect 30104 36722 30156 36728
rect 30012 36168 30064 36174
rect 30012 36110 30064 36116
rect 29828 36032 29880 36038
rect 29828 35974 29880 35980
rect 29736 35692 29788 35698
rect 29736 35634 29788 35640
rect 29368 35216 29420 35222
rect 29368 35158 29420 35164
rect 29840 35018 29868 35974
rect 30024 35894 30052 36110
rect 30116 36106 30144 36722
rect 30104 36100 30156 36106
rect 30104 36042 30156 36048
rect 30196 36032 30248 36038
rect 30196 35974 30248 35980
rect 30024 35866 30144 35894
rect 29920 35828 29972 35834
rect 29920 35770 29972 35776
rect 29644 35012 29696 35018
rect 29644 34954 29696 34960
rect 29828 35012 29880 35018
rect 29828 34954 29880 34960
rect 29552 34944 29604 34950
rect 29552 34886 29604 34892
rect 28908 34536 28960 34542
rect 28908 34478 28960 34484
rect 28816 33516 28868 33522
rect 28920 33504 28948 34478
rect 28868 33476 28948 33504
rect 28816 33458 28868 33464
rect 29368 32836 29420 32842
rect 29368 32778 29420 32784
rect 28816 32768 28868 32774
rect 28816 32710 28868 32716
rect 28724 32428 28776 32434
rect 28724 32370 28776 32376
rect 28736 32230 28764 32370
rect 28724 32224 28776 32230
rect 28724 32166 28776 32172
rect 28632 31476 28684 31482
rect 28632 31418 28684 31424
rect 28540 31340 28592 31346
rect 28540 31282 28592 31288
rect 28724 31340 28776 31346
rect 28724 31282 28776 31288
rect 28552 27690 28580 31282
rect 28736 30054 28764 31282
rect 28724 30048 28776 30054
rect 28724 29990 28776 29996
rect 28736 28626 28764 29990
rect 28724 28620 28776 28626
rect 28724 28562 28776 28568
rect 28828 28558 28856 32710
rect 29380 32570 29408 32778
rect 29368 32564 29420 32570
rect 29368 32506 29420 32512
rect 29460 32224 29512 32230
rect 29460 32166 29512 32172
rect 28908 31884 28960 31890
rect 28908 31826 28960 31832
rect 28920 31210 28948 31826
rect 29366 31784 29422 31793
rect 29366 31719 29368 31728
rect 29420 31719 29422 31728
rect 29368 31690 29420 31696
rect 28908 31204 28960 31210
rect 28908 31146 28960 31152
rect 29472 30326 29500 32166
rect 29564 31958 29592 34886
rect 29656 34610 29684 34954
rect 29932 34950 29960 35770
rect 30116 35766 30144 35866
rect 30104 35760 30156 35766
rect 30104 35702 30156 35708
rect 30208 35630 30236 35974
rect 30196 35624 30248 35630
rect 30196 35566 30248 35572
rect 29920 34944 29972 34950
rect 29920 34886 29972 34892
rect 29644 34604 29696 34610
rect 29644 34546 29696 34552
rect 29644 33924 29696 33930
rect 29644 33866 29696 33872
rect 29656 33658 29684 33866
rect 29920 33856 29972 33862
rect 29920 33798 29972 33804
rect 29644 33652 29696 33658
rect 29644 33594 29696 33600
rect 29734 33144 29790 33153
rect 29734 33079 29790 33088
rect 29748 32570 29776 33079
rect 29932 32570 29960 33798
rect 30392 33658 30420 38150
rect 30564 36168 30616 36174
rect 30564 36110 30616 36116
rect 30472 35624 30524 35630
rect 30472 35566 30524 35572
rect 30484 34406 30512 35566
rect 30576 35562 30604 36110
rect 30564 35556 30616 35562
rect 30564 35498 30616 35504
rect 30576 34474 30604 35498
rect 30564 34468 30616 34474
rect 30564 34410 30616 34416
rect 30472 34400 30524 34406
rect 30472 34342 30524 34348
rect 30484 34202 30512 34342
rect 30472 34196 30524 34202
rect 30472 34138 30524 34144
rect 30380 33652 30432 33658
rect 30380 33594 30432 33600
rect 30484 33454 30512 34138
rect 30472 33448 30524 33454
rect 30472 33390 30524 33396
rect 30380 33108 30432 33114
rect 30380 33050 30432 33056
rect 30392 32994 30420 33050
rect 30392 32966 30512 32994
rect 29736 32564 29788 32570
rect 29736 32506 29788 32512
rect 29920 32564 29972 32570
rect 29920 32506 29972 32512
rect 30196 32360 30248 32366
rect 30196 32302 30248 32308
rect 29644 32020 29696 32026
rect 29644 31962 29696 31968
rect 29552 31952 29604 31958
rect 29552 31894 29604 31900
rect 29656 31822 29684 31962
rect 30208 31822 30236 32302
rect 30288 32224 30340 32230
rect 30288 32166 30340 32172
rect 30300 31890 30328 32166
rect 30288 31884 30340 31890
rect 30288 31826 30340 31832
rect 29644 31816 29696 31822
rect 29644 31758 29696 31764
rect 30196 31816 30248 31822
rect 30196 31758 30248 31764
rect 30380 31748 30432 31754
rect 30380 31690 30432 31696
rect 29828 31680 29880 31686
rect 29828 31622 29880 31628
rect 29840 30734 29868 31622
rect 30392 31482 30420 31690
rect 30380 31476 30432 31482
rect 30380 31418 30432 31424
rect 30012 31340 30064 31346
rect 30012 31282 30064 31288
rect 29736 30728 29788 30734
rect 29736 30670 29788 30676
rect 29828 30728 29880 30734
rect 29828 30670 29880 30676
rect 29748 30394 29776 30670
rect 30024 30598 30052 31282
rect 30012 30592 30064 30598
rect 30012 30534 30064 30540
rect 29736 30388 29788 30394
rect 29736 30330 29788 30336
rect 29460 30320 29512 30326
rect 29460 30262 29512 30268
rect 28908 29640 28960 29646
rect 28908 29582 28960 29588
rect 28816 28552 28868 28558
rect 28816 28494 28868 28500
rect 28632 28416 28684 28422
rect 28632 28358 28684 28364
rect 28644 27878 28672 28358
rect 28632 27872 28684 27878
rect 28632 27814 28684 27820
rect 28552 27662 28672 27690
rect 28540 26988 28592 26994
rect 28540 26930 28592 26936
rect 28552 26586 28580 26930
rect 28540 26580 28592 26586
rect 28540 26522 28592 26528
rect 28644 26466 28672 27662
rect 28920 27402 28948 29582
rect 29828 28416 29880 28422
rect 29828 28358 29880 28364
rect 29840 27470 29868 28358
rect 29828 27464 29880 27470
rect 29828 27406 29880 27412
rect 28908 27396 28960 27402
rect 28908 27338 28960 27344
rect 28920 27062 28948 27338
rect 28908 27056 28960 27062
rect 28908 26998 28960 27004
rect 28552 26438 28672 26466
rect 29000 26512 29052 26518
rect 29000 26454 29052 26460
rect 28552 24614 28580 26438
rect 28632 25968 28684 25974
rect 28632 25910 28684 25916
rect 28644 25294 28672 25910
rect 28816 25696 28868 25702
rect 28816 25638 28868 25644
rect 28632 25288 28684 25294
rect 28632 25230 28684 25236
rect 28828 24970 28856 25638
rect 28736 24942 28856 24970
rect 28632 24812 28684 24818
rect 28632 24754 28684 24760
rect 28540 24608 28592 24614
rect 28540 24550 28592 24556
rect 28644 24070 28672 24754
rect 28736 24206 28764 24942
rect 29012 24818 29040 26454
rect 30024 26450 30052 30534
rect 30196 29232 30248 29238
rect 30196 29174 30248 29180
rect 30208 27606 30236 29174
rect 30196 27600 30248 27606
rect 30196 27542 30248 27548
rect 30012 26444 30064 26450
rect 30012 26386 30064 26392
rect 29276 26240 29328 26246
rect 29276 26182 29328 26188
rect 29288 26042 29316 26182
rect 29276 26036 29328 26042
rect 29276 25978 29328 25984
rect 29288 25362 29316 25978
rect 29552 25968 29604 25974
rect 29552 25910 29604 25916
rect 29276 25356 29328 25362
rect 29276 25298 29328 25304
rect 29368 25220 29420 25226
rect 29368 25162 29420 25168
rect 29000 24812 29052 24818
rect 29000 24754 29052 24760
rect 28908 24676 28960 24682
rect 28908 24618 28960 24624
rect 28920 24274 28948 24618
rect 28908 24268 28960 24274
rect 28908 24210 28960 24216
rect 28724 24200 28776 24206
rect 28724 24142 28776 24148
rect 28908 24132 28960 24138
rect 28908 24074 28960 24080
rect 28632 24064 28684 24070
rect 28632 24006 28684 24012
rect 28644 23662 28672 24006
rect 28920 23866 28948 24074
rect 28908 23860 28960 23866
rect 28908 23802 28960 23808
rect 29012 23730 29040 24754
rect 29380 24410 29408 25162
rect 29460 25152 29512 25158
rect 29460 25094 29512 25100
rect 29472 24818 29500 25094
rect 29564 24954 29592 25910
rect 30012 25492 30064 25498
rect 30012 25434 30064 25440
rect 29642 25256 29698 25265
rect 29642 25191 29644 25200
rect 29696 25191 29698 25200
rect 29644 25162 29696 25168
rect 29552 24948 29604 24954
rect 29552 24890 29604 24896
rect 30024 24818 30052 25434
rect 30380 25288 30432 25294
rect 30380 25230 30432 25236
rect 30392 25158 30420 25230
rect 30380 25152 30432 25158
rect 30380 25094 30432 25100
rect 30392 24954 30420 25094
rect 30380 24948 30432 24954
rect 30380 24890 30432 24896
rect 29460 24812 29512 24818
rect 29460 24754 29512 24760
rect 30012 24812 30064 24818
rect 30012 24754 30064 24760
rect 29368 24404 29420 24410
rect 29368 24346 29420 24352
rect 29642 24032 29698 24041
rect 29642 23967 29698 23976
rect 29656 23866 29684 23967
rect 29644 23860 29696 23866
rect 29644 23802 29696 23808
rect 30024 23730 30052 24754
rect 30380 24744 30432 24750
rect 30380 24686 30432 24692
rect 30104 24404 30156 24410
rect 30104 24346 30156 24352
rect 30116 24070 30144 24346
rect 30104 24064 30156 24070
rect 30104 24006 30156 24012
rect 29000 23724 29052 23730
rect 29000 23666 29052 23672
rect 30012 23724 30064 23730
rect 30012 23666 30064 23672
rect 30392 23662 30420 24686
rect 30484 23662 30512 32966
rect 30564 26784 30616 26790
rect 30564 26726 30616 26732
rect 30576 25362 30604 26726
rect 30564 25356 30616 25362
rect 30564 25298 30616 25304
rect 30668 24410 30696 41386
rect 30944 41138 30972 41414
rect 31864 41386 32076 41414
rect 30932 41132 30984 41138
rect 30932 41074 30984 41080
rect 31116 40520 31168 40526
rect 31114 40488 31116 40497
rect 31168 40488 31170 40497
rect 30748 40452 30800 40458
rect 31772 40458 31984 40474
rect 31114 40423 31170 40432
rect 31760 40452 31984 40458
rect 30748 40394 30800 40400
rect 31812 40446 31984 40452
rect 31760 40394 31812 40400
rect 30760 40050 30788 40394
rect 30840 40384 30892 40390
rect 30840 40326 30892 40332
rect 31668 40384 31720 40390
rect 31668 40326 31720 40332
rect 30748 40044 30800 40050
rect 30748 39986 30800 39992
rect 30852 38962 30880 40326
rect 31680 40118 31708 40326
rect 31024 40112 31076 40118
rect 31024 40054 31076 40060
rect 31668 40112 31720 40118
rect 31668 40054 31720 40060
rect 31036 39302 31064 40054
rect 31852 39636 31904 39642
rect 31852 39578 31904 39584
rect 30932 39296 30984 39302
rect 30930 39264 30932 39273
rect 31024 39296 31076 39302
rect 30984 39264 30986 39273
rect 31024 39238 31076 39244
rect 31668 39296 31720 39302
rect 31668 39238 31720 39244
rect 30930 39199 30986 39208
rect 30840 38956 30892 38962
rect 30840 38898 30892 38904
rect 31300 38956 31352 38962
rect 31300 38898 31352 38904
rect 31312 37466 31340 38898
rect 31300 37460 31352 37466
rect 31300 37402 31352 37408
rect 30748 37120 30800 37126
rect 30748 37062 30800 37068
rect 30760 36582 30788 37062
rect 30748 36576 30800 36582
rect 30748 36518 30800 36524
rect 30760 36292 30788 36518
rect 30760 36264 30880 36292
rect 30748 36100 30800 36106
rect 30748 36042 30800 36048
rect 30760 34678 30788 36042
rect 30748 34672 30800 34678
rect 30748 34614 30800 34620
rect 30760 32502 30788 34614
rect 30748 32496 30800 32502
rect 30748 32438 30800 32444
rect 30746 31784 30802 31793
rect 30746 31719 30748 31728
rect 30800 31719 30802 31728
rect 30748 31690 30800 31696
rect 30760 31346 30788 31690
rect 30852 31482 30880 36264
rect 31312 35766 31340 37402
rect 31392 36780 31444 36786
rect 31392 36722 31444 36728
rect 31404 35766 31432 36722
rect 31300 35760 31352 35766
rect 31300 35702 31352 35708
rect 31392 35760 31444 35766
rect 31392 35702 31444 35708
rect 31484 35692 31536 35698
rect 31484 35634 31536 35640
rect 31496 34746 31524 35634
rect 31576 35012 31628 35018
rect 31576 34954 31628 34960
rect 31588 34746 31616 34954
rect 31484 34740 31536 34746
rect 31484 34682 31536 34688
rect 31576 34740 31628 34746
rect 31576 34682 31628 34688
rect 31484 34128 31536 34134
rect 31484 34070 31536 34076
rect 31392 33516 31444 33522
rect 31392 33458 31444 33464
rect 31404 33114 31432 33458
rect 31496 33153 31524 34070
rect 31680 34066 31708 39238
rect 31864 39098 31892 39578
rect 31852 39092 31904 39098
rect 31852 39034 31904 39040
rect 31760 37868 31812 37874
rect 31760 37810 31812 37816
rect 31772 36718 31800 37810
rect 31956 36786 31984 40446
rect 31944 36780 31996 36786
rect 31944 36722 31996 36728
rect 31760 36712 31812 36718
rect 31760 36654 31812 36660
rect 31772 36310 31800 36654
rect 32048 36530 32076 41386
rect 32128 41132 32180 41138
rect 32128 41074 32180 41080
rect 32140 39642 32168 41074
rect 32312 41064 32364 41070
rect 32312 41006 32364 41012
rect 32220 40724 32272 40730
rect 32220 40666 32272 40672
rect 32232 40186 32260 40666
rect 32220 40180 32272 40186
rect 32220 40122 32272 40128
rect 32324 39982 32352 41006
rect 32404 40588 32456 40594
rect 32404 40530 32456 40536
rect 32956 40588 33008 40594
rect 32956 40530 33008 40536
rect 32416 40497 32444 40530
rect 32402 40488 32458 40497
rect 32402 40423 32458 40432
rect 32312 39976 32364 39982
rect 32312 39918 32364 39924
rect 32404 39840 32456 39846
rect 32404 39782 32456 39788
rect 32496 39840 32548 39846
rect 32496 39782 32548 39788
rect 32128 39636 32180 39642
rect 32128 39578 32180 39584
rect 32312 39432 32364 39438
rect 32310 39400 32312 39409
rect 32364 39400 32366 39409
rect 32310 39335 32366 39344
rect 32416 37398 32444 39782
rect 32508 39574 32536 39782
rect 32496 39568 32548 39574
rect 32496 39510 32548 39516
rect 32772 39432 32824 39438
rect 32772 39374 32824 39380
rect 32784 38962 32812 39374
rect 32772 38956 32824 38962
rect 32772 38898 32824 38904
rect 32864 38344 32916 38350
rect 32864 38286 32916 38292
rect 32496 38208 32548 38214
rect 32496 38150 32548 38156
rect 32508 37874 32536 38150
rect 32496 37868 32548 37874
rect 32496 37810 32548 37816
rect 32680 37664 32732 37670
rect 32680 37606 32732 37612
rect 32404 37392 32456 37398
rect 32404 37334 32456 37340
rect 32692 37262 32720 37606
rect 32876 37466 32904 38286
rect 32864 37460 32916 37466
rect 32864 37402 32916 37408
rect 32404 37256 32456 37262
rect 32404 37198 32456 37204
rect 32680 37256 32732 37262
rect 32680 37198 32732 37204
rect 32416 36786 32444 37198
rect 32312 36780 32364 36786
rect 32312 36722 32364 36728
rect 32404 36780 32456 36786
rect 32404 36722 32456 36728
rect 31864 36502 32076 36530
rect 31760 36304 31812 36310
rect 31760 36246 31812 36252
rect 31772 35154 31800 36246
rect 31760 35148 31812 35154
rect 31760 35090 31812 35096
rect 31668 34060 31720 34066
rect 31668 34002 31720 34008
rect 31576 33992 31628 33998
rect 31576 33934 31628 33940
rect 31588 33658 31616 33934
rect 31576 33652 31628 33658
rect 31576 33594 31628 33600
rect 31482 33144 31538 33153
rect 31392 33108 31444 33114
rect 31482 33079 31538 33088
rect 31392 33050 31444 33056
rect 30840 31476 30892 31482
rect 30840 31418 30892 31424
rect 30748 31340 30800 31346
rect 30748 31282 30800 31288
rect 30840 31272 30892 31278
rect 30840 31214 30892 31220
rect 30852 30802 30880 31214
rect 30840 30796 30892 30802
rect 30840 30738 30892 30744
rect 31208 29572 31260 29578
rect 31208 29514 31260 29520
rect 31116 29028 31168 29034
rect 31116 28970 31168 28976
rect 30748 28960 30800 28966
rect 30748 28902 30800 28908
rect 30760 28082 30788 28902
rect 30748 28076 30800 28082
rect 30748 28018 30800 28024
rect 31128 27334 31156 28970
rect 31220 28762 31248 29514
rect 31208 28756 31260 28762
rect 31208 28698 31260 28704
rect 31404 28626 31432 33050
rect 31496 32978 31524 33079
rect 31484 32972 31536 32978
rect 31484 32914 31536 32920
rect 31760 32904 31812 32910
rect 31760 32846 31812 32852
rect 31772 32230 31800 32846
rect 31760 32224 31812 32230
rect 31760 32166 31812 32172
rect 31772 31958 31800 32166
rect 31760 31952 31812 31958
rect 31760 31894 31812 31900
rect 31864 31754 31892 36502
rect 32036 35624 32088 35630
rect 32036 35566 32088 35572
rect 32048 35290 32076 35566
rect 32128 35488 32180 35494
rect 32128 35430 32180 35436
rect 32036 35284 32088 35290
rect 32036 35226 32088 35232
rect 32140 35086 32168 35430
rect 32128 35080 32180 35086
rect 32128 35022 32180 35028
rect 32036 35012 32088 35018
rect 32036 34954 32088 34960
rect 32048 33862 32076 34954
rect 32220 34536 32272 34542
rect 32220 34478 32272 34484
rect 32036 33856 32088 33862
rect 32036 33798 32088 33804
rect 32128 33856 32180 33862
rect 32128 33798 32180 33804
rect 32048 33522 32076 33798
rect 32140 33590 32168 33798
rect 32128 33584 32180 33590
rect 32128 33526 32180 33532
rect 32036 33516 32088 33522
rect 32036 33458 32088 33464
rect 32232 32910 32260 34478
rect 32220 32904 32272 32910
rect 32220 32846 32272 32852
rect 31864 31726 32168 31754
rect 31944 31340 31996 31346
rect 31944 31282 31996 31288
rect 31956 30734 31984 31282
rect 31944 30728 31996 30734
rect 31944 30670 31996 30676
rect 31484 29504 31536 29510
rect 31484 29446 31536 29452
rect 31392 28620 31444 28626
rect 31392 28562 31444 28568
rect 31496 27470 31524 29446
rect 31760 29164 31812 29170
rect 31760 29106 31812 29112
rect 31772 29073 31800 29106
rect 31758 29064 31814 29073
rect 31758 28999 31814 29008
rect 31576 28416 31628 28422
rect 31576 28358 31628 28364
rect 31588 27878 31616 28358
rect 31576 27872 31628 27878
rect 31576 27814 31628 27820
rect 31484 27464 31536 27470
rect 31484 27406 31536 27412
rect 31116 27328 31168 27334
rect 31116 27270 31168 27276
rect 31128 27130 31156 27270
rect 31116 27124 31168 27130
rect 31116 27066 31168 27072
rect 31208 26988 31260 26994
rect 31208 26930 31260 26936
rect 31220 26586 31248 26930
rect 31208 26580 31260 26586
rect 31208 26522 31260 26528
rect 31392 26376 31444 26382
rect 31392 26318 31444 26324
rect 31116 26308 31168 26314
rect 31116 26250 31168 26256
rect 30932 25832 30984 25838
rect 30932 25774 30984 25780
rect 30944 25430 30972 25774
rect 31128 25770 31156 26250
rect 31404 25906 31432 26318
rect 31392 25900 31444 25906
rect 31392 25842 31444 25848
rect 31116 25764 31168 25770
rect 31116 25706 31168 25712
rect 30932 25424 30984 25430
rect 30932 25366 30984 25372
rect 31128 25226 31156 25706
rect 31116 25220 31168 25226
rect 31116 25162 31168 25168
rect 31404 24954 31432 25842
rect 31392 24948 31444 24954
rect 31392 24890 31444 24896
rect 30656 24404 30708 24410
rect 30656 24346 30708 24352
rect 31300 24268 31352 24274
rect 31300 24210 31352 24216
rect 31312 23746 31340 24210
rect 31404 24138 31432 24890
rect 31588 24274 31616 27814
rect 31772 27470 31800 28999
rect 31944 28076 31996 28082
rect 31944 28018 31996 28024
rect 31956 27606 31984 28018
rect 31944 27600 31996 27606
rect 31944 27542 31996 27548
rect 31760 27464 31812 27470
rect 31760 27406 31812 27412
rect 31760 26920 31812 26926
rect 31760 26862 31812 26868
rect 31772 25362 31800 26862
rect 31760 25356 31812 25362
rect 31760 25298 31812 25304
rect 31852 24404 31904 24410
rect 31852 24346 31904 24352
rect 31576 24268 31628 24274
rect 31576 24210 31628 24216
rect 31392 24132 31444 24138
rect 31392 24074 31444 24080
rect 31576 23860 31628 23866
rect 31576 23802 31628 23808
rect 31588 23746 31616 23802
rect 30656 23724 30708 23730
rect 31312 23718 31616 23746
rect 31666 23760 31722 23769
rect 31666 23695 31668 23704
rect 30656 23666 30708 23672
rect 31720 23695 31722 23704
rect 31668 23666 31720 23672
rect 28632 23656 28684 23662
rect 28632 23598 28684 23604
rect 30380 23656 30432 23662
rect 30380 23598 30432 23604
rect 30472 23656 30524 23662
rect 30472 23598 30524 23604
rect 29920 23588 29972 23594
rect 29920 23530 29972 23536
rect 29368 23248 29420 23254
rect 29368 23190 29420 23196
rect 29460 23248 29512 23254
rect 29460 23190 29512 23196
rect 28632 23112 28684 23118
rect 28632 23054 28684 23060
rect 28540 22092 28592 22098
rect 28540 22034 28592 22040
rect 28448 21616 28500 21622
rect 28448 21558 28500 21564
rect 28552 21554 28580 22034
rect 28540 21548 28592 21554
rect 28540 21490 28592 21496
rect 28552 21457 28580 21490
rect 28538 21448 28594 21457
rect 28538 21383 28594 21392
rect 28264 21344 28316 21350
rect 28264 21286 28316 21292
rect 28170 21176 28226 21185
rect 28170 21111 28226 21120
rect 28172 20936 28224 20942
rect 28172 20878 28224 20884
rect 28184 20777 28212 20878
rect 28170 20768 28226 20777
rect 28170 20703 28226 20712
rect 28276 20618 28304 21286
rect 28448 21140 28500 21146
rect 28448 21082 28500 21088
rect 28276 20590 28396 20618
rect 28264 20460 28316 20466
rect 28264 20402 28316 20408
rect 28276 20058 28304 20402
rect 28264 20052 28316 20058
rect 28264 19994 28316 20000
rect 28172 18760 28224 18766
rect 28172 18702 28224 18708
rect 28184 18426 28212 18702
rect 28172 18420 28224 18426
rect 28172 18362 28224 18368
rect 28172 18284 28224 18290
rect 28172 18226 28224 18232
rect 28000 10118 28120 10146
rect 27896 9920 27948 9926
rect 27896 9862 27948 9868
rect 28000 9738 28028 10118
rect 28080 10056 28132 10062
rect 28080 9998 28132 10004
rect 27816 9710 28028 9738
rect 27816 9081 27844 9710
rect 27988 9580 28040 9586
rect 27988 9522 28040 9528
rect 27896 9172 27948 9178
rect 27896 9114 27948 9120
rect 27802 9072 27858 9081
rect 27802 9007 27858 9016
rect 27712 8968 27764 8974
rect 27712 8910 27764 8916
rect 27804 8900 27856 8906
rect 27804 8842 27856 8848
rect 27620 8424 27672 8430
rect 27620 8366 27672 8372
rect 27816 8294 27844 8842
rect 27908 8498 27936 9114
rect 28000 8906 28028 9522
rect 28092 9178 28120 9998
rect 28080 9172 28132 9178
rect 28080 9114 28132 9120
rect 27988 8900 28040 8906
rect 27988 8842 28040 8848
rect 27896 8492 27948 8498
rect 27896 8434 27948 8440
rect 27894 8392 27950 8401
rect 27894 8327 27950 8336
rect 27620 8288 27672 8294
rect 27620 8230 27672 8236
rect 27804 8288 27856 8294
rect 27804 8230 27856 8236
rect 27528 8084 27580 8090
rect 27528 8026 27580 8032
rect 27528 7812 27580 7818
rect 27528 7754 27580 7760
rect 27436 7336 27488 7342
rect 27436 7278 27488 7284
rect 27448 6798 27476 7278
rect 26240 6792 26292 6798
rect 26240 6734 26292 6740
rect 27068 6792 27120 6798
rect 27068 6734 27120 6740
rect 27160 6792 27212 6798
rect 27160 6734 27212 6740
rect 27436 6792 27488 6798
rect 27436 6734 27488 6740
rect 26148 6248 26200 6254
rect 26148 6190 26200 6196
rect 25964 3936 26016 3942
rect 25964 3878 26016 3884
rect 25976 3602 26004 3878
rect 25964 3596 26016 3602
rect 25964 3538 26016 3544
rect 25780 3528 25832 3534
rect 25780 3470 25832 3476
rect 25688 3460 25740 3466
rect 25688 3402 25740 3408
rect 25504 3392 25556 3398
rect 25504 3334 25556 3340
rect 25792 3058 25820 3470
rect 26160 3194 26188 6190
rect 27540 3670 27568 7754
rect 27632 7206 27660 8230
rect 27804 7744 27856 7750
rect 27804 7686 27856 7692
rect 27816 7274 27844 7686
rect 27804 7268 27856 7274
rect 27804 7210 27856 7216
rect 27620 7200 27672 7206
rect 27620 7142 27672 7148
rect 27712 6656 27764 6662
rect 27712 6598 27764 6604
rect 27724 6322 27752 6598
rect 27712 6316 27764 6322
rect 27712 6258 27764 6264
rect 27908 4690 27936 8327
rect 28000 7886 28028 8842
rect 28080 8356 28132 8362
rect 28080 8298 28132 8304
rect 28092 7954 28120 8298
rect 28080 7948 28132 7954
rect 28080 7890 28132 7896
rect 27988 7880 28040 7886
rect 27988 7822 28040 7828
rect 27896 4684 27948 4690
rect 27896 4626 27948 4632
rect 26884 3664 26936 3670
rect 26884 3606 26936 3612
rect 27528 3664 27580 3670
rect 27528 3606 27580 3612
rect 26424 3596 26476 3602
rect 26424 3538 26476 3544
rect 26148 3188 26200 3194
rect 26148 3130 26200 3136
rect 25780 3052 25832 3058
rect 25780 2994 25832 3000
rect 24676 2508 24728 2514
rect 24676 2450 24728 2456
rect 26148 2508 26200 2514
rect 26148 2450 26200 2456
rect 25136 2372 25188 2378
rect 25136 2314 25188 2320
rect 24492 2304 24544 2310
rect 24492 2246 24544 2252
rect 24308 2032 24360 2038
rect 24308 1974 24360 1980
rect 24504 800 24532 2246
rect 25148 800 25176 2314
rect 26160 2310 26188 2450
rect 26148 2304 26200 2310
rect 26148 2246 26200 2252
rect 26436 800 26464 3538
rect 26896 2854 26924 3606
rect 26884 2848 26936 2854
rect 26884 2790 26936 2796
rect 28184 2774 28212 18226
rect 28276 12102 28304 19994
rect 28368 18290 28396 20590
rect 28460 19854 28488 21082
rect 28540 20936 28592 20942
rect 28540 20878 28592 20884
rect 28552 19922 28580 20878
rect 28540 19916 28592 19922
rect 28540 19858 28592 19864
rect 28448 19848 28500 19854
rect 28448 19790 28500 19796
rect 28448 19440 28500 19446
rect 28448 19382 28500 19388
rect 28356 18284 28408 18290
rect 28356 18226 28408 18232
rect 28356 16108 28408 16114
rect 28356 16050 28408 16056
rect 28368 14074 28396 16050
rect 28356 14068 28408 14074
rect 28356 14010 28408 14016
rect 28354 13968 28410 13977
rect 28354 13903 28410 13912
rect 28368 12782 28396 13903
rect 28356 12776 28408 12782
rect 28356 12718 28408 12724
rect 28460 12628 28488 19382
rect 28368 12600 28488 12628
rect 28264 12096 28316 12102
rect 28264 12038 28316 12044
rect 28264 11688 28316 11694
rect 28264 11630 28316 11636
rect 28276 11286 28304 11630
rect 28264 11280 28316 11286
rect 28264 11222 28316 11228
rect 28264 11144 28316 11150
rect 28264 11086 28316 11092
rect 28276 8809 28304 11086
rect 28262 8800 28318 8809
rect 28262 8735 28318 8744
rect 28264 8560 28316 8566
rect 28264 8502 28316 8508
rect 28276 7546 28304 8502
rect 28264 7540 28316 7546
rect 28264 7482 28316 7488
rect 28368 2774 28396 12600
rect 28552 12209 28580 19858
rect 28644 17785 28672 23054
rect 29380 23050 29408 23190
rect 29368 23044 29420 23050
rect 29368 22986 29420 22992
rect 29380 22438 29408 22986
rect 29472 22642 29500 23190
rect 29644 23180 29696 23186
rect 29644 23122 29696 23128
rect 29656 22642 29684 23122
rect 29460 22636 29512 22642
rect 29460 22578 29512 22584
rect 29644 22636 29696 22642
rect 29644 22578 29696 22584
rect 29368 22432 29420 22438
rect 29368 22374 29420 22380
rect 29472 22234 29500 22578
rect 29552 22568 29604 22574
rect 29552 22510 29604 22516
rect 29460 22228 29512 22234
rect 29460 22170 29512 22176
rect 28722 22128 28778 22137
rect 28722 22063 28724 22072
rect 28776 22063 28778 22072
rect 28724 22034 28776 22040
rect 28816 22024 28868 22030
rect 28814 21992 28816 22001
rect 29564 22001 29592 22510
rect 29736 22228 29788 22234
rect 29788 22188 29868 22216
rect 29736 22170 29788 22176
rect 29642 22128 29698 22137
rect 29642 22063 29644 22072
rect 29696 22063 29698 22072
rect 29644 22034 29696 22040
rect 29736 22024 29788 22030
rect 28868 21992 28870 22001
rect 29550 21992 29606 22001
rect 28814 21927 28870 21936
rect 29184 21956 29236 21962
rect 29184 21898 29236 21904
rect 29460 21956 29512 21962
rect 29550 21927 29606 21936
rect 29734 21992 29736 22001
rect 29788 21992 29790 22001
rect 29734 21927 29790 21936
rect 29460 21898 29512 21904
rect 29092 21888 29144 21894
rect 29092 21830 29144 21836
rect 29104 21729 29132 21830
rect 29090 21720 29146 21729
rect 29090 21655 29146 21664
rect 28724 21616 28776 21622
rect 29196 21570 29224 21898
rect 28724 21558 28776 21564
rect 28736 21010 28764 21558
rect 29012 21542 29224 21570
rect 29368 21548 29420 21554
rect 28908 21344 28960 21350
rect 28908 21286 28960 21292
rect 28816 21140 28868 21146
rect 28816 21082 28868 21088
rect 28724 21004 28776 21010
rect 28724 20946 28776 20952
rect 28828 20942 28856 21082
rect 28816 20936 28868 20942
rect 28816 20878 28868 20884
rect 28920 20874 28948 21286
rect 28908 20868 28960 20874
rect 28908 20810 28960 20816
rect 28908 20460 28960 20466
rect 28908 20402 28960 20408
rect 28816 20392 28868 20398
rect 28816 20334 28868 20340
rect 28828 19854 28856 20334
rect 28816 19848 28868 19854
rect 28816 19790 28868 19796
rect 28724 18692 28776 18698
rect 28724 18634 28776 18640
rect 28736 18222 28764 18634
rect 28724 18216 28776 18222
rect 28724 18158 28776 18164
rect 28724 18080 28776 18086
rect 28724 18022 28776 18028
rect 28630 17776 28686 17785
rect 28630 17711 28686 17720
rect 28632 17672 28684 17678
rect 28632 17614 28684 17620
rect 28644 17134 28672 17614
rect 28632 17128 28684 17134
rect 28632 17070 28684 17076
rect 28644 15638 28672 17070
rect 28632 15632 28684 15638
rect 28632 15574 28684 15580
rect 28644 14958 28672 15574
rect 28736 15094 28764 18022
rect 28724 15088 28776 15094
rect 28724 15030 28776 15036
rect 28632 14952 28684 14958
rect 28632 14894 28684 14900
rect 28724 14340 28776 14346
rect 28724 14282 28776 14288
rect 28736 13938 28764 14282
rect 28724 13932 28776 13938
rect 28724 13874 28776 13880
rect 28736 12434 28764 13874
rect 28644 12406 28764 12434
rect 28538 12200 28594 12209
rect 28538 12135 28594 12144
rect 28540 12096 28592 12102
rect 28540 12038 28592 12044
rect 28448 11756 28500 11762
rect 28448 11698 28500 11704
rect 28460 11354 28488 11698
rect 28448 11348 28500 11354
rect 28448 11290 28500 11296
rect 28552 11234 28580 12038
rect 28644 11762 28672 12406
rect 28828 12322 28856 19790
rect 28920 19446 28948 20402
rect 29012 19854 29040 21542
rect 29368 21490 29420 21496
rect 29184 21344 29236 21350
rect 29184 21286 29236 21292
rect 29276 21344 29328 21350
rect 29276 21286 29328 21292
rect 29092 21004 29144 21010
rect 29092 20946 29144 20952
rect 29104 20330 29132 20946
rect 29092 20324 29144 20330
rect 29196 20312 29224 21286
rect 29288 20777 29316 21286
rect 29274 20768 29330 20777
rect 29274 20703 29330 20712
rect 29276 20324 29328 20330
rect 29196 20284 29276 20312
rect 29092 20266 29144 20272
rect 29276 20266 29328 20272
rect 29000 19848 29052 19854
rect 29000 19790 29052 19796
rect 28908 19440 28960 19446
rect 28908 19382 28960 19388
rect 29000 17264 29052 17270
rect 28998 17232 29000 17241
rect 29052 17232 29054 17241
rect 28908 17196 28960 17202
rect 28998 17167 29054 17176
rect 29092 17196 29144 17202
rect 28908 17138 28960 17144
rect 29092 17138 29144 17144
rect 28920 16794 28948 17138
rect 29000 17128 29052 17134
rect 28998 17096 29000 17105
rect 29052 17096 29054 17105
rect 28998 17031 29054 17040
rect 28908 16788 28960 16794
rect 28908 16730 28960 16736
rect 28908 16584 28960 16590
rect 28908 16526 28960 16532
rect 28920 15162 28948 16526
rect 29104 16114 29132 17138
rect 29000 16108 29052 16114
rect 29000 16050 29052 16056
rect 29092 16108 29144 16114
rect 29092 16050 29144 16056
rect 28908 15156 28960 15162
rect 28908 15098 28960 15104
rect 29012 14618 29040 16050
rect 29104 14958 29132 16050
rect 29182 15056 29238 15065
rect 29182 14991 29184 15000
rect 29236 14991 29238 15000
rect 29184 14962 29236 14968
rect 29092 14952 29144 14958
rect 29288 14906 29316 20266
rect 29380 20058 29408 21490
rect 29472 21486 29500 21898
rect 29840 21690 29868 22188
rect 29932 21894 29960 23530
rect 30564 23520 30616 23526
rect 30564 23462 30616 23468
rect 30576 23118 30604 23462
rect 30564 23112 30616 23118
rect 30564 23054 30616 23060
rect 30472 23044 30524 23050
rect 30472 22986 30524 22992
rect 30288 22976 30340 22982
rect 30288 22918 30340 22924
rect 30196 22228 30248 22234
rect 30196 22170 30248 22176
rect 30208 22137 30236 22170
rect 30194 22128 30250 22137
rect 30194 22063 30250 22072
rect 30012 22024 30064 22030
rect 30012 21966 30064 21972
rect 29920 21888 29972 21894
rect 29920 21830 29972 21836
rect 29828 21684 29880 21690
rect 29828 21626 29880 21632
rect 30024 21622 30052 21966
rect 30012 21616 30064 21622
rect 30012 21558 30064 21564
rect 29460 21480 29512 21486
rect 29460 21422 29512 21428
rect 29460 21344 29512 21350
rect 29458 21312 29460 21321
rect 29512 21312 29514 21321
rect 29458 21247 29514 21256
rect 29458 21176 29514 21185
rect 29458 21111 29514 21120
rect 29472 20262 29500 21111
rect 29918 21040 29974 21049
rect 29918 20975 29974 20984
rect 29932 20806 29960 20975
rect 30010 20904 30066 20913
rect 30010 20839 30066 20848
rect 30024 20806 30052 20839
rect 29920 20800 29972 20806
rect 29920 20742 29972 20748
rect 30012 20800 30064 20806
rect 30012 20742 30064 20748
rect 29460 20256 29512 20262
rect 29460 20198 29512 20204
rect 30196 20256 30248 20262
rect 30196 20198 30248 20204
rect 29368 20052 29420 20058
rect 29368 19994 29420 20000
rect 29472 17610 29500 20198
rect 30208 19922 30236 20198
rect 30196 19916 30248 19922
rect 30196 19858 30248 19864
rect 30300 19854 30328 22918
rect 30484 21865 30512 22986
rect 30668 22094 30696 23666
rect 30748 23656 30800 23662
rect 30748 23598 30800 23604
rect 30760 23526 30788 23598
rect 30748 23520 30800 23526
rect 30748 23462 30800 23468
rect 31024 23520 31076 23526
rect 31024 23462 31076 23468
rect 30932 22976 30984 22982
rect 30932 22918 30984 22924
rect 30840 22772 30892 22778
rect 30840 22714 30892 22720
rect 30748 22704 30800 22710
rect 30746 22672 30748 22681
rect 30800 22672 30802 22681
rect 30852 22642 30880 22714
rect 30746 22607 30802 22616
rect 30840 22636 30892 22642
rect 30840 22578 30892 22584
rect 30840 22228 30892 22234
rect 30840 22170 30892 22176
rect 30576 22066 30696 22094
rect 30470 21856 30526 21865
rect 30470 21791 30526 21800
rect 30380 20324 30432 20330
rect 30380 20266 30432 20272
rect 30392 20058 30420 20266
rect 30576 20058 30604 22066
rect 30748 21548 30800 21554
rect 30748 21490 30800 21496
rect 30656 21004 30708 21010
rect 30656 20946 30708 20952
rect 30380 20052 30432 20058
rect 30380 19994 30432 20000
rect 30564 20052 30616 20058
rect 30564 19994 30616 20000
rect 30668 19922 30696 20946
rect 30760 20262 30788 21490
rect 30852 20534 30880 22170
rect 30944 22098 30972 22918
rect 30932 22092 30984 22098
rect 30932 22034 30984 22040
rect 30932 21480 30984 21486
rect 30932 21422 30984 21428
rect 30944 21350 30972 21422
rect 30932 21344 30984 21350
rect 30932 21286 30984 21292
rect 30840 20528 30892 20534
rect 30840 20470 30892 20476
rect 30748 20256 30800 20262
rect 30748 20198 30800 20204
rect 30656 19916 30708 19922
rect 30656 19858 30708 19864
rect 30288 19848 30340 19854
rect 30288 19790 30340 19796
rect 29644 18692 29696 18698
rect 29644 18634 29696 18640
rect 29552 18624 29604 18630
rect 29552 18566 29604 18572
rect 29564 18358 29592 18566
rect 29552 18352 29604 18358
rect 29552 18294 29604 18300
rect 29656 18170 29684 18634
rect 29564 18142 29684 18170
rect 29564 18086 29592 18142
rect 29552 18080 29604 18086
rect 29552 18022 29604 18028
rect 29564 17678 29592 18022
rect 29920 17876 29972 17882
rect 29920 17818 29972 17824
rect 29552 17672 29604 17678
rect 29552 17614 29604 17620
rect 29460 17604 29512 17610
rect 29460 17546 29512 17552
rect 29564 17218 29592 17614
rect 29932 17610 29960 17818
rect 29828 17604 29880 17610
rect 29828 17546 29880 17552
rect 29920 17604 29972 17610
rect 29920 17546 29972 17552
rect 29840 17338 29868 17546
rect 29828 17332 29880 17338
rect 29828 17274 29880 17280
rect 29460 17196 29512 17202
rect 29564 17190 29868 17218
rect 29460 17138 29512 17144
rect 29472 17105 29500 17138
rect 29644 17128 29696 17134
rect 29458 17096 29514 17105
rect 29644 17070 29696 17076
rect 29458 17031 29514 17040
rect 29552 16108 29604 16114
rect 29552 16050 29604 16056
rect 29460 15564 29512 15570
rect 29460 15506 29512 15512
rect 29092 14894 29144 14900
rect 29000 14612 29052 14618
rect 29000 14554 29052 14560
rect 28908 14408 28960 14414
rect 28908 14350 28960 14356
rect 28920 14226 28948 14350
rect 28920 14198 29040 14226
rect 28908 14068 28960 14074
rect 28908 14010 28960 14016
rect 28736 12294 28856 12322
rect 28632 11756 28684 11762
rect 28632 11698 28684 11704
rect 28092 2746 28212 2774
rect 28276 2746 28396 2774
rect 28460 11206 28580 11234
rect 28092 2582 28120 2746
rect 28080 2576 28132 2582
rect 28080 2518 28132 2524
rect 28276 2446 28304 2746
rect 27068 2440 27120 2446
rect 27068 2382 27120 2388
rect 28264 2440 28316 2446
rect 28264 2382 28316 2388
rect 27080 800 27108 2382
rect 28460 2378 28488 11206
rect 28540 11076 28592 11082
rect 28540 11018 28592 11024
rect 28552 10146 28580 11018
rect 28644 10810 28672 11698
rect 28736 11150 28764 12294
rect 28814 12200 28870 12209
rect 28814 12135 28870 12144
rect 28724 11144 28776 11150
rect 28724 11086 28776 11092
rect 28724 11008 28776 11014
rect 28724 10950 28776 10956
rect 28632 10804 28684 10810
rect 28632 10746 28684 10752
rect 28736 10266 28764 10950
rect 28724 10260 28776 10266
rect 28724 10202 28776 10208
rect 28552 10118 28764 10146
rect 28540 9580 28592 9586
rect 28540 9522 28592 9528
rect 28552 9382 28580 9522
rect 28540 9376 28592 9382
rect 28540 9318 28592 9324
rect 28552 8974 28580 9318
rect 28540 8968 28592 8974
rect 28540 8910 28592 8916
rect 28632 8900 28684 8906
rect 28632 8842 28684 8848
rect 28538 8800 28594 8809
rect 28538 8735 28594 8744
rect 28552 8514 28580 8735
rect 28644 8634 28672 8842
rect 28632 8628 28684 8634
rect 28632 8570 28684 8576
rect 28552 8486 28672 8514
rect 28540 7404 28592 7410
rect 28540 7346 28592 7352
rect 28552 7206 28580 7346
rect 28540 7200 28592 7206
rect 28540 7142 28592 7148
rect 28552 6730 28580 7142
rect 28540 6724 28592 6730
rect 28540 6666 28592 6672
rect 28644 5574 28672 8486
rect 28736 6866 28764 10118
rect 28724 6860 28776 6866
rect 28724 6802 28776 6808
rect 28632 5568 28684 5574
rect 28632 5510 28684 5516
rect 28828 2774 28856 12135
rect 28920 11830 28948 14010
rect 29012 13802 29040 14198
rect 29000 13796 29052 13802
rect 29000 13738 29052 13744
rect 29000 13320 29052 13326
rect 29000 13262 29052 13268
rect 28908 11824 28960 11830
rect 28908 11766 28960 11772
rect 29012 11626 29040 13262
rect 29104 12986 29132 14894
rect 29196 14878 29316 14906
rect 29092 12980 29144 12986
rect 29092 12922 29144 12928
rect 29000 11620 29052 11626
rect 29000 11562 29052 11568
rect 28908 10124 28960 10130
rect 28908 10066 28960 10072
rect 28920 8838 28948 10066
rect 28998 9480 29054 9489
rect 28998 9415 29000 9424
rect 29052 9415 29054 9424
rect 29000 9386 29052 9392
rect 28908 8832 28960 8838
rect 28908 8774 28960 8780
rect 28908 8288 28960 8294
rect 28908 8230 28960 8236
rect 28920 6798 28948 8230
rect 28908 6792 28960 6798
rect 28908 6734 28960 6740
rect 28920 6458 28948 6734
rect 28908 6452 28960 6458
rect 28908 6394 28960 6400
rect 29196 4146 29224 14878
rect 29276 14816 29328 14822
rect 29276 14758 29328 14764
rect 29288 13938 29316 14758
rect 29276 13932 29328 13938
rect 29276 13874 29328 13880
rect 29472 13870 29500 15506
rect 29564 15434 29592 16050
rect 29656 16046 29684 17070
rect 29644 16040 29696 16046
rect 29644 15982 29696 15988
rect 29552 15428 29604 15434
rect 29552 15370 29604 15376
rect 29656 14958 29684 15982
rect 29840 15910 29868 17190
rect 30380 16176 30432 16182
rect 30380 16118 30432 16124
rect 29736 15904 29788 15910
rect 29736 15846 29788 15852
rect 29828 15904 29880 15910
rect 29828 15846 29880 15852
rect 29748 15570 29776 15846
rect 29736 15564 29788 15570
rect 29736 15506 29788 15512
rect 29840 15502 29868 15846
rect 30012 15700 30064 15706
rect 30012 15642 30064 15648
rect 29828 15496 29880 15502
rect 29828 15438 29880 15444
rect 29552 14952 29604 14958
rect 29552 14894 29604 14900
rect 29644 14952 29696 14958
rect 29644 14894 29696 14900
rect 29564 14618 29592 14894
rect 29552 14612 29604 14618
rect 29552 14554 29604 14560
rect 29564 13938 29592 14554
rect 29552 13932 29604 13938
rect 29552 13874 29604 13880
rect 29460 13864 29512 13870
rect 29460 13806 29512 13812
rect 29472 13530 29500 13806
rect 29460 13524 29512 13530
rect 29460 13466 29512 13472
rect 29460 13252 29512 13258
rect 29460 13194 29512 13200
rect 29276 12844 29328 12850
rect 29276 12786 29328 12792
rect 29288 12730 29316 12786
rect 29472 12782 29500 13194
rect 29656 13190 29684 14894
rect 29736 14884 29788 14890
rect 29736 14826 29788 14832
rect 29748 14521 29776 14826
rect 29734 14512 29790 14521
rect 29840 14482 29868 15438
rect 30024 14550 30052 15642
rect 30392 15502 30420 16118
rect 30472 15972 30524 15978
rect 30472 15914 30524 15920
rect 30380 15496 30432 15502
rect 30380 15438 30432 15444
rect 30484 15366 30512 15914
rect 30472 15360 30524 15366
rect 30472 15302 30524 15308
rect 30484 15094 30512 15302
rect 30472 15088 30524 15094
rect 30286 15056 30342 15065
rect 30472 15030 30524 15036
rect 30286 14991 30342 15000
rect 30656 15020 30708 15026
rect 30300 14958 30328 14991
rect 30656 14962 30708 14968
rect 30288 14952 30340 14958
rect 30288 14894 30340 14900
rect 30104 14816 30156 14822
rect 30104 14758 30156 14764
rect 30380 14816 30432 14822
rect 30380 14758 30432 14764
rect 30012 14544 30064 14550
rect 30012 14486 30064 14492
rect 29734 14447 29790 14456
rect 29828 14476 29880 14482
rect 29828 14418 29880 14424
rect 30116 14414 30144 14758
rect 30012 14408 30064 14414
rect 29932 14368 30012 14396
rect 29932 13530 29960 14368
rect 30012 14350 30064 14356
rect 30104 14408 30156 14414
rect 30104 14350 30156 14356
rect 29920 13524 29972 13530
rect 29920 13466 29972 13472
rect 29736 13320 29788 13326
rect 29736 13262 29788 13268
rect 29644 13184 29696 13190
rect 29644 13126 29696 13132
rect 29748 12918 29776 13262
rect 29736 12912 29788 12918
rect 29736 12854 29788 12860
rect 29460 12776 29512 12782
rect 29288 12702 29408 12730
rect 29460 12718 29512 12724
rect 29380 12238 29408 12702
rect 29368 12232 29420 12238
rect 29368 12174 29420 12180
rect 29472 10130 29500 12718
rect 29932 12306 29960 13466
rect 30392 13394 30420 14758
rect 30668 14618 30696 14962
rect 30656 14612 30708 14618
rect 30656 14554 30708 14560
rect 30564 14408 30616 14414
rect 30564 14350 30616 14356
rect 30380 13388 30432 13394
rect 30380 13330 30432 13336
rect 30012 13320 30064 13326
rect 30064 13268 30328 13274
rect 30012 13262 30328 13268
rect 30024 13246 30328 13262
rect 30012 13184 30064 13190
rect 30012 13126 30064 13132
rect 30196 13184 30248 13190
rect 30196 13126 30248 13132
rect 30024 12986 30052 13126
rect 30012 12980 30064 12986
rect 30012 12922 30064 12928
rect 29920 12300 29972 12306
rect 29920 12242 29972 12248
rect 30208 12238 30236 13126
rect 30012 12232 30064 12238
rect 30196 12232 30248 12238
rect 30064 12180 30144 12186
rect 30012 12174 30144 12180
rect 30196 12174 30248 12180
rect 30024 12158 30144 12174
rect 29644 12096 29696 12102
rect 29644 12038 29696 12044
rect 29656 11694 29684 12038
rect 29828 11756 29880 11762
rect 29828 11698 29880 11704
rect 29644 11688 29696 11694
rect 29644 11630 29696 11636
rect 29840 11370 29868 11698
rect 30012 11552 30064 11558
rect 30012 11494 30064 11500
rect 29840 11354 29960 11370
rect 29840 11348 29972 11354
rect 29840 11342 29920 11348
rect 29460 10124 29512 10130
rect 29460 10066 29512 10072
rect 29472 9518 29500 10066
rect 29840 9926 29868 11342
rect 29920 11290 29972 11296
rect 30024 11150 30052 11494
rect 30012 11144 30064 11150
rect 30012 11086 30064 11092
rect 29920 11076 29972 11082
rect 29920 11018 29972 11024
rect 29932 10062 29960 11018
rect 30012 11008 30064 11014
rect 30012 10950 30064 10956
rect 30024 10538 30052 10950
rect 30012 10532 30064 10538
rect 30012 10474 30064 10480
rect 30024 10062 30052 10474
rect 29920 10056 29972 10062
rect 29920 9998 29972 10004
rect 30012 10056 30064 10062
rect 30012 9998 30064 10004
rect 29828 9920 29880 9926
rect 29828 9862 29880 9868
rect 29460 9512 29512 9518
rect 29460 9454 29512 9460
rect 29552 8968 29604 8974
rect 29552 8910 29604 8916
rect 29460 8900 29512 8906
rect 29460 8842 29512 8848
rect 29368 7744 29420 7750
rect 29368 7686 29420 7692
rect 29380 7410 29408 7686
rect 29472 7410 29500 8842
rect 29564 8498 29592 8910
rect 29552 8492 29604 8498
rect 29552 8434 29604 8440
rect 29564 7954 29592 8434
rect 29644 8424 29696 8430
rect 29644 8366 29696 8372
rect 29552 7948 29604 7954
rect 29552 7890 29604 7896
rect 29368 7404 29420 7410
rect 29368 7346 29420 7352
rect 29460 7404 29512 7410
rect 29460 7346 29512 7352
rect 29472 7290 29500 7346
rect 29380 7262 29500 7290
rect 29276 6996 29328 7002
rect 29276 6938 29328 6944
rect 28908 4140 28960 4146
rect 28908 4082 28960 4088
rect 29184 4140 29236 4146
rect 29184 4082 29236 4088
rect 28920 3194 28948 4082
rect 29288 3534 29316 6938
rect 29380 6934 29408 7262
rect 29368 6928 29420 6934
rect 29368 6870 29420 6876
rect 29564 6798 29592 7890
rect 29656 7342 29684 8366
rect 29840 8362 29868 9862
rect 29932 9722 29960 9998
rect 29920 9716 29972 9722
rect 29920 9658 29972 9664
rect 29920 9580 29972 9586
rect 29920 9522 29972 9528
rect 29932 9110 29960 9522
rect 29920 9104 29972 9110
rect 29920 9046 29972 9052
rect 30024 8974 30052 9998
rect 30116 9586 30144 12158
rect 30300 9586 30328 13246
rect 30392 12850 30420 13330
rect 30576 13326 30604 14350
rect 30564 13320 30616 13326
rect 30564 13262 30616 13268
rect 30380 12844 30432 12850
rect 30380 12786 30432 12792
rect 30104 9580 30156 9586
rect 30104 9522 30156 9528
rect 30288 9580 30340 9586
rect 30288 9522 30340 9528
rect 30012 8968 30064 8974
rect 30012 8910 30064 8916
rect 30116 8906 30144 9522
rect 30196 9512 30248 9518
rect 30196 9454 30248 9460
rect 30208 9178 30236 9454
rect 30656 9376 30708 9382
rect 30656 9318 30708 9324
rect 30196 9172 30248 9178
rect 30196 9114 30248 9120
rect 30104 8900 30156 8906
rect 30104 8842 30156 8848
rect 30208 8566 30236 9114
rect 30668 8974 30696 9318
rect 30656 8968 30708 8974
rect 30656 8910 30708 8916
rect 30196 8560 30248 8566
rect 30196 8502 30248 8508
rect 29828 8356 29880 8362
rect 29828 8298 29880 8304
rect 29644 7336 29696 7342
rect 29644 7278 29696 7284
rect 29552 6792 29604 6798
rect 29552 6734 29604 6740
rect 29564 6390 29592 6734
rect 29656 6662 29684 7278
rect 29920 7268 29972 7274
rect 29920 7210 29972 7216
rect 29644 6656 29696 6662
rect 29644 6598 29696 6604
rect 29552 6384 29604 6390
rect 29552 6326 29604 6332
rect 29932 5114 29960 7210
rect 30104 7200 30156 7206
rect 30104 7142 30156 7148
rect 30116 6798 30144 7142
rect 30104 6792 30156 6798
rect 30104 6734 30156 6740
rect 29564 5086 29960 5114
rect 29460 4208 29512 4214
rect 29460 4150 29512 4156
rect 29000 3528 29052 3534
rect 29000 3470 29052 3476
rect 29276 3528 29328 3534
rect 29276 3470 29328 3476
rect 28908 3188 28960 3194
rect 28908 3130 28960 3136
rect 28736 2746 28856 2774
rect 28736 2514 28764 2746
rect 29012 2514 29040 3470
rect 29472 3398 29500 4150
rect 29460 3392 29512 3398
rect 29460 3334 29512 3340
rect 29564 2774 29592 5086
rect 29828 4140 29880 4146
rect 29828 4082 29880 4088
rect 29736 3936 29788 3942
rect 29736 3878 29788 3884
rect 29644 3460 29696 3466
rect 29644 3402 29696 3408
rect 29656 2836 29684 3402
rect 29748 3058 29776 3878
rect 29840 3466 29868 4082
rect 29828 3460 29880 3466
rect 29828 3402 29880 3408
rect 29920 3392 29972 3398
rect 29920 3334 29972 3340
rect 29932 3126 29960 3334
rect 29920 3120 29972 3126
rect 29920 3062 29972 3068
rect 29736 3052 29788 3058
rect 29736 2994 29788 3000
rect 30288 2984 30340 2990
rect 30288 2926 30340 2932
rect 29656 2808 29776 2836
rect 29564 2746 29684 2774
rect 28724 2508 28776 2514
rect 28724 2450 28776 2456
rect 29000 2508 29052 2514
rect 29000 2450 29052 2456
rect 27712 2372 27764 2378
rect 27712 2314 27764 2320
rect 28448 2372 28500 2378
rect 28448 2314 28500 2320
rect 27724 800 27752 2314
rect 29656 800 29684 2746
rect 29748 2514 29776 2808
rect 29736 2508 29788 2514
rect 29736 2450 29788 2456
rect 30300 800 30328 2926
rect 30760 2922 30788 20198
rect 30852 20058 30880 20470
rect 30944 20466 30972 21286
rect 31036 21146 31064 23462
rect 31116 23316 31168 23322
rect 31116 23258 31168 23264
rect 31128 23050 31156 23258
rect 31116 23044 31168 23050
rect 31116 22986 31168 22992
rect 31128 22794 31156 22986
rect 31128 22766 31248 22794
rect 31116 22704 31168 22710
rect 31116 22646 31168 22652
rect 31024 21140 31076 21146
rect 31024 21082 31076 21088
rect 31128 20806 31156 22646
rect 31220 21962 31248 22766
rect 31484 22636 31536 22642
rect 31484 22578 31536 22584
rect 31392 22500 31444 22506
rect 31392 22442 31444 22448
rect 31404 22094 31432 22442
rect 31496 22234 31524 22578
rect 31576 22568 31628 22574
rect 31576 22510 31628 22516
rect 31484 22228 31536 22234
rect 31484 22170 31536 22176
rect 31404 22066 31524 22094
rect 31392 22024 31444 22030
rect 31392 21966 31444 21972
rect 31208 21956 31260 21962
rect 31208 21898 31260 21904
rect 31300 21956 31352 21962
rect 31300 21898 31352 21904
rect 31312 21690 31340 21898
rect 31300 21684 31352 21690
rect 31300 21626 31352 21632
rect 31404 21468 31432 21966
rect 31496 21593 31524 22066
rect 31588 21690 31616 22510
rect 31576 21684 31628 21690
rect 31576 21626 31628 21632
rect 31482 21584 31538 21593
rect 31482 21519 31538 21528
rect 31404 21440 31524 21468
rect 31392 20936 31444 20942
rect 31392 20878 31444 20884
rect 31208 20868 31260 20874
rect 31208 20810 31260 20816
rect 31116 20800 31168 20806
rect 31116 20742 31168 20748
rect 30932 20460 30984 20466
rect 30932 20402 30984 20408
rect 30840 20052 30892 20058
rect 30840 19994 30892 20000
rect 31114 18456 31170 18465
rect 31114 18391 31170 18400
rect 30840 18284 30892 18290
rect 30840 18226 30892 18232
rect 30852 16114 30880 18226
rect 30932 17536 30984 17542
rect 30932 17478 30984 17484
rect 30944 17066 30972 17478
rect 31022 17096 31078 17105
rect 30932 17060 30984 17066
rect 31022 17031 31078 17040
rect 30932 17002 30984 17008
rect 31036 16998 31064 17031
rect 31024 16992 31076 16998
rect 31024 16934 31076 16940
rect 31024 16244 31076 16250
rect 31024 16186 31076 16192
rect 30840 16108 30892 16114
rect 30840 16050 30892 16056
rect 31036 15434 31064 16186
rect 31024 15428 31076 15434
rect 31024 15370 31076 15376
rect 30930 15328 30986 15337
rect 30930 15263 30986 15272
rect 30944 15162 30972 15263
rect 31128 15162 31156 18391
rect 30840 15156 30892 15162
rect 30840 15098 30892 15104
rect 30932 15156 30984 15162
rect 30932 15098 30984 15104
rect 31116 15156 31168 15162
rect 31116 15098 31168 15104
rect 30852 13462 30880 15098
rect 30932 14272 30984 14278
rect 30932 14214 30984 14220
rect 30840 13456 30892 13462
rect 30840 13398 30892 13404
rect 30944 13326 30972 14214
rect 31220 13802 31248 20810
rect 31404 20534 31432 20878
rect 31392 20528 31444 20534
rect 31392 20470 31444 20476
rect 31496 20398 31524 21440
rect 31576 21072 31628 21078
rect 31574 21040 31576 21049
rect 31628 21040 31630 21049
rect 31574 20975 31630 20984
rect 31680 20942 31708 23666
rect 31760 21344 31812 21350
rect 31760 21286 31812 21292
rect 31668 20936 31720 20942
rect 31668 20878 31720 20884
rect 31772 20874 31800 21286
rect 31760 20868 31812 20874
rect 31760 20810 31812 20816
rect 31484 20392 31536 20398
rect 31484 20334 31536 20340
rect 31392 20324 31444 20330
rect 31392 20266 31444 20272
rect 31404 19990 31432 20266
rect 31392 19984 31444 19990
rect 31392 19926 31444 19932
rect 31300 16992 31352 16998
rect 31300 16934 31352 16940
rect 31312 16658 31340 16934
rect 31300 16652 31352 16658
rect 31300 16594 31352 16600
rect 31208 13796 31260 13802
rect 31208 13738 31260 13744
rect 30932 13320 30984 13326
rect 30932 13262 30984 13268
rect 31300 12844 31352 12850
rect 31300 12786 31352 12792
rect 31312 12442 31340 12786
rect 31300 12436 31352 12442
rect 31300 12378 31352 12384
rect 31392 9580 31444 9586
rect 31392 9522 31444 9528
rect 30840 9444 30892 9450
rect 30840 9386 30892 9392
rect 30852 3194 30880 9386
rect 31404 9382 31432 9522
rect 31392 9376 31444 9382
rect 31392 9318 31444 9324
rect 31496 9110 31524 20334
rect 31760 19712 31812 19718
rect 31760 19654 31812 19660
rect 31772 17678 31800 19654
rect 31668 17672 31720 17678
rect 31668 17614 31720 17620
rect 31760 17672 31812 17678
rect 31760 17614 31812 17620
rect 31680 17134 31708 17614
rect 31668 17128 31720 17134
rect 31668 17070 31720 17076
rect 31668 14952 31720 14958
rect 31668 14894 31720 14900
rect 31576 13796 31628 13802
rect 31576 13738 31628 13744
rect 31588 12434 31616 13738
rect 31680 13138 31708 14894
rect 31772 13326 31800 17614
rect 31760 13320 31812 13326
rect 31760 13262 31812 13268
rect 31680 13110 31800 13138
rect 31772 12782 31800 13110
rect 31760 12776 31812 12782
rect 31760 12718 31812 12724
rect 31864 12434 31892 24346
rect 32140 23882 32168 31726
rect 32220 31340 32272 31346
rect 32220 31282 32272 31288
rect 32232 30938 32260 31282
rect 32220 30932 32272 30938
rect 32220 30874 32272 30880
rect 32324 27470 32352 36722
rect 32588 35556 32640 35562
rect 32588 35498 32640 35504
rect 32496 33992 32548 33998
rect 32600 33980 32628 35498
rect 32548 33952 32628 33980
rect 32496 33934 32548 33940
rect 32496 33516 32548 33522
rect 32496 33458 32548 33464
rect 32508 32842 32536 33458
rect 32600 32910 32628 33952
rect 32588 32904 32640 32910
rect 32588 32846 32640 32852
rect 32496 32836 32548 32842
rect 32496 32778 32548 32784
rect 32496 31816 32548 31822
rect 32496 31758 32548 31764
rect 32772 31816 32824 31822
rect 32772 31758 32824 31764
rect 32404 31748 32456 31754
rect 32404 31690 32456 31696
rect 32416 30122 32444 31690
rect 32508 31414 32536 31758
rect 32784 31482 32812 31758
rect 32968 31754 32996 40530
rect 33336 40526 33364 41414
rect 33324 40520 33376 40526
rect 33324 40462 33376 40468
rect 33416 40384 33468 40390
rect 33416 40326 33468 40332
rect 33428 40186 33456 40326
rect 33416 40180 33468 40186
rect 33416 40122 33468 40128
rect 33232 40044 33284 40050
rect 33232 39986 33284 39992
rect 33244 39506 33272 39986
rect 33232 39500 33284 39506
rect 33232 39442 33284 39448
rect 33324 39500 33376 39506
rect 33324 39442 33376 39448
rect 33336 39370 33364 39442
rect 33324 39364 33376 39370
rect 33324 39306 33376 39312
rect 33336 39030 33364 39306
rect 33324 39024 33376 39030
rect 33324 38966 33376 38972
rect 33140 38344 33192 38350
rect 33140 38286 33192 38292
rect 33152 38214 33180 38286
rect 33140 38208 33192 38214
rect 33140 38150 33192 38156
rect 33336 37330 33364 38966
rect 33324 37324 33376 37330
rect 33324 37266 33376 37272
rect 33232 37188 33284 37194
rect 33232 37130 33284 37136
rect 33140 37120 33192 37126
rect 33140 37062 33192 37068
rect 33152 36854 33180 37062
rect 33140 36848 33192 36854
rect 33140 36790 33192 36796
rect 33244 36786 33272 37130
rect 33232 36780 33284 36786
rect 33232 36722 33284 36728
rect 33324 36780 33376 36786
rect 33324 36722 33376 36728
rect 33244 36650 33272 36722
rect 33232 36644 33284 36650
rect 33232 36586 33284 36592
rect 33244 36378 33272 36586
rect 33336 36582 33364 36722
rect 33324 36576 33376 36582
rect 33324 36518 33376 36524
rect 33232 36372 33284 36378
rect 33232 36314 33284 36320
rect 33336 36038 33364 36518
rect 33324 36032 33376 36038
rect 33324 35974 33376 35980
rect 33232 34944 33284 34950
rect 33232 34886 33284 34892
rect 33244 34678 33272 34886
rect 33232 34672 33284 34678
rect 33232 34614 33284 34620
rect 33140 33856 33192 33862
rect 33140 33798 33192 33804
rect 33048 33516 33100 33522
rect 33048 33458 33100 33464
rect 33060 32230 33088 33458
rect 33152 32910 33180 33798
rect 33140 32904 33192 32910
rect 33140 32846 33192 32852
rect 33048 32224 33100 32230
rect 33048 32166 33100 32172
rect 32876 31726 32996 31754
rect 32772 31476 32824 31482
rect 32772 31418 32824 31424
rect 32496 31408 32548 31414
rect 32496 31350 32548 31356
rect 32876 30274 32904 31726
rect 33060 31346 33088 32166
rect 33048 31340 33100 31346
rect 33048 31282 33100 31288
rect 32956 30660 33008 30666
rect 32956 30602 33008 30608
rect 32784 30246 32904 30274
rect 32968 30258 32996 30602
rect 32956 30252 33008 30258
rect 32404 30116 32456 30122
rect 32404 30058 32456 30064
rect 32784 30002 32812 30246
rect 32956 30194 33008 30200
rect 33060 30190 33088 31282
rect 33244 30734 33272 34614
rect 33324 34536 33376 34542
rect 33428 34524 33456 40122
rect 33508 39432 33560 39438
rect 33508 39374 33560 39380
rect 33598 39400 33654 39409
rect 33520 39137 33548 39374
rect 33598 39335 33654 39344
rect 33612 39302 33640 39335
rect 33600 39296 33652 39302
rect 33600 39238 33652 39244
rect 33506 39128 33562 39137
rect 33506 39063 33562 39072
rect 33612 39030 33640 39238
rect 33600 39024 33652 39030
rect 33600 38966 33652 38972
rect 33600 37256 33652 37262
rect 33600 37198 33652 37204
rect 33612 36922 33640 37198
rect 33600 36916 33652 36922
rect 33600 36858 33652 36864
rect 33376 34496 33456 34524
rect 33508 34536 33560 34542
rect 33324 34478 33376 34484
rect 33508 34478 33560 34484
rect 33520 34066 33548 34478
rect 33508 34060 33560 34066
rect 33508 34002 33560 34008
rect 33324 33924 33376 33930
rect 33324 33866 33376 33872
rect 33336 33522 33364 33866
rect 33324 33516 33376 33522
rect 33324 33458 33376 33464
rect 33508 31816 33560 31822
rect 33508 31758 33560 31764
rect 33324 31680 33376 31686
rect 33324 31622 33376 31628
rect 33336 31414 33364 31622
rect 33324 31408 33376 31414
rect 33324 31350 33376 31356
rect 33416 31136 33468 31142
rect 33416 31078 33468 31084
rect 33232 30728 33284 30734
rect 33232 30670 33284 30676
rect 33428 30598 33456 31078
rect 33140 30592 33192 30598
rect 33140 30534 33192 30540
rect 33416 30592 33468 30598
rect 33416 30534 33468 30540
rect 33048 30184 33100 30190
rect 33048 30126 33100 30132
rect 32864 30116 32916 30122
rect 32864 30058 32916 30064
rect 32692 29974 32812 30002
rect 32692 29866 32720 29974
rect 32404 29844 32456 29850
rect 32404 29786 32456 29792
rect 32600 29838 32720 29866
rect 32416 29170 32444 29786
rect 32496 29232 32548 29238
rect 32494 29200 32496 29209
rect 32548 29200 32550 29209
rect 32404 29164 32456 29170
rect 32494 29135 32550 29144
rect 32404 29106 32456 29112
rect 32496 29096 32548 29102
rect 32496 29038 32548 29044
rect 32508 28150 32536 29038
rect 32600 28490 32628 29838
rect 32680 29708 32732 29714
rect 32680 29650 32732 29656
rect 32692 29306 32720 29650
rect 32680 29300 32732 29306
rect 32680 29242 32732 29248
rect 32876 29170 32904 30058
rect 33152 29850 33180 30534
rect 33140 29844 33192 29850
rect 33140 29786 33192 29792
rect 33324 29572 33376 29578
rect 33324 29514 33376 29520
rect 33048 29504 33100 29510
rect 33048 29446 33100 29452
rect 33060 29238 33088 29446
rect 33048 29232 33100 29238
rect 33048 29174 33100 29180
rect 32864 29164 32916 29170
rect 32864 29106 32916 29112
rect 33336 28762 33364 29514
rect 33324 28756 33376 28762
rect 33324 28698 33376 28704
rect 32588 28484 32640 28490
rect 32588 28426 32640 28432
rect 32496 28144 32548 28150
rect 32496 28086 32548 28092
rect 32508 28014 32536 28086
rect 32496 28008 32548 28014
rect 32496 27950 32548 27956
rect 32404 27872 32456 27878
rect 32404 27814 32456 27820
rect 32312 27464 32364 27470
rect 32312 27406 32364 27412
rect 32416 27062 32444 27814
rect 32404 27056 32456 27062
rect 32404 26998 32456 27004
rect 32600 25702 32628 28426
rect 32772 27872 32824 27878
rect 32772 27814 32824 27820
rect 32784 26382 32812 27814
rect 32864 27328 32916 27334
rect 32864 27270 32916 27276
rect 32876 26994 32904 27270
rect 32864 26988 32916 26994
rect 32864 26930 32916 26936
rect 33232 26988 33284 26994
rect 33232 26930 33284 26936
rect 32876 26874 32904 26930
rect 32876 26846 32996 26874
rect 32864 26784 32916 26790
rect 32864 26726 32916 26732
rect 32876 26382 32904 26726
rect 32772 26376 32824 26382
rect 32772 26318 32824 26324
rect 32864 26376 32916 26382
rect 32864 26318 32916 26324
rect 32588 25696 32640 25702
rect 32588 25638 32640 25644
rect 32784 25294 32812 26318
rect 32968 26042 32996 26846
rect 33244 26042 33272 26930
rect 32956 26036 33008 26042
rect 32956 25978 33008 25984
rect 33232 26036 33284 26042
rect 33232 25978 33284 25984
rect 32772 25288 32824 25294
rect 32772 25230 32824 25236
rect 32864 24200 32916 24206
rect 32968 24188 32996 25978
rect 33048 25900 33100 25906
rect 33048 25842 33100 25848
rect 33060 25702 33088 25842
rect 33048 25696 33100 25702
rect 33048 25638 33100 25644
rect 33324 25220 33376 25226
rect 33324 25162 33376 25168
rect 33048 24608 33100 24614
rect 33048 24550 33100 24556
rect 33232 24608 33284 24614
rect 33232 24550 33284 24556
rect 32916 24160 32996 24188
rect 32864 24142 32916 24148
rect 32140 23854 32352 23882
rect 32128 23724 32180 23730
rect 32128 23666 32180 23672
rect 32220 23724 32272 23730
rect 32220 23666 32272 23672
rect 32140 23118 32168 23666
rect 32128 23112 32180 23118
rect 32128 23054 32180 23060
rect 32140 22642 32168 23054
rect 32128 22636 32180 22642
rect 32128 22578 32180 22584
rect 32140 22030 32168 22578
rect 32128 22024 32180 22030
rect 32128 21966 32180 21972
rect 31944 21684 31996 21690
rect 31944 21626 31996 21632
rect 31956 21554 31984 21626
rect 31944 21548 31996 21554
rect 31944 21490 31996 21496
rect 32036 21480 32088 21486
rect 32036 21422 32088 21428
rect 32048 20874 32076 21422
rect 32036 20868 32088 20874
rect 32036 20810 32088 20816
rect 31944 20528 31996 20534
rect 31944 20470 31996 20476
rect 31956 18408 31984 20470
rect 32128 19780 32180 19786
rect 32128 19722 32180 19728
rect 32140 19378 32168 19722
rect 32128 19372 32180 19378
rect 32128 19314 32180 19320
rect 32232 18816 32260 23666
rect 32324 23118 32352 23854
rect 32588 23656 32640 23662
rect 32588 23598 32640 23604
rect 32312 23112 32364 23118
rect 32312 23054 32364 23060
rect 32600 21690 32628 23598
rect 32876 22098 32904 24142
rect 33060 23730 33088 24550
rect 33244 24138 33272 24550
rect 33336 24410 33364 25162
rect 33324 24404 33376 24410
rect 33324 24346 33376 24352
rect 33232 24132 33284 24138
rect 33232 24074 33284 24080
rect 33048 23724 33100 23730
rect 33048 23666 33100 23672
rect 32956 23248 33008 23254
rect 32956 23190 33008 23196
rect 32968 22982 32996 23190
rect 33048 23112 33100 23118
rect 33048 23054 33100 23060
rect 33060 22982 33088 23054
rect 32956 22976 33008 22982
rect 32956 22918 33008 22924
rect 33048 22976 33100 22982
rect 33048 22918 33100 22924
rect 32864 22092 32916 22098
rect 32864 22034 32916 22040
rect 32770 21992 32826 22001
rect 32680 21956 32732 21962
rect 32770 21927 32826 21936
rect 32680 21898 32732 21904
rect 32312 21684 32364 21690
rect 32312 21626 32364 21632
rect 32588 21684 32640 21690
rect 32588 21626 32640 21632
rect 32324 21486 32352 21626
rect 32496 21548 32548 21554
rect 32496 21490 32548 21496
rect 32312 21480 32364 21486
rect 32312 21422 32364 21428
rect 32324 21026 32352 21422
rect 32324 20998 32444 21026
rect 32312 19916 32364 19922
rect 32312 19858 32364 19864
rect 32140 18788 32260 18816
rect 32140 18601 32168 18788
rect 32220 18692 32272 18698
rect 32220 18634 32272 18640
rect 32126 18592 32182 18601
rect 32126 18527 32182 18536
rect 32232 18426 32260 18634
rect 32220 18420 32272 18426
rect 31956 18380 32168 18408
rect 32034 18320 32090 18329
rect 32140 18306 32168 18380
rect 32220 18362 32272 18368
rect 32140 18278 32260 18306
rect 32034 18255 32090 18264
rect 31944 17672 31996 17678
rect 31944 17614 31996 17620
rect 31956 17202 31984 17614
rect 31944 17196 31996 17202
rect 31944 17138 31996 17144
rect 31944 16448 31996 16454
rect 31944 16390 31996 16396
rect 31956 16182 31984 16390
rect 31944 16176 31996 16182
rect 31944 16118 31996 16124
rect 31944 14544 31996 14550
rect 31944 14486 31996 14492
rect 31588 12406 31708 12434
rect 31484 9104 31536 9110
rect 31484 9046 31536 9052
rect 30932 7812 30984 7818
rect 30932 7754 30984 7760
rect 30944 7546 30972 7754
rect 30932 7540 30984 7546
rect 30932 7482 30984 7488
rect 31576 7540 31628 7546
rect 31576 7482 31628 7488
rect 31588 7410 31616 7482
rect 31576 7404 31628 7410
rect 31576 7346 31628 7352
rect 31208 4616 31260 4622
rect 31208 4558 31260 4564
rect 30932 4140 30984 4146
rect 30932 4082 30984 4088
rect 30944 4010 30972 4082
rect 30932 4004 30984 4010
rect 30932 3946 30984 3952
rect 31116 4004 31168 4010
rect 31116 3946 31168 3952
rect 31128 3670 31156 3946
rect 31116 3664 31168 3670
rect 31116 3606 31168 3612
rect 31220 3534 31248 4558
rect 31392 3936 31444 3942
rect 31392 3878 31444 3884
rect 31208 3528 31260 3534
rect 31208 3470 31260 3476
rect 31404 3466 31432 3878
rect 31576 3596 31628 3602
rect 31576 3538 31628 3544
rect 31392 3460 31444 3466
rect 31392 3402 31444 3408
rect 30840 3188 30892 3194
rect 30840 3130 30892 3136
rect 30748 2916 30800 2922
rect 30748 2858 30800 2864
rect 30932 2508 30984 2514
rect 30932 2450 30984 2456
rect 30944 800 30972 2450
rect 31588 800 31616 3538
rect 31680 1902 31708 12406
rect 31772 12406 31892 12434
rect 31772 4146 31800 12406
rect 31956 8906 31984 14486
rect 31944 8900 31996 8906
rect 31944 8842 31996 8848
rect 31852 7200 31904 7206
rect 31852 7142 31904 7148
rect 31864 6866 31892 7142
rect 31852 6860 31904 6866
rect 31852 6802 31904 6808
rect 32048 5642 32076 18255
rect 32232 15314 32260 18278
rect 32324 17202 32352 19858
rect 32312 17196 32364 17202
rect 32312 17138 32364 17144
rect 32140 15286 32260 15314
rect 32140 13802 32168 15286
rect 32324 15042 32352 17138
rect 32232 15014 32352 15042
rect 32232 14958 32260 15014
rect 32220 14952 32272 14958
rect 32220 14894 32272 14900
rect 32312 14884 32364 14890
rect 32312 14826 32364 14832
rect 32324 14074 32352 14826
rect 32312 14068 32364 14074
rect 32312 14010 32364 14016
rect 32416 13954 32444 20998
rect 32508 20534 32536 21490
rect 32496 20528 32548 20534
rect 32496 20470 32548 20476
rect 32588 19712 32640 19718
rect 32588 19654 32640 19660
rect 32496 18148 32548 18154
rect 32496 18090 32548 18096
rect 32508 17746 32536 18090
rect 32496 17740 32548 17746
rect 32496 17682 32548 17688
rect 32508 16658 32536 17682
rect 32496 16652 32548 16658
rect 32496 16594 32548 16600
rect 32600 15201 32628 19654
rect 32586 15192 32642 15201
rect 32586 15127 32642 15136
rect 32496 15020 32548 15026
rect 32496 14962 32548 14968
rect 32508 14929 32536 14962
rect 32588 14952 32640 14958
rect 32494 14920 32550 14929
rect 32588 14894 32640 14900
rect 32494 14855 32550 14864
rect 32496 14816 32548 14822
rect 32496 14758 32548 14764
rect 32232 13926 32444 13954
rect 32128 13796 32180 13802
rect 32128 13738 32180 13744
rect 32128 9716 32180 9722
rect 32128 9658 32180 9664
rect 32140 8974 32168 9658
rect 32232 9178 32260 13926
rect 32404 13864 32456 13870
rect 32404 13806 32456 13812
rect 32312 13796 32364 13802
rect 32312 13738 32364 13744
rect 32220 9172 32272 9178
rect 32220 9114 32272 9120
rect 32128 8968 32180 8974
rect 32128 8910 32180 8916
rect 32220 8832 32272 8838
rect 32220 8774 32272 8780
rect 32232 8566 32260 8774
rect 32220 8560 32272 8566
rect 32220 8502 32272 8508
rect 32220 7812 32272 7818
rect 32220 7754 32272 7760
rect 32128 6860 32180 6866
rect 32128 6802 32180 6808
rect 32140 5914 32168 6802
rect 32232 6390 32260 7754
rect 32220 6384 32272 6390
rect 32220 6326 32272 6332
rect 32128 5908 32180 5914
rect 32128 5850 32180 5856
rect 32036 5636 32088 5642
rect 32036 5578 32088 5584
rect 32220 4752 32272 4758
rect 32220 4694 32272 4700
rect 31760 4140 31812 4146
rect 31760 4082 31812 4088
rect 31668 1896 31720 1902
rect 31668 1838 31720 1844
rect 32232 800 32260 4694
rect 32324 2774 32352 13738
rect 32416 13394 32444 13806
rect 32404 13388 32456 13394
rect 32404 13330 32456 13336
rect 32508 13326 32536 14758
rect 32600 14346 32628 14894
rect 32692 14550 32720 21898
rect 32784 21350 32812 21927
rect 32968 21554 32996 22918
rect 32956 21548 33008 21554
rect 32956 21490 33008 21496
rect 32772 21344 32824 21350
rect 32772 21286 32824 21292
rect 32772 18284 32824 18290
rect 32772 18226 32824 18232
rect 32784 16590 32812 18226
rect 32772 16584 32824 16590
rect 32772 16526 32824 16532
rect 32864 16584 32916 16590
rect 32864 16526 32916 16532
rect 32784 15366 32812 16526
rect 32876 15910 32904 16526
rect 32956 16108 33008 16114
rect 32956 16050 33008 16056
rect 32864 15904 32916 15910
rect 32864 15846 32916 15852
rect 32772 15360 32824 15366
rect 32772 15302 32824 15308
rect 32680 14544 32732 14550
rect 32680 14486 32732 14492
rect 32588 14340 32640 14346
rect 32588 14282 32640 14288
rect 32496 13320 32548 13326
rect 32496 13262 32548 13268
rect 32496 13184 32548 13190
rect 32600 13172 32628 14282
rect 32680 14272 32732 14278
rect 32680 14214 32732 14220
rect 32772 14272 32824 14278
rect 32772 14214 32824 14220
rect 32692 13938 32720 14214
rect 32784 14074 32812 14214
rect 32772 14068 32824 14074
rect 32772 14010 32824 14016
rect 32680 13932 32732 13938
rect 32680 13874 32732 13880
rect 32678 13832 32734 13841
rect 32678 13767 32734 13776
rect 32548 13144 32628 13172
rect 32496 13126 32548 13132
rect 32404 12844 32456 12850
rect 32404 12786 32456 12792
rect 32416 11150 32444 12786
rect 32404 11144 32456 11150
rect 32404 11086 32456 11092
rect 32508 10810 32536 13126
rect 32588 12096 32640 12102
rect 32588 12038 32640 12044
rect 32600 11286 32628 12038
rect 32588 11280 32640 11286
rect 32588 11222 32640 11228
rect 32588 11008 32640 11014
rect 32588 10950 32640 10956
rect 32600 10810 32628 10950
rect 32404 10804 32456 10810
rect 32404 10746 32456 10752
rect 32496 10804 32548 10810
rect 32496 10746 32548 10752
rect 32588 10804 32640 10810
rect 32588 10746 32640 10752
rect 32416 9518 32444 10746
rect 32508 10690 32536 10746
rect 32508 10662 32628 10690
rect 32496 10464 32548 10470
rect 32496 10406 32548 10412
rect 32508 10062 32536 10406
rect 32496 10056 32548 10062
rect 32496 9998 32548 10004
rect 32600 9636 32628 10662
rect 32508 9608 32628 9636
rect 32404 9512 32456 9518
rect 32404 9454 32456 9460
rect 32508 8956 32536 9608
rect 32692 9450 32720 13767
rect 32784 12850 32812 14010
rect 32772 12844 32824 12850
rect 32772 12786 32824 12792
rect 32772 10668 32824 10674
rect 32772 10610 32824 10616
rect 32680 9444 32732 9450
rect 32680 9386 32732 9392
rect 32680 9172 32732 9178
rect 32680 9114 32732 9120
rect 32588 8968 32640 8974
rect 32508 8928 32588 8956
rect 32508 7478 32536 8928
rect 32588 8910 32640 8916
rect 32588 7744 32640 7750
rect 32588 7686 32640 7692
rect 32496 7472 32548 7478
rect 32496 7414 32548 7420
rect 32496 7336 32548 7342
rect 32496 7278 32548 7284
rect 32508 6390 32536 7278
rect 32600 6730 32628 7686
rect 32588 6724 32640 6730
rect 32588 6666 32640 6672
rect 32496 6384 32548 6390
rect 32496 6326 32548 6332
rect 32600 6322 32628 6666
rect 32588 6316 32640 6322
rect 32588 6258 32640 6264
rect 32404 3936 32456 3942
rect 32404 3878 32456 3884
rect 32416 3126 32444 3878
rect 32404 3120 32456 3126
rect 32404 3062 32456 3068
rect 32324 2746 32536 2774
rect 32508 2514 32536 2746
rect 32692 2582 32720 9114
rect 32784 8906 32812 10610
rect 32876 9518 32904 15846
rect 32968 15434 32996 16050
rect 32956 15428 33008 15434
rect 32956 15370 33008 15376
rect 32968 14006 32996 15370
rect 32956 14000 33008 14006
rect 32956 13942 33008 13948
rect 33060 11218 33088 22918
rect 33140 22772 33192 22778
rect 33140 22714 33192 22720
rect 33152 22642 33180 22714
rect 33140 22636 33192 22642
rect 33140 22578 33192 22584
rect 33428 22030 33456 30534
rect 33520 30258 33548 31758
rect 33508 30252 33560 30258
rect 33508 30194 33560 30200
rect 33520 29170 33548 30194
rect 33600 30184 33652 30190
rect 33600 30126 33652 30132
rect 33612 29170 33640 30126
rect 33508 29164 33560 29170
rect 33508 29106 33560 29112
rect 33600 29164 33652 29170
rect 33600 29106 33652 29112
rect 33520 29073 33548 29106
rect 33506 29064 33562 29073
rect 33506 28999 33562 29008
rect 33508 24404 33560 24410
rect 33508 24346 33560 24352
rect 33416 22024 33468 22030
rect 33416 21966 33468 21972
rect 33416 21480 33468 21486
rect 33416 21422 33468 21428
rect 33232 20936 33284 20942
rect 33232 20878 33284 20884
rect 33244 20466 33272 20878
rect 33232 20460 33284 20466
rect 33232 20402 33284 20408
rect 33244 19854 33272 20402
rect 33324 20256 33376 20262
rect 33324 20198 33376 20204
rect 33232 19848 33284 19854
rect 33232 19790 33284 19796
rect 33140 19440 33192 19446
rect 33244 19394 33272 19790
rect 33336 19446 33364 20198
rect 33192 19388 33272 19394
rect 33140 19382 33272 19388
rect 33324 19440 33376 19446
rect 33324 19382 33376 19388
rect 33152 19366 33272 19382
rect 33140 18692 33192 18698
rect 33140 18634 33192 18640
rect 33152 18290 33180 18634
rect 33140 18284 33192 18290
rect 33140 18226 33192 18232
rect 33152 16998 33180 18226
rect 33140 16992 33192 16998
rect 33140 16934 33192 16940
rect 33152 16522 33180 16934
rect 33140 16516 33192 16522
rect 33140 16458 33192 16464
rect 33140 15360 33192 15366
rect 33140 15302 33192 15308
rect 33152 15026 33180 15302
rect 33140 15020 33192 15026
rect 33140 14962 33192 14968
rect 33152 14414 33180 14962
rect 33140 14408 33192 14414
rect 33140 14350 33192 14356
rect 33140 11280 33192 11286
rect 33140 11222 33192 11228
rect 33048 11212 33100 11218
rect 33048 11154 33100 11160
rect 33152 11150 33180 11222
rect 32956 11144 33008 11150
rect 33140 11144 33192 11150
rect 32956 11086 33008 11092
rect 33060 11092 33140 11098
rect 33060 11086 33192 11092
rect 32864 9512 32916 9518
rect 32864 9454 32916 9460
rect 32772 8900 32824 8906
rect 32772 8842 32824 8848
rect 32784 7546 32812 8842
rect 32968 7818 32996 11086
rect 33060 11070 33180 11086
rect 32956 7812 33008 7818
rect 32956 7754 33008 7760
rect 33060 7698 33088 11070
rect 33140 9512 33192 9518
rect 33138 9480 33140 9489
rect 33192 9480 33194 9489
rect 33138 9415 33194 9424
rect 33244 9382 33272 19366
rect 33428 18970 33456 21422
rect 33416 18964 33468 18970
rect 33416 18906 33468 18912
rect 33428 18290 33456 18906
rect 33416 18284 33468 18290
rect 33416 18226 33468 18232
rect 33414 14920 33470 14929
rect 33414 14855 33470 14864
rect 33428 12306 33456 14855
rect 33416 12300 33468 12306
rect 33416 12242 33468 12248
rect 33416 11076 33468 11082
rect 33416 11018 33468 11024
rect 33428 10674 33456 11018
rect 33416 10668 33468 10674
rect 33416 10610 33468 10616
rect 33428 10266 33456 10610
rect 33416 10260 33468 10266
rect 33416 10202 33468 10208
rect 33232 9376 33284 9382
rect 33232 9318 33284 9324
rect 33244 9042 33272 9318
rect 33140 9036 33192 9042
rect 33140 8978 33192 8984
rect 33232 9036 33284 9042
rect 33232 8978 33284 8984
rect 33152 8090 33180 8978
rect 33416 8968 33468 8974
rect 33416 8910 33468 8916
rect 33140 8084 33192 8090
rect 33140 8026 33192 8032
rect 33232 7880 33284 7886
rect 33232 7822 33284 7828
rect 32968 7670 33088 7698
rect 32968 7546 32996 7670
rect 32772 7540 32824 7546
rect 32772 7482 32824 7488
rect 32956 7540 33008 7546
rect 32956 7482 33008 7488
rect 33244 7342 33272 7822
rect 33428 7478 33456 8910
rect 33416 7472 33468 7478
rect 33416 7414 33468 7420
rect 33232 7336 33284 7342
rect 33232 7278 33284 7284
rect 33048 5636 33100 5642
rect 33048 5578 33100 5584
rect 32956 3936 33008 3942
rect 32956 3878 33008 3884
rect 32968 2990 32996 3878
rect 33060 3126 33088 5578
rect 33048 3120 33100 3126
rect 33520 3074 33548 24346
rect 33704 23254 33732 47058
rect 33784 40928 33836 40934
rect 33784 40870 33836 40876
rect 33796 40458 33824 40870
rect 33784 40452 33836 40458
rect 33784 40394 33836 40400
rect 33796 37074 33824 40394
rect 33968 39840 34020 39846
rect 33968 39782 34020 39788
rect 33876 39432 33928 39438
rect 33876 39374 33928 39380
rect 33888 38350 33916 39374
rect 33980 39370 34008 39782
rect 33968 39364 34020 39370
rect 33968 39306 34020 39312
rect 33876 38344 33928 38350
rect 33876 38286 33928 38292
rect 33888 37262 33916 38286
rect 33876 37256 33928 37262
rect 33876 37198 33928 37204
rect 33796 37046 33916 37074
rect 33888 33930 33916 37046
rect 33876 33924 33928 33930
rect 33876 33866 33928 33872
rect 33784 33856 33836 33862
rect 33784 33798 33836 33804
rect 33796 33658 33824 33798
rect 33784 33652 33836 33658
rect 33784 33594 33836 33600
rect 33796 29714 33824 33594
rect 33784 29708 33836 29714
rect 33784 29650 33836 29656
rect 33968 29708 34020 29714
rect 33968 29650 34020 29656
rect 33782 29200 33838 29209
rect 33782 29135 33784 29144
rect 33836 29135 33838 29144
rect 33784 29106 33836 29112
rect 33980 28626 34008 29650
rect 33968 28620 34020 28626
rect 33968 28562 34020 28568
rect 33784 28552 33836 28558
rect 33784 28494 33836 28500
rect 33796 28218 33824 28494
rect 33784 28212 33836 28218
rect 33784 28154 33836 28160
rect 33796 26314 33824 28154
rect 33968 26444 34020 26450
rect 33968 26386 34020 26392
rect 33784 26308 33836 26314
rect 33784 26250 33836 26256
rect 33980 25974 34008 26386
rect 33968 25968 34020 25974
rect 33968 25910 34020 25916
rect 33784 24948 33836 24954
rect 33784 24890 33836 24896
rect 33796 24206 33824 24890
rect 33784 24200 33836 24206
rect 33784 24142 33836 24148
rect 33966 23896 34022 23905
rect 33966 23831 34022 23840
rect 33784 23792 33836 23798
rect 33784 23734 33836 23740
rect 33796 23594 33824 23734
rect 33784 23588 33836 23594
rect 33784 23530 33836 23536
rect 33692 23248 33744 23254
rect 33692 23190 33744 23196
rect 33980 23186 34008 23831
rect 33968 23180 34020 23186
rect 33968 23122 34020 23128
rect 33600 22704 33652 22710
rect 33598 22672 33600 22681
rect 33652 22672 33654 22681
rect 33598 22607 33654 22616
rect 33600 22568 33652 22574
rect 33600 22510 33652 22516
rect 33612 21690 33640 22510
rect 33980 22030 34008 23122
rect 33968 22024 34020 22030
rect 33968 21966 34020 21972
rect 33600 21684 33652 21690
rect 33600 21626 33652 21632
rect 33876 21480 33928 21486
rect 33876 21422 33928 21428
rect 33692 20800 33744 20806
rect 33692 20742 33744 20748
rect 33704 20534 33732 20742
rect 33692 20528 33744 20534
rect 33692 20470 33744 20476
rect 33784 20392 33836 20398
rect 33784 20334 33836 20340
rect 33600 19304 33652 19310
rect 33600 19246 33652 19252
rect 33612 13734 33640 19246
rect 33692 18216 33744 18222
rect 33692 18158 33744 18164
rect 33704 17678 33732 18158
rect 33692 17672 33744 17678
rect 33692 17614 33744 17620
rect 33796 14414 33824 20334
rect 33888 20058 33916 21422
rect 34072 20398 34100 51326
rect 34150 51200 34206 51326
rect 34794 51200 34850 52000
rect 35438 51200 35494 52000
rect 36082 51200 36138 52000
rect 36726 51200 36782 52000
rect 37370 51354 37426 52000
rect 38014 51354 38070 52000
rect 37370 51326 37872 51354
rect 37370 51200 37426 51326
rect 34152 48544 34204 48550
rect 34152 48486 34204 48492
rect 34060 20392 34112 20398
rect 34060 20334 34112 20340
rect 33876 20052 33928 20058
rect 33876 19994 33928 20000
rect 34164 19310 34192 48486
rect 34808 47598 34836 51200
rect 34934 49532 35242 49552
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49456 35242 49476
rect 34888 49224 34940 49230
rect 34888 49166 34940 49172
rect 34900 48754 34928 49166
rect 34888 48748 34940 48754
rect 34888 48690 34940 48696
rect 36096 48686 36124 51200
rect 36084 48680 36136 48686
rect 36084 48622 36136 48628
rect 36176 48612 36228 48618
rect 36176 48554 36228 48560
rect 34934 48444 35242 48464
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48368 35242 48388
rect 35716 48136 35768 48142
rect 35438 48104 35494 48113
rect 35438 48039 35494 48048
rect 35714 48104 35716 48113
rect 35768 48104 35770 48113
rect 35714 48039 35770 48048
rect 34796 47592 34848 47598
rect 34796 47534 34848 47540
rect 34934 47356 35242 47376
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47280 35242 47300
rect 34934 46268 35242 46288
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46192 35242 46212
rect 34934 45180 35242 45200
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45104 35242 45124
rect 34934 44092 35242 44112
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44016 35242 44036
rect 34934 43004 35242 43024
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42928 35242 42948
rect 34934 41916 35242 41936
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41840 35242 41860
rect 34934 40828 35242 40848
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40752 35242 40772
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 34244 39364 34296 39370
rect 34244 39306 34296 39312
rect 34256 39030 34284 39306
rect 34334 39264 34390 39273
rect 34334 39199 34390 39208
rect 34348 39030 34376 39199
rect 34244 39024 34296 39030
rect 34244 38966 34296 38972
rect 34336 39024 34388 39030
rect 35452 39001 35480 48039
rect 36188 47802 36216 48554
rect 36740 48278 36768 51200
rect 37464 48544 37516 48550
rect 37464 48486 37516 48492
rect 36728 48272 36780 48278
rect 36728 48214 36780 48220
rect 37476 48210 37504 48486
rect 37464 48204 37516 48210
rect 37464 48146 37516 48152
rect 36176 47796 36228 47802
rect 36176 47738 36228 47744
rect 36084 47660 36136 47666
rect 36084 47602 36136 47608
rect 36096 47258 36124 47602
rect 36084 47252 36136 47258
rect 36084 47194 36136 47200
rect 37188 47252 37240 47258
rect 37188 47194 37240 47200
rect 37200 40050 37228 47194
rect 37844 45554 37872 51326
rect 38014 51326 38148 51354
rect 38014 51200 38070 51326
rect 38120 49230 38148 51326
rect 38658 51200 38714 52000
rect 39302 51354 39358 52000
rect 39132 51326 39358 51354
rect 38108 49224 38160 49230
rect 38108 49166 38160 49172
rect 38292 49088 38344 49094
rect 38292 49030 38344 49036
rect 37844 45526 38056 45554
rect 35900 40044 35952 40050
rect 35900 39986 35952 39992
rect 37188 40044 37240 40050
rect 37188 39986 37240 39992
rect 35912 39438 35940 39986
rect 35900 39432 35952 39438
rect 35900 39374 35952 39380
rect 34336 38966 34388 38972
rect 35438 38992 35494 39001
rect 34428 38956 34480 38962
rect 34480 38916 34560 38944
rect 35438 38927 35494 38936
rect 34428 38898 34480 38904
rect 34532 38758 34560 38916
rect 34428 38752 34480 38758
rect 34428 38694 34480 38700
rect 34520 38752 34572 38758
rect 34520 38694 34572 38700
rect 34440 38570 34468 38694
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 34440 38542 34560 38570
rect 34532 38214 34560 38542
rect 34520 38208 34572 38214
rect 34520 38150 34572 38156
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 34704 36372 34756 36378
rect 34704 36314 34756 36320
rect 34428 33992 34480 33998
rect 34428 33934 34480 33940
rect 34244 33448 34296 33454
rect 34244 33390 34296 33396
rect 34256 33114 34284 33390
rect 34440 33386 34468 33934
rect 34428 33380 34480 33386
rect 34428 33322 34480 33328
rect 34244 33108 34296 33114
rect 34244 33050 34296 33056
rect 34440 28558 34468 33322
rect 34612 30048 34664 30054
rect 34612 29990 34664 29996
rect 34624 29510 34652 29990
rect 34612 29504 34664 29510
rect 34612 29446 34664 29452
rect 34428 28552 34480 28558
rect 34428 28494 34480 28500
rect 34624 25430 34652 29446
rect 34716 26382 34744 36314
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 35348 26920 35400 26926
rect 35348 26862 35400 26868
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 34704 26376 34756 26382
rect 35256 26376 35308 26382
rect 34756 26336 34836 26364
rect 34704 26318 34756 26324
rect 34704 26240 34756 26246
rect 34704 26182 34756 26188
rect 34716 25974 34744 26182
rect 34704 25968 34756 25974
rect 34704 25910 34756 25916
rect 34704 25832 34756 25838
rect 34704 25774 34756 25780
rect 34612 25424 34664 25430
rect 34612 25366 34664 25372
rect 34716 25294 34744 25774
rect 34808 25294 34836 26336
rect 35360 26364 35388 26862
rect 35308 26336 35388 26364
rect 35256 26318 35308 26324
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 34888 25424 34940 25430
rect 34888 25366 34940 25372
rect 34704 25288 34756 25294
rect 34704 25230 34756 25236
rect 34796 25288 34848 25294
rect 34796 25230 34848 25236
rect 34612 25220 34664 25226
rect 34612 25162 34664 25168
rect 34520 25152 34572 25158
rect 34520 25094 34572 25100
rect 34244 24744 34296 24750
rect 34244 24686 34296 24692
rect 34256 24410 34284 24686
rect 34244 24404 34296 24410
rect 34244 24346 34296 24352
rect 34532 24138 34560 25094
rect 34520 24132 34572 24138
rect 34520 24074 34572 24080
rect 34624 23730 34652 25162
rect 34716 24750 34744 25230
rect 34900 25140 34928 25366
rect 35164 25288 35216 25294
rect 35360 25276 35388 26336
rect 35216 25248 35388 25276
rect 35164 25230 35216 25236
rect 34808 25112 34928 25140
rect 34704 24744 34756 24750
rect 34704 24686 34756 24692
rect 34520 23724 34572 23730
rect 34520 23666 34572 23672
rect 34612 23724 34664 23730
rect 34612 23666 34664 23672
rect 34532 23633 34560 23666
rect 34518 23624 34574 23633
rect 34518 23559 34574 23568
rect 34716 23186 34744 24686
rect 34808 23714 34836 25112
rect 35176 24954 35204 25230
rect 35164 24948 35216 24954
rect 35164 24890 35216 24896
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 34888 24132 34940 24138
rect 34888 24074 34940 24080
rect 34900 24041 34928 24074
rect 34886 24032 34942 24041
rect 34886 23967 34942 23976
rect 34978 23896 35034 23905
rect 34978 23831 35034 23840
rect 34992 23730 35020 23831
rect 35348 23792 35400 23798
rect 35348 23734 35400 23740
rect 34949 23724 35020 23730
rect 34796 23708 34848 23714
rect 35001 23684 35020 23724
rect 34949 23666 35001 23672
rect 34796 23650 34848 23656
rect 35360 23594 35388 23734
rect 35348 23588 35400 23594
rect 35348 23530 35400 23536
rect 34796 23520 34848 23526
rect 34796 23462 34848 23468
rect 34704 23180 34756 23186
rect 34704 23122 34756 23128
rect 34520 23044 34572 23050
rect 34520 22986 34572 22992
rect 34532 21962 34560 22986
rect 34612 22432 34664 22438
rect 34612 22374 34664 22380
rect 34624 22030 34652 22374
rect 34612 22024 34664 22030
rect 34612 21966 34664 21972
rect 34704 22024 34756 22030
rect 34704 21966 34756 21972
rect 34520 21956 34572 21962
rect 34520 21898 34572 21904
rect 34152 19304 34204 19310
rect 34152 19246 34204 19252
rect 34716 18834 34744 21966
rect 34808 21962 34836 23462
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 35452 22094 35480 38927
rect 35636 38814 35848 38842
rect 35636 38214 35664 38814
rect 35820 38758 35848 38814
rect 35716 38752 35768 38758
rect 35716 38694 35768 38700
rect 35808 38752 35860 38758
rect 35808 38694 35860 38700
rect 35624 38208 35676 38214
rect 35624 38150 35676 38156
rect 35532 37188 35584 37194
rect 35532 37130 35584 37136
rect 35544 36854 35572 37130
rect 35532 36848 35584 36854
rect 35532 36790 35584 36796
rect 35636 36786 35664 38150
rect 35728 37210 35756 38694
rect 35912 38350 35940 39374
rect 35992 39364 36044 39370
rect 35992 39306 36044 39312
rect 36004 39098 36032 39306
rect 35992 39092 36044 39098
rect 35992 39034 36044 39040
rect 36084 39092 36136 39098
rect 36084 39034 36136 39040
rect 36096 38876 36124 39034
rect 36176 39024 36228 39030
rect 36228 38984 36492 39012
rect 36176 38966 36228 38972
rect 36464 38944 36492 38984
rect 36636 38956 36688 38962
rect 36464 38916 36636 38944
rect 36636 38898 36688 38904
rect 36096 38848 36216 38876
rect 35900 38344 35952 38350
rect 35900 38286 35952 38292
rect 35808 38208 35860 38214
rect 35808 38150 35860 38156
rect 35820 37738 35848 38150
rect 35808 37732 35860 37738
rect 35808 37674 35860 37680
rect 35728 37182 35848 37210
rect 35716 37120 35768 37126
rect 35716 37062 35768 37068
rect 35624 36780 35676 36786
rect 35624 36722 35676 36728
rect 35728 36174 35756 37062
rect 35716 36168 35768 36174
rect 35716 36110 35768 36116
rect 35532 29028 35584 29034
rect 35532 28970 35584 28976
rect 35544 28422 35572 28970
rect 35532 28416 35584 28422
rect 35532 28358 35584 28364
rect 35544 25362 35572 28358
rect 35716 26988 35768 26994
rect 35716 26930 35768 26936
rect 35624 26784 35676 26790
rect 35624 26726 35676 26732
rect 35636 26382 35664 26726
rect 35624 26376 35676 26382
rect 35624 26318 35676 26324
rect 35532 25356 35584 25362
rect 35532 25298 35584 25304
rect 35624 25152 35676 25158
rect 35624 25094 35676 25100
rect 35636 24886 35664 25094
rect 35624 24880 35676 24886
rect 35624 24822 35676 24828
rect 35532 24404 35584 24410
rect 35532 24346 35584 24352
rect 35544 23526 35572 24346
rect 35728 24138 35756 26930
rect 35716 24132 35768 24138
rect 35716 24074 35768 24080
rect 35624 23724 35676 23730
rect 35624 23666 35676 23672
rect 35532 23520 35584 23526
rect 35532 23462 35584 23468
rect 35636 22506 35664 23666
rect 35728 22642 35756 24074
rect 35716 22636 35768 22642
rect 35716 22578 35768 22584
rect 35624 22500 35676 22506
rect 35624 22442 35676 22448
rect 35452 22066 35664 22094
rect 34796 21956 34848 21962
rect 34796 21898 34848 21904
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 35636 19718 35664 22066
rect 35624 19712 35676 19718
rect 35624 19654 35676 19660
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 34704 18828 34756 18834
rect 34704 18770 34756 18776
rect 34520 18624 34572 18630
rect 34520 18566 34572 18572
rect 34428 17808 34480 17814
rect 34428 17750 34480 17756
rect 33968 17604 34020 17610
rect 33968 17546 34020 17552
rect 33980 17338 34008 17546
rect 33968 17332 34020 17338
rect 33968 17274 34020 17280
rect 34440 17134 34468 17750
rect 34532 17746 34560 18566
rect 34612 18080 34664 18086
rect 34612 18022 34664 18028
rect 34520 17740 34572 17746
rect 34520 17682 34572 17688
rect 34624 17678 34652 18022
rect 34612 17672 34664 17678
rect 34612 17614 34664 17620
rect 34520 17196 34572 17202
rect 34520 17138 34572 17144
rect 34428 17128 34480 17134
rect 34532 17105 34560 17138
rect 34428 17070 34480 17076
rect 34518 17096 34574 17105
rect 34518 17031 34574 17040
rect 34520 15496 34572 15502
rect 34520 15438 34572 15444
rect 33784 14408 33836 14414
rect 33784 14350 33836 14356
rect 33796 14074 33824 14350
rect 33784 14068 33836 14074
rect 33784 14010 33836 14016
rect 33600 13728 33652 13734
rect 33600 13670 33652 13676
rect 33612 13530 33640 13670
rect 33600 13524 33652 13530
rect 33600 13466 33652 13472
rect 34532 13258 34560 15438
rect 34624 14958 34652 17614
rect 34716 16658 34744 18770
rect 35624 18760 35676 18766
rect 35624 18702 35676 18708
rect 35636 18426 35664 18702
rect 35624 18420 35676 18426
rect 35624 18362 35676 18368
rect 34796 18284 34848 18290
rect 34796 18226 34848 18232
rect 34808 17882 34836 18226
rect 35348 18080 35400 18086
rect 35348 18022 35400 18028
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 34796 17876 34848 17882
rect 34796 17818 34848 17824
rect 35360 17338 35388 18022
rect 35348 17332 35400 17338
rect 35348 17274 35400 17280
rect 35254 17232 35310 17241
rect 35254 17167 35256 17176
rect 35308 17167 35310 17176
rect 35624 17196 35676 17202
rect 35256 17138 35308 17144
rect 35624 17138 35676 17144
rect 35636 17105 35664 17138
rect 35622 17096 35678 17105
rect 35622 17031 35678 17040
rect 34796 16992 34848 16998
rect 34796 16934 34848 16940
rect 34704 16652 34756 16658
rect 34704 16594 34756 16600
rect 34808 16590 34836 16934
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 34796 16584 34848 16590
rect 34796 16526 34848 16532
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 35624 15360 35676 15366
rect 35624 15302 35676 15308
rect 35440 15020 35492 15026
rect 35440 14962 35492 14968
rect 34612 14952 34664 14958
rect 34612 14894 34664 14900
rect 34624 14006 34652 14894
rect 34794 14784 34850 14793
rect 34794 14719 34850 14728
rect 34704 14544 34756 14550
rect 34704 14486 34756 14492
rect 34612 14000 34664 14006
rect 34612 13942 34664 13948
rect 34716 13734 34744 14486
rect 34808 14482 34836 14719
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 35452 14618 35480 14962
rect 35440 14612 35492 14618
rect 35440 14554 35492 14560
rect 35532 14612 35584 14618
rect 35532 14554 35584 14560
rect 35544 14521 35572 14554
rect 35530 14512 35586 14521
rect 34796 14476 34848 14482
rect 35530 14447 35586 14456
rect 34796 14418 34848 14424
rect 35544 14414 35572 14447
rect 35636 14414 35664 15302
rect 35348 14408 35400 14414
rect 35346 14376 35348 14385
rect 35532 14408 35584 14414
rect 35400 14376 35402 14385
rect 35532 14350 35584 14356
rect 35624 14408 35676 14414
rect 35624 14350 35676 14356
rect 35346 14311 35402 14320
rect 34796 14000 34848 14006
rect 34796 13942 34848 13948
rect 34704 13728 34756 13734
rect 34704 13670 34756 13676
rect 34520 13252 34572 13258
rect 34520 13194 34572 13200
rect 34532 12238 34560 13194
rect 34808 12850 34836 13942
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 35544 13462 35572 14350
rect 35716 14340 35768 14346
rect 35716 14282 35768 14288
rect 35532 13456 35584 13462
rect 35532 13398 35584 13404
rect 35728 13326 35756 14282
rect 35348 13320 35400 13326
rect 35348 13262 35400 13268
rect 35532 13320 35584 13326
rect 35532 13262 35584 13268
rect 35716 13320 35768 13326
rect 35716 13262 35768 13268
rect 35072 13184 35124 13190
rect 35072 13126 35124 13132
rect 35084 12918 35112 13126
rect 35072 12912 35124 12918
rect 35072 12854 35124 12860
rect 34796 12844 34848 12850
rect 34796 12786 34848 12792
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 34520 12232 34572 12238
rect 34520 12174 34572 12180
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 33784 11008 33836 11014
rect 33784 10950 33836 10956
rect 33796 10606 33824 10950
rect 33784 10600 33836 10606
rect 33784 10542 33836 10548
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 33784 8288 33836 8294
rect 33784 8230 33836 8236
rect 33796 7886 33824 8230
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 33784 7880 33836 7886
rect 33784 7822 33836 7828
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 35360 4078 35388 13262
rect 35544 12442 35572 13262
rect 35532 12436 35584 12442
rect 35532 12378 35584 12384
rect 35820 8362 35848 37182
rect 35912 36378 35940 38286
rect 36084 38276 36136 38282
rect 36084 38218 36136 38224
rect 36096 38010 36124 38218
rect 36084 38004 36136 38010
rect 36084 37946 36136 37952
rect 36188 37806 36216 38848
rect 36648 37856 36676 38898
rect 36728 37868 36780 37874
rect 36648 37828 36728 37856
rect 36176 37800 36228 37806
rect 36176 37742 36228 37748
rect 36188 37398 36216 37742
rect 36176 37392 36228 37398
rect 36176 37334 36228 37340
rect 36648 37262 36676 37828
rect 36728 37810 36780 37816
rect 36084 37256 36136 37262
rect 36636 37256 36688 37262
rect 36136 37204 36400 37210
rect 36084 37198 36400 37204
rect 36636 37198 36688 37204
rect 36096 37194 36400 37198
rect 36096 37188 36412 37194
rect 36096 37182 36360 37188
rect 36360 37130 36412 37136
rect 35992 37120 36044 37126
rect 35992 37062 36044 37068
rect 36004 36922 36032 37062
rect 35992 36916 36044 36922
rect 35992 36858 36044 36864
rect 37004 36848 37056 36854
rect 37004 36790 37056 36796
rect 37016 36378 37044 36790
rect 35900 36372 35952 36378
rect 35900 36314 35952 36320
rect 37004 36372 37056 36378
rect 37004 36314 37056 36320
rect 36452 29572 36504 29578
rect 36452 29514 36504 29520
rect 36464 29306 36492 29514
rect 36452 29300 36504 29306
rect 36452 29242 36504 29248
rect 36360 29164 36412 29170
rect 36360 29106 36412 29112
rect 35900 25288 35952 25294
rect 35900 25230 35952 25236
rect 35912 24410 35940 25230
rect 35900 24404 35952 24410
rect 35900 24346 35952 24352
rect 35992 24132 36044 24138
rect 35992 24074 36044 24080
rect 36004 23730 36032 24074
rect 35992 23724 36044 23730
rect 35992 23666 36044 23672
rect 36082 23624 36138 23633
rect 36082 23559 36084 23568
rect 36136 23559 36138 23568
rect 36084 23530 36136 23536
rect 35900 22976 35952 22982
rect 35900 22918 35952 22924
rect 35912 22642 35940 22918
rect 36372 22778 36400 29106
rect 36452 27056 36504 27062
rect 36452 26998 36504 27004
rect 36464 25770 36492 26998
rect 36544 26240 36596 26246
rect 36544 26182 36596 26188
rect 36556 26042 36584 26182
rect 36544 26036 36596 26042
rect 36544 25978 36596 25984
rect 36452 25764 36504 25770
rect 36452 25706 36504 25712
rect 36464 25362 36492 25706
rect 36452 25356 36504 25362
rect 36452 25298 36504 25304
rect 36728 24608 36780 24614
rect 36728 24550 36780 24556
rect 36452 24336 36504 24342
rect 36452 24278 36504 24284
rect 36464 23769 36492 24278
rect 36740 24206 36768 24550
rect 36728 24200 36780 24206
rect 36728 24142 36780 24148
rect 36450 23760 36506 23769
rect 36740 23730 36768 24142
rect 36450 23695 36506 23704
rect 36728 23724 36780 23730
rect 36728 23666 36780 23672
rect 36360 22772 36412 22778
rect 36360 22714 36412 22720
rect 35900 22636 35952 22642
rect 35900 22578 35952 22584
rect 36084 22636 36136 22642
rect 36084 22578 36136 22584
rect 36096 21010 36124 22578
rect 36268 22500 36320 22506
rect 36268 22442 36320 22448
rect 36280 22166 36308 22442
rect 36268 22160 36320 22166
rect 36268 22102 36320 22108
rect 36280 22030 36308 22102
rect 36268 22024 36320 22030
rect 36268 21966 36320 21972
rect 36176 21888 36228 21894
rect 36176 21830 36228 21836
rect 36188 21146 36216 21830
rect 36268 21684 36320 21690
rect 36268 21626 36320 21632
rect 36176 21140 36228 21146
rect 36176 21082 36228 21088
rect 36280 21010 36308 21626
rect 36372 21554 36400 22714
rect 36360 21548 36412 21554
rect 36360 21490 36412 21496
rect 36372 21010 36400 21490
rect 36084 21004 36136 21010
rect 36084 20946 36136 20952
rect 36268 21004 36320 21010
rect 36268 20946 36320 20952
rect 36360 21004 36412 21010
rect 36360 20946 36412 20952
rect 36544 20324 36596 20330
rect 36544 20266 36596 20272
rect 36556 19990 36584 20266
rect 36544 19984 36596 19990
rect 36544 19926 36596 19932
rect 36636 19372 36688 19378
rect 36636 19314 36688 19320
rect 36544 19168 36596 19174
rect 36544 19110 36596 19116
rect 36556 18834 36584 19110
rect 36544 18828 36596 18834
rect 36544 18770 36596 18776
rect 36084 18692 36136 18698
rect 36084 18634 36136 18640
rect 36096 18290 36124 18634
rect 36648 18358 36676 19314
rect 36636 18352 36688 18358
rect 36636 18294 36688 18300
rect 36084 18284 36136 18290
rect 36084 18226 36136 18232
rect 36176 18284 36228 18290
rect 36176 18226 36228 18232
rect 35900 17740 35952 17746
rect 35900 17682 35952 17688
rect 35912 16794 35940 17682
rect 36096 17202 36124 18226
rect 36188 17882 36216 18226
rect 36176 17876 36228 17882
rect 36176 17818 36228 17824
rect 36648 17678 36676 18294
rect 36636 17672 36688 17678
rect 36636 17614 36688 17620
rect 36648 17202 36676 17614
rect 36084 17196 36136 17202
rect 36084 17138 36136 17144
rect 36268 17196 36320 17202
rect 36268 17138 36320 17144
rect 36636 17196 36688 17202
rect 36636 17138 36688 17144
rect 36280 16794 36308 17138
rect 35900 16788 35952 16794
rect 35900 16730 35952 16736
rect 36268 16788 36320 16794
rect 36268 16730 36320 16736
rect 36544 15428 36596 15434
rect 36544 15370 36596 15376
rect 36556 14822 36584 15370
rect 36544 14816 36596 14822
rect 36544 14758 36596 14764
rect 36268 14272 36320 14278
rect 36268 14214 36320 14220
rect 36280 14006 36308 14214
rect 36268 14000 36320 14006
rect 36268 13942 36320 13948
rect 36360 13728 36412 13734
rect 36360 13670 36412 13676
rect 36372 13326 36400 13670
rect 36360 13320 36412 13326
rect 36360 13262 36412 13268
rect 36360 12640 36412 12646
rect 36360 12582 36412 12588
rect 36372 12238 36400 12582
rect 36360 12232 36412 12238
rect 36360 12174 36412 12180
rect 36556 9654 36584 14758
rect 36728 14408 36780 14414
rect 36728 14350 36780 14356
rect 36912 14408 36964 14414
rect 36912 14350 36964 14356
rect 37002 14376 37058 14385
rect 36740 13530 36768 14350
rect 36924 14278 36952 14350
rect 37002 14311 37058 14320
rect 37016 14278 37044 14311
rect 36912 14272 36964 14278
rect 36912 14214 36964 14220
rect 37004 14272 37056 14278
rect 37004 14214 37056 14220
rect 36728 13524 36780 13530
rect 36728 13466 36780 13472
rect 36544 9648 36596 9654
rect 36544 9590 36596 9596
rect 35808 8356 35860 8362
rect 35808 8298 35860 8304
rect 36176 4140 36228 4146
rect 36176 4082 36228 4088
rect 35348 4072 35400 4078
rect 35348 4014 35400 4020
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 36188 3194 36216 4082
rect 36452 3936 36504 3942
rect 36452 3878 36504 3884
rect 36464 3602 36492 3878
rect 37200 3602 37228 39986
rect 37464 39296 37516 39302
rect 37464 39238 37516 39244
rect 37476 39137 37504 39238
rect 37462 39128 37518 39137
rect 37462 39063 37518 39072
rect 37476 39030 37504 39063
rect 37464 39024 37516 39030
rect 37370 38992 37426 39001
rect 37280 38956 37332 38962
rect 37464 38966 37516 38972
rect 37370 38927 37372 38936
rect 37280 38898 37332 38904
rect 37424 38927 37426 38936
rect 37372 38898 37424 38904
rect 37292 38758 37320 38898
rect 37280 38752 37332 38758
rect 37280 38694 37332 38700
rect 38028 29714 38056 45526
rect 38016 29708 38068 29714
rect 38016 29650 38068 29656
rect 37280 26580 37332 26586
rect 37280 26522 37332 26528
rect 37292 25906 37320 26522
rect 37372 26308 37424 26314
rect 37372 26250 37424 26256
rect 37384 26042 37412 26250
rect 37372 26036 37424 26042
rect 37372 25978 37424 25984
rect 37280 25900 37332 25906
rect 37280 25842 37332 25848
rect 37292 25294 37320 25842
rect 37372 25764 37424 25770
rect 37372 25706 37424 25712
rect 37280 25288 37332 25294
rect 37280 25230 37332 25236
rect 37292 24818 37320 25230
rect 37280 24812 37332 24818
rect 37280 24754 37332 24760
rect 37384 22094 37412 25706
rect 37648 24608 37700 24614
rect 37648 24550 37700 24556
rect 38200 24608 38252 24614
rect 38200 24550 38252 24556
rect 37660 24274 37688 24550
rect 37648 24268 37700 24274
rect 37648 24210 37700 24216
rect 38212 23662 38240 24550
rect 38200 23656 38252 23662
rect 38200 23598 38252 23604
rect 38304 23118 38332 49030
rect 38672 48226 38700 51200
rect 38752 48816 38804 48822
rect 38752 48758 38804 48764
rect 38764 48346 38792 48758
rect 38752 48340 38804 48346
rect 38752 48282 38804 48288
rect 38672 48198 39068 48226
rect 38660 48136 38712 48142
rect 38660 48078 38712 48084
rect 38672 44742 38700 48078
rect 38660 44736 38712 44742
rect 38660 44678 38712 44684
rect 38292 23112 38344 23118
rect 38292 23054 38344 23060
rect 37292 22066 37412 22094
rect 37292 21554 37320 22066
rect 37372 21956 37424 21962
rect 37372 21898 37424 21904
rect 37384 21690 37412 21898
rect 37372 21684 37424 21690
rect 37372 21626 37424 21632
rect 37280 21548 37332 21554
rect 37280 21490 37332 21496
rect 37292 4282 37320 21490
rect 37832 21004 37884 21010
rect 37832 20946 37884 20952
rect 37464 20800 37516 20806
rect 37464 20742 37516 20748
rect 37476 20534 37504 20742
rect 37464 20528 37516 20534
rect 37464 20470 37516 20476
rect 37464 19168 37516 19174
rect 37464 19110 37516 19116
rect 37476 18358 37504 19110
rect 37464 18352 37516 18358
rect 37464 18294 37516 18300
rect 37372 16992 37424 16998
rect 37372 16934 37424 16940
rect 37384 16522 37412 16934
rect 37372 16516 37424 16522
rect 37372 16458 37424 16464
rect 37280 4276 37332 4282
rect 37280 4218 37332 4224
rect 37740 4276 37792 4282
rect 37740 4218 37792 4224
rect 36452 3596 36504 3602
rect 36452 3538 36504 3544
rect 36728 3596 36780 3602
rect 36728 3538 36780 3544
rect 37188 3596 37240 3602
rect 37188 3538 37240 3544
rect 36268 3528 36320 3534
rect 36268 3470 36320 3476
rect 36176 3188 36228 3194
rect 36176 3130 36228 3136
rect 33048 3062 33100 3068
rect 33428 3046 33548 3074
rect 36280 3058 36308 3470
rect 36268 3052 36320 3058
rect 32956 2984 33008 2990
rect 32956 2926 33008 2932
rect 33428 2854 33456 3046
rect 36268 2994 36320 3000
rect 33508 2916 33560 2922
rect 33508 2858 33560 2864
rect 33416 2848 33468 2854
rect 33416 2790 33468 2796
rect 32680 2576 32732 2582
rect 32680 2518 32732 2524
rect 32496 2508 32548 2514
rect 32496 2450 32548 2456
rect 32864 2440 32916 2446
rect 32864 2382 32916 2388
rect 32876 800 32904 2382
rect 33520 800 33548 2858
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 34152 2372 34204 2378
rect 34152 2314 34204 2320
rect 34796 2372 34848 2378
rect 34796 2314 34848 2320
rect 36084 2372 36136 2378
rect 36084 2314 36136 2320
rect 34164 800 34192 2314
rect 34808 800 34836 2314
rect 36096 800 36124 2314
rect 36740 800 36768 3538
rect 37752 2990 37780 4218
rect 37844 4146 37872 20946
rect 37924 20868 37976 20874
rect 37924 20810 37976 20816
rect 37832 4140 37884 4146
rect 37832 4082 37884 4088
rect 37740 2984 37792 2990
rect 37740 2926 37792 2932
rect 37936 898 37964 20810
rect 39040 20534 39068 48198
rect 39028 20528 39080 20534
rect 39028 20470 39080 20476
rect 39132 17746 39160 51326
rect 39302 51200 39358 51326
rect 39946 51200 40002 52000
rect 40590 51200 40646 52000
rect 41234 51200 41290 52000
rect 41878 51200 41934 52000
rect 42522 51200 42578 52000
rect 43166 51200 43222 52000
rect 43810 51354 43866 52000
rect 43810 51326 43944 51354
rect 43810 51200 43866 51326
rect 39960 49450 39988 51200
rect 39960 49422 40080 49450
rect 40052 49366 40080 49422
rect 40040 49360 40092 49366
rect 40040 49302 40092 49308
rect 40604 49298 40632 51200
rect 40592 49292 40644 49298
rect 40592 49234 40644 49240
rect 39764 49224 39816 49230
rect 39764 49166 39816 49172
rect 39212 49088 39264 49094
rect 39212 49030 39264 49036
rect 39224 32298 39252 49030
rect 39776 47666 39804 49166
rect 40040 49156 40092 49162
rect 40040 49098 40092 49104
rect 40052 48278 40080 49098
rect 41248 48498 41276 51200
rect 41420 50244 41472 50250
rect 41420 50186 41472 50192
rect 41432 48822 41460 50186
rect 41892 48822 41920 51200
rect 41972 49224 42024 49230
rect 41972 49166 42024 49172
rect 41420 48816 41472 48822
rect 41420 48758 41472 48764
rect 41880 48816 41932 48822
rect 41880 48758 41932 48764
rect 40144 48470 41276 48498
rect 41604 48544 41656 48550
rect 41604 48486 41656 48492
rect 40040 48272 40092 48278
rect 40040 48214 40092 48220
rect 39856 48136 39908 48142
rect 39856 48078 39908 48084
rect 39764 47660 39816 47666
rect 39764 47602 39816 47608
rect 39868 34678 39896 48078
rect 39856 34672 39908 34678
rect 39856 34614 39908 34620
rect 39212 32292 39264 32298
rect 39212 32234 39264 32240
rect 39948 25152 40000 25158
rect 39948 25094 40000 25100
rect 39304 24132 39356 24138
rect 39304 24074 39356 24080
rect 39120 17740 39172 17746
rect 39120 17682 39172 17688
rect 38568 16652 38620 16658
rect 38568 16594 38620 16600
rect 38580 5370 38608 16594
rect 39316 9178 39344 24074
rect 39960 21350 39988 25094
rect 39948 21344 40000 21350
rect 39948 21286 40000 21292
rect 40144 18358 40172 48470
rect 41052 48136 41104 48142
rect 41052 48078 41104 48084
rect 40408 48068 40460 48074
rect 40408 48010 40460 48016
rect 40420 47802 40448 48010
rect 40408 47796 40460 47802
rect 40408 47738 40460 47744
rect 41064 47666 41092 48078
rect 40316 47660 40368 47666
rect 40316 47602 40368 47608
rect 41052 47660 41104 47666
rect 41052 47602 41104 47608
rect 40328 43246 40356 47602
rect 40316 43240 40368 43246
rect 40316 43182 40368 43188
rect 40684 37324 40736 37330
rect 40684 37266 40736 37272
rect 40132 18352 40184 18358
rect 40132 18294 40184 18300
rect 40696 10674 40724 37266
rect 40776 21956 40828 21962
rect 40776 21898 40828 21904
rect 40788 12442 40816 21898
rect 41616 20602 41644 48486
rect 41984 47666 42012 49166
rect 42536 48210 42564 51200
rect 43180 48686 43208 51200
rect 43720 49156 43772 49162
rect 43720 49098 43772 49104
rect 42800 48680 42852 48686
rect 42800 48622 42852 48628
rect 43168 48680 43220 48686
rect 43168 48622 43220 48628
rect 42524 48204 42576 48210
rect 42524 48146 42576 48152
rect 42812 47802 42840 48622
rect 42984 48612 43036 48618
rect 42984 48554 43036 48560
rect 42800 47796 42852 47802
rect 42800 47738 42852 47744
rect 41972 47660 42024 47666
rect 41972 47602 42024 47608
rect 42996 47258 43024 48554
rect 43536 47660 43588 47666
rect 43536 47602 43588 47608
rect 42984 47252 43036 47258
rect 42984 47194 43036 47200
rect 42800 37256 42852 37262
rect 42800 37198 42852 37204
rect 42812 33454 42840 37198
rect 42800 33448 42852 33454
rect 42800 33390 42852 33396
rect 43444 23656 43496 23662
rect 43444 23598 43496 23604
rect 42064 22568 42116 22574
rect 42064 22510 42116 22516
rect 41604 20596 41656 20602
rect 41604 20538 41656 20544
rect 40776 12436 40828 12442
rect 40776 12378 40828 12384
rect 40684 10668 40736 10674
rect 40684 10610 40736 10616
rect 39304 9172 39356 9178
rect 39304 9114 39356 9120
rect 38568 5364 38620 5370
rect 38568 5306 38620 5312
rect 40224 4480 40276 4486
rect 40224 4422 40276 4428
rect 40500 4480 40552 4486
rect 40500 4422 40552 4428
rect 38660 4072 38712 4078
rect 38660 4014 38712 4020
rect 38016 3936 38068 3942
rect 38016 3878 38068 3884
rect 37384 870 37504 898
rect 37384 800 37412 870
rect 9140 734 9444 762
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 23846 0 23902 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 25778 0 25834 800
rect 26422 0 26478 800
rect 27066 0 27122 800
rect 27710 0 27766 800
rect 28354 0 28410 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30286 0 30342 800
rect 30930 0 30986 800
rect 31574 0 31630 800
rect 32218 0 32274 800
rect 32862 0 32918 800
rect 33506 0 33562 800
rect 34150 0 34206 800
rect 34794 0 34850 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 36726 0 36782 800
rect 37370 0 37426 800
rect 37476 762 37504 870
rect 37752 870 37964 898
rect 37752 762 37780 870
rect 38028 800 38056 3878
rect 38672 3738 38700 4014
rect 38660 3732 38712 3738
rect 38660 3674 38712 3680
rect 40040 3392 40092 3398
rect 40040 3334 40092 3340
rect 39580 2848 39632 2854
rect 39580 2790 39632 2796
rect 39592 2514 39620 2790
rect 39948 2576 40000 2582
rect 39948 2518 40000 2524
rect 39580 2508 39632 2514
rect 39580 2450 39632 2456
rect 38660 2440 38712 2446
rect 38660 2382 38712 2388
rect 38752 2440 38804 2446
rect 38752 2382 38804 2388
rect 38672 800 38700 2382
rect 38764 1970 38792 2382
rect 38752 1964 38804 1970
rect 38752 1906 38804 1912
rect 39960 800 39988 2518
rect 40052 2514 40080 3334
rect 40236 3126 40264 4422
rect 40408 3188 40460 3194
rect 40408 3130 40460 3136
rect 40224 3120 40276 3126
rect 40224 3062 40276 3068
rect 40420 2922 40448 3130
rect 40512 2990 40540 4422
rect 41604 3936 41656 3942
rect 41604 3878 41656 3884
rect 41616 3602 41644 3878
rect 42076 3602 42104 22510
rect 42432 3936 42484 3942
rect 42432 3878 42484 3884
rect 41604 3596 41656 3602
rect 41604 3538 41656 3544
rect 41880 3596 41932 3602
rect 41880 3538 41932 3544
rect 42064 3596 42116 3602
rect 42064 3538 42116 3544
rect 40500 2984 40552 2990
rect 40500 2926 40552 2932
rect 41236 2984 41288 2990
rect 41236 2926 41288 2932
rect 40408 2916 40460 2922
rect 40408 2858 40460 2864
rect 40040 2508 40092 2514
rect 40040 2450 40092 2456
rect 41248 800 41276 2926
rect 41892 800 41920 3538
rect 42444 2514 42472 3878
rect 43456 3738 43484 23598
rect 43548 15026 43576 47602
rect 43732 46714 43760 49098
rect 43916 48142 43944 51326
rect 44454 51200 44510 52000
rect 45098 51200 45154 52000
rect 45742 51200 45798 52000
rect 46386 51200 46442 52000
rect 46662 51776 46718 51785
rect 46662 51711 46718 51720
rect 44088 49224 44140 49230
rect 44088 49166 44140 49172
rect 43904 48136 43956 48142
rect 43904 48078 43956 48084
rect 43812 48068 43864 48074
rect 43812 48010 43864 48016
rect 43824 47258 43852 48010
rect 43996 48000 44048 48006
rect 43996 47942 44048 47948
rect 43812 47252 43864 47258
rect 43812 47194 43864 47200
rect 43720 46708 43772 46714
rect 43720 46650 43772 46656
rect 43536 15020 43588 15026
rect 43536 14962 43588 14968
rect 44008 14278 44036 47942
rect 44100 46578 44128 49166
rect 44468 48142 44496 51200
rect 45112 49450 45140 51200
rect 45020 49422 45140 49450
rect 44916 48680 44968 48686
rect 44916 48622 44968 48628
rect 44456 48136 44508 48142
rect 44456 48078 44508 48084
rect 44180 47592 44232 47598
rect 44180 47534 44232 47540
rect 44364 47592 44416 47598
rect 44364 47534 44416 47540
rect 44088 46572 44140 46578
rect 44088 46514 44140 46520
rect 44192 46170 44220 47534
rect 44376 47258 44404 47534
rect 44364 47252 44416 47258
rect 44364 47194 44416 47200
rect 44548 46980 44600 46986
rect 44548 46922 44600 46928
rect 44560 46578 44588 46922
rect 44548 46572 44600 46578
rect 44548 46514 44600 46520
rect 44928 46170 44956 48622
rect 45020 47598 45048 49422
rect 45376 49156 45428 49162
rect 45376 49098 45428 49104
rect 45100 48680 45152 48686
rect 45100 48622 45152 48628
rect 45008 47592 45060 47598
rect 45008 47534 45060 47540
rect 45112 47258 45140 48622
rect 45192 48000 45244 48006
rect 45192 47942 45244 47948
rect 45100 47252 45152 47258
rect 45100 47194 45152 47200
rect 45204 46730 45232 47942
rect 45388 47802 45416 49098
rect 45756 48686 45784 51200
rect 46676 49298 46704 51711
rect 47030 51200 47086 52000
rect 47674 51354 47730 52000
rect 47674 51326 47808 51354
rect 47674 51200 47730 51326
rect 46754 51096 46810 51105
rect 46754 51031 46810 51040
rect 46768 49774 46796 51031
rect 46846 50416 46902 50425
rect 46846 50351 46902 50360
rect 46860 50250 46888 50351
rect 46848 50244 46900 50250
rect 46848 50186 46900 50192
rect 46756 49768 46808 49774
rect 46756 49710 46808 49716
rect 46846 49736 46902 49745
rect 46846 49671 46902 49680
rect 46860 49298 46888 49671
rect 46664 49292 46716 49298
rect 46664 49234 46716 49240
rect 46848 49292 46900 49298
rect 46848 49234 46900 49240
rect 47780 48822 47808 51326
rect 48318 51200 48374 52000
rect 48962 51200 49018 52000
rect 49606 51200 49662 52000
rect 47952 49088 48004 49094
rect 47858 49056 47914 49065
rect 47952 49030 48004 49036
rect 47858 48991 47914 49000
rect 47768 48816 47820 48822
rect 47768 48758 47820 48764
rect 45744 48680 45796 48686
rect 45744 48622 45796 48628
rect 46662 48376 46718 48385
rect 46662 48311 46718 48320
rect 45376 47796 45428 47802
rect 45376 47738 45428 47744
rect 46676 47734 46704 48311
rect 47032 48272 47084 48278
rect 47032 48214 47084 48220
rect 46664 47728 46716 47734
rect 46664 47670 46716 47676
rect 45560 47048 45612 47054
rect 45560 46990 45612 46996
rect 46296 47048 46348 47054
rect 46296 46990 46348 46996
rect 45020 46702 45232 46730
rect 44180 46164 44232 46170
rect 44180 46106 44232 46112
rect 44916 46164 44968 46170
rect 44916 46106 44968 46112
rect 44180 27872 44232 27878
rect 44180 27814 44232 27820
rect 44192 23322 44220 27814
rect 45020 24342 45048 46702
rect 45192 46504 45244 46510
rect 45192 46446 45244 46452
rect 45204 45490 45232 46446
rect 45192 45484 45244 45490
rect 45192 45426 45244 45432
rect 45572 35086 45600 46990
rect 46112 46504 46164 46510
rect 46112 46446 46164 46452
rect 45652 45960 45704 45966
rect 45652 45902 45704 45908
rect 45836 45960 45888 45966
rect 45836 45902 45888 45908
rect 45560 35080 45612 35086
rect 45560 35022 45612 35028
rect 45468 30388 45520 30394
rect 45468 30330 45520 30336
rect 45480 29209 45508 30330
rect 45466 29200 45522 29209
rect 45466 29135 45522 29144
rect 45466 26344 45522 26353
rect 45466 26279 45522 26288
rect 45008 24336 45060 24342
rect 45008 24278 45060 24284
rect 44180 23316 44232 23322
rect 44180 23258 44232 23264
rect 45480 21486 45508 26279
rect 45572 23526 45600 35022
rect 45664 25770 45692 45902
rect 45848 45490 45876 45902
rect 46124 45558 46152 46446
rect 46112 45552 46164 45558
rect 46112 45494 46164 45500
rect 45836 45484 45888 45490
rect 45836 45426 45888 45432
rect 46204 45484 46256 45490
rect 46204 45426 46256 45432
rect 45744 45348 45796 45354
rect 45744 45290 45796 45296
rect 45652 25764 45704 25770
rect 45652 25706 45704 25712
rect 45560 23520 45612 23526
rect 45560 23462 45612 23468
rect 45468 21480 45520 21486
rect 45468 21422 45520 21428
rect 43996 14272 44048 14278
rect 43996 14214 44048 14220
rect 45756 6914 45784 45290
rect 46018 44296 46074 44305
rect 46018 44231 46074 44240
rect 45836 43716 45888 43722
rect 45836 43658 45888 43664
rect 45848 43314 45876 43658
rect 45836 43308 45888 43314
rect 45836 43250 45888 43256
rect 45848 20466 45876 43250
rect 45928 38888 45980 38894
rect 45928 38830 45980 38836
rect 45940 31890 45968 38830
rect 45928 31884 45980 31890
rect 45928 31826 45980 31832
rect 46032 26314 46060 44231
rect 46112 34604 46164 34610
rect 46112 34546 46164 34552
rect 46020 26308 46072 26314
rect 46020 26250 46072 26256
rect 46124 22982 46152 34546
rect 46216 33538 46244 45426
rect 46308 45082 46336 46990
rect 46480 46980 46532 46986
rect 46480 46922 46532 46928
rect 46492 45558 46520 46922
rect 47044 46646 47072 48214
rect 47676 48068 47728 48074
rect 47676 48010 47728 48016
rect 47584 47524 47636 47530
rect 47584 47466 47636 47472
rect 47124 47456 47176 47462
rect 47124 47398 47176 47404
rect 47032 46640 47084 46646
rect 47032 46582 47084 46588
rect 46480 45552 46532 45558
rect 46480 45494 46532 45500
rect 46480 45280 46532 45286
rect 46480 45222 46532 45228
rect 46296 45076 46348 45082
rect 46296 45018 46348 45024
rect 46386 44976 46442 44985
rect 46492 44946 46520 45222
rect 46386 44911 46442 44920
rect 46480 44940 46532 44946
rect 46296 44872 46348 44878
rect 46296 44814 46348 44820
rect 46308 44402 46336 44814
rect 46296 44396 46348 44402
rect 46296 44338 46348 44344
rect 46296 42016 46348 42022
rect 46296 41958 46348 41964
rect 46308 41682 46336 41958
rect 46296 41676 46348 41682
rect 46296 41618 46348 41624
rect 46296 39840 46348 39846
rect 46296 39782 46348 39788
rect 46308 39506 46336 39782
rect 46296 39500 46348 39506
rect 46296 39442 46348 39448
rect 46296 36576 46348 36582
rect 46296 36518 46348 36524
rect 46308 36242 46336 36518
rect 46296 36236 46348 36242
rect 46296 36178 46348 36184
rect 46296 35488 46348 35494
rect 46296 35430 46348 35436
rect 46308 35154 46336 35430
rect 46296 35148 46348 35154
rect 46296 35090 46348 35096
rect 46216 33510 46336 33538
rect 46204 33448 46256 33454
rect 46202 33416 46204 33425
rect 46256 33416 46258 33425
rect 46202 33351 46258 33360
rect 46308 29170 46336 33510
rect 46296 29164 46348 29170
rect 46296 29106 46348 29112
rect 46296 24608 46348 24614
rect 46296 24550 46348 24556
rect 46308 24274 46336 24550
rect 46296 24268 46348 24274
rect 46296 24210 46348 24216
rect 46112 22976 46164 22982
rect 46112 22918 46164 22924
rect 45836 20460 45888 20466
rect 45836 20402 45888 20408
rect 46112 20324 46164 20330
rect 46112 20266 46164 20272
rect 45664 6886 45784 6914
rect 45664 5234 45692 6886
rect 45652 5228 45704 5234
rect 45652 5170 45704 5176
rect 43996 3936 44048 3942
rect 43996 3878 44048 3884
rect 44916 3936 44968 3942
rect 44916 3878 44968 3884
rect 43444 3732 43496 3738
rect 43444 3674 43496 3680
rect 43904 3528 43956 3534
rect 43904 3470 43956 3476
rect 43444 3460 43496 3466
rect 43444 3402 43496 3408
rect 43168 3052 43220 3058
rect 43168 2994 43220 3000
rect 42616 2848 42668 2854
rect 42616 2790 42668 2796
rect 42628 2514 42656 2790
rect 42432 2508 42484 2514
rect 42432 2450 42484 2456
rect 42616 2508 42668 2514
rect 42616 2450 42668 2456
rect 42708 2508 42760 2514
rect 42708 2450 42760 2456
rect 42720 1170 42748 2450
rect 42536 1142 42748 1170
rect 42536 800 42564 1142
rect 43180 800 43208 2994
rect 43456 2922 43484 3402
rect 43916 3194 43944 3470
rect 43904 3188 43956 3194
rect 43904 3130 43956 3136
rect 44008 3058 44036 3878
rect 44180 3392 44232 3398
rect 44180 3334 44232 3340
rect 44192 3126 44220 3334
rect 44180 3120 44232 3126
rect 44180 3062 44232 3068
rect 43996 3052 44048 3058
rect 43996 2994 44048 3000
rect 44456 2984 44508 2990
rect 44456 2926 44508 2932
rect 43444 2916 43496 2922
rect 43444 2858 43496 2864
rect 44468 800 44496 2926
rect 44928 2514 44956 3878
rect 45192 3392 45244 3398
rect 45192 3334 45244 3340
rect 45204 2514 45232 3334
rect 45664 2854 45692 5170
rect 46124 3194 46152 20266
rect 46400 18698 46428 44911
rect 46480 44882 46532 44888
rect 47032 44192 47084 44198
rect 47032 44134 47084 44140
rect 47044 43858 47072 44134
rect 47032 43852 47084 43858
rect 47032 43794 47084 43800
rect 46940 43716 46992 43722
rect 46940 43658 46992 43664
rect 46952 43450 46980 43658
rect 46940 43444 46992 43450
rect 46940 43386 46992 43392
rect 46480 41540 46532 41546
rect 46480 41482 46532 41488
rect 46492 41274 46520 41482
rect 46480 41268 46532 41274
rect 46480 41210 46532 41216
rect 46664 41132 46716 41138
rect 46664 41074 46716 41080
rect 46480 40452 46532 40458
rect 46480 40394 46532 40400
rect 46492 40186 46520 40394
rect 46480 40180 46532 40186
rect 46480 40122 46532 40128
rect 46572 34604 46624 34610
rect 46572 34546 46624 34552
rect 46480 34400 46532 34406
rect 46480 34342 46532 34348
rect 46492 34066 46520 34342
rect 46480 34060 46532 34066
rect 46480 34002 46532 34008
rect 46584 26246 46612 34546
rect 46572 26240 46624 26246
rect 46572 26182 46624 26188
rect 46676 23594 46704 41074
rect 47136 40746 47164 47398
rect 47596 46578 47624 47466
rect 47688 46714 47716 48010
rect 47872 47734 47900 48991
rect 47860 47728 47912 47734
rect 47860 47670 47912 47676
rect 47768 47456 47820 47462
rect 47768 47398 47820 47404
rect 47676 46708 47728 46714
rect 47676 46650 47728 46656
rect 47584 46572 47636 46578
rect 47584 46514 47636 46520
rect 47596 45490 47624 46514
rect 47584 45484 47636 45490
rect 47584 45426 47636 45432
rect 47216 43104 47268 43110
rect 47216 43046 47268 43052
rect 46952 40718 47164 40746
rect 46756 39364 46808 39370
rect 46756 39306 46808 39312
rect 46768 39098 46796 39306
rect 46756 39092 46808 39098
rect 46756 39034 46808 39040
rect 46756 38752 46808 38758
rect 46756 38694 46808 38700
rect 46768 37874 46796 38694
rect 46756 37868 46808 37874
rect 46756 37810 46808 37816
rect 46846 37496 46902 37505
rect 46846 37431 46902 37440
rect 46860 37330 46888 37431
rect 46848 37324 46900 37330
rect 46848 37266 46900 37272
rect 46848 34536 46900 34542
rect 46848 34478 46900 34484
rect 46860 32842 46888 34478
rect 46848 32836 46900 32842
rect 46848 32778 46900 32784
rect 46664 23588 46716 23594
rect 46664 23530 46716 23536
rect 46952 22234 46980 40718
rect 47124 38208 47176 38214
rect 47124 38150 47176 38156
rect 47032 35488 47084 35494
rect 47032 35430 47084 35436
rect 47044 34134 47072 35430
rect 47032 34128 47084 34134
rect 47032 34070 47084 34076
rect 47136 22710 47164 38150
rect 47124 22704 47176 22710
rect 47124 22646 47176 22652
rect 46940 22228 46992 22234
rect 46940 22170 46992 22176
rect 46480 20256 46532 20262
rect 46480 20198 46532 20204
rect 46492 19922 46520 20198
rect 46480 19916 46532 19922
rect 46480 19858 46532 19864
rect 46388 18692 46440 18698
rect 46388 18634 46440 18640
rect 46846 17776 46902 17785
rect 46846 17711 46902 17720
rect 46860 17542 46888 17711
rect 47124 17672 47176 17678
rect 47124 17614 47176 17620
rect 46848 17536 46900 17542
rect 46848 17478 46900 17484
rect 46480 16992 46532 16998
rect 46480 16934 46532 16940
rect 46492 16658 46520 16934
rect 46480 16652 46532 16658
rect 46480 16594 46532 16600
rect 47032 15904 47084 15910
rect 47032 15846 47084 15852
rect 46480 14816 46532 14822
rect 46480 14758 46532 14764
rect 46492 14482 46520 14758
rect 47044 14550 47072 15846
rect 47136 15638 47164 17614
rect 47124 15632 47176 15638
rect 47124 15574 47176 15580
rect 47032 14544 47084 14550
rect 47032 14486 47084 14492
rect 46480 14476 46532 14482
rect 46480 14418 46532 14424
rect 47228 14346 47256 43046
rect 47400 40928 47452 40934
rect 47400 40870 47452 40876
rect 47308 31816 47360 31822
rect 47308 31758 47360 31764
rect 47320 31385 47348 31758
rect 47306 31376 47362 31385
rect 47306 31311 47362 31320
rect 47308 29300 47360 29306
rect 47308 29242 47360 29248
rect 47320 24818 47348 29242
rect 47308 24812 47360 24818
rect 47308 24754 47360 24760
rect 47412 22710 47440 40870
rect 47676 36100 47728 36106
rect 47676 36042 47728 36048
rect 47688 34746 47716 36042
rect 47676 34740 47728 34746
rect 47676 34682 47728 34688
rect 47584 34604 47636 34610
rect 47584 34546 47636 34552
rect 47492 32360 47544 32366
rect 47492 32302 47544 32308
rect 47504 29306 47532 32302
rect 47492 29300 47544 29306
rect 47492 29242 47544 29248
rect 47492 29096 47544 29102
rect 47492 29038 47544 29044
rect 47504 23798 47532 29038
rect 47596 24818 47624 34546
rect 47676 34536 47728 34542
rect 47676 34478 47728 34484
rect 47688 32586 47716 34478
rect 47780 33402 47808 47398
rect 47860 43308 47912 43314
rect 47860 43250 47912 43256
rect 47872 42945 47900 43250
rect 47858 42936 47914 42945
rect 47858 42871 47914 42880
rect 47964 42786 47992 49030
rect 48228 48544 48280 48550
rect 48228 48486 48280 48492
rect 48136 47048 48188 47054
rect 48134 47016 48136 47025
rect 48188 47016 48190 47025
rect 48134 46951 48190 46960
rect 48134 46336 48190 46345
rect 48134 46271 48190 46280
rect 48148 46034 48176 46271
rect 48136 46028 48188 46034
rect 48136 45970 48188 45976
rect 48134 45656 48190 45665
rect 48134 45591 48190 45600
rect 48148 44946 48176 45591
rect 48136 44940 48188 44946
rect 48136 44882 48188 44888
rect 48136 43716 48188 43722
rect 48136 43658 48188 43664
rect 48148 43625 48176 43658
rect 48134 43616 48190 43625
rect 48134 43551 48190 43560
rect 47872 42758 47992 42786
rect 47872 40746 47900 42758
rect 47952 42628 48004 42634
rect 47952 42570 48004 42576
rect 47964 42265 47992 42570
rect 48044 42560 48096 42566
rect 48044 42502 48096 42508
rect 48056 42362 48084 42502
rect 48044 42356 48096 42362
rect 48044 42298 48096 42304
rect 47950 42256 48006 42265
rect 47950 42191 48006 42200
rect 48136 41608 48188 41614
rect 48134 41576 48136 41585
rect 48188 41576 48190 41585
rect 48134 41511 48190 41520
rect 47952 41132 48004 41138
rect 47952 41074 48004 41080
rect 47964 40905 47992 41074
rect 47950 40896 48006 40905
rect 47950 40831 48006 40840
rect 47872 40718 47992 40746
rect 47860 38344 47912 38350
rect 47860 38286 47912 38292
rect 47872 38185 47900 38286
rect 47858 38176 47914 38185
rect 47858 38111 47914 38120
rect 47858 36136 47914 36145
rect 47858 36071 47914 36080
rect 47872 35698 47900 36071
rect 47860 35692 47912 35698
rect 47860 35634 47912 35640
rect 47780 33374 47900 33402
rect 47768 33312 47820 33318
rect 47768 33254 47820 33260
rect 47780 32978 47808 33254
rect 47768 32972 47820 32978
rect 47768 32914 47820 32920
rect 47688 32558 47808 32586
rect 47676 32428 47728 32434
rect 47676 32370 47728 32376
rect 47688 32065 47716 32370
rect 47674 32056 47730 32065
rect 47674 31991 47730 32000
rect 47780 29102 47808 32558
rect 47768 29096 47820 29102
rect 47768 29038 47820 29044
rect 47676 28960 47728 28966
rect 47676 28902 47728 28908
rect 47688 28626 47716 28902
rect 47676 28620 47728 28626
rect 47676 28562 47728 28568
rect 47676 28484 47728 28490
rect 47676 28426 47728 28432
rect 47688 27606 47716 28426
rect 47676 27600 47728 27606
rect 47676 27542 47728 27548
rect 47872 26234 47900 33374
rect 47964 31090 47992 40718
rect 48136 40452 48188 40458
rect 48136 40394 48188 40400
rect 48148 40225 48176 40394
rect 48134 40216 48190 40225
rect 48134 40151 48190 40160
rect 48134 39536 48190 39545
rect 48134 39471 48136 39480
rect 48188 39471 48190 39480
rect 48136 39442 48188 39448
rect 48136 38956 48188 38962
rect 48136 38898 48188 38904
rect 48148 38865 48176 38898
rect 48134 38856 48190 38865
rect 48134 38791 48190 38800
rect 48134 36816 48190 36825
rect 48134 36751 48190 36760
rect 48148 36242 48176 36751
rect 48136 36236 48188 36242
rect 48136 36178 48188 36184
rect 48044 35488 48096 35494
rect 48044 35430 48096 35436
rect 48134 35456 48190 35465
rect 48056 34542 48084 35430
rect 48134 35391 48190 35400
rect 48148 35154 48176 35391
rect 48136 35148 48188 35154
rect 48136 35090 48188 35096
rect 48134 34776 48190 34785
rect 48134 34711 48190 34720
rect 48044 34536 48096 34542
rect 48044 34478 48096 34484
rect 48042 34096 48098 34105
rect 48148 34066 48176 34711
rect 48042 34031 48098 34040
rect 48136 34060 48188 34066
rect 48056 32978 48084 34031
rect 48136 34002 48188 34008
rect 48044 32972 48096 32978
rect 48044 32914 48096 32920
rect 47964 31062 48176 31090
rect 47952 30252 48004 30258
rect 47952 30194 48004 30200
rect 47964 30025 47992 30194
rect 48044 30048 48096 30054
rect 47950 30016 48006 30025
rect 48044 29990 48096 29996
rect 47950 29951 48006 29960
rect 48056 29782 48084 29990
rect 48044 29776 48096 29782
rect 48044 29718 48096 29724
rect 48148 29594 48176 31062
rect 48056 29566 48176 29594
rect 47952 28076 48004 28082
rect 47952 28018 48004 28024
rect 47964 27985 47992 28018
rect 47950 27976 48006 27985
rect 47950 27911 48006 27920
rect 47952 26308 48004 26314
rect 47952 26250 48004 26256
rect 47780 26206 47900 26234
rect 47584 24812 47636 24818
rect 47584 24754 47636 24760
rect 47676 24608 47728 24614
rect 47676 24550 47728 24556
rect 47688 24274 47716 24550
rect 47676 24268 47728 24274
rect 47676 24210 47728 24216
rect 47492 23792 47544 23798
rect 47492 23734 47544 23740
rect 47584 22976 47636 22982
rect 47584 22918 47636 22924
rect 47400 22704 47452 22710
rect 47400 22646 47452 22652
rect 47412 22098 47440 22646
rect 47596 22642 47624 22918
rect 47584 22636 47636 22642
rect 47584 22578 47636 22584
rect 47400 22092 47452 22098
rect 47400 22034 47452 22040
rect 47596 22030 47624 22578
rect 47676 22432 47728 22438
rect 47676 22374 47728 22380
rect 47584 22024 47636 22030
rect 47584 21966 47636 21972
rect 47688 20874 47716 22374
rect 47676 20868 47728 20874
rect 47676 20810 47728 20816
rect 47492 20460 47544 20466
rect 47492 20402 47544 20408
rect 47216 14340 47268 14346
rect 47216 14282 47268 14288
rect 46754 13016 46810 13025
rect 46754 12951 46810 12960
rect 46768 11898 46796 12951
rect 46848 12436 46900 12442
rect 46848 12378 46900 12384
rect 46860 12345 46888 12378
rect 46846 12336 46902 12345
rect 46846 12271 46902 12280
rect 46756 11892 46808 11898
rect 46756 11834 46808 11840
rect 47216 11144 47268 11150
rect 47216 11086 47268 11092
rect 46846 9616 46902 9625
rect 46846 9551 46902 9560
rect 46860 9178 46888 9551
rect 46848 9172 46900 9178
rect 46848 9114 46900 9120
rect 46480 8832 46532 8838
rect 46480 8774 46532 8780
rect 46492 7818 46520 8774
rect 47032 8288 47084 8294
rect 47032 8230 47084 8236
rect 47044 7954 47072 8230
rect 47032 7948 47084 7954
rect 47032 7890 47084 7896
rect 46480 7812 46532 7818
rect 46480 7754 46532 7760
rect 46846 6896 46902 6905
rect 46846 6831 46902 6840
rect 46860 6458 46888 6831
rect 46848 6452 46900 6458
rect 46848 6394 46900 6400
rect 46754 6216 46810 6225
rect 46754 6151 46810 6160
rect 46768 5302 46796 6151
rect 46848 5364 46900 5370
rect 46848 5306 46900 5312
rect 46756 5296 46808 5302
rect 46756 5238 46808 5244
rect 46296 5024 46348 5030
rect 46296 4966 46348 4972
rect 46308 4690 46336 4966
rect 46296 4684 46348 4690
rect 46296 4626 46348 4632
rect 46756 4208 46808 4214
rect 46860 4185 46888 5306
rect 46756 4150 46808 4156
rect 46846 4176 46902 4185
rect 46388 4140 46440 4146
rect 46388 4082 46440 4088
rect 46204 3596 46256 3602
rect 46204 3538 46256 3544
rect 46216 3505 46244 3538
rect 46202 3496 46258 3505
rect 46202 3431 46258 3440
rect 46112 3188 46164 3194
rect 46112 3130 46164 3136
rect 45744 3052 45796 3058
rect 45744 2994 45796 3000
rect 45652 2848 45704 2854
rect 45652 2790 45704 2796
rect 44916 2508 44968 2514
rect 44916 2450 44968 2456
rect 45192 2508 45244 2514
rect 45192 2450 45244 2456
rect 45376 2508 45428 2514
rect 45376 2450 45428 2456
rect 45112 870 45232 898
rect 45112 800 45140 870
rect 37476 734 37780 762
rect 38014 0 38070 800
rect 38658 0 38714 800
rect 39946 0 40002 800
rect 40590 0 40646 800
rect 41234 0 41290 800
rect 41878 0 41934 800
rect 42522 0 42578 800
rect 43166 0 43222 800
rect 43810 0 43866 800
rect 44454 0 44510 800
rect 45098 0 45154 800
rect 45204 762 45232 870
rect 45388 762 45416 2450
rect 45756 800 45784 2994
rect 45836 2644 45888 2650
rect 45836 2586 45888 2592
rect 45848 1465 45876 2586
rect 45834 1456 45890 1465
rect 45834 1391 45890 1400
rect 46400 800 46428 4082
rect 46480 3936 46532 3942
rect 46480 3878 46532 3884
rect 46492 3602 46520 3878
rect 46480 3596 46532 3602
rect 46480 3538 46532 3544
rect 45204 734 45416 762
rect 45742 0 45798 800
rect 46386 0 46442 800
rect 46768 105 46796 4150
rect 46846 4111 46902 4120
rect 46940 4140 46992 4146
rect 46940 4082 46992 4088
rect 46952 3466 46980 4082
rect 47228 4078 47256 11086
rect 47308 11008 47360 11014
rect 47308 10950 47360 10956
rect 47320 10130 47348 10950
rect 47308 10124 47360 10130
rect 47308 10066 47360 10072
rect 47504 4146 47532 20402
rect 47676 19780 47728 19786
rect 47676 19722 47728 19728
rect 47688 18970 47716 19722
rect 47780 19514 47808 26206
rect 47964 25945 47992 26250
rect 47950 25936 48006 25945
rect 47950 25871 48006 25880
rect 47860 25288 47912 25294
rect 47858 25256 47860 25265
rect 47912 25256 47914 25265
rect 47858 25191 47914 25200
rect 48056 24834 48084 29566
rect 48134 28656 48190 28665
rect 48134 28591 48136 28600
rect 48188 28591 48190 28600
rect 48136 28562 48188 28568
rect 48136 26308 48188 26314
rect 48136 26250 48188 26256
rect 47872 24806 48084 24834
rect 47872 22234 47900 24806
rect 48148 24698 48176 26250
rect 48056 24670 48176 24698
rect 48056 24410 48084 24670
rect 48134 24576 48190 24585
rect 48134 24511 48190 24520
rect 48044 24404 48096 24410
rect 48044 24346 48096 24352
rect 48148 24274 48176 24511
rect 48136 24268 48188 24274
rect 48136 24210 48188 24216
rect 47950 23896 48006 23905
rect 47950 23831 48006 23840
rect 47964 23798 47992 23831
rect 47952 23792 48004 23798
rect 47952 23734 48004 23740
rect 48136 23112 48188 23118
rect 48136 23054 48188 23060
rect 48148 22545 48176 23054
rect 48134 22536 48190 22545
rect 48134 22471 48190 22480
rect 47860 22228 47912 22234
rect 47860 22170 47912 22176
rect 47860 22024 47912 22030
rect 47860 21966 47912 21972
rect 47872 21690 47900 21966
rect 47950 21856 48006 21865
rect 47950 21791 48006 21800
rect 47860 21684 47912 21690
rect 47860 21626 47912 21632
rect 47872 20074 47900 21626
rect 47964 21622 47992 21791
rect 47952 21616 48004 21622
rect 47952 21558 48004 21564
rect 48240 21418 48268 48486
rect 48332 48210 48360 51200
rect 48976 49230 49004 51200
rect 48964 49224 49016 49230
rect 48964 49166 49016 49172
rect 49620 48278 49648 51200
rect 49608 48272 49660 48278
rect 49608 48214 49660 48220
rect 48320 48204 48372 48210
rect 48320 48146 48372 48152
rect 48504 25220 48556 25226
rect 48504 25162 48556 25168
rect 48228 21412 48280 21418
rect 48228 21354 48280 21360
rect 48044 21344 48096 21350
rect 48044 21286 48096 21292
rect 48056 21078 48084 21286
rect 48044 21072 48096 21078
rect 48044 21014 48096 21020
rect 47872 20046 47992 20074
rect 47768 19508 47820 19514
rect 47768 19450 47820 19456
rect 47860 19372 47912 19378
rect 47860 19314 47912 19320
rect 47872 19145 47900 19314
rect 47858 19136 47914 19145
rect 47858 19071 47914 19080
rect 47676 18964 47728 18970
rect 47676 18906 47728 18912
rect 47768 16992 47820 16998
rect 47768 16934 47820 16940
rect 47780 16726 47808 16934
rect 47768 16720 47820 16726
rect 47768 16662 47820 16668
rect 47584 16108 47636 16114
rect 47584 16050 47636 16056
rect 47596 15026 47624 16050
rect 47676 15904 47728 15910
rect 47676 15846 47728 15852
rect 47688 15570 47716 15846
rect 47676 15564 47728 15570
rect 47676 15506 47728 15512
rect 47964 15162 47992 20046
rect 48134 19816 48190 19825
rect 48134 19751 48136 19760
rect 48188 19751 48190 19760
rect 48136 19722 48188 19728
rect 48044 19168 48096 19174
rect 48044 19110 48096 19116
rect 47952 15156 48004 15162
rect 47952 15098 48004 15104
rect 47860 15088 47912 15094
rect 47860 15030 47912 15036
rect 47950 15056 48006 15065
rect 47584 15020 47636 15026
rect 47584 14962 47636 14968
rect 47872 14074 47900 15030
rect 47950 14991 47952 15000
rect 48004 14991 48006 15000
rect 47952 14962 48004 14968
rect 47860 14068 47912 14074
rect 47860 14010 47912 14016
rect 47860 13932 47912 13938
rect 47860 13874 47912 13880
rect 47872 13705 47900 13874
rect 47858 13696 47914 13705
rect 47858 13631 47914 13640
rect 48056 11234 48084 19110
rect 48134 17096 48190 17105
rect 48134 17031 48190 17040
rect 48148 16658 48176 17031
rect 48136 16652 48188 16658
rect 48136 16594 48188 16600
rect 48134 16416 48190 16425
rect 48134 16351 48190 16360
rect 48148 15570 48176 16351
rect 48136 15564 48188 15570
rect 48136 15506 48188 15512
rect 48134 14376 48190 14385
rect 48134 14311 48136 14320
rect 48188 14311 48190 14320
rect 48136 14282 48188 14288
rect 47964 11206 48084 11234
rect 47964 10742 47992 11206
rect 48044 11144 48096 11150
rect 48044 11086 48096 11092
rect 47952 10736 48004 10742
rect 47952 10678 48004 10684
rect 47768 10668 47820 10674
rect 47768 10610 47820 10616
rect 47780 10305 47808 10610
rect 47766 10296 47822 10305
rect 47766 10231 47822 10240
rect 48056 10198 48084 11086
rect 48134 10976 48190 10985
rect 48134 10911 48190 10920
rect 48044 10192 48096 10198
rect 48044 10134 48096 10140
rect 48148 10130 48176 10911
rect 48136 10124 48188 10130
rect 48136 10066 48188 10072
rect 47950 8936 48006 8945
rect 47950 8871 47952 8880
rect 48004 8871 48006 8880
rect 47952 8842 48004 8848
rect 47860 8492 47912 8498
rect 47860 8434 47912 8440
rect 47872 8265 47900 8434
rect 47858 8256 47914 8265
rect 47858 8191 47914 8200
rect 48136 7812 48188 7818
rect 48136 7754 48188 7760
rect 48148 7585 48176 7754
rect 48134 7576 48190 7585
rect 48134 7511 48190 7520
rect 47860 5704 47912 5710
rect 47860 5646 47912 5652
rect 47872 5545 47900 5646
rect 47858 5536 47914 5545
rect 47858 5471 47914 5480
rect 47676 5024 47728 5030
rect 47676 4966 47728 4972
rect 47688 4690 47716 4966
rect 48134 4856 48190 4865
rect 48134 4791 48190 4800
rect 48148 4690 48176 4791
rect 47676 4684 47728 4690
rect 47676 4626 47728 4632
rect 48136 4684 48188 4690
rect 48136 4626 48188 4632
rect 47492 4140 47544 4146
rect 47492 4082 47544 4088
rect 47216 4072 47268 4078
rect 47216 4014 47268 4020
rect 47032 3732 47084 3738
rect 47032 3674 47084 3680
rect 46940 3460 46992 3466
rect 46940 3402 46992 3408
rect 47044 800 47072 3674
rect 48044 3664 48096 3670
rect 48044 3606 48096 3612
rect 48056 3194 48084 3606
rect 48320 3460 48372 3466
rect 48320 3402 48372 3408
rect 48044 3188 48096 3194
rect 48044 3130 48096 3136
rect 47768 2372 47820 2378
rect 47768 2314 47820 2320
rect 46754 96 46810 105
rect 46754 31 46810 40
rect 47030 0 47086 800
rect 47674 0 47730 800
rect 47780 785 47808 2314
rect 47860 2304 47912 2310
rect 47860 2246 47912 2252
rect 47872 2038 47900 2246
rect 47860 2032 47912 2038
rect 47860 1974 47912 1980
rect 48332 800 48360 3402
rect 47766 776 47822 785
rect 47766 711 47822 720
rect 48318 0 48374 800
rect 48516 762 48544 25162
rect 49608 3052 49660 3058
rect 49608 2994 49660 3000
rect 48884 870 49004 898
rect 48884 762 48912 870
rect 48976 800 49004 870
rect 49620 800 49648 2994
rect 48516 734 48912 762
rect 48962 0 49018 800
rect 49606 0 49662 800
<< via2 >>
rect 1398 47640 1454 47696
rect 1398 34720 1454 34776
rect 1398 31320 1454 31376
rect 1398 25900 1454 25936
rect 1398 25880 1400 25900
rect 1400 25880 1452 25900
rect 1452 25880 1454 25900
rect 2870 51720 2926 51776
rect 3422 51040 3478 51096
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 1858 46960 1914 47016
rect 1858 45600 1914 45656
rect 1858 44240 1914 44296
rect 1858 43560 1914 43616
rect 1858 41520 1914 41576
rect 1858 40840 1914 40896
rect 1858 40160 1914 40216
rect 1858 37440 1914 37496
rect 1858 36760 1914 36816
rect 2318 31184 2374 31240
rect 1858 23840 1914 23896
rect 1858 22480 1914 22536
rect 1398 12280 1454 12336
rect 2410 30912 2466 30968
rect 2962 46280 3018 46336
rect 2778 44920 2834 44976
rect 2778 39480 2834 39536
rect 2778 36080 2834 36136
rect 2778 34060 2834 34096
rect 2778 34040 2780 34060
rect 2780 34040 2832 34060
rect 2832 34040 2834 34060
rect 2778 33396 2780 33416
rect 2780 33396 2832 33416
rect 2832 33396 2834 33416
rect 2778 33360 2834 33396
rect 3054 32680 3110 32736
rect 3054 32000 3110 32056
rect 2778 29960 2834 30016
rect 2778 28620 2834 28656
rect 2778 28600 2780 28620
rect 2780 28600 2832 28620
rect 2832 28600 2834 28620
rect 2778 27240 2834 27296
rect 2778 26560 2834 26616
rect 2226 19080 2282 19136
rect 1858 17040 1914 17096
rect 1858 10920 1914 10976
rect 1858 8200 1914 8256
rect 1858 7520 1914 7576
rect 1858 3440 1914 3496
rect 2778 23180 2834 23216
rect 2778 23160 2780 23180
rect 2780 23160 2832 23180
rect 2832 23160 2834 23180
rect 2778 17740 2834 17776
rect 2778 17720 2780 17740
rect 2780 17720 2832 17740
rect 2832 17720 2834 17740
rect 2778 16360 2834 16416
rect 3330 48320 3386 48376
rect 4066 49000 4122 49056
rect 3422 38120 3478 38176
rect 2778 13640 2834 13696
rect 2778 10240 2834 10296
rect 2778 9560 2834 9616
rect 2778 6860 2834 6896
rect 2778 6840 2780 6860
rect 2780 6840 2832 6860
rect 2832 6840 2834 6860
rect 2778 5480 2834 5536
rect 2778 4800 2834 4856
rect 2226 2372 2282 2408
rect 2226 2352 2228 2372
rect 2228 2352 2280 2372
rect 2280 2352 2282 2372
rect 3146 2080 3202 2136
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 4710 50360 4766 50416
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4066 29280 4122 29336
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 3974 21800 4030 21856
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4066 21120 4122 21176
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4066 19760 4122 19816
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 3422 8880 3478 8936
rect 3422 6160 3478 6216
rect 3422 4120 3478 4176
rect 4066 18400 4122 18456
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4066 12960 4122 13016
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4802 2524 4804 2544
rect 4804 2524 4856 2544
rect 4856 2524 4858 2544
rect 4802 2488 4858 2524
rect 1858 720 1914 776
rect 11702 24012 11704 24032
rect 11704 24012 11756 24032
rect 11756 24012 11758 24032
rect 11702 23976 11758 24012
rect 10782 22636 10838 22672
rect 10782 22616 10784 22636
rect 10784 22616 10836 22636
rect 10836 22616 10838 22636
rect 10966 19352 11022 19408
rect 12162 30812 12164 30832
rect 12164 30812 12216 30832
rect 12216 30812 12218 30832
rect 12162 30776 12218 30812
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 13266 30812 13268 30832
rect 13268 30812 13320 30832
rect 13320 30812 13322 30832
rect 13266 30776 13322 30812
rect 12530 19352 12586 19408
rect 12162 3304 12218 3360
rect 13726 22516 13728 22536
rect 13728 22516 13780 22536
rect 13780 22516 13782 22536
rect 13726 22480 13782 22516
rect 14922 22500 14978 22536
rect 14922 22480 14924 22500
rect 14924 22480 14976 22500
rect 14976 22480 14978 22500
rect 15474 29180 15476 29200
rect 15476 29180 15528 29200
rect 15528 29180 15530 29200
rect 15474 29144 15530 29180
rect 15750 20576 15806 20632
rect 16946 29164 17002 29200
rect 16946 29144 16948 29164
rect 16948 29144 17000 29164
rect 17000 29144 17002 29164
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 16578 23976 16634 24032
rect 17406 24012 17408 24032
rect 17408 24012 17460 24032
rect 17460 24012 17462 24032
rect 17406 23976 17462 24012
rect 16670 20440 16726 20496
rect 12622 3304 12678 3360
rect 18326 31864 18382 31920
rect 18418 22616 18474 22672
rect 17958 20596 18014 20632
rect 17958 20576 17960 20596
rect 17960 20576 18012 20596
rect 18012 20576 18014 20596
rect 18142 20460 18198 20496
rect 18142 20440 18144 20460
rect 18144 20440 18196 20460
rect 18196 20440 18198 20460
rect 18326 8372 18328 8392
rect 18328 8372 18380 8392
rect 18380 8372 18382 8392
rect 18326 8336 18382 8372
rect 19154 31864 19210 31920
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19890 22480 19946 22536
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19798 19352 19854 19408
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19890 17176 19946 17232
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 20258 13232 20314 13288
rect 20166 12552 20222 12608
rect 20350 12552 20406 12608
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19430 11076 19486 11112
rect 19430 11056 19432 11076
rect 19432 11056 19484 11076
rect 19484 11056 19486 11076
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19430 10376 19486 10432
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 21270 31728 21326 31784
rect 22742 31764 22744 31784
rect 22744 31764 22796 31784
rect 22796 31764 22798 31784
rect 22742 31728 22798 31764
rect 23202 32544 23258 32600
rect 20810 22380 20812 22400
rect 20812 22380 20864 22400
rect 20864 22380 20866 22400
rect 20810 22344 20866 22380
rect 20994 17176 21050 17232
rect 21086 8336 21142 8392
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 21270 18028 21272 18048
rect 21272 18028 21324 18048
rect 21324 18028 21326 18048
rect 21270 17992 21326 18028
rect 21454 19760 21510 19816
rect 21546 18672 21602 18728
rect 21730 18264 21786 18320
rect 22190 21956 22246 21992
rect 22190 21936 22192 21956
rect 22192 21936 22244 21956
rect 22244 21936 22246 21956
rect 22374 21428 22376 21448
rect 22376 21428 22428 21448
rect 22428 21428 22430 21448
rect 22374 21392 22430 21428
rect 22374 21140 22430 21176
rect 22374 21120 22376 21140
rect 22376 21120 22428 21140
rect 22428 21120 22430 21140
rect 22466 19372 22522 19408
rect 22466 19352 22468 19372
rect 22468 19352 22520 19372
rect 22520 19352 22522 19372
rect 23478 32408 23534 32464
rect 23478 32000 23534 32056
rect 23662 39888 23718 39944
rect 23846 39888 23902 39944
rect 23478 29588 23480 29608
rect 23480 29588 23532 29608
rect 23532 29588 23534 29608
rect 23478 29552 23534 29588
rect 23018 21392 23074 21448
rect 23110 21120 23166 21176
rect 22926 19760 22982 19816
rect 22926 18572 22928 18592
rect 22928 18572 22980 18592
rect 22980 18572 22982 18592
rect 22926 18536 22982 18572
rect 23018 17040 23074 17096
rect 24122 32408 24178 32464
rect 23478 21936 23534 21992
rect 23662 21936 23718 21992
rect 23386 17448 23442 17504
rect 23386 16768 23442 16824
rect 24030 18808 24086 18864
rect 24214 18400 24270 18456
rect 24030 16904 24086 16960
rect 23570 12688 23626 12744
rect 24214 16788 24270 16824
rect 24214 16768 24216 16788
rect 24216 16768 24268 16788
rect 24268 16768 24270 16788
rect 23938 12280 23994 12336
rect 24030 11076 24086 11112
rect 24030 11056 24032 11076
rect 24032 11056 24084 11076
rect 24084 11056 24086 11076
rect 25134 29588 25136 29608
rect 25136 29588 25188 29608
rect 25188 29588 25190 29608
rect 25134 29552 25190 29588
rect 24398 17040 24454 17096
rect 24490 16768 24546 16824
rect 24398 16516 24454 16552
rect 24398 16496 24400 16516
rect 24400 16496 24452 16516
rect 24452 16496 24454 16516
rect 24490 16360 24546 16416
rect 25226 22344 25282 22400
rect 25318 21800 25374 21856
rect 24950 18572 24952 18592
rect 24952 18572 25004 18592
rect 25004 18572 25006 18592
rect 24950 18536 25006 18572
rect 24858 18128 24914 18184
rect 24950 17584 25006 17640
rect 24858 16768 24914 16824
rect 25134 12708 25190 12744
rect 25134 12688 25136 12708
rect 25136 12688 25188 12708
rect 25188 12688 25190 12708
rect 25686 32544 25742 32600
rect 25778 32000 25834 32056
rect 25594 26988 25650 27024
rect 25594 26968 25596 26988
rect 25596 26968 25648 26988
rect 25648 26968 25650 26988
rect 25502 22072 25558 22128
rect 25594 17196 25650 17232
rect 25594 17176 25596 17196
rect 25596 17176 25648 17196
rect 25648 17176 25650 17196
rect 26882 33088 26938 33144
rect 26054 21548 26110 21584
rect 26054 21528 26056 21548
rect 26056 21528 26108 21548
rect 26108 21528 26110 21548
rect 26606 21664 26662 21720
rect 26514 21528 26570 21584
rect 26698 21392 26754 21448
rect 26882 22480 26938 22536
rect 26974 21256 27030 21312
rect 27434 26968 27490 27024
rect 27986 26988 28042 27024
rect 27986 26968 27988 26988
rect 27988 26968 28040 26988
rect 28040 26968 28042 26988
rect 27342 21528 27398 21584
rect 27434 20848 27490 20904
rect 28354 25236 28356 25256
rect 28356 25236 28408 25256
rect 28408 25236 28410 25256
rect 28354 25200 28410 25236
rect 26054 18264 26110 18320
rect 26146 18164 26148 18184
rect 26148 18164 26200 18184
rect 26200 18164 26202 18184
rect 26146 18128 26202 18164
rect 26422 18672 26478 18728
rect 26238 17620 26240 17640
rect 26240 17620 26292 17640
rect 26292 17620 26294 17640
rect 26238 17584 26294 17620
rect 26974 17448 27030 17504
rect 27066 17196 27122 17232
rect 27066 17176 27068 17196
rect 27068 17176 27120 17196
rect 27120 17176 27122 17196
rect 25870 16360 25926 16416
rect 27158 16496 27214 16552
rect 26790 14764 26792 14784
rect 26792 14764 26844 14784
rect 26844 14764 26846 14784
rect 26790 14728 26846 14764
rect 27250 14184 27306 14240
rect 27526 17992 27582 18048
rect 27710 18264 27766 18320
rect 27986 16652 28042 16688
rect 27986 16632 27988 16652
rect 27988 16632 28040 16652
rect 28040 16632 28042 16652
rect 27802 15272 27858 15328
rect 27894 14220 27896 14240
rect 27896 14220 27948 14240
rect 27948 14220 27950 14240
rect 27894 14184 27950 14220
rect 29182 42356 29238 42392
rect 29182 42336 29184 42356
rect 29184 42336 29236 42356
rect 29236 42336 29238 42356
rect 29550 48048 29606 48104
rect 30838 42356 30894 42392
rect 30838 42336 30840 42356
rect 30840 42336 30892 42356
rect 30892 42336 30894 42356
rect 29366 31748 29422 31784
rect 29366 31728 29368 31748
rect 29368 31728 29420 31748
rect 29420 31728 29422 31748
rect 29734 33088 29790 33144
rect 29642 25220 29698 25256
rect 29642 25200 29644 25220
rect 29644 25200 29696 25220
rect 29696 25200 29698 25220
rect 29642 23976 29698 24032
rect 31114 40468 31116 40488
rect 31116 40468 31168 40488
rect 31168 40468 31170 40488
rect 31114 40432 31170 40468
rect 30930 39244 30932 39264
rect 30932 39244 30984 39264
rect 30984 39244 30986 39264
rect 30930 39208 30986 39244
rect 30746 31748 30802 31784
rect 30746 31728 30748 31748
rect 30748 31728 30800 31748
rect 30800 31728 30802 31748
rect 32402 40432 32458 40488
rect 32310 39380 32312 39400
rect 32312 39380 32364 39400
rect 32364 39380 32366 39400
rect 32310 39344 32366 39380
rect 31482 33088 31538 33144
rect 31758 29008 31814 29064
rect 31666 23724 31722 23760
rect 31666 23704 31668 23724
rect 31668 23704 31720 23724
rect 31720 23704 31722 23724
rect 28538 21392 28594 21448
rect 28170 21120 28226 21176
rect 28170 20712 28226 20768
rect 27802 9016 27858 9072
rect 27894 8336 27950 8392
rect 28354 13912 28410 13968
rect 28262 8744 28318 8800
rect 28722 22092 28778 22128
rect 28722 22072 28724 22092
rect 28724 22072 28776 22092
rect 28776 22072 28778 22092
rect 29642 22092 29698 22128
rect 29642 22072 29644 22092
rect 29644 22072 29696 22092
rect 29696 22072 29698 22092
rect 28814 21972 28816 21992
rect 28816 21972 28868 21992
rect 28868 21972 28870 21992
rect 28814 21936 28870 21972
rect 29550 21936 29606 21992
rect 29734 21972 29736 21992
rect 29736 21972 29788 21992
rect 29788 21972 29790 21992
rect 29734 21936 29790 21972
rect 29090 21664 29146 21720
rect 28630 17720 28686 17776
rect 28538 12144 28594 12200
rect 29274 20712 29330 20768
rect 28998 17212 29000 17232
rect 29000 17212 29052 17232
rect 29052 17212 29054 17232
rect 28998 17176 29054 17212
rect 28998 17076 29000 17096
rect 29000 17076 29052 17096
rect 29052 17076 29054 17096
rect 28998 17040 29054 17076
rect 29182 15020 29238 15056
rect 29182 15000 29184 15020
rect 29184 15000 29236 15020
rect 29236 15000 29238 15020
rect 30194 22072 30250 22128
rect 29458 21292 29460 21312
rect 29460 21292 29512 21312
rect 29512 21292 29514 21312
rect 29458 21256 29514 21292
rect 29458 21120 29514 21176
rect 29918 20984 29974 21040
rect 30010 20848 30066 20904
rect 30746 22652 30748 22672
rect 30748 22652 30800 22672
rect 30800 22652 30802 22672
rect 30746 22616 30802 22652
rect 30470 21800 30526 21856
rect 29458 17040 29514 17096
rect 28814 12144 28870 12200
rect 28538 8744 28594 8800
rect 28998 9444 29054 9480
rect 28998 9424 29000 9444
rect 29000 9424 29052 9444
rect 29052 9424 29054 9444
rect 29734 14456 29790 14512
rect 30286 15000 30342 15056
rect 31482 21528 31538 21584
rect 31114 18400 31170 18456
rect 31022 17040 31078 17096
rect 30930 15272 30986 15328
rect 31574 21020 31576 21040
rect 31576 21020 31628 21040
rect 31628 21020 31630 21040
rect 31574 20984 31630 21020
rect 33598 39344 33654 39400
rect 33506 39072 33562 39128
rect 32494 29180 32496 29200
rect 32496 29180 32548 29200
rect 32548 29180 32550 29200
rect 32494 29144 32550 29180
rect 32770 21936 32826 21992
rect 32126 18536 32182 18592
rect 32034 18264 32090 18320
rect 32586 15136 32642 15192
rect 32494 14864 32550 14920
rect 32678 13776 32734 13832
rect 33506 29008 33562 29064
rect 33138 9460 33140 9480
rect 33140 9460 33192 9480
rect 33192 9460 33194 9480
rect 33138 9424 33194 9460
rect 33414 14864 33470 14920
rect 33782 29164 33838 29200
rect 33782 29144 33784 29164
rect 33784 29144 33836 29164
rect 33836 29144 33838 29164
rect 33966 23840 34022 23896
rect 33598 22652 33600 22672
rect 33600 22652 33652 22672
rect 33652 22652 33654 22672
rect 33598 22616 33654 22652
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 35438 48048 35494 48104
rect 35714 48084 35716 48104
rect 35716 48084 35768 48104
rect 35768 48084 35770 48104
rect 35714 48048 35770 48084
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34334 39208 34390 39264
rect 35438 38936 35494 38992
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34518 23568 34574 23624
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34886 23976 34942 24032
rect 34978 23840 35034 23896
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34518 17040 34574 17096
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 35254 17196 35310 17232
rect 35254 17176 35256 17196
rect 35256 17176 35308 17196
rect 35308 17176 35310 17196
rect 35622 17040 35678 17096
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34794 14728 34850 14784
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 35530 14456 35586 14512
rect 35346 14356 35348 14376
rect 35348 14356 35400 14376
rect 35400 14356 35402 14376
rect 35346 14320 35402 14356
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 36082 23588 36138 23624
rect 36082 23568 36084 23588
rect 36084 23568 36136 23588
rect 36136 23568 36138 23588
rect 36450 23704 36506 23760
rect 37002 14320 37058 14376
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 37462 39072 37518 39128
rect 37370 38956 37426 38992
rect 37370 38936 37372 38956
rect 37372 38936 37424 38956
rect 37424 38936 37426 38956
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 46662 51720 46718 51776
rect 46754 51040 46810 51096
rect 46846 50360 46902 50416
rect 46846 49680 46902 49736
rect 47858 49000 47914 49056
rect 46662 48320 46718 48376
rect 45466 29144 45522 29200
rect 45466 26288 45522 26344
rect 46018 44240 46074 44296
rect 46386 44920 46442 44976
rect 46202 33396 46204 33416
rect 46204 33396 46256 33416
rect 46256 33396 46258 33416
rect 46202 33360 46258 33396
rect 46846 37440 46902 37496
rect 46846 17720 46902 17776
rect 47306 31320 47362 31376
rect 47858 42880 47914 42936
rect 48134 46996 48136 47016
rect 48136 46996 48188 47016
rect 48188 46996 48190 47016
rect 48134 46960 48190 46996
rect 48134 46280 48190 46336
rect 48134 45600 48190 45656
rect 48134 43560 48190 43616
rect 47950 42200 48006 42256
rect 48134 41556 48136 41576
rect 48136 41556 48188 41576
rect 48188 41556 48190 41576
rect 48134 41520 48190 41556
rect 47950 40840 48006 40896
rect 47858 38120 47914 38176
rect 47858 36080 47914 36136
rect 47674 32000 47730 32056
rect 48134 40160 48190 40216
rect 48134 39500 48190 39536
rect 48134 39480 48136 39500
rect 48136 39480 48188 39500
rect 48188 39480 48190 39500
rect 48134 38800 48190 38856
rect 48134 36760 48190 36816
rect 48134 35400 48190 35456
rect 48134 34720 48190 34776
rect 48042 34040 48098 34096
rect 47950 29960 48006 30016
rect 47950 27920 48006 27976
rect 46754 12960 46810 13016
rect 46846 12280 46902 12336
rect 46846 9560 46902 9616
rect 46846 6840 46902 6896
rect 46754 6160 46810 6216
rect 46202 3440 46258 3496
rect 45834 1400 45890 1456
rect 46846 4120 46902 4176
rect 47950 25880 48006 25936
rect 47858 25236 47860 25256
rect 47860 25236 47912 25256
rect 47912 25236 47914 25256
rect 47858 25200 47914 25236
rect 48134 28620 48190 28656
rect 48134 28600 48136 28620
rect 48136 28600 48188 28620
rect 48188 28600 48190 28620
rect 48134 24520 48190 24576
rect 47950 23840 48006 23896
rect 48134 22480 48190 22536
rect 47950 21800 48006 21856
rect 47858 19080 47914 19136
rect 48134 19780 48190 19816
rect 48134 19760 48136 19780
rect 48136 19760 48188 19780
rect 48188 19760 48190 19780
rect 47950 15020 48006 15056
rect 47950 15000 47952 15020
rect 47952 15000 48004 15020
rect 48004 15000 48006 15020
rect 47858 13640 47914 13696
rect 48134 17040 48190 17096
rect 48134 16360 48190 16416
rect 48134 14340 48190 14376
rect 48134 14320 48136 14340
rect 48136 14320 48188 14340
rect 48188 14320 48190 14340
rect 47766 10240 47822 10296
rect 48134 10920 48190 10976
rect 47950 8900 48006 8936
rect 47950 8880 47952 8900
rect 47952 8880 48004 8900
rect 48004 8880 48006 8900
rect 47858 8200 47914 8256
rect 48134 7520 48190 7576
rect 47858 5480 47914 5536
rect 48134 4800 48190 4856
rect 46754 40 46810 96
rect 47766 720 47822 776
<< metal3 >>
rect 0 51778 800 51808
rect 2865 51778 2931 51781
rect 0 51776 2931 51778
rect 0 51720 2870 51776
rect 2926 51720 2931 51776
rect 0 51718 2931 51720
rect 0 51688 800 51718
rect 2865 51715 2931 51718
rect 46657 51778 46723 51781
rect 49200 51778 50000 51808
rect 46657 51776 50000 51778
rect 46657 51720 46662 51776
rect 46718 51720 50000 51776
rect 46657 51718 50000 51720
rect 46657 51715 46723 51718
rect 49200 51688 50000 51718
rect 0 51098 800 51128
rect 3417 51098 3483 51101
rect 0 51096 3483 51098
rect 0 51040 3422 51096
rect 3478 51040 3483 51096
rect 0 51038 3483 51040
rect 0 51008 800 51038
rect 3417 51035 3483 51038
rect 46749 51098 46815 51101
rect 49200 51098 50000 51128
rect 46749 51096 50000 51098
rect 46749 51040 46754 51096
rect 46810 51040 50000 51096
rect 46749 51038 50000 51040
rect 46749 51035 46815 51038
rect 49200 51008 50000 51038
rect 0 50418 800 50448
rect 4705 50418 4771 50421
rect 0 50416 4771 50418
rect 0 50360 4710 50416
rect 4766 50360 4771 50416
rect 0 50358 4771 50360
rect 0 50328 800 50358
rect 4705 50355 4771 50358
rect 46841 50418 46907 50421
rect 49200 50418 50000 50448
rect 46841 50416 50000 50418
rect 46841 50360 46846 50416
rect 46902 50360 50000 50416
rect 46841 50358 50000 50360
rect 46841 50355 46907 50358
rect 49200 50328 50000 50358
rect 0 49648 800 49768
rect 46841 49738 46907 49741
rect 49200 49738 50000 49768
rect 46841 49736 50000 49738
rect 46841 49680 46846 49736
rect 46902 49680 50000 49736
rect 46841 49678 50000 49680
rect 46841 49675 46907 49678
rect 49200 49648 50000 49678
rect 4208 49536 4528 49537
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 49471 4528 49472
rect 34928 49536 35248 49537
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 49471 35248 49472
rect 0 49058 800 49088
rect 4061 49058 4127 49061
rect 0 49056 4127 49058
rect 0 49000 4066 49056
rect 4122 49000 4127 49056
rect 0 48998 4127 49000
rect 0 48968 800 48998
rect 4061 48995 4127 48998
rect 47853 49058 47919 49061
rect 49200 49058 50000 49088
rect 47853 49056 50000 49058
rect 47853 49000 47858 49056
rect 47914 49000 50000 49056
rect 47853 48998 50000 49000
rect 47853 48995 47919 48998
rect 19568 48992 19888 48993
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 49200 48968 50000 48998
rect 19568 48927 19888 48928
rect 4208 48448 4528 48449
rect 0 48378 800 48408
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 48383 4528 48384
rect 34928 48448 35248 48449
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 48383 35248 48384
rect 3325 48378 3391 48381
rect 0 48376 3391 48378
rect 0 48320 3330 48376
rect 3386 48320 3391 48376
rect 0 48318 3391 48320
rect 0 48288 800 48318
rect 3325 48315 3391 48318
rect 46657 48378 46723 48381
rect 49200 48378 50000 48408
rect 46657 48376 50000 48378
rect 46657 48320 46662 48376
rect 46718 48320 50000 48376
rect 46657 48318 50000 48320
rect 46657 48315 46723 48318
rect 49200 48288 50000 48318
rect 29545 48106 29611 48109
rect 35433 48106 35499 48109
rect 35709 48106 35775 48109
rect 29545 48104 35775 48106
rect 29545 48048 29550 48104
rect 29606 48048 35438 48104
rect 35494 48048 35714 48104
rect 35770 48048 35775 48104
rect 29545 48046 35775 48048
rect 29545 48043 29611 48046
rect 35433 48043 35499 48046
rect 35709 48043 35775 48046
rect 19568 47904 19888 47905
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 47839 19888 47840
rect 0 47698 800 47728
rect 1393 47698 1459 47701
rect 0 47696 1459 47698
rect 0 47640 1398 47696
rect 1454 47640 1459 47696
rect 0 47638 1459 47640
rect 0 47608 800 47638
rect 1393 47635 1459 47638
rect 49200 47608 50000 47728
rect 4208 47360 4528 47361
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 47295 4528 47296
rect 34928 47360 35248 47361
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 47295 35248 47296
rect 0 47018 800 47048
rect 1853 47018 1919 47021
rect 0 47016 1919 47018
rect 0 46960 1858 47016
rect 1914 46960 1919 47016
rect 0 46958 1919 46960
rect 0 46928 800 46958
rect 1853 46955 1919 46958
rect 48129 47018 48195 47021
rect 49200 47018 50000 47048
rect 48129 47016 50000 47018
rect 48129 46960 48134 47016
rect 48190 46960 50000 47016
rect 48129 46958 50000 46960
rect 48129 46955 48195 46958
rect 49200 46928 50000 46958
rect 19568 46816 19888 46817
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 46751 19888 46752
rect 0 46338 800 46368
rect 2957 46338 3023 46341
rect 0 46336 3023 46338
rect 0 46280 2962 46336
rect 3018 46280 3023 46336
rect 0 46278 3023 46280
rect 0 46248 800 46278
rect 2957 46275 3023 46278
rect 48129 46338 48195 46341
rect 49200 46338 50000 46368
rect 48129 46336 50000 46338
rect 48129 46280 48134 46336
rect 48190 46280 50000 46336
rect 48129 46278 50000 46280
rect 48129 46275 48195 46278
rect 4208 46272 4528 46273
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 46207 4528 46208
rect 34928 46272 35248 46273
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 49200 46248 50000 46278
rect 34928 46207 35248 46208
rect 19568 45728 19888 45729
rect 0 45658 800 45688
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 45663 19888 45664
rect 1853 45658 1919 45661
rect 0 45656 1919 45658
rect 0 45600 1858 45656
rect 1914 45600 1919 45656
rect 0 45598 1919 45600
rect 0 45568 800 45598
rect 1853 45595 1919 45598
rect 48129 45658 48195 45661
rect 49200 45658 50000 45688
rect 48129 45656 50000 45658
rect 48129 45600 48134 45656
rect 48190 45600 50000 45656
rect 48129 45598 50000 45600
rect 48129 45595 48195 45598
rect 49200 45568 50000 45598
rect 4208 45184 4528 45185
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 45119 4528 45120
rect 34928 45184 35248 45185
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 45119 35248 45120
rect 0 44978 800 45008
rect 2773 44978 2839 44981
rect 0 44976 2839 44978
rect 0 44920 2778 44976
rect 2834 44920 2839 44976
rect 0 44918 2839 44920
rect 0 44888 800 44918
rect 2773 44915 2839 44918
rect 46381 44978 46447 44981
rect 49200 44978 50000 45008
rect 46381 44976 50000 44978
rect 46381 44920 46386 44976
rect 46442 44920 50000 44976
rect 46381 44918 50000 44920
rect 46381 44915 46447 44918
rect 49200 44888 50000 44918
rect 19568 44640 19888 44641
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 44575 19888 44576
rect 0 44298 800 44328
rect 1853 44298 1919 44301
rect 0 44296 1919 44298
rect 0 44240 1858 44296
rect 1914 44240 1919 44296
rect 0 44238 1919 44240
rect 0 44208 800 44238
rect 1853 44235 1919 44238
rect 46013 44298 46079 44301
rect 49200 44298 50000 44328
rect 46013 44296 50000 44298
rect 46013 44240 46018 44296
rect 46074 44240 50000 44296
rect 46013 44238 50000 44240
rect 46013 44235 46079 44238
rect 49200 44208 50000 44238
rect 4208 44096 4528 44097
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 44031 4528 44032
rect 34928 44096 35248 44097
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 44031 35248 44032
rect 0 43618 800 43648
rect 1853 43618 1919 43621
rect 0 43616 1919 43618
rect 0 43560 1858 43616
rect 1914 43560 1919 43616
rect 0 43558 1919 43560
rect 0 43528 800 43558
rect 1853 43555 1919 43558
rect 48129 43618 48195 43621
rect 49200 43618 50000 43648
rect 48129 43616 50000 43618
rect 48129 43560 48134 43616
rect 48190 43560 50000 43616
rect 48129 43558 50000 43560
rect 48129 43555 48195 43558
rect 19568 43552 19888 43553
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 49200 43528 50000 43558
rect 19568 43487 19888 43488
rect 4208 43008 4528 43009
rect 0 42848 800 42968
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 42943 4528 42944
rect 34928 43008 35248 43009
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 42943 35248 42944
rect 47853 42938 47919 42941
rect 49200 42938 50000 42968
rect 47853 42936 50000 42938
rect 47853 42880 47858 42936
rect 47914 42880 50000 42936
rect 47853 42878 50000 42880
rect 47853 42875 47919 42878
rect 49200 42848 50000 42878
rect 19568 42464 19888 42465
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 42399 19888 42400
rect 29177 42394 29243 42397
rect 30833 42394 30899 42397
rect 29177 42392 30899 42394
rect 29177 42336 29182 42392
rect 29238 42336 30838 42392
rect 30894 42336 30899 42392
rect 29177 42334 30899 42336
rect 29177 42331 29243 42334
rect 30833 42331 30899 42334
rect 47945 42258 48011 42261
rect 49200 42258 50000 42288
rect 47945 42256 50000 42258
rect 47945 42200 47950 42256
rect 48006 42200 50000 42256
rect 47945 42198 50000 42200
rect 47945 42195 48011 42198
rect 49200 42168 50000 42198
rect 4208 41920 4528 41921
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 41855 4528 41856
rect 34928 41920 35248 41921
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 41855 35248 41856
rect 0 41578 800 41608
rect 1853 41578 1919 41581
rect 0 41576 1919 41578
rect 0 41520 1858 41576
rect 1914 41520 1919 41576
rect 0 41518 1919 41520
rect 0 41488 800 41518
rect 1853 41515 1919 41518
rect 48129 41578 48195 41581
rect 49200 41578 50000 41608
rect 48129 41576 50000 41578
rect 48129 41520 48134 41576
rect 48190 41520 50000 41576
rect 48129 41518 50000 41520
rect 48129 41515 48195 41518
rect 49200 41488 50000 41518
rect 19568 41376 19888 41377
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 41311 19888 41312
rect 0 40898 800 40928
rect 1853 40898 1919 40901
rect 0 40896 1919 40898
rect 0 40840 1858 40896
rect 1914 40840 1919 40896
rect 0 40838 1919 40840
rect 0 40808 800 40838
rect 1853 40835 1919 40838
rect 47945 40898 48011 40901
rect 49200 40898 50000 40928
rect 47945 40896 50000 40898
rect 47945 40840 47950 40896
rect 48006 40840 50000 40896
rect 47945 40838 50000 40840
rect 47945 40835 48011 40838
rect 4208 40832 4528 40833
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 40767 4528 40768
rect 34928 40832 35248 40833
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 49200 40808 50000 40838
rect 34928 40767 35248 40768
rect 31109 40490 31175 40493
rect 32397 40490 32463 40493
rect 31109 40488 32463 40490
rect 31109 40432 31114 40488
rect 31170 40432 32402 40488
rect 32458 40432 32463 40488
rect 31109 40430 32463 40432
rect 31109 40427 31175 40430
rect 32397 40427 32463 40430
rect 19568 40288 19888 40289
rect 0 40218 800 40248
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 40223 19888 40224
rect 1853 40218 1919 40221
rect 0 40216 1919 40218
rect 0 40160 1858 40216
rect 1914 40160 1919 40216
rect 0 40158 1919 40160
rect 0 40128 800 40158
rect 1853 40155 1919 40158
rect 48129 40218 48195 40221
rect 49200 40218 50000 40248
rect 48129 40216 50000 40218
rect 48129 40160 48134 40216
rect 48190 40160 50000 40216
rect 48129 40158 50000 40160
rect 48129 40155 48195 40158
rect 49200 40128 50000 40158
rect 23657 39946 23723 39949
rect 23841 39946 23907 39949
rect 23657 39944 23907 39946
rect 23657 39888 23662 39944
rect 23718 39888 23846 39944
rect 23902 39888 23907 39944
rect 23657 39886 23907 39888
rect 23657 39883 23723 39886
rect 23841 39883 23907 39886
rect 4208 39744 4528 39745
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 0 39538 800 39568
rect 2773 39538 2839 39541
rect 0 39536 2839 39538
rect 0 39480 2778 39536
rect 2834 39480 2839 39536
rect 0 39478 2839 39480
rect 0 39448 800 39478
rect 2773 39475 2839 39478
rect 48129 39538 48195 39541
rect 49200 39538 50000 39568
rect 48129 39536 50000 39538
rect 48129 39480 48134 39536
rect 48190 39480 50000 39536
rect 48129 39478 50000 39480
rect 48129 39475 48195 39478
rect 49200 39448 50000 39478
rect 32305 39402 32371 39405
rect 33593 39402 33659 39405
rect 32305 39400 33659 39402
rect 32305 39344 32310 39400
rect 32366 39344 33598 39400
rect 33654 39344 33659 39400
rect 32305 39342 33659 39344
rect 32305 39339 32371 39342
rect 33593 39339 33659 39342
rect 30925 39266 30991 39269
rect 34329 39266 34395 39269
rect 30925 39264 34395 39266
rect 30925 39208 30930 39264
rect 30986 39208 34334 39264
rect 34390 39208 34395 39264
rect 30925 39206 34395 39208
rect 30925 39203 30991 39206
rect 34329 39203 34395 39206
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 39135 19888 39136
rect 33501 39130 33567 39133
rect 37457 39130 37523 39133
rect 33501 39128 37523 39130
rect 33501 39072 33506 39128
rect 33562 39072 37462 39128
rect 37518 39072 37523 39128
rect 33501 39070 37523 39072
rect 33501 39067 33567 39070
rect 37457 39067 37523 39070
rect 35433 38994 35499 38997
rect 37365 38994 37431 38997
rect 35433 38992 37431 38994
rect 35433 38936 35438 38992
rect 35494 38936 37370 38992
rect 37426 38936 37431 38992
rect 35433 38934 37431 38936
rect 35433 38931 35499 38934
rect 37365 38931 37431 38934
rect 0 38768 800 38888
rect 48129 38858 48195 38861
rect 49200 38858 50000 38888
rect 48129 38856 50000 38858
rect 48129 38800 48134 38856
rect 48190 38800 50000 38856
rect 48129 38798 50000 38800
rect 48129 38795 48195 38798
rect 49200 38768 50000 38798
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 38591 35248 38592
rect 0 38178 800 38208
rect 3417 38178 3483 38181
rect 0 38176 3483 38178
rect 0 38120 3422 38176
rect 3478 38120 3483 38176
rect 0 38118 3483 38120
rect 0 38088 800 38118
rect 3417 38115 3483 38118
rect 47853 38178 47919 38181
rect 49200 38178 50000 38208
rect 47853 38176 50000 38178
rect 47853 38120 47858 38176
rect 47914 38120 50000 38176
rect 47853 38118 50000 38120
rect 47853 38115 47919 38118
rect 19568 38112 19888 38113
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 49200 38088 50000 38118
rect 19568 38047 19888 38048
rect 4208 37568 4528 37569
rect 0 37498 800 37528
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 1853 37498 1919 37501
rect 0 37496 1919 37498
rect 0 37440 1858 37496
rect 1914 37440 1919 37496
rect 0 37438 1919 37440
rect 0 37408 800 37438
rect 1853 37435 1919 37438
rect 46841 37498 46907 37501
rect 49200 37498 50000 37528
rect 46841 37496 50000 37498
rect 46841 37440 46846 37496
rect 46902 37440 50000 37496
rect 46841 37438 50000 37440
rect 46841 37435 46907 37438
rect 49200 37408 50000 37438
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 0 36818 800 36848
rect 1853 36818 1919 36821
rect 0 36816 1919 36818
rect 0 36760 1858 36816
rect 1914 36760 1919 36816
rect 0 36758 1919 36760
rect 0 36728 800 36758
rect 1853 36755 1919 36758
rect 48129 36818 48195 36821
rect 49200 36818 50000 36848
rect 48129 36816 50000 36818
rect 48129 36760 48134 36816
rect 48190 36760 50000 36816
rect 48129 36758 50000 36760
rect 48129 36755 48195 36758
rect 49200 36728 50000 36758
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 0 36138 800 36168
rect 2773 36138 2839 36141
rect 0 36136 2839 36138
rect 0 36080 2778 36136
rect 2834 36080 2839 36136
rect 0 36078 2839 36080
rect 0 36048 800 36078
rect 2773 36075 2839 36078
rect 47853 36138 47919 36141
rect 49200 36138 50000 36168
rect 47853 36136 50000 36138
rect 47853 36080 47858 36136
rect 47914 36080 50000 36136
rect 47853 36078 50000 36080
rect 47853 36075 47919 36078
rect 49200 36048 50000 36078
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 0 35368 800 35488
rect 48129 35458 48195 35461
rect 49200 35458 50000 35488
rect 48129 35456 50000 35458
rect 48129 35400 48134 35456
rect 48190 35400 50000 35456
rect 48129 35398 50000 35400
rect 48129 35395 48195 35398
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 49200 35368 50000 35398
rect 34928 35327 35248 35328
rect 19568 34848 19888 34849
rect 0 34778 800 34808
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 1393 34778 1459 34781
rect 0 34776 1459 34778
rect 0 34720 1398 34776
rect 1454 34720 1459 34776
rect 0 34718 1459 34720
rect 0 34688 800 34718
rect 1393 34715 1459 34718
rect 48129 34778 48195 34781
rect 49200 34778 50000 34808
rect 48129 34776 50000 34778
rect 48129 34720 48134 34776
rect 48190 34720 50000 34776
rect 48129 34718 50000 34720
rect 48129 34715 48195 34718
rect 49200 34688 50000 34718
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 0 34098 800 34128
rect 2773 34098 2839 34101
rect 0 34096 2839 34098
rect 0 34040 2778 34096
rect 2834 34040 2839 34096
rect 0 34038 2839 34040
rect 0 34008 800 34038
rect 2773 34035 2839 34038
rect 48037 34098 48103 34101
rect 49200 34098 50000 34128
rect 48037 34096 50000 34098
rect 48037 34040 48042 34096
rect 48098 34040 50000 34096
rect 48037 34038 50000 34040
rect 48037 34035 48103 34038
rect 49200 34008 50000 34038
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 0 33418 800 33448
rect 2773 33418 2839 33421
rect 0 33416 2839 33418
rect 0 33360 2778 33416
rect 2834 33360 2839 33416
rect 0 33358 2839 33360
rect 0 33328 800 33358
rect 2773 33355 2839 33358
rect 46197 33418 46263 33421
rect 49200 33418 50000 33448
rect 46197 33416 50000 33418
rect 46197 33360 46202 33416
rect 46258 33360 50000 33416
rect 46197 33358 50000 33360
rect 46197 33355 46263 33358
rect 49200 33328 50000 33358
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 26877 33146 26943 33149
rect 29729 33146 29795 33149
rect 31477 33146 31543 33149
rect 26877 33144 31543 33146
rect 26877 33088 26882 33144
rect 26938 33088 29734 33144
rect 29790 33088 31482 33144
rect 31538 33088 31543 33144
rect 26877 33086 31543 33088
rect 26877 33083 26943 33086
rect 29729 33083 29795 33086
rect 31477 33083 31543 33086
rect 0 32738 800 32768
rect 3049 32738 3115 32741
rect 0 32736 3115 32738
rect 0 32680 3054 32736
rect 3110 32680 3115 32736
rect 0 32678 3115 32680
rect 0 32648 800 32678
rect 3049 32675 3115 32678
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 49200 32648 50000 32768
rect 19568 32607 19888 32608
rect 23197 32602 23263 32605
rect 25681 32602 25747 32605
rect 23197 32600 25747 32602
rect 23197 32544 23202 32600
rect 23258 32544 25686 32600
rect 25742 32544 25747 32600
rect 23197 32542 25747 32544
rect 23197 32539 23263 32542
rect 25681 32539 25747 32542
rect 23473 32466 23539 32469
rect 24117 32466 24183 32469
rect 23473 32464 24183 32466
rect 23473 32408 23478 32464
rect 23534 32408 24122 32464
rect 24178 32408 24183 32464
rect 23473 32406 24183 32408
rect 23473 32403 23539 32406
rect 24117 32403 24183 32406
rect 4208 32128 4528 32129
rect 0 32058 800 32088
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 3049 32058 3115 32061
rect 0 32056 3115 32058
rect 0 32000 3054 32056
rect 3110 32000 3115 32056
rect 0 31998 3115 32000
rect 0 31968 800 31998
rect 3049 31995 3115 31998
rect 23473 32058 23539 32061
rect 25773 32058 25839 32061
rect 23473 32056 25839 32058
rect 23473 32000 23478 32056
rect 23534 32000 25778 32056
rect 25834 32000 25839 32056
rect 23473 31998 25839 32000
rect 23473 31995 23539 31998
rect 25773 31995 25839 31998
rect 47669 32058 47735 32061
rect 49200 32058 50000 32088
rect 47669 32056 50000 32058
rect 47669 32000 47674 32056
rect 47730 32000 50000 32056
rect 47669 31998 50000 32000
rect 47669 31995 47735 31998
rect 49200 31968 50000 31998
rect 18321 31922 18387 31925
rect 19149 31922 19215 31925
rect 18321 31920 19215 31922
rect 18321 31864 18326 31920
rect 18382 31864 19154 31920
rect 19210 31864 19215 31920
rect 18321 31862 19215 31864
rect 18321 31859 18387 31862
rect 19149 31859 19215 31862
rect 21265 31786 21331 31789
rect 22737 31786 22803 31789
rect 21265 31784 22803 31786
rect 21265 31728 21270 31784
rect 21326 31728 22742 31784
rect 22798 31728 22803 31784
rect 21265 31726 22803 31728
rect 21265 31723 21331 31726
rect 22737 31723 22803 31726
rect 29361 31786 29427 31789
rect 30741 31786 30807 31789
rect 29361 31784 30807 31786
rect 29361 31728 29366 31784
rect 29422 31728 30746 31784
rect 30802 31728 30807 31784
rect 29361 31726 30807 31728
rect 29361 31723 29427 31726
rect 30741 31723 30807 31726
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 0 31378 800 31408
rect 1393 31378 1459 31381
rect 0 31376 1459 31378
rect 0 31320 1398 31376
rect 1454 31320 1459 31376
rect 0 31318 1459 31320
rect 0 31288 800 31318
rect 1393 31315 1459 31318
rect 47301 31378 47367 31381
rect 49200 31378 50000 31408
rect 47301 31376 50000 31378
rect 47301 31320 47306 31376
rect 47362 31320 50000 31376
rect 47301 31318 50000 31320
rect 47301 31315 47367 31318
rect 49200 31288 50000 31318
rect 2313 31242 2379 31245
rect 2270 31240 2379 31242
rect 2270 31184 2318 31240
rect 2374 31184 2379 31240
rect 2270 31179 2379 31184
rect 2270 30970 2330 31179
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 2405 30970 2471 30973
rect 2270 30968 2471 30970
rect 2270 30912 2410 30968
rect 2466 30912 2471 30968
rect 2270 30910 2471 30912
rect 2405 30907 2471 30910
rect 12157 30834 12223 30837
rect 13261 30834 13327 30837
rect 12157 30832 13327 30834
rect 12157 30776 12162 30832
rect 12218 30776 13266 30832
rect 13322 30776 13327 30832
rect 12157 30774 13327 30776
rect 12157 30771 12223 30774
rect 13261 30771 13327 30774
rect 0 30608 800 30728
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 0 30018 800 30048
rect 2773 30018 2839 30021
rect 0 30016 2839 30018
rect 0 29960 2778 30016
rect 2834 29960 2839 30016
rect 0 29958 2839 29960
rect 0 29928 800 29958
rect 2773 29955 2839 29958
rect 47945 30018 48011 30021
rect 49200 30018 50000 30048
rect 47945 30016 50000 30018
rect 47945 29960 47950 30016
rect 48006 29960 50000 30016
rect 47945 29958 50000 29960
rect 47945 29955 48011 29958
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 49200 29928 50000 29958
rect 34928 29887 35248 29888
rect 23473 29610 23539 29613
rect 25129 29610 25195 29613
rect 23473 29608 25195 29610
rect 23473 29552 23478 29608
rect 23534 29552 25134 29608
rect 25190 29552 25195 29608
rect 23473 29550 25195 29552
rect 23473 29547 23539 29550
rect 25129 29547 25195 29550
rect 19568 29408 19888 29409
rect 0 29338 800 29368
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 4061 29338 4127 29341
rect 49200 29338 50000 29368
rect 0 29336 4127 29338
rect 0 29280 4066 29336
rect 4122 29280 4127 29336
rect 0 29278 4127 29280
rect 0 29248 800 29278
rect 4061 29275 4127 29278
rect 45510 29278 50000 29338
rect 45510 29205 45570 29278
rect 49200 29248 50000 29278
rect 15469 29202 15535 29205
rect 16941 29202 17007 29205
rect 15469 29200 17007 29202
rect 15469 29144 15474 29200
rect 15530 29144 16946 29200
rect 17002 29144 17007 29200
rect 15469 29142 17007 29144
rect 15469 29139 15535 29142
rect 16941 29139 17007 29142
rect 32489 29202 32555 29205
rect 33777 29202 33843 29205
rect 32489 29200 33843 29202
rect 32489 29144 32494 29200
rect 32550 29144 33782 29200
rect 33838 29144 33843 29200
rect 32489 29142 33843 29144
rect 32489 29139 32555 29142
rect 33777 29139 33843 29142
rect 45461 29200 45570 29205
rect 45461 29144 45466 29200
rect 45522 29144 45570 29200
rect 45461 29142 45570 29144
rect 45461 29139 45527 29142
rect 31753 29066 31819 29069
rect 33501 29066 33567 29069
rect 31753 29064 33567 29066
rect 31753 29008 31758 29064
rect 31814 29008 33506 29064
rect 33562 29008 33567 29064
rect 31753 29006 33567 29008
rect 31753 29003 31819 29006
rect 33501 29003 33567 29006
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 0 28658 800 28688
rect 2773 28658 2839 28661
rect 0 28656 2839 28658
rect 0 28600 2778 28656
rect 2834 28600 2839 28656
rect 0 28598 2839 28600
rect 0 28568 800 28598
rect 2773 28595 2839 28598
rect 48129 28658 48195 28661
rect 49200 28658 50000 28688
rect 48129 28656 50000 28658
rect 48129 28600 48134 28656
rect 48190 28600 50000 28656
rect 48129 28598 50000 28600
rect 48129 28595 48195 28598
rect 49200 28568 50000 28598
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 0 27888 800 28008
rect 47945 27978 48011 27981
rect 49200 27978 50000 28008
rect 47945 27976 50000 27978
rect 47945 27920 47950 27976
rect 48006 27920 50000 27976
rect 47945 27918 50000 27920
rect 47945 27915 48011 27918
rect 49200 27888 50000 27918
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 0 27298 800 27328
rect 2773 27298 2839 27301
rect 0 27296 2839 27298
rect 0 27240 2778 27296
rect 2834 27240 2839 27296
rect 0 27238 2839 27240
rect 0 27208 800 27238
rect 2773 27235 2839 27238
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 49200 27208 50000 27328
rect 19568 27167 19888 27168
rect 25589 27026 25655 27029
rect 27429 27026 27495 27029
rect 27981 27026 28047 27029
rect 25589 27024 28047 27026
rect 25589 26968 25594 27024
rect 25650 26968 27434 27024
rect 27490 26968 27986 27024
rect 28042 26968 28047 27024
rect 25589 26966 28047 26968
rect 25589 26963 25655 26966
rect 27429 26963 27495 26966
rect 27981 26963 28047 26966
rect 4208 26688 4528 26689
rect 0 26618 800 26648
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 2773 26618 2839 26621
rect 49200 26618 50000 26648
rect 0 26616 2839 26618
rect 0 26560 2778 26616
rect 2834 26560 2839 26616
rect 0 26558 2839 26560
rect 0 26528 800 26558
rect 2773 26555 2839 26558
rect 45510 26558 50000 26618
rect 45510 26349 45570 26558
rect 49200 26528 50000 26558
rect 45461 26344 45570 26349
rect 45461 26288 45466 26344
rect 45522 26288 45570 26344
rect 45461 26286 45570 26288
rect 45461 26283 45527 26286
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 0 25938 800 25968
rect 1393 25938 1459 25941
rect 0 25936 1459 25938
rect 0 25880 1398 25936
rect 1454 25880 1459 25936
rect 0 25878 1459 25880
rect 0 25848 800 25878
rect 1393 25875 1459 25878
rect 47945 25938 48011 25941
rect 49200 25938 50000 25968
rect 47945 25936 50000 25938
rect 47945 25880 47950 25936
rect 48006 25880 50000 25936
rect 47945 25878 50000 25880
rect 47945 25875 48011 25878
rect 49200 25848 50000 25878
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 0 25168 800 25288
rect 28349 25258 28415 25261
rect 29637 25258 29703 25261
rect 28349 25256 29703 25258
rect 28349 25200 28354 25256
rect 28410 25200 29642 25256
rect 29698 25200 29703 25256
rect 28349 25198 29703 25200
rect 28349 25195 28415 25198
rect 29637 25195 29703 25198
rect 47853 25258 47919 25261
rect 49200 25258 50000 25288
rect 47853 25256 50000 25258
rect 47853 25200 47858 25256
rect 47914 25200 50000 25256
rect 47853 25198 50000 25200
rect 47853 25195 47919 25198
rect 49200 25168 50000 25198
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 0 24488 800 24608
rect 48129 24578 48195 24581
rect 49200 24578 50000 24608
rect 48129 24576 50000 24578
rect 48129 24520 48134 24576
rect 48190 24520 50000 24576
rect 48129 24518 50000 24520
rect 48129 24515 48195 24518
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 49200 24488 50000 24518
rect 34928 24447 35248 24448
rect 11697 24034 11763 24037
rect 16573 24034 16639 24037
rect 17401 24034 17467 24037
rect 11697 24032 17467 24034
rect 11697 23976 11702 24032
rect 11758 23976 16578 24032
rect 16634 23976 17406 24032
rect 17462 23976 17467 24032
rect 11697 23974 17467 23976
rect 11697 23971 11763 23974
rect 16573 23971 16639 23974
rect 17401 23971 17467 23974
rect 29637 24034 29703 24037
rect 34881 24034 34947 24037
rect 29637 24032 34947 24034
rect 29637 23976 29642 24032
rect 29698 23976 34886 24032
rect 34942 23976 34947 24032
rect 29637 23974 34947 23976
rect 29637 23971 29703 23974
rect 34881 23971 34947 23974
rect 19568 23968 19888 23969
rect 0 23898 800 23928
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 1853 23898 1919 23901
rect 0 23896 1919 23898
rect 0 23840 1858 23896
rect 1914 23840 1919 23896
rect 0 23838 1919 23840
rect 0 23808 800 23838
rect 1853 23835 1919 23838
rect 33961 23898 34027 23901
rect 34973 23898 35039 23901
rect 33961 23896 35039 23898
rect 33961 23840 33966 23896
rect 34022 23840 34978 23896
rect 35034 23840 35039 23896
rect 33961 23838 35039 23840
rect 33961 23835 34027 23838
rect 34973 23835 35039 23838
rect 47945 23898 48011 23901
rect 49200 23898 50000 23928
rect 47945 23896 50000 23898
rect 47945 23840 47950 23896
rect 48006 23840 50000 23896
rect 47945 23838 50000 23840
rect 47945 23835 48011 23838
rect 49200 23808 50000 23838
rect 31661 23762 31727 23765
rect 36445 23762 36511 23765
rect 31661 23760 36511 23762
rect 31661 23704 31666 23760
rect 31722 23704 36450 23760
rect 36506 23704 36511 23760
rect 31661 23702 36511 23704
rect 31661 23699 31727 23702
rect 36445 23699 36511 23702
rect 34513 23626 34579 23629
rect 36077 23626 36143 23629
rect 34513 23624 36143 23626
rect 34513 23568 34518 23624
rect 34574 23568 36082 23624
rect 36138 23568 36143 23624
rect 34513 23566 36143 23568
rect 34513 23563 34579 23566
rect 36077 23563 36143 23566
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 0 23218 800 23248
rect 2773 23218 2839 23221
rect 0 23216 2839 23218
rect 0 23160 2778 23216
rect 2834 23160 2839 23216
rect 0 23158 2839 23160
rect 0 23128 800 23158
rect 2773 23155 2839 23158
rect 49200 23128 50000 23248
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 10777 22674 10843 22677
rect 18413 22674 18479 22677
rect 10777 22672 18479 22674
rect 10777 22616 10782 22672
rect 10838 22616 18418 22672
rect 18474 22616 18479 22672
rect 10777 22614 18479 22616
rect 10777 22611 10843 22614
rect 18413 22611 18479 22614
rect 30741 22674 30807 22677
rect 33593 22674 33659 22677
rect 30741 22672 33659 22674
rect 30741 22616 30746 22672
rect 30802 22616 33598 22672
rect 33654 22616 33659 22672
rect 30741 22614 33659 22616
rect 30741 22611 30807 22614
rect 33593 22611 33659 22614
rect 0 22538 800 22568
rect 1853 22538 1919 22541
rect 0 22536 1919 22538
rect 0 22480 1858 22536
rect 1914 22480 1919 22536
rect 0 22478 1919 22480
rect 0 22448 800 22478
rect 1853 22475 1919 22478
rect 13721 22538 13787 22541
rect 14917 22538 14983 22541
rect 13721 22536 14983 22538
rect 13721 22480 13726 22536
rect 13782 22480 14922 22536
rect 14978 22480 14983 22536
rect 13721 22478 14983 22480
rect 13721 22475 13787 22478
rect 14917 22475 14983 22478
rect 19885 22538 19951 22541
rect 26877 22538 26943 22541
rect 19885 22536 26943 22538
rect 19885 22480 19890 22536
rect 19946 22480 26882 22536
rect 26938 22480 26943 22536
rect 19885 22478 26943 22480
rect 19885 22475 19951 22478
rect 26877 22475 26943 22478
rect 48129 22538 48195 22541
rect 49200 22538 50000 22568
rect 48129 22536 50000 22538
rect 48129 22480 48134 22536
rect 48190 22480 50000 22536
rect 48129 22478 50000 22480
rect 48129 22475 48195 22478
rect 49200 22448 50000 22478
rect 20805 22402 20871 22405
rect 25221 22402 25287 22405
rect 20805 22400 25287 22402
rect 20805 22344 20810 22400
rect 20866 22344 25226 22400
rect 25282 22344 25287 22400
rect 20805 22342 25287 22344
rect 20805 22339 20871 22342
rect 25221 22339 25287 22342
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 25497 22130 25563 22133
rect 28717 22130 28783 22133
rect 25497 22128 28783 22130
rect 25497 22072 25502 22128
rect 25558 22072 28722 22128
rect 28778 22072 28783 22128
rect 25497 22070 28783 22072
rect 25497 22067 25563 22070
rect 28717 22067 28783 22070
rect 29637 22130 29703 22133
rect 30189 22130 30255 22133
rect 29637 22128 30255 22130
rect 29637 22072 29642 22128
rect 29698 22072 30194 22128
rect 30250 22072 30255 22128
rect 29637 22070 30255 22072
rect 29637 22067 29703 22070
rect 30189 22067 30255 22070
rect 22185 21994 22251 21997
rect 23473 21994 23539 21997
rect 23657 21994 23723 21997
rect 28809 21996 28875 21997
rect 28758 21994 28764 21996
rect 22185 21992 23723 21994
rect 22185 21936 22190 21992
rect 22246 21936 23478 21992
rect 23534 21936 23662 21992
rect 23718 21936 23723 21992
rect 22185 21934 23723 21936
rect 28682 21934 28764 21994
rect 28828 21994 28875 21996
rect 29545 21994 29611 21997
rect 28828 21992 29611 21994
rect 28870 21936 29550 21992
rect 29606 21936 29611 21992
rect 22185 21931 22251 21934
rect 23473 21931 23539 21934
rect 23657 21931 23723 21934
rect 28758 21932 28764 21934
rect 28828 21934 29611 21936
rect 28828 21932 28875 21934
rect 28809 21931 28875 21932
rect 29545 21931 29611 21934
rect 29729 21994 29795 21997
rect 32765 21994 32831 21997
rect 29729 21992 32831 21994
rect 29729 21936 29734 21992
rect 29790 21936 32770 21992
rect 32826 21936 32831 21992
rect 29729 21934 32831 21936
rect 29729 21931 29795 21934
rect 32765 21931 32831 21934
rect 0 21858 800 21888
rect 3969 21858 4035 21861
rect 0 21856 4035 21858
rect 0 21800 3974 21856
rect 4030 21800 4035 21856
rect 0 21798 4035 21800
rect 0 21768 800 21798
rect 3969 21795 4035 21798
rect 25313 21858 25379 21861
rect 30465 21858 30531 21861
rect 25313 21856 30531 21858
rect 25313 21800 25318 21856
rect 25374 21800 30470 21856
rect 30526 21800 30531 21856
rect 25313 21798 30531 21800
rect 25313 21795 25379 21798
rect 30465 21795 30531 21798
rect 47945 21858 48011 21861
rect 49200 21858 50000 21888
rect 47945 21856 50000 21858
rect 47945 21800 47950 21856
rect 48006 21800 50000 21856
rect 47945 21798 50000 21800
rect 47945 21795 48011 21798
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 49200 21768 50000 21798
rect 19568 21727 19888 21728
rect 26601 21722 26667 21725
rect 29085 21722 29151 21725
rect 26601 21720 29151 21722
rect 26601 21664 26606 21720
rect 26662 21664 29090 21720
rect 29146 21664 29151 21720
rect 26601 21662 29151 21664
rect 26601 21659 26667 21662
rect 29085 21659 29151 21662
rect 26049 21586 26115 21589
rect 26509 21586 26575 21589
rect 26049 21584 26575 21586
rect 26049 21528 26054 21584
rect 26110 21528 26514 21584
rect 26570 21528 26575 21584
rect 26049 21526 26575 21528
rect 26049 21523 26115 21526
rect 26509 21523 26575 21526
rect 27337 21586 27403 21589
rect 31477 21586 31543 21589
rect 27337 21584 31543 21586
rect 27337 21528 27342 21584
rect 27398 21528 31482 21584
rect 31538 21528 31543 21584
rect 27337 21526 31543 21528
rect 27337 21523 27403 21526
rect 31477 21523 31543 21526
rect 22369 21450 22435 21453
rect 23013 21450 23079 21453
rect 22369 21448 23079 21450
rect 22369 21392 22374 21448
rect 22430 21392 23018 21448
rect 23074 21392 23079 21448
rect 22369 21390 23079 21392
rect 22369 21387 22435 21390
rect 23013 21387 23079 21390
rect 26693 21450 26759 21453
rect 28533 21450 28599 21453
rect 26693 21448 28599 21450
rect 26693 21392 26698 21448
rect 26754 21392 28538 21448
rect 28594 21392 28599 21448
rect 26693 21390 28599 21392
rect 26693 21387 26759 21390
rect 28533 21387 28599 21390
rect 26969 21314 27035 21317
rect 29453 21314 29519 21317
rect 26969 21312 29519 21314
rect 26969 21256 26974 21312
rect 27030 21256 29458 21312
rect 29514 21256 29519 21312
rect 26969 21254 29519 21256
rect 26969 21251 27035 21254
rect 29453 21251 29519 21254
rect 4208 21248 4528 21249
rect 0 21178 800 21208
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 4061 21178 4127 21181
rect 0 21176 4127 21178
rect 0 21120 4066 21176
rect 4122 21120 4127 21176
rect 0 21118 4127 21120
rect 0 21088 800 21118
rect 4061 21115 4127 21118
rect 22369 21178 22435 21181
rect 23105 21178 23171 21181
rect 22369 21176 23171 21178
rect 22369 21120 22374 21176
rect 22430 21120 23110 21176
rect 23166 21120 23171 21176
rect 22369 21118 23171 21120
rect 22369 21115 22435 21118
rect 23105 21115 23171 21118
rect 28165 21178 28231 21181
rect 29453 21178 29519 21181
rect 28165 21176 29519 21178
rect 28165 21120 28170 21176
rect 28226 21120 29458 21176
rect 29514 21120 29519 21176
rect 28165 21118 29519 21120
rect 28165 21115 28231 21118
rect 29453 21115 29519 21118
rect 49200 21088 50000 21208
rect 29913 21042 29979 21045
rect 31569 21042 31635 21045
rect 29913 21040 31635 21042
rect 29913 20984 29918 21040
rect 29974 20984 31574 21040
rect 31630 20984 31635 21040
rect 29913 20982 31635 20984
rect 29913 20979 29979 20982
rect 31569 20979 31635 20982
rect 27429 20906 27495 20909
rect 30005 20906 30071 20909
rect 27429 20904 30071 20906
rect 27429 20848 27434 20904
rect 27490 20848 30010 20904
rect 30066 20848 30071 20904
rect 27429 20846 30071 20848
rect 27429 20843 27495 20846
rect 30005 20843 30071 20846
rect 28165 20770 28231 20773
rect 28390 20770 28396 20772
rect 28165 20768 28396 20770
rect 28165 20712 28170 20768
rect 28226 20712 28396 20768
rect 28165 20710 28396 20712
rect 28165 20707 28231 20710
rect 28390 20708 28396 20710
rect 28460 20770 28466 20772
rect 29269 20770 29335 20773
rect 28460 20768 29335 20770
rect 28460 20712 29274 20768
rect 29330 20712 29335 20768
rect 28460 20710 29335 20712
rect 28460 20708 28466 20710
rect 29269 20707 29335 20710
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 15745 20634 15811 20637
rect 17953 20634 18019 20637
rect 15745 20632 18019 20634
rect 15745 20576 15750 20632
rect 15806 20576 17958 20632
rect 18014 20576 18019 20632
rect 15745 20574 18019 20576
rect 15745 20571 15811 20574
rect 17953 20571 18019 20574
rect 0 20408 800 20528
rect 16665 20498 16731 20501
rect 18137 20498 18203 20501
rect 16665 20496 18203 20498
rect 16665 20440 16670 20496
rect 16726 20440 18142 20496
rect 18198 20440 18203 20496
rect 16665 20438 18203 20440
rect 16665 20435 16731 20438
rect 18137 20435 18203 20438
rect 49200 20408 50000 20528
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 0 19818 800 19848
rect 4061 19818 4127 19821
rect 0 19816 4127 19818
rect 0 19760 4066 19816
rect 4122 19760 4127 19816
rect 0 19758 4127 19760
rect 0 19728 800 19758
rect 4061 19755 4127 19758
rect 21449 19818 21515 19821
rect 22921 19818 22987 19821
rect 21449 19816 22987 19818
rect 21449 19760 21454 19816
rect 21510 19760 22926 19816
rect 22982 19760 22987 19816
rect 21449 19758 22987 19760
rect 21449 19755 21515 19758
rect 22921 19755 22987 19758
rect 48129 19818 48195 19821
rect 49200 19818 50000 19848
rect 48129 19816 50000 19818
rect 48129 19760 48134 19816
rect 48190 19760 50000 19816
rect 48129 19758 50000 19760
rect 48129 19755 48195 19758
rect 49200 19728 50000 19758
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 10961 19410 11027 19413
rect 12525 19410 12591 19413
rect 10961 19408 12591 19410
rect 10961 19352 10966 19408
rect 11022 19352 12530 19408
rect 12586 19352 12591 19408
rect 10961 19350 12591 19352
rect 10961 19347 11027 19350
rect 12525 19347 12591 19350
rect 19793 19410 19859 19413
rect 22461 19410 22527 19413
rect 19793 19408 22527 19410
rect 19793 19352 19798 19408
rect 19854 19352 22466 19408
rect 22522 19352 22527 19408
rect 19793 19350 22527 19352
rect 19793 19347 19859 19350
rect 22461 19347 22527 19350
rect 0 19138 800 19168
rect 2221 19138 2287 19141
rect 0 19136 2287 19138
rect 0 19080 2226 19136
rect 2282 19080 2287 19136
rect 0 19078 2287 19080
rect 0 19048 800 19078
rect 2221 19075 2287 19078
rect 47853 19138 47919 19141
rect 49200 19138 50000 19168
rect 47853 19136 50000 19138
rect 47853 19080 47858 19136
rect 47914 19080 50000 19136
rect 47853 19078 50000 19080
rect 47853 19075 47919 19078
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 49200 19048 50000 19078
rect 34928 19007 35248 19008
rect 23790 18804 23796 18868
rect 23860 18866 23866 18868
rect 24025 18866 24091 18869
rect 23860 18864 24091 18866
rect 23860 18808 24030 18864
rect 24086 18808 24091 18864
rect 23860 18806 24091 18808
rect 23860 18804 23866 18806
rect 24025 18803 24091 18806
rect 21541 18730 21607 18733
rect 26417 18730 26483 18733
rect 21541 18728 26483 18730
rect 21541 18672 21546 18728
rect 21602 18672 26422 18728
rect 26478 18672 26483 18728
rect 21541 18670 26483 18672
rect 21541 18667 21607 18670
rect 26417 18667 26483 18670
rect 22921 18594 22987 18597
rect 24945 18594 25011 18597
rect 32121 18594 32187 18597
rect 22921 18592 25011 18594
rect 22921 18536 22926 18592
rect 22982 18536 24950 18592
rect 25006 18536 25011 18592
rect 22921 18534 25011 18536
rect 22921 18531 22987 18534
rect 24945 18531 25011 18534
rect 32078 18592 32187 18594
rect 32078 18536 32126 18592
rect 32182 18536 32187 18592
rect 32078 18531 32187 18536
rect 19568 18528 19888 18529
rect 0 18458 800 18488
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 4061 18458 4127 18461
rect 0 18456 4127 18458
rect 0 18400 4066 18456
rect 4122 18400 4127 18456
rect 0 18398 4127 18400
rect 0 18368 800 18398
rect 4061 18395 4127 18398
rect 24209 18458 24275 18461
rect 31109 18458 31175 18461
rect 24209 18456 31175 18458
rect 24209 18400 24214 18456
rect 24270 18400 31114 18456
rect 31170 18400 31175 18456
rect 24209 18398 31175 18400
rect 24209 18395 24275 18398
rect 31109 18395 31175 18398
rect 32078 18325 32138 18531
rect 49200 18368 50000 18488
rect 21725 18322 21791 18325
rect 26049 18322 26115 18325
rect 27705 18322 27771 18325
rect 21725 18320 27771 18322
rect 21725 18264 21730 18320
rect 21786 18264 26054 18320
rect 26110 18264 27710 18320
rect 27766 18264 27771 18320
rect 21725 18262 27771 18264
rect 21725 18259 21791 18262
rect 26049 18259 26115 18262
rect 27705 18259 27771 18262
rect 32029 18320 32138 18325
rect 32029 18264 32034 18320
rect 32090 18264 32138 18320
rect 32029 18262 32138 18264
rect 32029 18259 32095 18262
rect 24853 18186 24919 18189
rect 26141 18186 26207 18189
rect 24853 18184 26207 18186
rect 24853 18128 24858 18184
rect 24914 18128 26146 18184
rect 26202 18128 26207 18184
rect 24853 18126 26207 18128
rect 24853 18123 24919 18126
rect 26141 18123 26207 18126
rect 21265 18050 21331 18053
rect 27521 18050 27587 18053
rect 21265 18048 27587 18050
rect 21265 17992 21270 18048
rect 21326 17992 27526 18048
rect 27582 17992 27587 18048
rect 21265 17990 27587 17992
rect 21265 17987 21331 17990
rect 27521 17987 27587 17990
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 0 17778 800 17808
rect 2773 17778 2839 17781
rect 28625 17780 28691 17781
rect 28574 17778 28580 17780
rect 0 17776 2839 17778
rect 0 17720 2778 17776
rect 2834 17720 2839 17776
rect 0 17718 2839 17720
rect 28534 17718 28580 17778
rect 28644 17776 28691 17780
rect 28686 17720 28691 17776
rect 0 17688 800 17718
rect 2773 17715 2839 17718
rect 28574 17716 28580 17718
rect 28644 17716 28691 17720
rect 28625 17715 28691 17716
rect 46841 17778 46907 17781
rect 49200 17778 50000 17808
rect 46841 17776 50000 17778
rect 46841 17720 46846 17776
rect 46902 17720 50000 17776
rect 46841 17718 50000 17720
rect 46841 17715 46907 17718
rect 49200 17688 50000 17718
rect 24945 17642 25011 17645
rect 26233 17642 26299 17645
rect 24945 17640 26299 17642
rect 24945 17584 24950 17640
rect 25006 17584 26238 17640
rect 26294 17584 26299 17640
rect 24945 17582 26299 17584
rect 24945 17579 25011 17582
rect 26233 17579 26299 17582
rect 23381 17506 23447 17509
rect 26969 17506 27035 17509
rect 23381 17504 27035 17506
rect 23381 17448 23386 17504
rect 23442 17448 26974 17504
rect 27030 17448 27035 17504
rect 23381 17446 27035 17448
rect 23381 17443 23447 17446
rect 26969 17443 27035 17446
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 19885 17234 19951 17237
rect 20989 17234 21055 17237
rect 19885 17232 21055 17234
rect 19885 17176 19890 17232
rect 19946 17176 20994 17232
rect 21050 17176 21055 17232
rect 19885 17174 21055 17176
rect 19885 17171 19951 17174
rect 20989 17171 21055 17174
rect 25589 17234 25655 17237
rect 27061 17234 27127 17237
rect 25589 17232 27127 17234
rect 25589 17176 25594 17232
rect 25650 17176 27066 17232
rect 27122 17176 27127 17232
rect 25589 17174 27127 17176
rect 25589 17171 25655 17174
rect 27061 17171 27127 17174
rect 28993 17234 29059 17237
rect 35249 17234 35315 17237
rect 28993 17232 35315 17234
rect 28993 17176 28998 17232
rect 29054 17176 35254 17232
rect 35310 17176 35315 17232
rect 28993 17174 35315 17176
rect 28993 17171 29059 17174
rect 35249 17171 35315 17174
rect 0 17098 800 17128
rect 1853 17098 1919 17101
rect 0 17096 1919 17098
rect 0 17040 1858 17096
rect 1914 17040 1919 17096
rect 0 17038 1919 17040
rect 0 17008 800 17038
rect 1853 17035 1919 17038
rect 23013 17098 23079 17101
rect 24393 17098 24459 17101
rect 23013 17096 24459 17098
rect 23013 17040 23018 17096
rect 23074 17040 24398 17096
rect 24454 17040 24459 17096
rect 23013 17038 24459 17040
rect 23013 17035 23079 17038
rect 24393 17035 24459 17038
rect 28993 17098 29059 17101
rect 29453 17098 29519 17101
rect 28993 17096 29519 17098
rect 28993 17040 28998 17096
rect 29054 17040 29458 17096
rect 29514 17040 29519 17096
rect 28993 17038 29519 17040
rect 28993 17035 29059 17038
rect 29453 17035 29519 17038
rect 31017 17098 31083 17101
rect 34513 17098 34579 17101
rect 35617 17098 35683 17101
rect 31017 17096 35683 17098
rect 31017 17040 31022 17096
rect 31078 17040 34518 17096
rect 34574 17040 35622 17096
rect 35678 17040 35683 17096
rect 31017 17038 35683 17040
rect 31017 17035 31083 17038
rect 34513 17035 34579 17038
rect 35617 17035 35683 17038
rect 48129 17098 48195 17101
rect 49200 17098 50000 17128
rect 48129 17096 50000 17098
rect 48129 17040 48134 17096
rect 48190 17040 50000 17096
rect 48129 17038 50000 17040
rect 48129 17035 48195 17038
rect 49200 17008 50000 17038
rect 24025 16962 24091 16965
rect 24025 16960 24778 16962
rect 24025 16904 24030 16960
rect 24086 16904 24778 16960
rect 24025 16902 24778 16904
rect 24025 16899 24091 16902
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 23381 16826 23447 16829
rect 24209 16826 24275 16829
rect 24485 16826 24551 16829
rect 23381 16824 24551 16826
rect 23381 16768 23386 16824
rect 23442 16768 24214 16824
rect 24270 16768 24490 16824
rect 24546 16768 24551 16824
rect 23381 16766 24551 16768
rect 24718 16826 24778 16902
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 24853 16826 24919 16829
rect 24718 16824 24919 16826
rect 24718 16768 24858 16824
rect 24914 16768 24919 16824
rect 24718 16766 24919 16768
rect 23381 16763 23447 16766
rect 24209 16763 24275 16766
rect 24485 16763 24551 16766
rect 24853 16763 24919 16766
rect 23790 16628 23796 16692
rect 23860 16690 23866 16692
rect 27981 16690 28047 16693
rect 23860 16688 28047 16690
rect 23860 16632 27986 16688
rect 28042 16632 28047 16688
rect 23860 16630 28047 16632
rect 23860 16628 23866 16630
rect 27981 16627 28047 16630
rect 24393 16554 24459 16557
rect 27153 16554 27219 16557
rect 24393 16552 27219 16554
rect 24393 16496 24398 16552
rect 24454 16496 27158 16552
rect 27214 16496 27219 16552
rect 24393 16494 27219 16496
rect 24393 16491 24459 16494
rect 27153 16491 27219 16494
rect 0 16418 800 16448
rect 2773 16418 2839 16421
rect 0 16416 2839 16418
rect 0 16360 2778 16416
rect 2834 16360 2839 16416
rect 0 16358 2839 16360
rect 0 16328 800 16358
rect 2773 16355 2839 16358
rect 24485 16418 24551 16421
rect 25865 16418 25931 16421
rect 24485 16416 25931 16418
rect 24485 16360 24490 16416
rect 24546 16360 25870 16416
rect 25926 16360 25931 16416
rect 24485 16358 25931 16360
rect 24485 16355 24551 16358
rect 25865 16355 25931 16358
rect 48129 16418 48195 16421
rect 49200 16418 50000 16448
rect 48129 16416 50000 16418
rect 48129 16360 48134 16416
rect 48190 16360 50000 16416
rect 48129 16358 50000 16360
rect 48129 16355 48195 16358
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 49200 16328 50000 16358
rect 19568 16287 19888 16288
rect 4208 15808 4528 15809
rect 0 15648 800 15768
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 49200 15648 50000 15768
rect 27797 15330 27863 15333
rect 30925 15330 30991 15333
rect 27797 15328 30991 15330
rect 27797 15272 27802 15328
rect 27858 15272 30930 15328
rect 30986 15272 30991 15328
rect 27797 15270 30991 15272
rect 27797 15267 27863 15270
rect 30925 15267 30991 15270
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 32581 15196 32647 15197
rect 32581 15194 32628 15196
rect 32536 15192 32628 15194
rect 32536 15136 32586 15192
rect 32536 15134 32628 15136
rect 32581 15132 32628 15134
rect 32692 15132 32698 15196
rect 32581 15131 32647 15132
rect 0 14968 800 15088
rect 29177 15058 29243 15061
rect 30281 15058 30347 15061
rect 29177 15056 30347 15058
rect 29177 15000 29182 15056
rect 29238 15000 30286 15056
rect 30342 15000 30347 15056
rect 29177 14998 30347 15000
rect 29177 14995 29243 14998
rect 30281 14995 30347 14998
rect 47945 15058 48011 15061
rect 49200 15058 50000 15088
rect 47945 15056 50000 15058
rect 47945 15000 47950 15056
rect 48006 15000 50000 15056
rect 47945 14998 50000 15000
rect 47945 14995 48011 14998
rect 49200 14968 50000 14998
rect 32489 14922 32555 14925
rect 33409 14922 33475 14925
rect 32489 14920 33475 14922
rect 32489 14864 32494 14920
rect 32550 14864 33414 14920
rect 33470 14864 33475 14920
rect 32489 14862 33475 14864
rect 32489 14859 32555 14862
rect 33409 14859 33475 14862
rect 26785 14786 26851 14789
rect 34789 14786 34855 14789
rect 26785 14784 34855 14786
rect 26785 14728 26790 14784
rect 26846 14728 34794 14784
rect 34850 14728 34855 14784
rect 26785 14726 34855 14728
rect 26785 14723 26851 14726
rect 34789 14723 34855 14726
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 29729 14514 29795 14517
rect 35525 14514 35591 14517
rect 29729 14512 35591 14514
rect 29729 14456 29734 14512
rect 29790 14456 35530 14512
rect 35586 14456 35591 14512
rect 29729 14454 35591 14456
rect 29729 14451 29795 14454
rect 35525 14451 35591 14454
rect 0 14288 800 14408
rect 35341 14378 35407 14381
rect 36997 14378 37063 14381
rect 35341 14376 37063 14378
rect 35341 14320 35346 14376
rect 35402 14320 37002 14376
rect 37058 14320 37063 14376
rect 35341 14318 37063 14320
rect 35341 14315 35407 14318
rect 36997 14315 37063 14318
rect 48129 14378 48195 14381
rect 49200 14378 50000 14408
rect 48129 14376 50000 14378
rect 48129 14320 48134 14376
rect 48190 14320 50000 14376
rect 48129 14318 50000 14320
rect 48129 14315 48195 14318
rect 49200 14288 50000 14318
rect 27245 14242 27311 14245
rect 27889 14242 27955 14245
rect 27245 14240 27955 14242
rect 27245 14184 27250 14240
rect 27306 14184 27894 14240
rect 27950 14184 27955 14240
rect 27245 14182 27955 14184
rect 27245 14179 27311 14182
rect 27889 14179 27955 14182
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 28349 13970 28415 13973
rect 28574 13970 28580 13972
rect 28349 13968 28580 13970
rect 28349 13912 28354 13968
rect 28410 13912 28580 13968
rect 28349 13910 28580 13912
rect 28349 13907 28415 13910
rect 28574 13908 28580 13910
rect 28644 13908 28650 13972
rect 32673 13836 32739 13837
rect 32622 13834 32628 13836
rect 32582 13774 32628 13834
rect 32692 13832 32739 13836
rect 32734 13776 32739 13832
rect 32622 13772 32628 13774
rect 32692 13772 32739 13776
rect 32673 13771 32739 13772
rect 0 13698 800 13728
rect 2773 13698 2839 13701
rect 0 13696 2839 13698
rect 0 13640 2778 13696
rect 2834 13640 2839 13696
rect 0 13638 2839 13640
rect 0 13608 800 13638
rect 2773 13635 2839 13638
rect 47853 13698 47919 13701
rect 49200 13698 50000 13728
rect 47853 13696 50000 13698
rect 47853 13640 47858 13696
rect 47914 13640 50000 13696
rect 47853 13638 50000 13640
rect 47853 13635 47919 13638
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 49200 13608 50000 13638
rect 34928 13567 35248 13568
rect 20110 13228 20116 13292
rect 20180 13290 20186 13292
rect 20253 13290 20319 13293
rect 20180 13288 20319 13290
rect 20180 13232 20258 13288
rect 20314 13232 20319 13288
rect 20180 13230 20319 13232
rect 20180 13228 20186 13230
rect 20253 13227 20319 13230
rect 19568 13088 19888 13089
rect 0 13018 800 13048
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 4061 13018 4127 13021
rect 0 13016 4127 13018
rect 0 12960 4066 13016
rect 4122 12960 4127 13016
rect 0 12958 4127 12960
rect 0 12928 800 12958
rect 4061 12955 4127 12958
rect 46749 13018 46815 13021
rect 49200 13018 50000 13048
rect 46749 13016 50000 13018
rect 46749 12960 46754 13016
rect 46810 12960 50000 13016
rect 46749 12958 50000 12960
rect 46749 12955 46815 12958
rect 49200 12928 50000 12958
rect 23565 12746 23631 12749
rect 25129 12746 25195 12749
rect 23565 12744 25195 12746
rect 23565 12688 23570 12744
rect 23626 12688 25134 12744
rect 25190 12688 25195 12744
rect 23565 12686 25195 12688
rect 23565 12683 23631 12686
rect 25129 12683 25195 12686
rect 20161 12610 20227 12613
rect 20345 12610 20411 12613
rect 20161 12608 20411 12610
rect 20161 12552 20166 12608
rect 20222 12552 20350 12608
rect 20406 12552 20411 12608
rect 20161 12550 20411 12552
rect 20161 12547 20227 12550
rect 20345 12547 20411 12550
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 0 12338 800 12368
rect 1393 12338 1459 12341
rect 0 12336 1459 12338
rect 0 12280 1398 12336
rect 1454 12280 1459 12336
rect 0 12278 1459 12280
rect 0 12248 800 12278
rect 1393 12275 1459 12278
rect 23790 12276 23796 12340
rect 23860 12338 23866 12340
rect 23933 12338 23999 12341
rect 23860 12336 23999 12338
rect 23860 12280 23938 12336
rect 23994 12280 23999 12336
rect 23860 12278 23999 12280
rect 23860 12276 23866 12278
rect 23933 12275 23999 12278
rect 46841 12338 46907 12341
rect 49200 12338 50000 12368
rect 46841 12336 50000 12338
rect 46841 12280 46846 12336
rect 46902 12280 50000 12336
rect 46841 12278 50000 12280
rect 46841 12275 46907 12278
rect 49200 12248 50000 12278
rect 28533 12202 28599 12205
rect 28809 12202 28875 12205
rect 28533 12200 28875 12202
rect 28533 12144 28538 12200
rect 28594 12144 28814 12200
rect 28870 12144 28875 12200
rect 28533 12142 28875 12144
rect 28533 12139 28599 12142
rect 28809 12139 28875 12142
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 0 11568 800 11688
rect 49200 11568 50000 11688
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 19425 11114 19491 11117
rect 24025 11114 24091 11117
rect 19425 11112 24091 11114
rect 19425 11056 19430 11112
rect 19486 11056 24030 11112
rect 24086 11056 24091 11112
rect 19425 11054 24091 11056
rect 19425 11051 19491 11054
rect 24025 11051 24091 11054
rect 0 10978 800 11008
rect 1853 10978 1919 10981
rect 0 10976 1919 10978
rect 0 10920 1858 10976
rect 1914 10920 1919 10976
rect 0 10918 1919 10920
rect 0 10888 800 10918
rect 1853 10915 1919 10918
rect 48129 10978 48195 10981
rect 49200 10978 50000 11008
rect 48129 10976 50000 10978
rect 48129 10920 48134 10976
rect 48190 10920 50000 10976
rect 48129 10918 50000 10920
rect 48129 10915 48195 10918
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 49200 10888 50000 10918
rect 19568 10847 19888 10848
rect 19425 10434 19491 10437
rect 20110 10434 20116 10436
rect 19425 10432 20116 10434
rect 19425 10376 19430 10432
rect 19486 10376 20116 10432
rect 19425 10374 20116 10376
rect 19425 10371 19491 10374
rect 20110 10372 20116 10374
rect 20180 10372 20186 10436
rect 4208 10368 4528 10369
rect 0 10298 800 10328
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 2773 10298 2839 10301
rect 0 10296 2839 10298
rect 0 10240 2778 10296
rect 2834 10240 2839 10296
rect 0 10238 2839 10240
rect 0 10208 800 10238
rect 2773 10235 2839 10238
rect 47761 10298 47827 10301
rect 49200 10298 50000 10328
rect 47761 10296 50000 10298
rect 47761 10240 47766 10296
rect 47822 10240 50000 10296
rect 47761 10238 50000 10240
rect 47761 10235 47827 10238
rect 49200 10208 50000 10238
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 0 9618 800 9648
rect 2773 9618 2839 9621
rect 0 9616 2839 9618
rect 0 9560 2778 9616
rect 2834 9560 2839 9616
rect 0 9558 2839 9560
rect 0 9528 800 9558
rect 2773 9555 2839 9558
rect 46841 9618 46907 9621
rect 49200 9618 50000 9648
rect 46841 9616 50000 9618
rect 46841 9560 46846 9616
rect 46902 9560 50000 9616
rect 46841 9558 50000 9560
rect 46841 9555 46907 9558
rect 49200 9528 50000 9558
rect 28993 9482 29059 9485
rect 33133 9482 33199 9485
rect 28993 9480 33199 9482
rect 28993 9424 28998 9480
rect 29054 9424 33138 9480
rect 33194 9424 33199 9480
rect 28993 9422 33199 9424
rect 28993 9419 29059 9422
rect 33133 9419 33199 9422
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 27797 9074 27863 9077
rect 27797 9072 27906 9074
rect 27797 9016 27802 9072
rect 27858 9016 27906 9072
rect 27797 9011 27906 9016
rect 0 8938 800 8968
rect 3417 8938 3483 8941
rect 0 8936 3483 8938
rect 0 8880 3422 8936
rect 3478 8880 3483 8936
rect 0 8878 3483 8880
rect 0 8848 800 8878
rect 3417 8875 3483 8878
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 27846 8397 27906 9011
rect 47945 8938 48011 8941
rect 49200 8938 50000 8968
rect 47945 8936 50000 8938
rect 47945 8880 47950 8936
rect 48006 8880 50000 8936
rect 47945 8878 50000 8880
rect 47945 8875 48011 8878
rect 49200 8848 50000 8878
rect 28257 8802 28323 8805
rect 28533 8802 28599 8805
rect 28257 8800 28599 8802
rect 28257 8744 28262 8800
rect 28318 8744 28538 8800
rect 28594 8744 28599 8800
rect 28257 8742 28599 8744
rect 28257 8739 28323 8742
rect 28533 8739 28599 8742
rect 18321 8394 18387 8397
rect 21081 8394 21147 8397
rect 18321 8392 21147 8394
rect 18321 8336 18326 8392
rect 18382 8336 21086 8392
rect 21142 8336 21147 8392
rect 18321 8334 21147 8336
rect 27846 8392 27955 8397
rect 27846 8336 27894 8392
rect 27950 8336 27955 8392
rect 27846 8334 27955 8336
rect 18321 8331 18387 8334
rect 21081 8331 21147 8334
rect 27889 8331 27955 8334
rect 0 8258 800 8288
rect 1853 8258 1919 8261
rect 0 8256 1919 8258
rect 0 8200 1858 8256
rect 1914 8200 1919 8256
rect 0 8198 1919 8200
rect 0 8168 800 8198
rect 1853 8195 1919 8198
rect 47853 8258 47919 8261
rect 49200 8258 50000 8288
rect 47853 8256 50000 8258
rect 47853 8200 47858 8256
rect 47914 8200 50000 8256
rect 47853 8198 50000 8200
rect 47853 8195 47919 8198
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 49200 8168 50000 8198
rect 34928 8127 35248 8128
rect 19568 7648 19888 7649
rect 0 7578 800 7608
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 1853 7578 1919 7581
rect 0 7576 1919 7578
rect 0 7520 1858 7576
rect 1914 7520 1919 7576
rect 0 7518 1919 7520
rect 0 7488 800 7518
rect 1853 7515 1919 7518
rect 48129 7578 48195 7581
rect 49200 7578 50000 7608
rect 48129 7576 50000 7578
rect 48129 7520 48134 7576
rect 48190 7520 50000 7576
rect 48129 7518 50000 7520
rect 48129 7515 48195 7518
rect 49200 7488 50000 7518
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 0 6898 800 6928
rect 2773 6898 2839 6901
rect 0 6896 2839 6898
rect 0 6840 2778 6896
rect 2834 6840 2839 6896
rect 0 6838 2839 6840
rect 0 6808 800 6838
rect 2773 6835 2839 6838
rect 46841 6898 46907 6901
rect 49200 6898 50000 6928
rect 46841 6896 50000 6898
rect 46841 6840 46846 6896
rect 46902 6840 50000 6896
rect 46841 6838 50000 6840
rect 46841 6835 46907 6838
rect 49200 6808 50000 6838
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 0 6218 800 6248
rect 3417 6218 3483 6221
rect 0 6216 3483 6218
rect 0 6160 3422 6216
rect 3478 6160 3483 6216
rect 0 6158 3483 6160
rect 0 6128 800 6158
rect 3417 6155 3483 6158
rect 46749 6218 46815 6221
rect 49200 6218 50000 6248
rect 46749 6216 50000 6218
rect 46749 6160 46754 6216
rect 46810 6160 50000 6216
rect 46749 6158 50000 6160
rect 46749 6155 46815 6158
rect 49200 6128 50000 6158
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 0 5538 800 5568
rect 2773 5538 2839 5541
rect 0 5536 2839 5538
rect 0 5480 2778 5536
rect 2834 5480 2839 5536
rect 0 5478 2839 5480
rect 0 5448 800 5478
rect 2773 5475 2839 5478
rect 47853 5538 47919 5541
rect 49200 5538 50000 5568
rect 47853 5536 50000 5538
rect 47853 5480 47858 5536
rect 47914 5480 50000 5536
rect 47853 5478 50000 5480
rect 47853 5475 47919 5478
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 49200 5448 50000 5478
rect 19568 5407 19888 5408
rect 4208 4928 4528 4929
rect 0 4858 800 4888
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 2773 4858 2839 4861
rect 0 4856 2839 4858
rect 0 4800 2778 4856
rect 2834 4800 2839 4856
rect 0 4798 2839 4800
rect 0 4768 800 4798
rect 2773 4795 2839 4798
rect 48129 4858 48195 4861
rect 49200 4858 50000 4888
rect 48129 4856 50000 4858
rect 48129 4800 48134 4856
rect 48190 4800 50000 4856
rect 48129 4798 50000 4800
rect 48129 4795 48195 4798
rect 49200 4768 50000 4798
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 0 4178 800 4208
rect 3417 4178 3483 4181
rect 0 4176 3483 4178
rect 0 4120 3422 4176
rect 3478 4120 3483 4176
rect 0 4118 3483 4120
rect 0 4088 800 4118
rect 3417 4115 3483 4118
rect 46841 4178 46907 4181
rect 49200 4178 50000 4208
rect 46841 4176 50000 4178
rect 46841 4120 46846 4176
rect 46902 4120 50000 4176
rect 46841 4118 50000 4120
rect 46841 4115 46907 4118
rect 49200 4088 50000 4118
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 0 3498 800 3528
rect 1853 3498 1919 3501
rect 0 3496 1919 3498
rect 0 3440 1858 3496
rect 1914 3440 1919 3496
rect 0 3438 1919 3440
rect 0 3408 800 3438
rect 1853 3435 1919 3438
rect 46197 3498 46263 3501
rect 49200 3498 50000 3528
rect 46197 3496 50000 3498
rect 46197 3440 46202 3496
rect 46258 3440 50000 3496
rect 46197 3438 50000 3440
rect 46197 3435 46263 3438
rect 49200 3408 50000 3438
rect 12157 3362 12223 3365
rect 12617 3362 12683 3365
rect 12157 3360 12683 3362
rect 12157 3304 12162 3360
rect 12218 3304 12622 3360
rect 12678 3304 12683 3360
rect 12157 3302 12683 3304
rect 12157 3299 12223 3302
rect 12617 3299 12683 3302
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 0 2728 800 2848
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 49200 2728 50000 2848
rect 34928 2687 35248 2688
rect 4797 2546 4863 2549
rect 28390 2546 28396 2548
rect 4797 2544 28396 2546
rect 4797 2488 4802 2544
rect 4858 2488 28396 2544
rect 4797 2486 28396 2488
rect 4797 2483 4863 2486
rect 28390 2484 28396 2486
rect 28460 2484 28466 2548
rect 2221 2410 2287 2413
rect 28758 2410 28764 2412
rect 2221 2408 28764 2410
rect 2221 2352 2226 2408
rect 2282 2352 28764 2408
rect 2221 2350 28764 2352
rect 2221 2347 2287 2350
rect 28758 2348 28764 2350
rect 28828 2348 28834 2412
rect 19568 2208 19888 2209
rect 0 2138 800 2168
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 3141 2138 3207 2141
rect 0 2136 3207 2138
rect 0 2080 3146 2136
rect 3202 2080 3207 2136
rect 0 2078 3207 2080
rect 0 2048 800 2078
rect 3141 2075 3207 2078
rect 49200 2048 50000 2168
rect 0 1368 800 1488
rect 45829 1458 45895 1461
rect 49200 1458 50000 1488
rect 45829 1456 50000 1458
rect 45829 1400 45834 1456
rect 45890 1400 50000 1456
rect 45829 1398 50000 1400
rect 45829 1395 45895 1398
rect 49200 1368 50000 1398
rect 0 778 800 808
rect 1853 778 1919 781
rect 0 776 1919 778
rect 0 720 1858 776
rect 1914 720 1919 776
rect 0 718 1919 720
rect 0 688 800 718
rect 1853 715 1919 718
rect 47761 778 47827 781
rect 49200 778 50000 808
rect 47761 776 50000 778
rect 47761 720 47766 776
rect 47822 720 50000 776
rect 47761 718 50000 720
rect 47761 715 47827 718
rect 49200 688 50000 718
rect 46749 98 46815 101
rect 49200 98 50000 128
rect 46749 96 50000 98
rect 46749 40 46754 96
rect 46810 40 50000 96
rect 46749 38 50000 40
rect 46749 35 46815 38
rect 49200 8 50000 38
<< via3 >>
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 28764 21992 28828 21996
rect 28764 21936 28814 21992
rect 28814 21936 28828 21992
rect 28764 21932 28828 21936
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 28396 20708 28460 20772
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 23796 18804 23860 18868
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 28580 17776 28644 17780
rect 28580 17720 28630 17776
rect 28630 17720 28644 17776
rect 28580 17716 28644 17720
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 23796 16628 23860 16692
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 32628 15192 32692 15196
rect 32628 15136 32642 15192
rect 32642 15136 32692 15192
rect 32628 15132 32692 15136
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 28580 13908 28644 13972
rect 32628 13832 32692 13836
rect 32628 13776 32678 13832
rect 32678 13776 32692 13832
rect 32628 13772 32692 13776
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 20116 13228 20180 13292
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 23796 12276 23860 12340
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 20116 10372 20180 10436
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 28396 2484 28460 2548
rect 28764 2348 28828 2412
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 49536 4528 49552
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 48992 19888 49552
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 34928 49536 35248 49552
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 28763 21996 28829 21997
rect 28763 21932 28764 21996
rect 28828 21932 28829 21996
rect 28763 21931 28829 21932
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 28395 20772 28461 20773
rect 28395 20708 28396 20772
rect 28460 20708 28461 20772
rect 28395 20707 28461 20708
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 23795 18868 23861 18869
rect 23795 18804 23796 18868
rect 23860 18804 23861 18868
rect 23795 18803 23861 18804
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 23798 16693 23858 18803
rect 23795 16692 23861 16693
rect 23795 16628 23796 16692
rect 23860 16628 23861 16692
rect 23795 16627 23861 16628
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 20115 13292 20181 13293
rect 20115 13228 20116 13292
rect 20180 13228 20181 13292
rect 20115 13227 20181 13228
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 20118 10437 20178 13227
rect 23798 12341 23858 16627
rect 23795 12340 23861 12341
rect 23795 12276 23796 12340
rect 23860 12276 23861 12340
rect 23795 12275 23861 12276
rect 20115 10436 20181 10437
rect 20115 10372 20116 10436
rect 20180 10372 20181 10436
rect 20115 10371 20181 10372
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 28398 2549 28458 20707
rect 28579 17780 28645 17781
rect 28579 17716 28580 17780
rect 28644 17716 28645 17780
rect 28579 17715 28645 17716
rect 28582 13973 28642 17715
rect 28579 13972 28645 13973
rect 28579 13908 28580 13972
rect 28644 13908 28645 13972
rect 28579 13907 28645 13908
rect 28395 2548 28461 2549
rect 28395 2484 28396 2548
rect 28460 2484 28461 2548
rect 28395 2483 28461 2484
rect 28766 2413 28826 21931
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 32627 15196 32693 15197
rect 32627 15132 32628 15196
rect 32692 15132 32693 15196
rect 32627 15131 32693 15132
rect 32630 13837 32690 15131
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 32627 13836 32693 13837
rect 32627 13772 32628 13836
rect 32692 13772 32693 13836
rect 32627 13771 32693 13772
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 28763 2412 28829 2413
rect 28763 2348 28764 2412
rect 28828 2348 28829 2412
rect 28763 2347 28829 2348
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28980 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1644511149
transform -1 0 30820 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1644511149
transform 1 0 30452 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1644511149
transform 1 0 17112 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1644511149
transform -1 0 17848 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1644511149
transform 1 0 17480 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1644511149
transform 1 0 11960 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1644511149
transform 1 0 30728 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1644511149
transform 1 0 30452 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13
timestamp 1644511149
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37
timestamp 1644511149
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_42 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4968 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79
timestamp 1644511149
transform 1 0 8372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1644511149
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_95
timestamp 1644511149
transform 1 0 9844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_103
timestamp 1644511149
transform 1 0 10580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1644511149
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_124
timestamp 1644511149
transform 1 0 12512 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_131
timestamp 1644511149
transform 1 0 13156 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1644511149
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_162
timestamp 1644511149
transform 1 0 16008 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177
timestamp 1644511149
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_182
timestamp 1644511149
transform 1 0 17848 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1644511149
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_205
timestamp 1644511149
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_210
timestamp 1644511149
transform 1 0 20424 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1644511149
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_246
timestamp 1644511149
transform 1 0 23736 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_261
timestamp 1644511149
transform 1 0 25116 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_266
timestamp 1644511149
transform 1 0 25576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_274
timestamp 1644511149
transform 1 0 26312 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_287
timestamp 1644511149
transform 1 0 27508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_295
timestamp 1644511149
transform 1 0 28244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1644511149
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_330
timestamp 1644511149
transform 1 0 31464 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_345
timestamp 1644511149
transform 1 0 32844 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_350
timestamp 1644511149
transform 1 0 33304 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_360
timestamp 1644511149
transform 1 0 34224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_373
timestamp 1644511149
transform 1 0 35420 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_385
timestamp 1644511149
transform 1 0 36524 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1644511149
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_393
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_405
timestamp 1644511149
transform 1 0 38364 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_416
timestamp 1644511149
transform 1 0 39376 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_442
timestamp 1644511149
transform 1 0 41768 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_470
timestamp 1644511149
transform 1 0 44344 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_498
timestamp 1644511149
transform 1 0 46920 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_505
timestamp 1644511149
transform 1 0 47564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_512
timestamp 1644511149
transform 1 0 48208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_9
timestamp 1644511149
transform 1 0 1932 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_13
timestamp 1644511149
transform 1 0 2300 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_25
timestamp 1644511149
transform 1 0 3404 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1644511149
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_78
timestamp 1644511149
transform 1 0 8280 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_92
timestamp 1644511149
transform 1 0 9568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_100
timestamp 1644511149
transform 1 0 10304 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_142
timestamp 1644511149
transform 1 0 14168 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_150
timestamp 1644511149
transform 1 0 14904 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_157
timestamp 1644511149
transform 1 0 15548 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1644511149
transform 1 0 17756 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_204
timestamp 1644511149
transform 1 0 19872 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_211
timestamp 1644511149
transform 1 0 20516 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_218
timestamp 1644511149
transform 1 0 21160 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_233
timestamp 1644511149
transform 1 0 22540 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_238
timestamp 1644511149
transform 1 0 23000 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_263
timestamp 1644511149
transform 1 0 25300 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_272
timestamp 1644511149
transform 1 0 26128 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_284
timestamp 1644511149
transform 1 0 27232 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_296
timestamp 1644511149
transform 1 0 28336 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_308
timestamp 1644511149
transform 1 0 29440 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_332
timestamp 1644511149
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_359
timestamp 1644511149
transform 1 0 34132 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_371
timestamp 1644511149
transform 1 0 35236 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_386
timestamp 1644511149
transform 1 0 36616 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_405
timestamp 1644511149
transform 1 0 38364 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_413
timestamp 1644511149
transform 1 0 39100 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_419
timestamp 1644511149
transform 1 0 39652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_444
timestamp 1644511149
transform 1 0 41952 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_452
timestamp 1644511149
transform 1 0 42688 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_462
timestamp 1644511149
transform 1 0 43608 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_487
timestamp 1644511149
transform 1 0 45908 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_495
timestamp 1644511149
transform 1 0 46644 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1644511149
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_505
timestamp 1644511149
transform 1 0 47564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_512
timestamp 1644511149
transform 1 0 48208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1644511149
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_50
timestamp 1644511149
transform 1 0 5704 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_57
timestamp 1644511149
transform 1 0 6348 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_64
timestamp 1644511149
transform 1 0 6992 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_68
timestamp 1644511149
transform 1 0 7360 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_72
timestamp 1644511149
transform 1 0 7728 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_91
timestamp 1644511149
transform 1 0 9476 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_103
timestamp 1644511149
transform 1 0 10580 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_110
timestamp 1644511149
transform 1 0 11224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_135
timestamp 1644511149
transform 1 0 13524 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1644511149
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_144
timestamp 1644511149
transform 1 0 14352 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_171
timestamp 1644511149
transform 1 0 16836 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_183
timestamp 1644511149
transform 1 0 17940 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1644511149
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_205
timestamp 1644511149
transform 1 0 19964 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_227
timestamp 1644511149
transform 1 0 21988 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_239
timestamp 1644511149
transform 1 0 23092 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_246
timestamp 1644511149
transform 1 0 23736 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_265
timestamp 1644511149
transform 1 0 25484 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_289
timestamp 1644511149
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_304
timestamp 1644511149
transform 1 0 29072 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_312
timestamp 1644511149
transform 1 0 29808 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_319
timestamp 1644511149
transform 1 0 30452 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_348
timestamp 1644511149
transform 1 0 33120 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_360
timestamp 1644511149
transform 1 0 34224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_381
timestamp 1644511149
transform 1 0 36156 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_403
timestamp 1644511149
transform 1 0 38180 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_407
timestamp 1644511149
transform 1 0 38548 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_411
timestamp 1644511149
transform 1 0 38916 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1644511149
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_424
timestamp 1644511149
transform 1 0 40112 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_430
timestamp 1644511149
transform 1 0 40664 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_434
timestamp 1644511149
transform 1 0 41032 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_459
timestamp 1644511149
transform 1 0 43332 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_468
timestamp 1644511149
transform 1 0 44160 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_480
timestamp 1644511149
transform 1 0 45264 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_487
timestamp 1644511149
transform 1 0 45908 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_512
timestamp 1644511149
transform 1 0 48208 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7
timestamp 1644511149
transform 1 0 1748 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_11
timestamp 1644511149
transform 1 0 2116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_23
timestamp 1644511149
transform 1 0 3220 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_28
timestamp 1644511149
transform 1 0 3680 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_32
timestamp 1644511149
transform 1 0 4048 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_36
timestamp 1644511149
transform 1 0 4416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_43
timestamp 1644511149
transform 1 0 5060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1644511149
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_61
timestamp 1644511149
transform 1 0 6716 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_73
timestamp 1644511149
transform 1 0 7820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_85
timestamp 1644511149
transform 1 0 8924 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1644511149
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_134
timestamp 1644511149
transform 1 0 13432 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_141
timestamp 1644511149
transform 1 0 14076 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_156
timestamp 1644511149
transform 1 0 15456 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_181
timestamp 1644511149
transform 1 0 17756 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_187
timestamp 1644511149
transform 1 0 18308 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_199
timestamp 1644511149
transform 1 0 19412 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_208
timestamp 1644511149
transform 1 0 20240 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_212
timestamp 1644511149
transform 1 0 20608 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_216
timestamp 1644511149
transform 1 0 20976 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_237
timestamp 1644511149
transform 1 0 22908 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_244
timestamp 1644511149
transform 1 0 23552 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_256
timestamp 1644511149
transform 1 0 24656 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_268
timestamp 1644511149
transform 1 0 25760 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_274
timestamp 1644511149
transform 1 0 26312 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_311
timestamp 1644511149
transform 1 0 29716 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_315
timestamp 1644511149
transform 1 0 30084 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_323
timestamp 1644511149
transform 1 0 30820 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_327
timestamp 1644511149
transform 1 0 31188 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_340
timestamp 1644511149
transform 1 0 32384 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_347
timestamp 1644511149
transform 1 0 33028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_359
timestamp 1644511149
transform 1 0 34132 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_371
timestamp 1644511149
transform 1 0 35236 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_379
timestamp 1644511149
transform 1 0 35972 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_384
timestamp 1644511149
transform 1 0 36432 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_402
timestamp 1644511149
transform 1 0 38088 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_429
timestamp 1644511149
transform 1 0 40572 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_440
timestamp 1644511149
transform 1 0 41584 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_452
timestamp 1644511149
transform 1 0 42688 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_464
timestamp 1644511149
transform 1 0 43792 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_470
timestamp 1644511149
transform 1 0 44344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_477
timestamp 1644511149
transform 1 0 44988 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_489
timestamp 1644511149
transform 1 0 46092 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_500
timestamp 1644511149
transform 1 0 47104 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_505
timestamp 1644511149
transform 1 0 47564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_512
timestamp 1644511149
transform 1 0 48208 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1644511149
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_35
timestamp 1644511149
transform 1 0 4324 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_39
timestamp 1644511149
transform 1 0 4692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_51
timestamp 1644511149
transform 1 0 5796 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_63
timestamp 1644511149
transform 1 0 6900 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_75
timestamp 1644511149
transform 1 0 8004 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_109
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_118
timestamp 1644511149
transform 1 0 11960 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_125
timestamp 1644511149
transform 1 0 12604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_137
timestamp 1644511149
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1644511149
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_221
timestamp 1644511149
transform 1 0 21436 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_225
timestamp 1644511149
transform 1 0 21804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_231
timestamp 1644511149
transform 1 0 22356 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_243
timestamp 1644511149
transform 1 0 23460 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1644511149
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1644511149
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_327
timestamp 1644511149
transform 1 0 31188 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_331
timestamp 1644511149
transform 1 0 31556 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_343
timestamp 1644511149
transform 1 0 32660 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_355
timestamp 1644511149
transform 1 0 33764 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_401
timestamp 1644511149
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1644511149
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1644511149
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_424
timestamp 1644511149
transform 1 0 40112 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_431
timestamp 1644511149
transform 1 0 40756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_443
timestamp 1644511149
transform 1 0 41860 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_455
timestamp 1644511149
transform 1 0 42964 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_467
timestamp 1644511149
transform 1 0 44068 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1644511149
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_477
timestamp 1644511149
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_489
timestamp 1644511149
transform 1 0 46092 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_512
timestamp 1644511149
transform 1 0 48208 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_7
timestamp 1644511149
transform 1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_32
timestamp 1644511149
transform 1 0 4048 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_44
timestamp 1644511149
transform 1 0 5152 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_208
timestamp 1644511149
transform 1 0 20240 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_220
timestamp 1644511149
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_236
timestamp 1644511149
transform 1 0 22816 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_258
timestamp 1644511149
transform 1 0 24840 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_270
timestamp 1644511149
transform 1 0 25944 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_278
timestamp 1644511149
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1644511149
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_405
timestamp 1644511149
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_417
timestamp 1644511149
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_429
timestamp 1644511149
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1644511149
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1644511149
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_449
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_461
timestamp 1644511149
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_473
timestamp 1644511149
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_485
timestamp 1644511149
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_500
timestamp 1644511149
transform 1 0 47104 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_508
timestamp 1644511149
transform 1 0 47840 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_14
timestamp 1644511149
transform 1 0 2392 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_21
timestamp 1644511149
transform 1 0 3036 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1644511149
transform 1 0 4048 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1644511149
transform 1 0 5152 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1644511149
transform 1 0 6256 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1644511149
transform 1 0 7360 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp 1644511149
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_200
timestamp 1644511149
transform 1 0 19504 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_224
timestamp 1644511149
transform 1 0 21712 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_248
timestamp 1644511149
transform 1 0 23920 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1644511149
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1644511149
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_433
timestamp 1644511149
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_445
timestamp 1644511149
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_457
timestamp 1644511149
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1644511149
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1644511149
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_477
timestamp 1644511149
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_489
timestamp 1644511149
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_501
timestamp 1644511149
transform 1 0 47196 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_507
timestamp 1644511149
transform 1 0 47748 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_512
timestamp 1644511149
transform 1 0 48208 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_14
timestamp 1644511149
transform 1 0 2392 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_26
timestamp 1644511149
transform 1 0 3496 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_38
timestamp 1644511149
transform 1 0 4600 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_50
timestamp 1644511149
transform 1 0 5704 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_206
timestamp 1644511149
transform 1 0 20056 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_218
timestamp 1644511149
transform 1 0 21160 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_230
timestamp 1644511149
transform 1 0 22264 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_234
timestamp 1644511149
transform 1 0 22632 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_243
timestamp 1644511149
transform 1 0 23460 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_255
timestamp 1644511149
transform 1 0 24564 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_267
timestamp 1644511149
transform 1 0 25668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_285
timestamp 1644511149
transform 1 0 27324 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_302
timestamp 1644511149
transform 1 0 28888 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_314
timestamp 1644511149
transform 1 0 29992 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_326
timestamp 1644511149
transform 1 0 31096 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_334
timestamp 1644511149
transform 1 0 31832 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_342
timestamp 1644511149
transform 1 0 32568 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_354
timestamp 1644511149
transform 1 0 33672 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_366
timestamp 1644511149
transform 1 0 34776 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_378
timestamp 1644511149
transform 1 0 35880 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_390
timestamp 1644511149
transform 1 0 36984 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1644511149
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1644511149
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_461
timestamp 1644511149
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_473
timestamp 1644511149
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_485
timestamp 1644511149
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1644511149
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1644511149
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_505
timestamp 1644511149
transform 1 0 47564 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_513
timestamp 1644511149
transform 1 0 48300 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1644511149
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_185
timestamp 1644511149
transform 1 0 18124 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_190
timestamp 1644511149
transform 1 0 18584 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_205
timestamp 1644511149
transform 1 0 19964 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_224
timestamp 1644511149
transform 1 0 21712 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_232
timestamp 1644511149
transform 1 0 22448 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_239
timestamp 1644511149
transform 1 0 23092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_276
timestamp 1644511149
transform 1 0 26496 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_325
timestamp 1644511149
transform 1 0 31004 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_331
timestamp 1644511149
transform 1 0 31556 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_353
timestamp 1644511149
transform 1 0 33580 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_361
timestamp 1644511149
transform 1 0 34316 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_401
timestamp 1644511149
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1644511149
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1644511149
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_433
timestamp 1644511149
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_445
timestamp 1644511149
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_457
timestamp 1644511149
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1644511149
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1644511149
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_477
timestamp 1644511149
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_489
timestamp 1644511149
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_501
timestamp 1644511149
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_513
timestamp 1644511149
transform 1 0 48300 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7
timestamp 1644511149
transform 1 0 1748 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_11
timestamp 1644511149
transform 1 0 2116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_23
timestamp 1644511149
transform 1 0 3220 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_35
timestamp 1644511149
transform 1 0 4324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_47
timestamp 1644511149
transform 1 0 5428 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_173
timestamp 1644511149
transform 1 0 17020 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_190
timestamp 1644511149
transform 1 0 18584 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_202
timestamp 1644511149
transform 1 0 19688 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_211
timestamp 1644511149
transform 1 0 20516 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_218
timestamp 1644511149
transform 1 0 21160 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_259
timestamp 1644511149
transform 1 0 24932 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_267
timestamp 1644511149
transform 1 0 25668 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_276
timestamp 1644511149
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_290
timestamp 1644511149
transform 1 0 27784 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_303
timestamp 1644511149
transform 1 0 28980 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_316
timestamp 1644511149
transform 1 0 30176 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_332
timestamp 1644511149
transform 1 0 31648 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_340
timestamp 1644511149
transform 1 0 32384 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_344
timestamp 1644511149
transform 1 0 32752 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_366
timestamp 1644511149
transform 1 0 34776 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_378
timestamp 1644511149
transform 1 0 35880 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_390
timestamp 1644511149
transform 1 0 36984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_417
timestamp 1644511149
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_429
timestamp 1644511149
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1644511149
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1644511149
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_461
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_473
timestamp 1644511149
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_485
timestamp 1644511149
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1644511149
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1644511149
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_505
timestamp 1644511149
transform 1 0 47564 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_513
timestamp 1644511149
transform 1 0 48300 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_13
timestamp 1644511149
transform 1 0 2300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1644511149
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_173
timestamp 1644511149
transform 1 0 17020 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_180
timestamp 1644511149
transform 1 0 17664 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_192
timestamp 1644511149
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_202
timestamp 1644511149
transform 1 0 19688 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_235
timestamp 1644511149
transform 1 0 22724 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_248
timestamp 1644511149
transform 1 0 23920 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_262
timestamp 1644511149
transform 1 0 25208 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_266
timestamp 1644511149
transform 1 0 25576 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_288
timestamp 1644511149
transform 1 0 27600 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_299
timestamp 1644511149
transform 1 0 28612 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_343
timestamp 1644511149
transform 1 0 32660 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_352
timestamp 1644511149
transform 1 0 33488 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1644511149
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1644511149
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1644511149
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_457
timestamp 1644511149
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1644511149
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1644511149
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_477
timestamp 1644511149
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_489
timestamp 1644511149
transform 1 0 46092 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_512
timestamp 1644511149
transform 1 0 48208 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_13
timestamp 1644511149
transform 1 0 2300 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_25
timestamp 1644511149
transform 1 0 3404 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_37
timestamp 1644511149
transform 1 0 4508 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_49
timestamp 1644511149
transform 1 0 5612 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_185
timestamp 1644511149
transform 1 0 18124 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_194
timestamp 1644511149
transform 1 0 18952 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_214
timestamp 1644511149
transform 1 0 20792 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1644511149
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_241
timestamp 1644511149
transform 1 0 23276 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_246
timestamp 1644511149
transform 1 0 23736 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_253
timestamp 1644511149
transform 1 0 24380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_265
timestamp 1644511149
transform 1 0 25484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_277
timestamp 1644511149
transform 1 0 26588 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_290
timestamp 1644511149
transform 1 0 27784 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_299
timestamp 1644511149
transform 1 0 28612 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_303
timestamp 1644511149
transform 1 0 28980 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_310
timestamp 1644511149
transform 1 0 29624 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_322
timestamp 1644511149
transform 1 0 30728 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp 1644511149
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_356
timestamp 1644511149
transform 1 0 33856 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_368
timestamp 1644511149
transform 1 0 34960 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_380
timestamp 1644511149
transform 1 0 36064 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_417
timestamp 1644511149
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1644511149
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1644511149
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_449
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_461
timestamp 1644511149
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_473
timestamp 1644511149
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_485
timestamp 1644511149
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_500
timestamp 1644511149
transform 1 0 47104 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_505
timestamp 1644511149
transform 1 0 47564 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_512
timestamp 1644511149
transform 1 0 48208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_186
timestamp 1644511149
transform 1 0 18216 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1644511149
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_209
timestamp 1644511149
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_221
timestamp 1644511149
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_233
timestamp 1644511149
transform 1 0 22540 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_241
timestamp 1644511149
transform 1 0 23276 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_248
timestamp 1644511149
transform 1 0 23920 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_259
timestamp 1644511149
transform 1 0 24932 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_271
timestamp 1644511149
transform 1 0 26036 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_279
timestamp 1644511149
transform 1 0 26772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_284
timestamp 1644511149
transform 1 0 27232 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_294
timestamp 1644511149
transform 1 0 28152 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_303
timestamp 1644511149
transform 1 0 28980 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_313
timestamp 1644511149
transform 1 0 29900 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_330
timestamp 1644511149
transform 1 0 31464 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_346
timestamp 1644511149
transform 1 0 32936 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_353
timestamp 1644511149
transform 1 0 33580 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_361
timestamp 1644511149
transform 1 0 34316 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_445
timestamp 1644511149
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_457
timestamp 1644511149
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1644511149
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1644511149
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_477
timestamp 1644511149
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_489
timestamp 1644511149
transform 1 0 46092 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_495
timestamp 1644511149
transform 1 0 46644 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_499
timestamp 1644511149
transform 1 0 47012 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_507
timestamp 1644511149
transform 1 0 47748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_512
timestamp 1644511149
transform 1 0 48208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_28
timestamp 1644511149
transform 1 0 3680 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_40
timestamp 1644511149
transform 1 0 4784 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_52
timestamp 1644511149
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_177
timestamp 1644511149
transform 1 0 17388 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_200
timestamp 1644511149
transform 1 0 19504 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_212
timestamp 1644511149
transform 1 0 20608 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_245
timestamp 1644511149
transform 1 0 23644 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_259
timestamp 1644511149
transform 1 0 24932 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_269
timestamp 1644511149
transform 1 0 25852 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_277
timestamp 1644511149
transform 1 0 26588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_289
timestamp 1644511149
transform 1 0 27692 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_294
timestamp 1644511149
transform 1 0 28152 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_309
timestamp 1644511149
transform 1 0 29532 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_322
timestamp 1644511149
transform 1 0 30728 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_328
timestamp 1644511149
transform 1 0 31280 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_332
timestamp 1644511149
transform 1 0 31648 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_341
timestamp 1644511149
transform 1 0 32476 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_363
timestamp 1644511149
transform 1 0 34500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_375
timestamp 1644511149
transform 1 0 35604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_387
timestamp 1644511149
transform 1 0 36708 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_417
timestamp 1644511149
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_429
timestamp 1644511149
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1644511149
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1644511149
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_461
timestamp 1644511149
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_473
timestamp 1644511149
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_485
timestamp 1644511149
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1644511149
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1644511149
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_505
timestamp 1644511149
transform 1 0 47564 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_513
timestamp 1644511149
transform 1 0 48300 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 1644511149
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_202
timestamp 1644511149
transform 1 0 19688 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_212
timestamp 1644511149
transform 1 0 20608 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_232
timestamp 1644511149
transform 1 0 22448 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_238
timestamp 1644511149
transform 1 0 23000 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_248
timestamp 1644511149
transform 1 0 23920 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_273
timestamp 1644511149
transform 1 0 26220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_282
timestamp 1644511149
transform 1 0 27048 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_291
timestamp 1644511149
transform 1 0 27876 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_303
timestamp 1644511149
transform 1 0 28980 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1644511149
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_318
timestamp 1644511149
transform 1 0 30360 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_330
timestamp 1644511149
transform 1 0 31464 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_338
timestamp 1644511149
transform 1 0 32200 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_356
timestamp 1644511149
transform 1 0 33856 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1644511149
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1644511149
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_433
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_445
timestamp 1644511149
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_457
timestamp 1644511149
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1644511149
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1644511149
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_477
timestamp 1644511149
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_489
timestamp 1644511149
transform 1 0 46092 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_512
timestamp 1644511149
transform 1 0 48208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_7
timestamp 1644511149
transform 1 0 1748 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_14
timestamp 1644511149
transform 1 0 2392 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_21
timestamp 1644511149
transform 1 0 3036 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_33
timestamp 1644511149
transform 1 0 4140 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_45
timestamp 1644511149
transform 1 0 5244 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 1644511149
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_195
timestamp 1644511149
transform 1 0 19044 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1644511149
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_233
timestamp 1644511149
transform 1 0 22540 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_254
timestamp 1644511149
transform 1 0 24472 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_263
timestamp 1644511149
transform 1 0 25300 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_276
timestamp 1644511149
transform 1 0 26496 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_284
timestamp 1644511149
transform 1 0 27232 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_301
timestamp 1644511149
transform 1 0 28796 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_306
timestamp 1644511149
transform 1 0 29256 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_318
timestamp 1644511149
transform 1 0 30360 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_330
timestamp 1644511149
transform 1 0 31464 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_345
timestamp 1644511149
transform 1 0 32844 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_374
timestamp 1644511149
transform 1 0 35512 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_386
timestamp 1644511149
transform 1 0 36616 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_417
timestamp 1644511149
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_429
timestamp 1644511149
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1644511149
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1644511149
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_461
timestamp 1644511149
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_473
timestamp 1644511149
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_485
timestamp 1644511149
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1644511149
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1644511149
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_505
timestamp 1644511149
transform 1 0 47564 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_512
timestamp 1644511149
transform 1 0 48208 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_11
timestamp 1644511149
transform 1 0 2116 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_18
timestamp 1644511149
transform 1 0 2760 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1644511149
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_185
timestamp 1644511149
transform 1 0 18124 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1644511149
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_205
timestamp 1644511149
transform 1 0 19964 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_217
timestamp 1644511149
transform 1 0 21068 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_230
timestamp 1644511149
transform 1 0 22264 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_238
timestamp 1644511149
transform 1 0 23000 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_248
timestamp 1644511149
transform 1 0 23920 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_256
timestamp 1644511149
transform 1 0 24656 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_278
timestamp 1644511149
transform 1 0 26680 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_286
timestamp 1644511149
transform 1 0 27416 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_291
timestamp 1644511149
transform 1 0 27876 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_304
timestamp 1644511149
transform 1 0 29072 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_315
timestamp 1644511149
transform 1 0 30084 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_335
timestamp 1644511149
transform 1 0 31924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_348
timestamp 1644511149
transform 1 0 33120 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_355
timestamp 1644511149
transform 1 0 33764 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1644511149
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1644511149
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_433
timestamp 1644511149
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_445
timestamp 1644511149
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_457
timestamp 1644511149
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1644511149
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1644511149
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_477
timestamp 1644511149
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_489
timestamp 1644511149
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_504
timestamp 1644511149
transform 1 0 47472 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_511
timestamp 1644511149
transform 1 0 48116 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_515
timestamp 1644511149
transform 1 0 48484 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1644511149
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_185
timestamp 1644511149
transform 1 0 18124 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_205
timestamp 1644511149
transform 1 0 19964 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_214
timestamp 1644511149
transform 1 0 20792 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1644511149
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_235
timestamp 1644511149
transform 1 0 22724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_247
timestamp 1644511149
transform 1 0 23828 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_259
timestamp 1644511149
transform 1 0 24932 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_265
timestamp 1644511149
transform 1 0 25484 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_272
timestamp 1644511149
transform 1 0 26128 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_285
timestamp 1644511149
transform 1 0 27324 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_300
timestamp 1644511149
transform 1 0 28704 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_313
timestamp 1644511149
transform 1 0 29900 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_325
timestamp 1644511149
transform 1 0 31004 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_333
timestamp 1644511149
transform 1 0 31740 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_417
timestamp 1644511149
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_429
timestamp 1644511149
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1644511149
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1644511149
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_449
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_461
timestamp 1644511149
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_473
timestamp 1644511149
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_485
timestamp 1644511149
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1644511149
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1644511149
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_505
timestamp 1644511149
transform 1 0 47564 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_513
timestamp 1644511149
transform 1 0 48300 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_145
timestamp 1644511149
transform 1 0 14444 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_158
timestamp 1644511149
transform 1 0 15640 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_183
timestamp 1644511149
transform 1 0 17940 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_192
timestamp 1644511149
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_202
timestamp 1644511149
transform 1 0 19688 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_227
timestamp 1644511149
transform 1 0 21988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_239
timestamp 1644511149
transform 1 0 23092 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_246
timestamp 1644511149
transform 1 0 23736 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_282
timestamp 1644511149
transform 1 0 27048 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_296
timestamp 1644511149
transform 1 0 28336 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_304
timestamp 1644511149
transform 1 0 29072 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_329
timestamp 1644511149
transform 1 0 31372 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_341
timestamp 1644511149
transform 1 0 32476 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_353
timestamp 1644511149
transform 1 0 33580 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_361
timestamp 1644511149
transform 1 0 34316 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_373
timestamp 1644511149
transform 1 0 35420 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_385
timestamp 1644511149
transform 1 0 36524 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_397
timestamp 1644511149
transform 1 0 37628 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_409
timestamp 1644511149
transform 1 0 38732 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_417
timestamp 1644511149
transform 1 0 39468 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_421
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_433
timestamp 1644511149
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_445
timestamp 1644511149
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_457
timestamp 1644511149
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1644511149
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1644511149
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_477
timestamp 1644511149
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_489
timestamp 1644511149
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_501
timestamp 1644511149
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_513
timestamp 1644511149
transform 1 0 48300 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_13
timestamp 1644511149
transform 1 0 2300 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_25
timestamp 1644511149
transform 1 0 3404 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_37
timestamp 1644511149
transform 1 0 4508 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_49
timestamp 1644511149
transform 1 0 5612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_162
timestamp 1644511149
transform 1 0 16008 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_185
timestamp 1644511149
transform 1 0 18124 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_199
timestamp 1644511149
transform 1 0 19412 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_207
timestamp 1644511149
transform 1 0 20148 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_211
timestamp 1644511149
transform 1 0 20516 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_216
timestamp 1644511149
transform 1 0 20976 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_237
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_250
timestamp 1644511149
transform 1 0 24104 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_263
timestamp 1644511149
transform 1 0 25300 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_275
timestamp 1644511149
transform 1 0 26404 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_301
timestamp 1644511149
transform 1 0 28796 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_311
timestamp 1644511149
transform 1 0 29716 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_323
timestamp 1644511149
transform 1 0 30820 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_347
timestamp 1644511149
transform 1 0 33028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_359
timestamp 1644511149
transform 1 0 34132 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_367
timestamp 1644511149
transform 1 0 34868 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_384
timestamp 1644511149
transform 1 0 36432 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_417
timestamp 1644511149
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_429
timestamp 1644511149
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1644511149
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1644511149
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_461
timestamp 1644511149
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_473
timestamp 1644511149
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_485
timestamp 1644511149
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1644511149
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1644511149
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_505
timestamp 1644511149
transform 1 0 47564 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_513
timestamp 1644511149
transform 1 0 48300 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_24
timestamp 1644511149
transform 1 0 3312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1644511149
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_164
timestamp 1644511149
transform 1 0 16192 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_172
timestamp 1644511149
transform 1 0 16928 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_178
timestamp 1644511149
transform 1 0 17480 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_190
timestamp 1644511149
transform 1 0 18584 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_205
timestamp 1644511149
transform 1 0 19964 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_212
timestamp 1644511149
transform 1 0 20608 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_224
timestamp 1644511149
transform 1 0 21712 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_248
timestamp 1644511149
transform 1 0 23920 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_265
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_273
timestamp 1644511149
transform 1 0 26220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_277
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_282
timestamp 1644511149
transform 1 0 27048 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_290
timestamp 1644511149
transform 1 0 27784 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_295
timestamp 1644511149
transform 1 0 28244 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_303
timestamp 1644511149
transform 1 0 28980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_318
timestamp 1644511149
transform 1 0 30360 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_325
timestamp 1644511149
transform 1 0 31004 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_331
timestamp 1644511149
transform 1 0 31556 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_336
timestamp 1644511149
transform 1 0 32016 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_356
timestamp 1644511149
transform 1 0 33856 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_386
timestamp 1644511149
transform 1 0 36616 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_398
timestamp 1644511149
transform 1 0 37720 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_410
timestamp 1644511149
transform 1 0 38824 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_418
timestamp 1644511149
transform 1 0 39560 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_433
timestamp 1644511149
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_445
timestamp 1644511149
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_457
timestamp 1644511149
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1644511149
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1644511149
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_477
timestamp 1644511149
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_489
timestamp 1644511149
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_501
timestamp 1644511149
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_513
timestamp 1644511149
transform 1 0 48300 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_9
timestamp 1644511149
transform 1 0 1932 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_13
timestamp 1644511149
transform 1 0 2300 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_20
timestamp 1644511149
transform 1 0 2944 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_32
timestamp 1644511149
transform 1 0 4048 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_44
timestamp 1644511149
transform 1 0 5152 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_75
timestamp 1644511149
transform 1 0 8004 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_97
timestamp 1644511149
transform 1 0 10028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_109
timestamp 1644511149
transform 1 0 11132 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_121
timestamp 1644511149
transform 1 0 12236 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_144
timestamp 1644511149
transform 1 0 14352 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_148
timestamp 1644511149
transform 1 0 14720 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_153
timestamp 1644511149
transform 1 0 15180 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_160
timestamp 1644511149
transform 1 0 15824 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_173
timestamp 1644511149
transform 1 0 17020 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_202
timestamp 1644511149
transform 1 0 19688 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_208
timestamp 1644511149
transform 1 0 20240 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_213
timestamp 1644511149
transform 1 0 20700 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_221
timestamp 1644511149
transform 1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_233
timestamp 1644511149
transform 1 0 22540 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_241
timestamp 1644511149
transform 1 0 23276 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_258
timestamp 1644511149
transform 1 0 24840 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_264
timestamp 1644511149
transform 1 0 25392 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1644511149
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1644511149
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_301
timestamp 1644511149
transform 1 0 28796 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_311
timestamp 1644511149
transform 1 0 29716 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_319
timestamp 1644511149
transform 1 0 30452 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_332
timestamp 1644511149
transform 1 0 31648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_341
timestamp 1644511149
transform 1 0 32476 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_358
timestamp 1644511149
transform 1 0 34040 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_366
timestamp 1644511149
transform 1 0 34776 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_417
timestamp 1644511149
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_429
timestamp 1644511149
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1644511149
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1644511149
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_461
timestamp 1644511149
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_473
timestamp 1644511149
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_485
timestamp 1644511149
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1644511149
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1644511149
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_505
timestamp 1644511149
transform 1 0 47564 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_512
timestamp 1644511149
transform 1 0 48208 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1644511149
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_126
timestamp 1644511149
transform 1 0 12696 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1644511149
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_147
timestamp 1644511149
transform 1 0 14628 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_151
timestamp 1644511149
transform 1 0 14996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_163
timestamp 1644511149
transform 1 0 16100 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_175
timestamp 1644511149
transform 1 0 17204 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_187
timestamp 1644511149
transform 1 0 18308 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_192
timestamp 1644511149
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_201
timestamp 1644511149
transform 1 0 19596 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_210
timestamp 1644511149
transform 1 0 20424 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_230
timestamp 1644511149
transform 1 0 22264 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_238
timestamp 1644511149
transform 1 0 23000 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1644511149
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_275
timestamp 1644511149
transform 1 0 26404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_285
timestamp 1644511149
transform 1 0 27324 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_295
timestamp 1644511149
transform 1 0 28244 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_304
timestamp 1644511149
transform 1 0 29072 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_313
timestamp 1644511149
transform 1 0 29900 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_330
timestamp 1644511149
transform 1 0 31464 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_338
timestamp 1644511149
transform 1 0 32200 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_349
timestamp 1644511149
transform 1 0 33212 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_358
timestamp 1644511149
transform 1 0 34040 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_369
timestamp 1644511149
transform 1 0 35052 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_378
timestamp 1644511149
transform 1 0 35880 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_390
timestamp 1644511149
transform 1 0 36984 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_402
timestamp 1644511149
transform 1 0 38088 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_414
timestamp 1644511149
transform 1 0 39192 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_433
timestamp 1644511149
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_445
timestamp 1644511149
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_457
timestamp 1644511149
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1644511149
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1644511149
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_477
timestamp 1644511149
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_489
timestamp 1644511149
transform 1 0 46092 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_512
timestamp 1644511149
transform 1 0 48208 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1644511149
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1644511149
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1644511149
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_89
timestamp 1644511149
transform 1 0 9292 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_94
timestamp 1644511149
transform 1 0 9752 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_121
timestamp 1644511149
transform 1 0 12236 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_138
timestamp 1644511149
transform 1 0 13800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_147
timestamp 1644511149
transform 1 0 14628 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_159
timestamp 1644511149
transform 1 0 15732 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_185
timestamp 1644511149
transform 1 0 18124 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_192
timestamp 1644511149
transform 1 0 18768 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1644511149
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_230
timestamp 1644511149
transform 1 0 22264 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_238
timestamp 1644511149
transform 1 0 23000 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_250
timestamp 1644511149
transform 1 0 24104 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_262
timestamp 1644511149
transform 1 0 25208 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_268
timestamp 1644511149
transform 1 0 25760 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_276
timestamp 1644511149
transform 1 0 26496 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_296
timestamp 1644511149
transform 1 0 28336 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_304
timestamp 1644511149
transform 1 0 29072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_315
timestamp 1644511149
transform 1 0 30084 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_325
timestamp 1644511149
transform 1 0 31004 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_333
timestamp 1644511149
transform 1 0 31740 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_348
timestamp 1644511149
transform 1 0 33120 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_360
timestamp 1644511149
transform 1 0 34224 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_368
timestamp 1644511149
transform 1 0 34960 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_386
timestamp 1644511149
transform 1 0 36616 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_417
timestamp 1644511149
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_429
timestamp 1644511149
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1644511149
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1644511149
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_461
timestamp 1644511149
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_473
timestamp 1644511149
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_485
timestamp 1644511149
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_500
timestamp 1644511149
transform 1 0 47104 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_505
timestamp 1644511149
transform 1 0 47564 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_512
timestamp 1644511149
transform 1 0 48208 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1644511149
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_134
timestamp 1644511149
transform 1 0 13432 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_149
timestamp 1644511149
transform 1 0 14812 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_156
timestamp 1644511149
transform 1 0 15456 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_172
timestamp 1644511149
transform 1 0 16928 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_181
timestamp 1644511149
transform 1 0 17756 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1644511149
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1644511149
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_207
timestamp 1644511149
transform 1 0 20148 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_219
timestamp 1644511149
transform 1 0 21252 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_228
timestamp 1644511149
transform 1 0 22080 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_240
timestamp 1644511149
transform 1 0 23184 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_262
timestamp 1644511149
transform 1 0 25208 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_270
timestamp 1644511149
transform 1 0 25944 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_276
timestamp 1644511149
transform 1 0 26496 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_290
timestamp 1644511149
transform 1 0 27784 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_294
timestamp 1644511149
transform 1 0 28152 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_304
timestamp 1644511149
transform 1 0 29072 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_328
timestamp 1644511149
transform 1 0 31280 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_336
timestamp 1644511149
transform 1 0 32016 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_344
timestamp 1644511149
transform 1 0 32752 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_356
timestamp 1644511149
transform 1 0 33856 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_373
timestamp 1644511149
transform 1 0 35420 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_385
timestamp 1644511149
transform 1 0 36524 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_397
timestamp 1644511149
transform 1 0 37628 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_409
timestamp 1644511149
transform 1 0 38732 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_417
timestamp 1644511149
transform 1 0 39468 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_433
timestamp 1644511149
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_445
timestamp 1644511149
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_457
timestamp 1644511149
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1644511149
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1644511149
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_477
timestamp 1644511149
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_489
timestamp 1644511149
transform 1 0 46092 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_512
timestamp 1644511149
transform 1 0 48208 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_9
timestamp 1644511149
transform 1 0 1932 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_31
timestamp 1644511149
transform 1 0 3956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_43
timestamp 1644511149
transform 1 0 5060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_100
timestamp 1644511149
transform 1 0 10304 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_121
timestamp 1644511149
transform 1 0 12236 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_138
timestamp 1644511149
transform 1 0 13800 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_152
timestamp 1644511149
transform 1 0 15088 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_164
timestamp 1644511149
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_176
timestamp 1644511149
transform 1 0 17296 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_184
timestamp 1644511149
transform 1 0 18032 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_192
timestamp 1644511149
transform 1 0 18768 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_202
timestamp 1644511149
transform 1 0 19688 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_210
timestamp 1644511149
transform 1 0 20424 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1644511149
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_237
timestamp 1644511149
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_249
timestamp 1644511149
transform 1 0 24012 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_258
timestamp 1644511149
transform 1 0 24840 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_270
timestamp 1644511149
transform 1 0 25944 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1644511149
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_288
timestamp 1644511149
transform 1 0 27600 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_294
timestamp 1644511149
transform 1 0 28152 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_299
timestamp 1644511149
transform 1 0 28612 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_312
timestamp 1644511149
transform 1 0 29808 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_320
timestamp 1644511149
transform 1 0 30544 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_332
timestamp 1644511149
transform 1 0 31648 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_353
timestamp 1644511149
transform 1 0 33580 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_365
timestamp 1644511149
transform 1 0 34684 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_377
timestamp 1644511149
transform 1 0 35788 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_389
timestamp 1644511149
transform 1 0 36892 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_417
timestamp 1644511149
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_429
timestamp 1644511149
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1644511149
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1644511149
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_461
timestamp 1644511149
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_473
timestamp 1644511149
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_485
timestamp 1644511149
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_500
timestamp 1644511149
transform 1 0 47104 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_508
timestamp 1644511149
transform 1 0 47840 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_9
timestamp 1644511149
transform 1 0 1932 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_13
timestamp 1644511149
transform 1 0 2300 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_22
timestamp 1644511149
transform 1 0 3128 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_93
timestamp 1644511149
transform 1 0 9660 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1644511149
transform 1 0 11868 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_129
timestamp 1644511149
transform 1 0 12972 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1644511149
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_145
timestamp 1644511149
transform 1 0 14444 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_154
timestamp 1644511149
transform 1 0 15272 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_166
timestamp 1644511149
transform 1 0 16376 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_170
timestamp 1644511149
transform 1 0 16744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_179
timestamp 1644511149
transform 1 0 17572 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_187
timestamp 1644511149
transform 1 0 18308 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1644511149
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_213
timestamp 1644511149
transform 1 0 20700 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_225
timestamp 1644511149
transform 1 0 21804 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_231
timestamp 1644511149
transform 1 0 22356 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_248
timestamp 1644511149
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_257
timestamp 1644511149
transform 1 0 24748 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_269
timestamp 1644511149
transform 1 0 25852 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_277
timestamp 1644511149
transform 1 0 26588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_284
timestamp 1644511149
transform 1 0 27232 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_288
timestamp 1644511149
transform 1 0 27600 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_293
timestamp 1644511149
transform 1 0 28060 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_305
timestamp 1644511149
transform 1 0 29164 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_321
timestamp 1644511149
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_333
timestamp 1644511149
transform 1 0 31740 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_343
timestamp 1644511149
transform 1 0 32660 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_352
timestamp 1644511149
transform 1 0 33488 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_381
timestamp 1644511149
transform 1 0 36156 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_410
timestamp 1644511149
transform 1 0 38824 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_418
timestamp 1644511149
transform 1 0 39560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_421
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_433
timestamp 1644511149
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_445
timestamp 1644511149
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_457
timestamp 1644511149
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1644511149
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1644511149
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_477
timestamp 1644511149
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_489
timestamp 1644511149
transform 1 0 46092 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_512
timestamp 1644511149
transform 1 0 48208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_11
timestamp 1644511149
transform 1 0 2116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_23
timestamp 1644511149
transform 1 0 3220 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_35
timestamp 1644511149
transform 1 0 4324 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_47
timestamp 1644511149
transform 1 0 5428 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_89
timestamp 1644511149
transform 1 0 9292 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_95
timestamp 1644511149
transform 1 0 9844 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_107
timestamp 1644511149
transform 1 0 10948 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_137
timestamp 1644511149
transform 1 0 13708 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_145
timestamp 1644511149
transform 1 0 14444 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_162
timestamp 1644511149
transform 1 0 16008 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_189
timestamp 1644511149
transform 1 0 18492 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_201
timestamp 1644511149
transform 1 0 19596 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_210
timestamp 1644511149
transform 1 0 20424 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_219
timestamp 1644511149
transform 1 0 21252 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1644511149
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_237
timestamp 1644511149
transform 1 0 22908 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_248
timestamp 1644511149
transform 1 0 23920 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_261
timestamp 1644511149
transform 1 0 25116 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_271
timestamp 1644511149
transform 1 0 26036 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_285
timestamp 1644511149
transform 1 0 27324 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_298
timestamp 1644511149
transform 1 0 28520 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_311
timestamp 1644511149
transform 1 0 29716 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_323
timestamp 1644511149
transform 1 0 30820 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1644511149
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_340
timestamp 1644511149
transform 1 0 32384 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_352
timestamp 1644511149
transform 1 0 33488 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_364
timestamp 1644511149
transform 1 0 34592 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_376
timestamp 1644511149
transform 1 0 35696 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1644511149
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1644511149
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_396
timestamp 1644511149
transform 1 0 37536 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_408
timestamp 1644511149
transform 1 0 38640 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_420
timestamp 1644511149
transform 1 0 39744 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_432
timestamp 1644511149
transform 1 0 40848 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_444
timestamp 1644511149
transform 1 0 41952 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_449
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_461
timestamp 1644511149
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_473
timestamp 1644511149
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_485
timestamp 1644511149
transform 1 0 45724 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_493
timestamp 1644511149
transform 1 0 46460 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_499
timestamp 1644511149
transform 1 0 47012 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1644511149
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_508
timestamp 1644511149
transform 1 0 47840 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1644511149
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_59
timestamp 1644511149
transform 1 0 6532 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_69
timestamp 1644511149
transform 1 0 7452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_81
timestamp 1644511149
transform 1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_101
timestamp 1644511149
transform 1 0 10396 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1644511149
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1644511149
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_147
timestamp 1644511149
transform 1 0 14628 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_153
timestamp 1644511149
transform 1 0 15180 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_178
timestamp 1644511149
transform 1 0 17480 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_186
timestamp 1644511149
transform 1 0 18216 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1644511149
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_205
timestamp 1644511149
transform 1 0 19964 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_225
timestamp 1644511149
transform 1 0 21804 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_237
timestamp 1644511149
transform 1 0 22908 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_249
timestamp 1644511149
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_260
timestamp 1644511149
transform 1 0 25024 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_264
timestamp 1644511149
transform 1 0 25392 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_269
timestamp 1644511149
transform 1 0 25852 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_280
timestamp 1644511149
transform 1 0 26864 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_294
timestamp 1644511149
transform 1 0 28152 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_302
timestamp 1644511149
transform 1 0 28888 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_325
timestamp 1644511149
transform 1 0 31004 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_333
timestamp 1644511149
transform 1 0 31740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_344
timestamp 1644511149
transform 1 0 32752 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_356
timestamp 1644511149
transform 1 0 33856 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_382
timestamp 1644511149
transform 1 0 36248 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_389
timestamp 1644511149
transform 1 0 36892 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_414
timestamp 1644511149
transform 1 0 39192 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_421
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_433
timestamp 1644511149
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_445
timestamp 1644511149
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_457
timestamp 1644511149
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1644511149
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1644511149
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_477
timestamp 1644511149
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_489
timestamp 1644511149
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_501
timestamp 1644511149
transform 1 0 47196 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_507
timestamp 1644511149
transform 1 0 47748 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_515
timestamp 1644511149
transform 1 0 48484 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_9
timestamp 1644511149
transform 1 0 1932 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_13
timestamp 1644511149
transform 1 0 2300 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_20
timestamp 1644511149
transform 1 0 2944 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_32
timestamp 1644511149
transform 1 0 4048 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_44
timestamp 1644511149
transform 1 0 5152 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_61
timestamp 1644511149
transform 1 0 6716 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_65
timestamp 1644511149
transform 1 0 7084 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_85
timestamp 1644511149
transform 1 0 8924 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_89
timestamp 1644511149
transform 1 0 9292 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_98
timestamp 1644511149
transform 1 0 10120 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_107
timestamp 1644511149
transform 1 0 10948 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_118
timestamp 1644511149
transform 1 0 11960 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_126
timestamp 1644511149
transform 1 0 12696 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_145
timestamp 1644511149
transform 1 0 14444 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_157
timestamp 1644511149
transform 1 0 15548 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_163
timestamp 1644511149
transform 1 0 16100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1644511149
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_179
timestamp 1644511149
transform 1 0 17572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_191
timestamp 1644511149
transform 1 0 18676 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_203
timestamp 1644511149
transform 1 0 19780 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1644511149
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_225
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_237
timestamp 1644511149
transform 1 0 22908 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_243
timestamp 1644511149
transform 1 0 23460 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_251
timestamp 1644511149
transform 1 0 24196 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_263
timestamp 1644511149
transform 1 0 25300 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_276
timestamp 1644511149
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_290
timestamp 1644511149
transform 1 0 27784 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_303
timestamp 1644511149
transform 1 0 28980 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_323
timestamp 1644511149
transform 1 0 30820 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1644511149
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_345
timestamp 1644511149
transform 1 0 32844 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_354
timestamp 1644511149
transform 1 0 33672 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_376
timestamp 1644511149
transform 1 0 35696 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1644511149
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1644511149
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_414
timestamp 1644511149
transform 1 0 39192 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_426
timestamp 1644511149
transform 1 0 40296 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_438
timestamp 1644511149
transform 1 0 41400 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_446
timestamp 1644511149
transform 1 0 42136 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_449
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_461
timestamp 1644511149
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_473
timestamp 1644511149
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_485
timestamp 1644511149
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1644511149
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1644511149
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_505
timestamp 1644511149
transform 1 0 47564 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_513
timestamp 1644511149
transform 1 0 48300 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_14
timestamp 1644511149
transform 1 0 2392 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1644511149
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_94
timestamp 1644511149
transform 1 0 9752 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_106
timestamp 1644511149
transform 1 0 10856 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_110
timestamp 1644511149
transform 1 0 11224 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_119
timestamp 1644511149
transform 1 0 12052 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_127
timestamp 1644511149
transform 1 0 12788 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_136
timestamp 1644511149
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_146
timestamp 1644511149
transform 1 0 14536 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_158
timestamp 1644511149
transform 1 0 15640 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_162
timestamp 1644511149
transform 1 0 16008 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_166
timestamp 1644511149
transform 1 0 16376 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_191
timestamp 1644511149
transform 1 0 18676 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1644511149
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_209
timestamp 1644511149
transform 1 0 20332 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_218
timestamp 1644511149
transform 1 0 21160 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_225
timestamp 1644511149
transform 1 0 21804 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_237
timestamp 1644511149
transform 1 0 22908 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_248
timestamp 1644511149
transform 1 0 23920 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_262
timestamp 1644511149
transform 1 0 25208 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_271
timestamp 1644511149
transform 1 0 26036 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_277
timestamp 1644511149
transform 1 0 26588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_282
timestamp 1644511149
transform 1 0 27048 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_291
timestamp 1644511149
transform 1 0 27876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_303
timestamp 1644511149
transform 1 0 28980 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1644511149
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_312
timestamp 1644511149
transform 1 0 29808 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_324
timestamp 1644511149
transform 1 0 30912 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_332
timestamp 1644511149
transform 1 0 31648 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_351
timestamp 1644511149
transform 1 0 33396 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1644511149
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_370
timestamp 1644511149
transform 1 0 35144 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_382
timestamp 1644511149
transform 1 0 36248 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_404
timestamp 1644511149
transform 1 0 38272 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_416
timestamp 1644511149
transform 1 0 39376 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_421
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_433
timestamp 1644511149
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_445
timestamp 1644511149
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_457
timestamp 1644511149
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1644511149
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1644511149
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_477
timestamp 1644511149
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_489
timestamp 1644511149
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_501
timestamp 1644511149
transform 1 0 47196 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_507
timestamp 1644511149
transform 1 0 47748 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_515
timestamp 1644511149
transform 1 0 48484 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_28
timestamp 1644511149
transform 1 0 3680 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_40
timestamp 1644511149
transform 1 0 4784 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1644511149
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_91
timestamp 1644511149
transform 1 0 9476 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_100
timestamp 1644511149
transform 1 0 10304 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_121
timestamp 1644511149
transform 1 0 12236 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_129
timestamp 1644511149
transform 1 0 12972 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_139
timestamp 1644511149
transform 1 0 13892 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_148
timestamp 1644511149
transform 1 0 14720 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_162
timestamp 1644511149
transform 1 0 16008 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_173
timestamp 1644511149
transform 1 0 17020 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_178
timestamp 1644511149
transform 1 0 17480 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_190
timestamp 1644511149
transform 1 0 18584 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_197
timestamp 1644511149
transform 1 0 19228 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_205
timestamp 1644511149
transform 1 0 19964 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_212
timestamp 1644511149
transform 1 0 20608 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_216
timestamp 1644511149
transform 1 0 20976 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1644511149
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_229
timestamp 1644511149
transform 1 0 22172 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_235
timestamp 1644511149
transform 1 0 22724 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_252
timestamp 1644511149
transform 1 0 24288 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_259
timestamp 1644511149
transform 1 0 24932 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_271
timestamp 1644511149
transform 1 0 26036 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1644511149
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_286
timestamp 1644511149
transform 1 0 27416 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_298
timestamp 1644511149
transform 1 0 28520 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_310
timestamp 1644511149
transform 1 0 29624 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_322
timestamp 1644511149
transform 1 0 30728 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_334
timestamp 1644511149
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_341
timestamp 1644511149
transform 1 0 32476 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_347
timestamp 1644511149
transform 1 0 33028 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_369
timestamp 1644511149
transform 1 0 35052 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_381
timestamp 1644511149
transform 1 0 36156 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_387
timestamp 1644511149
transform 1 0 36708 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1644511149
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_396
timestamp 1644511149
transform 1 0 37536 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_408
timestamp 1644511149
transform 1 0 38640 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_420
timestamp 1644511149
transform 1 0 39744 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_432
timestamp 1644511149
transform 1 0 40848 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_444
timestamp 1644511149
transform 1 0 41952 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_449
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_461
timestamp 1644511149
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_473
timestamp 1644511149
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_485
timestamp 1644511149
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1644511149
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1644511149
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_505
timestamp 1644511149
transform 1 0 47564 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_512
timestamp 1644511149
transform 1 0 48208 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_7
timestamp 1644511149
transform 1 0 1748 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_11
timestamp 1644511149
transform 1 0 2116 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_23
timestamp 1644511149
transform 1 0 3220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_37
timestamp 1644511149
transform 1 0 4508 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_60
timestamp 1644511149
transform 1 0 6624 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_72
timestamp 1644511149
transform 1 0 7728 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_76
timestamp 1644511149
transform 1 0 8096 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_80
timestamp 1644511149
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_96
timestamp 1644511149
transform 1 0 9936 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_116
timestamp 1644511149
transform 1 0 11776 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_120
timestamp 1644511149
transform 1 0 12144 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_132
timestamp 1644511149
transform 1 0 13248 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_149
timestamp 1644511149
transform 1 0 14812 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_169
timestamp 1644511149
transform 1 0 16652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_174
timestamp 1644511149
transform 1 0 17112 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_181
timestamp 1644511149
transform 1 0 17756 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_191
timestamp 1644511149
transform 1 0 18676 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1644511149
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_201
timestamp 1644511149
transform 1 0 19596 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_208
timestamp 1644511149
transform 1 0 20240 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_212
timestamp 1644511149
transform 1 0 20608 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_217
timestamp 1644511149
transform 1 0 21068 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_221
timestamp 1644511149
transform 1 0 21436 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_226
timestamp 1644511149
transform 1 0 21896 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_234
timestamp 1644511149
transform 1 0 22632 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_246
timestamp 1644511149
transform 1 0 23736 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_265
timestamp 1644511149
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_277
timestamp 1644511149
transform 1 0 26588 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_288
timestamp 1644511149
transform 1 0 27600 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_296
timestamp 1644511149
transform 1 0 28336 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_303
timestamp 1644511149
transform 1 0 28980 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1644511149
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_321
timestamp 1644511149
transform 1 0 30636 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_329
timestamp 1644511149
transform 1 0 31372 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_351
timestamp 1644511149
transform 1 0 33396 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_358
timestamp 1644511149
transform 1 0 34040 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_389
timestamp 1644511149
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_401
timestamp 1644511149
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1644511149
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1644511149
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_421
timestamp 1644511149
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_433
timestamp 1644511149
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_445
timestamp 1644511149
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_457
timestamp 1644511149
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1644511149
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1644511149
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_477
timestamp 1644511149
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_489
timestamp 1644511149
transform 1 0 46092 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_512
timestamp 1644511149
transform 1 0 48208 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_43
timestamp 1644511149
transform 1 0 5060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_104
timestamp 1644511149
transform 1 0 10672 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_118
timestamp 1644511149
transform 1 0 11960 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_146
timestamp 1644511149
transform 1 0 14536 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_154
timestamp 1644511149
transform 1 0 15272 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_164
timestamp 1644511149
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_173
timestamp 1644511149
transform 1 0 17020 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_176
timestamp 1644511149
transform 1 0 17296 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_186
timestamp 1644511149
transform 1 0 18216 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_196
timestamp 1644511149
transform 1 0 19136 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_216
timestamp 1644511149
transform 1 0 20976 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_229
timestamp 1644511149
transform 1 0 22172 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_237
timestamp 1644511149
transform 1 0 22908 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_245
timestamp 1644511149
transform 1 0 23644 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_253
timestamp 1644511149
transform 1 0 24380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_265
timestamp 1644511149
transform 1 0 25484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_277
timestamp 1644511149
transform 1 0 26588 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_291
timestamp 1644511149
transform 1 0 27876 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_305
timestamp 1644511149
transform 1 0 29164 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_315
timestamp 1644511149
transform 1 0 30084 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_321
timestamp 1644511149
transform 1 0 30636 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1644511149
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1644511149
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_348
timestamp 1644511149
transform 1 0 33120 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_373
timestamp 1644511149
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1644511149
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1644511149
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_414
timestamp 1644511149
transform 1 0 39192 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_426
timestamp 1644511149
transform 1 0 40296 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_438
timestamp 1644511149
transform 1 0 41400 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_446
timestamp 1644511149
transform 1 0 42136 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_449
timestamp 1644511149
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_461
timestamp 1644511149
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_473
timestamp 1644511149
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_485
timestamp 1644511149
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1644511149
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1644511149
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_508
timestamp 1644511149
transform 1 0 47840 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_72
timestamp 1644511149
transform 1 0 7728 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_109
timestamp 1644511149
transform 1 0 11132 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_117
timestamp 1644511149
transform 1 0 11868 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_122
timestamp 1644511149
transform 1 0 12328 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 1644511149
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_146
timestamp 1644511149
transform 1 0 14536 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_158
timestamp 1644511149
transform 1 0 15640 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_170
timestamp 1644511149
transform 1 0 16744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_187
timestamp 1644511149
transform 1 0 18308 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1644511149
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_207
timestamp 1644511149
transform 1 0 20148 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_215
timestamp 1644511149
transform 1 0 20884 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_226
timestamp 1644511149
transform 1 0 21896 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_240
timestamp 1644511149
transform 1 0 23184 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_268
timestamp 1644511149
transform 1 0 25760 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_282
timestamp 1644511149
transform 1 0 27048 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_292
timestamp 1644511149
transform 1 0 27968 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_302
timestamp 1644511149
transform 1 0 28888 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_315
timestamp 1644511149
transform 1 0 30084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_333
timestamp 1644511149
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_345
timestamp 1644511149
transform 1 0 32844 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_354
timestamp 1644511149
transform 1 0 33672 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_362
timestamp 1644511149
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_377
timestamp 1644511149
transform 1 0 35788 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_401
timestamp 1644511149
transform 1 0 37996 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_408
timestamp 1644511149
transform 1 0 38640 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_421
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_433
timestamp 1644511149
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_445
timestamp 1644511149
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_457
timestamp 1644511149
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1644511149
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1644511149
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_477
timestamp 1644511149
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_489
timestamp 1644511149
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_501
timestamp 1644511149
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_513
timestamp 1644511149
transform 1 0 48300 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_65
timestamp 1644511149
transform 1 0 7084 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_88
timestamp 1644511149
transform 1 0 9200 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_100
timestamp 1644511149
transform 1 0 10304 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_134
timestamp 1644511149
transform 1 0 13432 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_149
timestamp 1644511149
transform 1 0 14812 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_160
timestamp 1644511149
transform 1 0 15824 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_181
timestamp 1644511149
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_193
timestamp 1644511149
transform 1 0 18860 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_199
timestamp 1644511149
transform 1 0 19412 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_203
timestamp 1644511149
transform 1 0 19780 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_211
timestamp 1644511149
transform 1 0 20516 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_215
timestamp 1644511149
transform 1 0 20884 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_220
timestamp 1644511149
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_230
timestamp 1644511149
transform 1 0 22264 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_250
timestamp 1644511149
transform 1 0 24104 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_258
timestamp 1644511149
transform 1 0 24840 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_262
timestamp 1644511149
transform 1 0 25208 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_276
timestamp 1644511149
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_287
timestamp 1644511149
transform 1 0 27508 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_301
timestamp 1644511149
transform 1 0 28796 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_305
timestamp 1644511149
transform 1 0 29164 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_313
timestamp 1644511149
transform 1 0 29900 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_321
timestamp 1644511149
transform 1 0 30636 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_324
timestamp 1644511149
transform 1 0 30912 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_332
timestamp 1644511149
transform 1 0 31648 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_343
timestamp 1644511149
transform 1 0 32660 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_350
timestamp 1644511149
transform 1 0 33304 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_375
timestamp 1644511149
transform 1 0 35604 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_381
timestamp 1644511149
transform 1 0 36156 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1644511149
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1644511149
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_396
timestamp 1644511149
transform 1 0 37536 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_408
timestamp 1644511149
transform 1 0 38640 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_420
timestamp 1644511149
transform 1 0 39744 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_432
timestamp 1644511149
transform 1 0 40848 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_444
timestamp 1644511149
transform 1 0 41952 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_449
timestamp 1644511149
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_461
timestamp 1644511149
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_473
timestamp 1644511149
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_485
timestamp 1644511149
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1644511149
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1644511149
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_505
timestamp 1644511149
transform 1 0 47564 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_512
timestamp 1644511149
transform 1 0 48208 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_61
timestamp 1644511149
transform 1 0 6716 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_78
timestamp 1644511149
transform 1 0 8280 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_93
timestamp 1644511149
transform 1 0 9660 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_100
timestamp 1644511149
transform 1 0 10304 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_112
timestamp 1644511149
transform 1 0 11408 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_124
timestamp 1644511149
transform 1 0 12512 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_136
timestamp 1644511149
transform 1 0 13616 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_146
timestamp 1644511149
transform 1 0 14536 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_158
timestamp 1644511149
transform 1 0 15640 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_170
timestamp 1644511149
transform 1 0 16744 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_178
timestamp 1644511149
transform 1 0 17480 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_186
timestamp 1644511149
transform 1 0 18216 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1644511149
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_197
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_207
timestamp 1644511149
transform 1 0 20148 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_216
timestamp 1644511149
transform 1 0 20976 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_228
timestamp 1644511149
transform 1 0 22080 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_240
timestamp 1644511149
transform 1 0 23184 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_269
timestamp 1644511149
transform 1 0 25852 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_276
timestamp 1644511149
transform 1 0 26496 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_283
timestamp 1644511149
transform 1 0 27140 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_295
timestamp 1644511149
transform 1 0 28244 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_304
timestamp 1644511149
transform 1 0 29072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_317
timestamp 1644511149
transform 1 0 30268 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_321
timestamp 1644511149
transform 1 0 30636 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_329
timestamp 1644511149
transform 1 0 31372 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_345
timestamp 1644511149
transform 1 0 32844 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_351
timestamp 1644511149
transform 1 0 33396 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_360
timestamp 1644511149
transform 1 0 34224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_384
timestamp 1644511149
transform 1 0 36432 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_388
timestamp 1644511149
transform 1 0 36800 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_410
timestamp 1644511149
transform 1 0 38824 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_418
timestamp 1644511149
transform 1 0 39560 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_421
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_433
timestamp 1644511149
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_445
timestamp 1644511149
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_457
timestamp 1644511149
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1644511149
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1644511149
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_477
timestamp 1644511149
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_489
timestamp 1644511149
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_501
timestamp 1644511149
transform 1 0 47196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_512
timestamp 1644511149
transform 1 0 48208 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_11
timestamp 1644511149
transform 1 0 2116 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_18
timestamp 1644511149
transform 1 0 2760 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_30
timestamp 1644511149
transform 1 0 3864 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_42
timestamp 1644511149
transform 1 0 4968 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1644511149
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_100
timestamp 1644511149
transform 1 0 10304 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_108
timestamp 1644511149
transform 1 0 11040 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_125
timestamp 1644511149
transform 1 0 12604 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_131
timestamp 1644511149
transform 1 0 13156 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_137
timestamp 1644511149
transform 1 0 13708 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_149
timestamp 1644511149
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1644511149
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_177
timestamp 1644511149
transform 1 0 17388 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_180
timestamp 1644511149
transform 1 0 17664 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_190
timestamp 1644511149
transform 1 0 18584 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_202
timestamp 1644511149
transform 1 0 19688 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_210
timestamp 1644511149
transform 1 0 20424 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_220
timestamp 1644511149
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_237
timestamp 1644511149
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_255
timestamp 1644511149
transform 1 0 24564 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_263
timestamp 1644511149
transform 1 0 25300 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_270
timestamp 1644511149
transform 1 0 25944 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1644511149
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_293
timestamp 1644511149
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_305
timestamp 1644511149
transform 1 0 29164 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_314
timestamp 1644511149
transform 1 0 29992 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_322
timestamp 1644511149
transform 1 0 30728 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_331
timestamp 1644511149
transform 1 0 31556 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1644511149
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_346
timestamp 1644511149
transform 1 0 32936 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_350
timestamp 1644511149
transform 1 0 33304 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_372
timestamp 1644511149
transform 1 0 35328 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_381
timestamp 1644511149
transform 1 0 36156 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_389
timestamp 1644511149
transform 1 0 36892 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_417
timestamp 1644511149
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_429
timestamp 1644511149
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1644511149
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1644511149
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_449
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_461
timestamp 1644511149
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_473
timestamp 1644511149
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_485
timestamp 1644511149
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1644511149
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1644511149
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_508
timestamp 1644511149
transform 1 0 47840 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_24
timestamp 1644511149
transform 1 0 3312 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_93
timestamp 1644511149
transform 1 0 9660 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_104
timestamp 1644511149
transform 1 0 10672 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_116
timestamp 1644511149
transform 1 0 11776 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_134
timestamp 1644511149
transform 1 0 13432 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_151
timestamp 1644511149
transform 1 0 14996 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_162
timestamp 1644511149
transform 1 0 16008 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_166
timestamp 1644511149
transform 1 0 16376 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_172
timestamp 1644511149
transform 1 0 16928 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_192
timestamp 1644511149
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_202
timestamp 1644511149
transform 1 0 19688 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_226
timestamp 1644511149
transform 1 0 21896 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_246
timestamp 1644511149
transform 1 0 23736 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_269
timestamp 1644511149
transform 1 0 25852 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_277
timestamp 1644511149
transform 1 0 26588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_282
timestamp 1644511149
transform 1 0 27048 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_289
timestamp 1644511149
transform 1 0 27692 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_299
timestamp 1644511149
transform 1 0 28612 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1644511149
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_316
timestamp 1644511149
transform 1 0 30176 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_329
timestamp 1644511149
transform 1 0 31372 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_353
timestamp 1644511149
transform 1 0 33580 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_361
timestamp 1644511149
transform 1 0 34316 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_381
timestamp 1644511149
transform 1 0 36156 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_393
timestamp 1644511149
transform 1 0 37260 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_405
timestamp 1644511149
transform 1 0 38364 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_417
timestamp 1644511149
transform 1 0 39468 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_421
timestamp 1644511149
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_433
timestamp 1644511149
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_445
timestamp 1644511149
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_457
timestamp 1644511149
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1644511149
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1644511149
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_477
timestamp 1644511149
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_489
timestamp 1644511149
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_501
timestamp 1644511149
transform 1 0 47196 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_512
timestamp 1644511149
transform 1 0 48208 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_7
timestamp 1644511149
transform 1 0 1748 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_11
timestamp 1644511149
transform 1 0 2116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_23
timestamp 1644511149
transform 1 0 3220 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_35
timestamp 1644511149
transform 1 0 4324 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_47
timestamp 1644511149
transform 1 0 5428 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_77
timestamp 1644511149
transform 1 0 8188 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_85
timestamp 1644511149
transform 1 0 8924 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_95
timestamp 1644511149
transform 1 0 9844 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_108
timestamp 1644511149
transform 1 0 11040 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_119
timestamp 1644511149
transform 1 0 12052 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_126
timestamp 1644511149
transform 1 0 12696 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_134
timestamp 1644511149
transform 1 0 13432 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_142
timestamp 1644511149
transform 1 0 14168 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_153
timestamp 1644511149
transform 1 0 15180 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_162
timestamp 1644511149
transform 1 0 16008 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_177
timestamp 1644511149
transform 1 0 17388 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_185
timestamp 1644511149
transform 1 0 18124 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_203
timestamp 1644511149
transform 1 0 19780 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_211
timestamp 1644511149
transform 1 0 20516 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_220
timestamp 1644511149
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_231
timestamp 1644511149
transform 1 0 22356 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_248
timestamp 1644511149
transform 1 0 23920 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_260
timestamp 1644511149
transform 1 0 25024 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_269
timestamp 1644511149
transform 1 0 25852 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_277
timestamp 1644511149
transform 1 0 26588 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_285
timestamp 1644511149
transform 1 0 27324 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_291
timestamp 1644511149
transform 1 0 27876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_303
timestamp 1644511149
transform 1 0 28980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_309
timestamp 1644511149
transform 1 0 29532 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_313
timestamp 1644511149
transform 1 0 29900 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_319
timestamp 1644511149
transform 1 0 30452 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_323
timestamp 1644511149
transform 1 0 30820 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_331
timestamp 1644511149
transform 1 0 31556 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1644511149
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_353
timestamp 1644511149
transform 1 0 33580 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_361
timestamp 1644511149
transform 1 0 34316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_370
timestamp 1644511149
transform 1 0 35144 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_379
timestamp 1644511149
transform 1 0 35972 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1644511149
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_415
timestamp 1644511149
transform 1 0 39284 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_427
timestamp 1644511149
transform 1 0 40388 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_439
timestamp 1644511149
transform 1 0 41492 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1644511149
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_449
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_461
timestamp 1644511149
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_473
timestamp 1644511149
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_485
timestamp 1644511149
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1644511149
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1644511149
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_505
timestamp 1644511149
transform 1 0 47564 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_512
timestamp 1644511149
transform 1 0 48208 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_11
timestamp 1644511149
transform 1 0 2116 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_23
timestamp 1644511149
transform 1 0 3220 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_91
timestamp 1644511149
transform 1 0 9476 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_102
timestamp 1644511149
transform 1 0 10488 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_110
timestamp 1644511149
transform 1 0 11224 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_114
timestamp 1644511149
transform 1 0 11592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_122
timestamp 1644511149
transform 1 0 12328 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1644511149
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_150
timestamp 1644511149
transform 1 0 14904 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_157
timestamp 1644511149
transform 1 0 15548 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_161
timestamp 1644511149
transform 1 0 15916 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_178
timestamp 1644511149
transform 1 0 17480 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_182
timestamp 1644511149
transform 1 0 17848 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1644511149
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_209
timestamp 1644511149
transform 1 0 20332 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_215
timestamp 1644511149
transform 1 0 20884 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_227
timestamp 1644511149
transform 1 0 21988 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_248
timestamp 1644511149
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_256
timestamp 1644511149
transform 1 0 24656 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_268
timestamp 1644511149
transform 1 0 25760 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_274
timestamp 1644511149
transform 1 0 26312 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_294
timestamp 1644511149
transform 1 0 28152 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1644511149
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1644511149
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_309
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_317
timestamp 1644511149
transform 1 0 30268 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_325
timestamp 1644511149
transform 1 0 31004 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_346
timestamp 1644511149
transform 1 0 32936 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_358
timestamp 1644511149
transform 1 0 34040 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_370
timestamp 1644511149
transform 1 0 35144 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_379
timestamp 1644511149
transform 1 0 35972 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_391
timestamp 1644511149
transform 1 0 37076 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_416
timestamp 1644511149
transform 1 0 39376 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_421
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_433
timestamp 1644511149
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_445
timestamp 1644511149
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_457
timestamp 1644511149
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1644511149
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1644511149
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_477
timestamp 1644511149
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_489
timestamp 1644511149
transform 1 0 46092 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_512
timestamp 1644511149
transform 1 0 48208 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_88
timestamp 1644511149
transform 1 0 9200 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_96
timestamp 1644511149
transform 1 0 9936 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_101
timestamp 1644511149
transform 1 0 10396 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_109
timestamp 1644511149
transform 1 0 11132 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_137
timestamp 1644511149
transform 1 0 13708 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_151
timestamp 1644511149
transform 1 0 14996 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_163
timestamp 1644511149
transform 1 0 16100 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_181
timestamp 1644511149
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_193
timestamp 1644511149
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_205
timestamp 1644511149
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1644511149
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1644511149
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_242
timestamp 1644511149
transform 1 0 23368 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_254
timestamp 1644511149
transform 1 0 24472 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_266
timestamp 1644511149
transform 1 0 25576 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_270
timestamp 1644511149
transform 1 0 25944 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_275
timestamp 1644511149
transform 1 0 26404 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1644511149
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_286
timestamp 1644511149
transform 1 0 27416 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_295
timestamp 1644511149
transform 1 0 28244 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_303
timestamp 1644511149
transform 1 0 28980 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_323
timestamp 1644511149
transform 1 0 30820 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_331
timestamp 1644511149
transform 1 0 31556 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1644511149
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_361
timestamp 1644511149
transform 1 0 34316 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_369
timestamp 1644511149
transform 1 0 35052 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_388
timestamp 1644511149
transform 1 0 36800 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_398
timestamp 1644511149
transform 1 0 37720 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_417
timestamp 1644511149
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_429
timestamp 1644511149
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1644511149
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1644511149
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_449
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_461
timestamp 1644511149
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_473
timestamp 1644511149
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_485
timestamp 1644511149
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_500
timestamp 1644511149
transform 1 0 47104 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_508
timestamp 1644511149
transform 1 0 47840 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1644511149
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_80
timestamp 1644511149
transform 1 0 8464 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_88
timestamp 1644511149
transform 1 0 9200 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_100
timestamp 1644511149
transform 1 0 10304 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_109
timestamp 1644511149
transform 1 0 11132 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_118
timestamp 1644511149
transform 1 0 11960 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_130
timestamp 1644511149
transform 1 0 13064 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1644511149
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_146
timestamp 1644511149
transform 1 0 14536 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_158
timestamp 1644511149
transform 1 0 15640 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_170
timestamp 1644511149
transform 1 0 16744 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_190
timestamp 1644511149
transform 1 0 18584 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_205
timestamp 1644511149
transform 1 0 19964 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_228
timestamp 1644511149
transform 1 0 22080 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_240
timestamp 1644511149
transform 1 0 23184 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_258
timestamp 1644511149
transform 1 0 24840 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_270
timestamp 1644511149
transform 1 0 25944 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_282
timestamp 1644511149
transform 1 0 27048 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_289
timestamp 1644511149
transform 1 0 27692 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_295
timestamp 1644511149
transform 1 0 28244 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_304
timestamp 1644511149
transform 1 0 29072 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_314
timestamp 1644511149
transform 1 0 29992 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_339
timestamp 1644511149
transform 1 0 32292 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_359
timestamp 1644511149
transform 1 0 34132 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1644511149
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_373
timestamp 1644511149
transform 1 0 35420 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_385
timestamp 1644511149
transform 1 0 36524 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_390
timestamp 1644511149
transform 1 0 36984 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_415
timestamp 1644511149
transform 1 0 39284 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1644511149
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_421
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_433
timestamp 1644511149
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_445
timestamp 1644511149
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_457
timestamp 1644511149
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1644511149
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1644511149
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_477
timestamp 1644511149
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_489
timestamp 1644511149
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_501
timestamp 1644511149
transform 1 0 47196 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_507
timestamp 1644511149
transform 1 0 47748 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_512
timestamp 1644511149
transform 1 0 48208 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_7
timestamp 1644511149
transform 1 0 1748 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_14
timestamp 1644511149
transform 1 0 2392 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_26
timestamp 1644511149
transform 1 0 3496 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_38
timestamp 1644511149
transform 1 0 4600 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_50
timestamp 1644511149
transform 1 0 5704 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_68
timestamp 1644511149
transform 1 0 7360 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_80
timestamp 1644511149
transform 1 0 8464 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_86
timestamp 1644511149
transform 1 0 9016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_90
timestamp 1644511149
transform 1 0 9384 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_103
timestamp 1644511149
transform 1 0 10580 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_122
timestamp 1644511149
transform 1 0 12328 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_126
timestamp 1644511149
transform 1 0 12696 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_131
timestamp 1644511149
transform 1 0 13156 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_143
timestamp 1644511149
transform 1 0 14260 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_147
timestamp 1644511149
transform 1 0 14628 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_155
timestamp 1644511149
transform 1 0 15364 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_162
timestamp 1644511149
transform 1 0 16008 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_180
timestamp 1644511149
transform 1 0 17664 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_184
timestamp 1644511149
transform 1 0 18032 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_201
timestamp 1644511149
transform 1 0 19596 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_205
timestamp 1644511149
transform 1 0 19964 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_210
timestamp 1644511149
transform 1 0 20424 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1644511149
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1644511149
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_235
timestamp 1644511149
transform 1 0 22724 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_259
timestamp 1644511149
transform 1 0 24932 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_271
timestamp 1644511149
transform 1 0 26036 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1644511149
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_281
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_287
timestamp 1644511149
transform 1 0 27508 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_307
timestamp 1644511149
transform 1 0 29348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_319
timestamp 1644511149
transform 1 0 30452 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_332
timestamp 1644511149
transform 1 0 31648 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_353
timestamp 1644511149
transform 1 0 33580 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_362
timestamp 1644511149
transform 1 0 34408 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_43_386
timestamp 1644511149
transform 1 0 36616 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_396
timestamp 1644511149
transform 1 0 37536 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_408
timestamp 1644511149
transform 1 0 38640 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_420
timestamp 1644511149
transform 1 0 39744 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_432
timestamp 1644511149
transform 1 0 40848 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_444
timestamp 1644511149
transform 1 0 41952 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_449
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_461
timestamp 1644511149
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_473
timestamp 1644511149
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_485
timestamp 1644511149
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1644511149
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1644511149
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_505
timestamp 1644511149
transform 1 0 47564 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_513
timestamp 1644511149
transform 1 0 48300 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_24
timestamp 1644511149
transform 1 0 3312 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_101
timestamp 1644511149
transform 1 0 10396 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_115
timestamp 1644511149
transform 1 0 11684 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_119
timestamp 1644511149
transform 1 0 12052 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_125
timestamp 1644511149
transform 1 0 12604 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_136
timestamp 1644511149
transform 1 0 13616 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_158
timestamp 1644511149
transform 1 0 15640 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_186
timestamp 1644511149
transform 1 0 18216 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 1644511149
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_213
timestamp 1644511149
transform 1 0 20700 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_225
timestamp 1644511149
transform 1 0 21804 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_237
timestamp 1644511149
transform 1 0 22908 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_249
timestamp 1644511149
transform 1 0 24012 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_257
timestamp 1644511149
transform 1 0 24748 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_274
timestamp 1644511149
transform 1 0 26312 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_287
timestamp 1644511149
transform 1 0 27508 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_299
timestamp 1644511149
transform 1 0 28612 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1644511149
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_318
timestamp 1644511149
transform 1 0 30360 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_322
timestamp 1644511149
transform 1 0 30728 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_327
timestamp 1644511149
transform 1 0 31188 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_335
timestamp 1644511149
transform 1 0 31924 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_343
timestamp 1644511149
transform 1 0 32660 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_360
timestamp 1644511149
transform 1 0 34224 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_373
timestamp 1644511149
transform 1 0 35420 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_385
timestamp 1644511149
transform 1 0 36524 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_389
timestamp 1644511149
transform 1 0 36892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_411
timestamp 1644511149
transform 1 0 38916 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1644511149
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_421
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_433
timestamp 1644511149
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_445
timestamp 1644511149
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_457
timestamp 1644511149
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1644511149
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1644511149
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_477
timestamp 1644511149
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_489
timestamp 1644511149
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_501
timestamp 1644511149
transform 1 0 47196 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_507
timestamp 1644511149
transform 1 0 47748 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_512
timestamp 1644511149
transform 1 0 48208 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_28
timestamp 1644511149
transform 1 0 3680 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_40
timestamp 1644511149
transform 1 0 4784 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_52
timestamp 1644511149
transform 1 0 5888 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_77
timestamp 1644511149
transform 1 0 8188 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_83
timestamp 1644511149
transform 1 0 8740 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_94
timestamp 1644511149
transform 1 0 9752 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_108
timestamp 1644511149
transform 1 0 11040 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_121
timestamp 1644511149
transform 1 0 12236 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_133
timestamp 1644511149
transform 1 0 13340 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_145
timestamp 1644511149
transform 1 0 14444 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_153
timestamp 1644511149
transform 1 0 15180 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_164
timestamp 1644511149
transform 1 0 16192 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_177
timestamp 1644511149
transform 1 0 17388 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_189
timestamp 1644511149
transform 1 0 18492 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_198
timestamp 1644511149
transform 1 0 19320 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_206
timestamp 1644511149
transform 1 0 20056 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_216
timestamp 1644511149
transform 1 0 20976 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_237
timestamp 1644511149
transform 1 0 22908 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_243
timestamp 1644511149
transform 1 0 23460 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_255
timestamp 1644511149
transform 1 0 24564 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_264
timestamp 1644511149
transform 1 0 25392 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_270
timestamp 1644511149
transform 1 0 25944 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_276
timestamp 1644511149
transform 1 0 26496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_293
timestamp 1644511149
transform 1 0 28060 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_302
timestamp 1644511149
transform 1 0 28888 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_314
timestamp 1644511149
transform 1 0 29992 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_326
timestamp 1644511149
transform 1 0 31096 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_330
timestamp 1644511149
transform 1 0 31464 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_341
timestamp 1644511149
transform 1 0 32476 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_350
timestamp 1644511149
transform 1 0 33304 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_362
timestamp 1644511149
transform 1 0 34408 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_366
timestamp 1644511149
transform 1 0 34776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_372
timestamp 1644511149
transform 1 0 35328 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_384
timestamp 1644511149
transform 1 0 36432 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_417
timestamp 1644511149
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_429
timestamp 1644511149
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1644511149
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1644511149
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_461
timestamp 1644511149
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_473
timestamp 1644511149
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_485
timestamp 1644511149
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1644511149
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1644511149
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_505
timestamp 1644511149
transform 1 0 47564 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_513
timestamp 1644511149
transform 1 0 48300 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_6
timestamp 1644511149
transform 1 0 1656 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_13
timestamp 1644511149
transform 1 0 2300 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_20
timestamp 1644511149
transform 1 0 2944 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_61
timestamp 1644511149
transform 1 0 6716 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_80
timestamp 1644511149
transform 1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_96
timestamp 1644511149
transform 1 0 9936 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_105
timestamp 1644511149
transform 1 0 10764 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_117
timestamp 1644511149
transform 1 0 11868 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_129
timestamp 1644511149
transform 1 0 12972 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_137
timestamp 1644511149
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_153
timestamp 1644511149
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_165
timestamp 1644511149
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_177
timestamp 1644511149
transform 1 0 17388 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_188
timestamp 1644511149
transform 1 0 18400 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_205
timestamp 1644511149
transform 1 0 19964 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_216
timestamp 1644511149
transform 1 0 20976 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_224
timestamp 1644511149
transform 1 0 21712 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_243
timestamp 1644511149
transform 1 0 23460 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1644511149
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_260
timestamp 1644511149
transform 1 0 25024 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_272
timestamp 1644511149
transform 1 0 26128 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_292
timestamp 1644511149
transform 1 0 27968 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_304
timestamp 1644511149
transform 1 0 29072 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_46_317
timestamp 1644511149
transform 1 0 30268 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_323
timestamp 1644511149
transform 1 0 30820 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_332
timestamp 1644511149
transform 1 0 31648 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_340
timestamp 1644511149
transform 1 0 32384 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_352
timestamp 1644511149
transform 1 0 33488 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_389
timestamp 1644511149
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_401
timestamp 1644511149
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1644511149
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1644511149
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_421
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_433
timestamp 1644511149
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_445
timestamp 1644511149
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_457
timestamp 1644511149
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1644511149
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1644511149
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_477
timestamp 1644511149
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_489
timestamp 1644511149
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_501
timestamp 1644511149
transform 1 0 47196 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_507
timestamp 1644511149
transform 1 0 47748 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_515
timestamp 1644511149
transform 1 0 48484 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_11
timestamp 1644511149
transform 1 0 2116 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_75
timestamp 1644511149
transform 1 0 8004 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_84
timestamp 1644511149
transform 1 0 8832 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_98
timestamp 1644511149
transform 1 0 10120 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_121
timestamp 1644511149
transform 1 0 12236 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_133
timestamp 1644511149
transform 1 0 13340 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_137
timestamp 1644511149
transform 1 0 13708 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_143
timestamp 1644511149
transform 1 0 14260 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_150
timestamp 1644511149
transform 1 0 14904 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_162
timestamp 1644511149
transform 1 0 16008 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_174
timestamp 1644511149
transform 1 0 17112 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_186
timestamp 1644511149
transform 1 0 18216 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_198
timestamp 1644511149
transform 1 0 19320 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_210
timestamp 1644511149
transform 1 0 20424 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_222
timestamp 1644511149
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_233
timestamp 1644511149
transform 1 0 22540 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_242
timestamp 1644511149
transform 1 0 23368 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_262
timestamp 1644511149
transform 1 0 25208 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_274
timestamp 1644511149
transform 1 0 26312 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_47_305
timestamp 1644511149
transform 1 0 29164 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_313
timestamp 1644511149
transform 1 0 29900 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_332
timestamp 1644511149
transform 1 0 31648 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_357
timestamp 1644511149
transform 1 0 33948 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_369
timestamp 1644511149
transform 1 0 35052 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_381
timestamp 1644511149
transform 1 0 36156 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_389
timestamp 1644511149
transform 1 0 36892 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_405
timestamp 1644511149
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_417
timestamp 1644511149
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_429
timestamp 1644511149
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1644511149
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1644511149
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_449
timestamp 1644511149
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_461
timestamp 1644511149
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_473
timestamp 1644511149
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_485
timestamp 1644511149
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1644511149
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1644511149
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_47_505
timestamp 1644511149
transform 1 0 47564 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_512
timestamp 1644511149
transform 1 0 48208 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_24
timestamp 1644511149
transform 1 0 3312 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_80
timestamp 1644511149
transform 1 0 8464 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_89
timestamp 1644511149
transform 1 0 9292 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_114
timestamp 1644511149
transform 1 0 11592 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_125
timestamp 1644511149
transform 1 0 12604 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_136
timestamp 1644511149
transform 1 0 13616 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_159
timestamp 1644511149
transform 1 0 15732 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_173
timestamp 1644511149
transform 1 0 17020 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_185
timestamp 1644511149
transform 1 0 18124 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_193
timestamp 1644511149
transform 1 0 18860 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_221
timestamp 1644511149
transform 1 0 21436 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_241
timestamp 1644511149
transform 1 0 23276 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_249
timestamp 1644511149
transform 1 0 24012 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_272
timestamp 1644511149
transform 1 0 26128 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_288
timestamp 1644511149
transform 1 0 27600 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_294
timestamp 1644511149
transform 1 0 28152 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_304
timestamp 1644511149
transform 1 0 29072 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_321
timestamp 1644511149
transform 1 0 30636 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_329
timestamp 1644511149
transform 1 0 31372 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_339
timestamp 1644511149
transform 1 0 32292 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_347
timestamp 1644511149
transform 1 0 33028 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_360
timestamp 1644511149
transform 1 0 34224 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_377
timestamp 1644511149
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_389
timestamp 1644511149
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_401
timestamp 1644511149
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1644511149
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1644511149
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_421
timestamp 1644511149
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_433
timestamp 1644511149
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_445
timestamp 1644511149
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_457
timestamp 1644511149
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1644511149
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1644511149
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_477
timestamp 1644511149
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_489
timestamp 1644511149
transform 1 0 46092 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_512
timestamp 1644511149
transform 1 0 48208 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_28
timestamp 1644511149
transform 1 0 3680 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_35
timestamp 1644511149
transform 1 0 4324 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_47
timestamp 1644511149
transform 1 0 5428 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_89
timestamp 1644511149
transform 1 0 9292 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_98
timestamp 1644511149
transform 1 0 10120 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_110
timestamp 1644511149
transform 1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_130
timestamp 1644511149
transform 1 0 13064 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_139
timestamp 1644511149
transform 1 0 13892 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_147
timestamp 1644511149
transform 1 0 14628 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_155
timestamp 1644511149
transform 1 0 15364 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_164
timestamp 1644511149
transform 1 0 16192 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_185
timestamp 1644511149
transform 1 0 18124 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_205
timestamp 1644511149
transform 1 0 19964 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1644511149
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1644511149
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_233
timestamp 1644511149
transform 1 0 22540 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_250
timestamp 1644511149
transform 1 0 24104 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_270
timestamp 1644511149
transform 1 0 25944 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_278
timestamp 1644511149
transform 1 0 26680 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_288
timestamp 1644511149
transform 1 0 27600 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_297
timestamp 1644511149
transform 1 0 28428 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_305
timestamp 1644511149
transform 1 0 29164 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_318
timestamp 1644511149
transform 1 0 30360 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_330
timestamp 1644511149
transform 1 0 31464 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_349
timestamp 1644511149
transform 1 0 33212 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_353
timestamp 1644511149
transform 1 0 33580 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_370
timestamp 1644511149
transform 1 0 35144 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_382
timestamp 1644511149
transform 1 0 36248 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_386
timestamp 1644511149
transform 1 0 36616 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_417
timestamp 1644511149
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_429
timestamp 1644511149
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1644511149
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1644511149
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_449
timestamp 1644511149
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_461
timestamp 1644511149
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_473
timestamp 1644511149
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_485
timestamp 1644511149
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1644511149
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1644511149
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_508
timestamp 1644511149
transform 1 0 47840 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_6
timestamp 1644511149
transform 1 0 1656 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_13
timestamp 1644511149
transform 1 0 2300 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_20
timestamp 1644511149
transform 1 0 2944 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_88
timestamp 1644511149
transform 1 0 9200 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_96
timestamp 1644511149
transform 1 0 9936 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_107
timestamp 1644511149
transform 1 0 10948 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_119
timestamp 1644511149
transform 1 0 12052 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_127
timestamp 1644511149
transform 1 0 12788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_148
timestamp 1644511149
transform 1 0 14720 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_156
timestamp 1644511149
transform 1 0 15456 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_161
timestamp 1644511149
transform 1 0 15916 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_175
timestamp 1644511149
transform 1 0 17204 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_50_188
timestamp 1644511149
transform 1 0 18400 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_209
timestamp 1644511149
transform 1 0 20332 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_218
timestamp 1644511149
transform 1 0 21160 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_230
timestamp 1644511149
transform 1 0 22264 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_248
timestamp 1644511149
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_261
timestamp 1644511149
transform 1 0 25116 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_269
timestamp 1644511149
transform 1 0 25852 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_281
timestamp 1644511149
transform 1 0 26956 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_297
timestamp 1644511149
transform 1 0 28428 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_305
timestamp 1644511149
transform 1 0 29164 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_321
timestamp 1644511149
transform 1 0 30636 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_332
timestamp 1644511149
transform 1 0 31648 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_340
timestamp 1644511149
transform 1 0 32384 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_347
timestamp 1644511149
transform 1 0 33028 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_360
timestamp 1644511149
transform 1 0 34224 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_402
timestamp 1644511149
transform 1 0 38088 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_414
timestamp 1644511149
transform 1 0 39192 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_421
timestamp 1644511149
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_433
timestamp 1644511149
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_445
timestamp 1644511149
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_457
timestamp 1644511149
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1644511149
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1644511149
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_477
timestamp 1644511149
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_489
timestamp 1644511149
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_501
timestamp 1644511149
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_513
timestamp 1644511149
transform 1 0 48300 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_28
timestamp 1644511149
transform 1 0 3680 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_36
timestamp 1644511149
transform 1 0 4416 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_42
timestamp 1644511149
transform 1 0 4968 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_54
timestamp 1644511149
transform 1 0 6072 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_77
timestamp 1644511149
transform 1 0 8188 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_97
timestamp 1644511149
transform 1 0 10028 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_106
timestamp 1644511149
transform 1 0 10856 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_149
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1644511149
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1644511149
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_177
timestamp 1644511149
transform 1 0 17388 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_183
timestamp 1644511149
transform 1 0 17940 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_191
timestamp 1644511149
transform 1 0 18676 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_211
timestamp 1644511149
transform 1 0 20516 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_215
timestamp 1644511149
transform 1 0 20884 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_220
timestamp 1644511149
transform 1 0 21344 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_235
timestamp 1644511149
transform 1 0 22724 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_243
timestamp 1644511149
transform 1 0 23460 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_255
timestamp 1644511149
transform 1 0 24564 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_267
timestamp 1644511149
transform 1 0 25668 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_303
timestamp 1644511149
transform 1 0 28980 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_311
timestamp 1644511149
transform 1 0 29716 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_323
timestamp 1644511149
transform 1 0 30820 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1644511149
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_349
timestamp 1644511149
transform 1 0 33212 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_369
timestamp 1644511149
transform 1 0 35052 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_381
timestamp 1644511149
transform 1 0 36156 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_389
timestamp 1644511149
transform 1 0 36892 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_417
timestamp 1644511149
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_429
timestamp 1644511149
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1644511149
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1644511149
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_449
timestamp 1644511149
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_461
timestamp 1644511149
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_473
timestamp 1644511149
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_485
timestamp 1644511149
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1644511149
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1644511149
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_505
timestamp 1644511149
transform 1 0 47564 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_512
timestamp 1644511149
transform 1 0 48208 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_7
timestamp 1644511149
transform 1 0 1748 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_11
timestamp 1644511149
transform 1 0 2116 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_17
timestamp 1644511149
transform 1 0 2668 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_21
timestamp 1644511149
transform 1 0 3036 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_91
timestamp 1644511149
transform 1 0 9476 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_115
timestamp 1644511149
transform 1 0 11684 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_124
timestamp 1644511149
transform 1 0 12512 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_135
timestamp 1644511149
transform 1 0 13524 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_162
timestamp 1644511149
transform 1 0 16008 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_170
timestamp 1644511149
transform 1 0 16744 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_182
timestamp 1644511149
transform 1 0 17848 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1644511149
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_205
timestamp 1644511149
transform 1 0 19964 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_214
timestamp 1644511149
transform 1 0 20792 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_225
timestamp 1644511149
transform 1 0 21804 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_234
timestamp 1644511149
transform 1 0 22632 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_248
timestamp 1644511149
transform 1 0 23920 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_265
timestamp 1644511149
transform 1 0 25484 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_273
timestamp 1644511149
transform 1 0 26220 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_290
timestamp 1644511149
transform 1 0 27784 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_299
timestamp 1644511149
transform 1 0 28612 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1644511149
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_327
timestamp 1644511149
transform 1 0 31188 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_335
timestamp 1644511149
transform 1 0 31924 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_341
timestamp 1644511149
transform 1 0 32476 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_354
timestamp 1644511149
transform 1 0 33672 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_362
timestamp 1644511149
transform 1 0 34408 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_377
timestamp 1644511149
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_389
timestamp 1644511149
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_401
timestamp 1644511149
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1644511149
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1644511149
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_421
timestamp 1644511149
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_433
timestamp 1644511149
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_445
timestamp 1644511149
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_457
timestamp 1644511149
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1644511149
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1644511149
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_477
timestamp 1644511149
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_489
timestamp 1644511149
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_501
timestamp 1644511149
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_513
timestamp 1644511149
transform 1 0 48300 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_30
timestamp 1644511149
transform 1 0 3864 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_42
timestamp 1644511149
transform 1 0 4968 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_54
timestamp 1644511149
transform 1 0 6072 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_89
timestamp 1644511149
transform 1 0 9292 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_108
timestamp 1644511149
transform 1 0 11040 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_132
timestamp 1644511149
transform 1 0 13248 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_144
timestamp 1644511149
transform 1 0 14352 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_156
timestamp 1644511149
transform 1 0 15456 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_164
timestamp 1644511149
transform 1 0 16192 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_174
timestamp 1644511149
transform 1 0 17112 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_186
timestamp 1644511149
transform 1 0 18216 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_190
timestamp 1644511149
transform 1 0 18584 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_194
timestamp 1644511149
transform 1 0 18952 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_208
timestamp 1644511149
transform 1 0 20240 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_220
timestamp 1644511149
transform 1 0 21344 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_241
timestamp 1644511149
transform 1 0 23276 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_261
timestamp 1644511149
transform 1 0 25116 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_267
timestamp 1644511149
transform 1 0 25668 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_276
timestamp 1644511149
transform 1 0 26496 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_294
timestamp 1644511149
transform 1 0 28152 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_307
timestamp 1644511149
transform 1 0 29348 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_315
timestamp 1644511149
transform 1 0 30084 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_326
timestamp 1644511149
transform 1 0 31096 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_334
timestamp 1644511149
transform 1 0 31832 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_343
timestamp 1644511149
transform 1 0 32660 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_363
timestamp 1644511149
transform 1 0 34500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_375
timestamp 1644511149
transform 1 0 35604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_387
timestamp 1644511149
transform 1 0 36708 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1644511149
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_405
timestamp 1644511149
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_417
timestamp 1644511149
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_429
timestamp 1644511149
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1644511149
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1644511149
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_449
timestamp 1644511149
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_461
timestamp 1644511149
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_473
timestamp 1644511149
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_485
timestamp 1644511149
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1644511149
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1644511149
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_505
timestamp 1644511149
transform 1 0 47564 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_513
timestamp 1644511149
transform 1 0 48300 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_7
timestamp 1644511149
transform 1 0 1748 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_14
timestamp 1644511149
transform 1 0 2392 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_18
timestamp 1644511149
transform 1 0 2760 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_22
timestamp 1644511149
transform 1 0 3128 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_126
timestamp 1644511149
transform 1 0 12696 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_138
timestamp 1644511149
transform 1 0 13800 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_147
timestamp 1644511149
transform 1 0 14628 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_171
timestamp 1644511149
transform 1 0 16836 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_179
timestamp 1644511149
transform 1 0 17572 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_192
timestamp 1644511149
transform 1 0 18768 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_213
timestamp 1644511149
transform 1 0 20700 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_219
timestamp 1644511149
transform 1 0 21252 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_224
timestamp 1644511149
transform 1 0 21712 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_236
timestamp 1644511149
transform 1 0 22816 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_248
timestamp 1644511149
transform 1 0 23920 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_269
timestamp 1644511149
transform 1 0 25852 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_277
timestamp 1644511149
transform 1 0 26588 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_284
timestamp 1644511149
transform 1 0 27232 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_297
timestamp 1644511149
transform 1 0 28428 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_305
timestamp 1644511149
transform 1 0 29164 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_317
timestamp 1644511149
transform 1 0 30268 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_326
timestamp 1644511149
transform 1 0 31096 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_334
timestamp 1644511149
transform 1 0 31832 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_338
timestamp 1644511149
transform 1 0 32200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_347
timestamp 1644511149
transform 1 0 33028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_359
timestamp 1644511149
transform 1 0 34132 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1644511149
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1644511149
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_389
timestamp 1644511149
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_401
timestamp 1644511149
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1644511149
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1644511149
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_421
timestamp 1644511149
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_433
timestamp 1644511149
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_445
timestamp 1644511149
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_457
timestamp 1644511149
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1644511149
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1644511149
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_477
timestamp 1644511149
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_489
timestamp 1644511149
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_501
timestamp 1644511149
transform 1 0 47196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_512
timestamp 1644511149
transform 1 0 48208 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_9
timestamp 1644511149
transform 1 0 1932 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_31
timestamp 1644511149
transform 1 0 3956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_43
timestamp 1644511149
transform 1 0 5060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_159
timestamp 1644511149
transform 1 0 15732 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_172
timestamp 1644511149
transform 1 0 16928 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_184
timestamp 1644511149
transform 1 0 18032 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_200
timestamp 1644511149
transform 1 0 19504 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_209
timestamp 1644511149
transform 1 0 20332 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1644511149
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1644511149
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_233
timestamp 1644511149
transform 1 0 22540 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_237
timestamp 1644511149
transform 1 0 22908 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_243
timestamp 1644511149
transform 1 0 23460 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_255
timestamp 1644511149
transform 1 0 24564 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_267
timestamp 1644511149
transform 1 0 25668 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_271
timestamp 1644511149
transform 1 0 26036 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_276
timestamp 1644511149
transform 1 0 26496 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_290
timestamp 1644511149
transform 1 0 27784 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_298
timestamp 1644511149
transform 1 0 28520 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_303
timestamp 1644511149
transform 1 0 28980 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_315
timestamp 1644511149
transform 1 0 30084 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_323
timestamp 1644511149
transform 1 0 30820 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1644511149
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_349
timestamp 1644511149
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_361
timestamp 1644511149
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_373
timestamp 1644511149
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1644511149
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1644511149
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_405
timestamp 1644511149
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_417
timestamp 1644511149
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_429
timestamp 1644511149
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1644511149
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1644511149
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_449
timestamp 1644511149
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_461
timestamp 1644511149
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_473
timestamp 1644511149
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_485
timestamp 1644511149
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1644511149
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1644511149
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_505
timestamp 1644511149
transform 1 0 47564 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_512
timestamp 1644511149
transform 1 0 48208 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_14
timestamp 1644511149
transform 1 0 2392 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_21
timestamp 1644511149
transform 1 0 3036 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_157
timestamp 1644511149
transform 1 0 15548 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_162
timestamp 1644511149
transform 1 0 16008 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_174
timestamp 1644511149
transform 1 0 17112 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_182
timestamp 1644511149
transform 1 0 17848 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_192
timestamp 1644511149
transform 1 0 18768 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_213
timestamp 1644511149
transform 1 0 20700 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_225
timestamp 1644511149
transform 1 0 21804 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_237
timestamp 1644511149
transform 1 0 22908 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_243
timestamp 1644511149
transform 1 0 23460 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_248
timestamp 1644511149
transform 1 0 23920 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_269
timestamp 1644511149
transform 1 0 25852 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_281
timestamp 1644511149
transform 1 0 26956 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_298
timestamp 1644511149
transform 1 0 28520 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_306
timestamp 1644511149
transform 1 0 29256 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_313
timestamp 1644511149
transform 1 0 29900 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_330
timestamp 1644511149
transform 1 0 31464 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_334
timestamp 1644511149
transform 1 0 31832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_343
timestamp 1644511149
transform 1 0 32660 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_352
timestamp 1644511149
transform 1 0 33488 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_377
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_389
timestamp 1644511149
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_401
timestamp 1644511149
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1644511149
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1644511149
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_421
timestamp 1644511149
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_433
timestamp 1644511149
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_445
timestamp 1644511149
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_457
timestamp 1644511149
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1644511149
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1644511149
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_477
timestamp 1644511149
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_489
timestamp 1644511149
transform 1 0 46092 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_512
timestamp 1644511149
transform 1 0 48208 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_28
timestamp 1644511149
transform 1 0 3680 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_40
timestamp 1644511149
transform 1 0 4784 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_52
timestamp 1644511149
transform 1 0 5888 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_119
timestamp 1644511149
transform 1 0 12052 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_131
timestamp 1644511149
transform 1 0 13156 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_143
timestamp 1644511149
transform 1 0 14260 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_150
timestamp 1644511149
transform 1 0 14904 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_162
timestamp 1644511149
transform 1 0 16008 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_173
timestamp 1644511149
transform 1 0 17020 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_177
timestamp 1644511149
transform 1 0 17388 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_188
timestamp 1644511149
transform 1 0 18400 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_194
timestamp 1644511149
transform 1 0 18952 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_205
timestamp 1644511149
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1644511149
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1644511149
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_237
timestamp 1644511149
transform 1 0 22908 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_242
timestamp 1644511149
transform 1 0 23368 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_248
timestamp 1644511149
transform 1 0 23920 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_254
timestamp 1644511149
transform 1 0 24472 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_266
timestamp 1644511149
transform 1 0 25576 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_276
timestamp 1644511149
transform 1 0 26496 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_285
timestamp 1644511149
transform 1 0 27324 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_295
timestamp 1644511149
transform 1 0 28244 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_303
timestamp 1644511149
transform 1 0 28980 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_311
timestamp 1644511149
transform 1 0 29716 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_322
timestamp 1644511149
transform 1 0 30728 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_334
timestamp 1644511149
transform 1 0 31832 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_342
timestamp 1644511149
transform 1 0 32568 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_346
timestamp 1644511149
transform 1 0 32936 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_363
timestamp 1644511149
transform 1 0 34500 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_383
timestamp 1644511149
transform 1 0 36340 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1644511149
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_417
timestamp 1644511149
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_429
timestamp 1644511149
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1644511149
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1644511149
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_449
timestamp 1644511149
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_461
timestamp 1644511149
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_473
timestamp 1644511149
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_485
timestamp 1644511149
transform 1 0 45724 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_489
timestamp 1644511149
transform 1 0 46092 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_500
timestamp 1644511149
transform 1 0 47104 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_508
timestamp 1644511149
transform 1 0 47840 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_24
timestamp 1644511149
transform 1 0 3312 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_136
timestamp 1644511149
transform 1 0 13616 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_173
timestamp 1644511149
transform 1 0 17020 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_183
timestamp 1644511149
transform 1 0 17940 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_191
timestamp 1644511149
transform 1 0 18676 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_201
timestamp 1644511149
transform 1 0 19596 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_206
timestamp 1644511149
transform 1 0 20056 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_218
timestamp 1644511149
transform 1 0 21160 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_229
timestamp 1644511149
transform 1 0 22172 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_237
timestamp 1644511149
transform 1 0 22908 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_248
timestamp 1644511149
transform 1 0 23920 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_261
timestamp 1644511149
transform 1 0 25116 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_273
timestamp 1644511149
transform 1 0 26220 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_279
timestamp 1644511149
transform 1 0 26772 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_288
timestamp 1644511149
transform 1 0 27600 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_297
timestamp 1644511149
transform 1 0 28428 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_305
timestamp 1644511149
transform 1 0 29164 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_315
timestamp 1644511149
transform 1 0 30084 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_323
timestamp 1644511149
transform 1 0 30820 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_334
timestamp 1644511149
transform 1 0 31832 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_347
timestamp 1644511149
transform 1 0 33028 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_360
timestamp 1644511149
transform 1 0 34224 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_377
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_389
timestamp 1644511149
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_401
timestamp 1644511149
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1644511149
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1644511149
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_421
timestamp 1644511149
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_433
timestamp 1644511149
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_445
timestamp 1644511149
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_457
timestamp 1644511149
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1644511149
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1644511149
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_477
timestamp 1644511149
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_489
timestamp 1644511149
transform 1 0 46092 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_512
timestamp 1644511149
transform 1 0 48208 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_6
timestamp 1644511149
transform 1 0 1656 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_13
timestamp 1644511149
transform 1 0 2300 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_20
timestamp 1644511149
transform 1 0 2944 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_32
timestamp 1644511149
transform 1 0 4048 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_44
timestamp 1644511149
transform 1 0 5152 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_141
timestamp 1644511149
transform 1 0 14076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_175
timestamp 1644511149
transform 1 0 17204 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_182
timestamp 1644511149
transform 1 0 17848 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_190
timestamp 1644511149
transform 1 0 18584 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_199
timestamp 1644511149
transform 1 0 19412 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_208
timestamp 1644511149
transform 1 0 20240 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_214
timestamp 1644511149
transform 1 0 20792 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_220
timestamp 1644511149
transform 1 0 21344 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_241
timestamp 1644511149
transform 1 0 23276 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_247
timestamp 1644511149
transform 1 0 23828 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_264
timestamp 1644511149
transform 1 0 25392 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_276
timestamp 1644511149
transform 1 0 26496 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_291
timestamp 1644511149
transform 1 0 27876 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_301
timestamp 1644511149
transform 1 0 28796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_315
timestamp 1644511149
transform 1 0 30084 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_323
timestamp 1644511149
transform 1 0 30820 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1644511149
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_343
timestamp 1644511149
transform 1 0 32660 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_353
timestamp 1644511149
transform 1 0 33580 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_365
timestamp 1644511149
transform 1 0 34684 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_377
timestamp 1644511149
transform 1 0 35788 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_389
timestamp 1644511149
transform 1 0 36892 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_417
timestamp 1644511149
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_429
timestamp 1644511149
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1644511149
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1644511149
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_449
timestamp 1644511149
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_461
timestamp 1644511149
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_473
timestamp 1644511149
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_485
timestamp 1644511149
transform 1 0 45724 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_492
timestamp 1644511149
transform 1 0 46368 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_499
timestamp 1644511149
transform 1 0 47012 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1644511149
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_508
timestamp 1644511149
transform 1 0 47840 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_13
timestamp 1644511149
transform 1 0 2300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_25
timestamp 1644511149
transform 1 0 3404 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_177
timestamp 1644511149
transform 1 0 17388 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_184
timestamp 1644511149
transform 1 0 18032 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_213
timestamp 1644511149
transform 1 0 20700 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_60_231
timestamp 1644511149
transform 1 0 22356 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_239
timestamp 1644511149
transform 1 0 23092 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_244
timestamp 1644511149
transform 1 0 23552 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_261
timestamp 1644511149
transform 1 0 25116 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_273
timestamp 1644511149
transform 1 0 26220 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_287
timestamp 1644511149
transform 1 0 27508 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_60_299
timestamp 1644511149
transform 1 0 28612 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1644511149
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_325
timestamp 1644511149
transform 1 0 31004 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_336
timestamp 1644511149
transform 1 0 32016 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_356
timestamp 1644511149
transform 1 0 33856 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_401
timestamp 1644511149
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1644511149
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1644511149
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_421
timestamp 1644511149
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_433
timestamp 1644511149
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_445
timestamp 1644511149
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_457
timestamp 1644511149
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1644511149
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1644511149
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_477
timestamp 1644511149
transform 1 0 44988 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_483
timestamp 1644511149
transform 1 0 45540 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_487
timestamp 1644511149
transform 1 0 45908 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_512
timestamp 1644511149
transform 1 0 48208 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_9
timestamp 1644511149
transform 1 0 1932 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_31
timestamp 1644511149
transform 1 0 3956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_43
timestamp 1644511149
transform 1 0 5060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1644511149
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_189
timestamp 1644511149
transform 1 0 18492 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_206
timestamp 1644511149
transform 1 0 20056 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_215
timestamp 1644511149
transform 1 0 20884 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_229
timestamp 1644511149
transform 1 0 22172 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_237
timestamp 1644511149
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_249
timestamp 1644511149
transform 1 0 24012 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_257
timestamp 1644511149
transform 1 0 24748 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_269
timestamp 1644511149
transform 1 0 25852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_276
timestamp 1644511149
transform 1 0 26496 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_297
timestamp 1644511149
transform 1 0 28428 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_308
timestamp 1644511149
transform 1 0 29440 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_321
timestamp 1644511149
transform 1 0 30636 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1644511149
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1644511149
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_345
timestamp 1644511149
transform 1 0 32844 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_357
timestamp 1644511149
transform 1 0 33948 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_369
timestamp 1644511149
transform 1 0 35052 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_381
timestamp 1644511149
transform 1 0 36156 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_389
timestamp 1644511149
transform 1 0 36892 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_417
timestamp 1644511149
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_429
timestamp 1644511149
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1644511149
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1644511149
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_449
timestamp 1644511149
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_461
timestamp 1644511149
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_473
timestamp 1644511149
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_485
timestamp 1644511149
transform 1 0 45724 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_489
timestamp 1644511149
transform 1 0 46092 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_493
timestamp 1644511149
transform 1 0 46460 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_500
timestamp 1644511149
transform 1 0 47104 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_61_505
timestamp 1644511149
transform 1 0 47564 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_512
timestamp 1644511149
transform 1 0 48208 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_9
timestamp 1644511149
transform 1 0 1932 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_13
timestamp 1644511149
transform 1 0 2300 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_62_22
timestamp 1644511149
transform 1 0 3128 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_165
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_177
timestamp 1644511149
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1644511149
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1644511149
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_205
timestamp 1644511149
transform 1 0 19964 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_213
timestamp 1644511149
transform 1 0 20700 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_219
timestamp 1644511149
transform 1 0 21252 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_227
timestamp 1644511149
transform 1 0 21988 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_231
timestamp 1644511149
transform 1 0 22356 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_240
timestamp 1644511149
transform 1 0 23184 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_261
timestamp 1644511149
transform 1 0 25116 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_275
timestamp 1644511149
transform 1 0 26404 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_288
timestamp 1644511149
transform 1 0 27600 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_297
timestamp 1644511149
transform 1 0 28428 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_305
timestamp 1644511149
transform 1 0 29164 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_317
timestamp 1644511149
transform 1 0 30268 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_325
timestamp 1644511149
transform 1 0 31004 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_333
timestamp 1644511149
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_345
timestamp 1644511149
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1644511149
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1644511149
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_373
timestamp 1644511149
transform 1 0 35420 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_391
timestamp 1644511149
transform 1 0 37076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_403
timestamp 1644511149
transform 1 0 38180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_415
timestamp 1644511149
transform 1 0 39284 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1644511149
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_421
timestamp 1644511149
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_433
timestamp 1644511149
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_445
timestamp 1644511149
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_457
timestamp 1644511149
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1644511149
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1644511149
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_477
timestamp 1644511149
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_489
timestamp 1644511149
transform 1 0 46092 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_512
timestamp 1644511149
transform 1 0 48208 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1644511149
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1644511149
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1644511149
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1644511149
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1644511149
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_189
timestamp 1644511149
transform 1 0 18492 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_206
timestamp 1644511149
transform 1 0 20056 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_215
timestamp 1644511149
transform 1 0 20884 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1644511149
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_242
timestamp 1644511149
transform 1 0 23368 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_246
timestamp 1644511149
transform 1 0 23736 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_263
timestamp 1644511149
transform 1 0 25300 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_275
timestamp 1644511149
transform 1 0 26404 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1644511149
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_289
timestamp 1644511149
transform 1 0 27692 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_297
timestamp 1644511149
transform 1 0 28428 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_301
timestamp 1644511149
transform 1 0 28796 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_310
timestamp 1644511149
transform 1 0 29624 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_330
timestamp 1644511149
transform 1 0 31464 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_341
timestamp 1644511149
transform 1 0 32476 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_351
timestamp 1644511149
transform 1 0 33396 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_371
timestamp 1644511149
transform 1 0 35236 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_380
timestamp 1644511149
transform 1 0 36064 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_417
timestamp 1644511149
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_429
timestamp 1644511149
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1644511149
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1644511149
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_449
timestamp 1644511149
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_461
timestamp 1644511149
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_473
timestamp 1644511149
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_485
timestamp 1644511149
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1644511149
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1644511149
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_508
timestamp 1644511149
transform 1 0 47840 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_11
timestamp 1644511149
transform 1 0 2116 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_23
timestamp 1644511149
transform 1 0 3220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1644511149
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1644511149
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_205
timestamp 1644511149
transform 1 0 19964 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_209
timestamp 1644511149
transform 1 0 20332 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_214
timestamp 1644511149
transform 1 0 20792 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_218
timestamp 1644511149
transform 1 0 21160 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_223
timestamp 1644511149
transform 1 0 21620 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_231
timestamp 1644511149
transform 1 0 22356 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_239
timestamp 1644511149
transform 1 0 23092 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1644511149
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_258
timestamp 1644511149
transform 1 0 24840 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_266
timestamp 1644511149
transform 1 0 25576 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_274
timestamp 1644511149
transform 1 0 26312 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_294
timestamp 1644511149
transform 1 0 28152 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_302
timestamp 1644511149
transform 1 0 28888 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_314
timestamp 1644511149
transform 1 0 29992 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_327
timestamp 1644511149
transform 1 0 31188 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_335
timestamp 1644511149
transform 1 0 31924 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_344
timestamp 1644511149
transform 1 0 32752 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_356
timestamp 1644511149
transform 1 0 33856 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_385
timestamp 1644511149
transform 1 0 36524 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_397
timestamp 1644511149
transform 1 0 37628 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_409
timestamp 1644511149
transform 1 0 38732 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_417
timestamp 1644511149
transform 1 0 39468 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_421
timestamp 1644511149
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_433
timestamp 1644511149
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_445
timestamp 1644511149
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_457
timestamp 1644511149
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1644511149
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1644511149
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_477
timestamp 1644511149
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_489
timestamp 1644511149
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_501
timestamp 1644511149
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_513
timestamp 1644511149
transform 1 0 48300 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_11
timestamp 1644511149
transform 1 0 2116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_23
timestamp 1644511149
transform 1 0 3220 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_35
timestamp 1644511149
transform 1 0 4324 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_47
timestamp 1644511149
transform 1 0 5428 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_149
timestamp 1644511149
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1644511149
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1644511149
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_181
timestamp 1644511149
transform 1 0 17756 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_189
timestamp 1644511149
transform 1 0 18492 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_198
timestamp 1644511149
transform 1 0 19320 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_207
timestamp 1644511149
transform 1 0 20148 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_211
timestamp 1644511149
transform 1 0 20516 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_216
timestamp 1644511149
transform 1 0 20976 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_65_229
timestamp 1644511149
transform 1 0 22172 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_241
timestamp 1644511149
transform 1 0 23276 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_255
timestamp 1644511149
transform 1 0 24564 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_263
timestamp 1644511149
transform 1 0 25300 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_269
timestamp 1644511149
transform 1 0 25852 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_277
timestamp 1644511149
transform 1 0 26588 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_65_281
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_291
timestamp 1644511149
transform 1 0 27876 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_299
timestamp 1644511149
transform 1 0 28612 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_65_306
timestamp 1644511149
transform 1 0 29256 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_318
timestamp 1644511149
transform 1 0 30360 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_330
timestamp 1644511149
transform 1 0 31464 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_65_337
timestamp 1644511149
transform 1 0 32108 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_356
timestamp 1644511149
transform 1 0 33856 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_368
timestamp 1644511149
transform 1 0 34960 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_388
timestamp 1644511149
transform 1 0 36800 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_393
timestamp 1644511149
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_405
timestamp 1644511149
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_417
timestamp 1644511149
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_429
timestamp 1644511149
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1644511149
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1644511149
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_449
timestamp 1644511149
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_461
timestamp 1644511149
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_473
timestamp 1644511149
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_485
timestamp 1644511149
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1644511149
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1644511149
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_505
timestamp 1644511149
transform 1 0 47564 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_513
timestamp 1644511149
transform 1 0 48300 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1644511149
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1644511149
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1644511149
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_165
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_177
timestamp 1644511149
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1644511149
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1644511149
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_213
timestamp 1644511149
transform 1 0 20700 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_221
timestamp 1644511149
transform 1 0 21436 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_232
timestamp 1644511149
transform 1 0 22448 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_240
timestamp 1644511149
transform 1 0 23184 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_263
timestamp 1644511149
transform 1 0 25300 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_275
timestamp 1644511149
transform 1 0 26404 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_287
timestamp 1644511149
transform 1 0 27508 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_295
timestamp 1644511149
transform 1 0 28244 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_304
timestamp 1644511149
transform 1 0 29072 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_325
timestamp 1644511149
transform 1 0 31004 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_337
timestamp 1644511149
transform 1 0 32108 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_348
timestamp 1644511149
transform 1 0 33120 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_360
timestamp 1644511149
transform 1 0 34224 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_365
timestamp 1644511149
transform 1 0 34684 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_378
timestamp 1644511149
transform 1 0 35880 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_398
timestamp 1644511149
transform 1 0 37720 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_410
timestamp 1644511149
transform 1 0 38824 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_418
timestamp 1644511149
transform 1 0 39560 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_421
timestamp 1644511149
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_433
timestamp 1644511149
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_445
timestamp 1644511149
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_457
timestamp 1644511149
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1644511149
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1644511149
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_477
timestamp 1644511149
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_489
timestamp 1644511149
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_501
timestamp 1644511149
transform 1 0 47196 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_507
timestamp 1644511149
transform 1 0 47748 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_512
timestamp 1644511149
transform 1 0 48208 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_9
timestamp 1644511149
transform 1 0 1932 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_31
timestamp 1644511149
transform 1 0 3956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_43
timestamp 1644511149
transform 1 0 5060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1644511149
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1644511149
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_149
timestamp 1644511149
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1644511149
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1644511149
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_181
timestamp 1644511149
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_193
timestamp 1644511149
transform 1 0 18860 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_201
timestamp 1644511149
transform 1 0 19596 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_212
timestamp 1644511149
transform 1 0 20608 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_241
timestamp 1644511149
transform 1 0 23276 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_67_253
timestamp 1644511149
transform 1 0 24380 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_259
timestamp 1644511149
transform 1 0 24932 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_276
timestamp 1644511149
transform 1 0 26496 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_287
timestamp 1644511149
transform 1 0 27508 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_299
timestamp 1644511149
transform 1 0 28612 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_314
timestamp 1644511149
transform 1 0 29992 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_326
timestamp 1644511149
transform 1 0 31096 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_334
timestamp 1644511149
transform 1 0 31832 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_67_337
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_349
timestamp 1644511149
transform 1 0 33212 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_356
timestamp 1644511149
transform 1 0 33856 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_368
timestamp 1644511149
transform 1 0 34960 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_376
timestamp 1644511149
transform 1 0 35696 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_387
timestamp 1644511149
transform 1 0 36708 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1644511149
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_398
timestamp 1644511149
transform 1 0 37720 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_410
timestamp 1644511149
transform 1 0 38824 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_422
timestamp 1644511149
transform 1 0 39928 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_434
timestamp 1644511149
transform 1 0 41032 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_446
timestamp 1644511149
transform 1 0 42136 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_67_449
timestamp 1644511149
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_461
timestamp 1644511149
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_473
timestamp 1644511149
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_485
timestamp 1644511149
transform 1 0 45724 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_493
timestamp 1644511149
transform 1 0 46460 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_67_498
timestamp 1644511149
transform 1 0 46920 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_505
timestamp 1644511149
transform 1 0 47564 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_512
timestamp 1644511149
transform 1 0 48208 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_15
timestamp 1644511149
transform 1 0 2484 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_22
timestamp 1644511149
transform 1 0 3128 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_41
timestamp 1644511149
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_53
timestamp 1644511149
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_65
timestamp 1644511149
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1644511149
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1644511149
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_109
timestamp 1644511149
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_121
timestamp 1644511149
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1644511149
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1644511149
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1644511149
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_165
timestamp 1644511149
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_177
timestamp 1644511149
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1644511149
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1644511149
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_197
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_203
timestamp 1644511149
transform 1 0 19780 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_220
timestamp 1644511149
transform 1 0 21344 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_68_233
timestamp 1644511149
transform 1 0 22540 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_239
timestamp 1644511149
transform 1 0 23092 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_248
timestamp 1644511149
transform 1 0 23920 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_253
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_259
timestamp 1644511149
transform 1 0 24932 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_267
timestamp 1644511149
transform 1 0 25668 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_285
timestamp 1644511149
transform 1 0 27324 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_295
timestamp 1644511149
transform 1 0 28244 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1644511149
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_333
timestamp 1644511149
transform 1 0 31740 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_345
timestamp 1644511149
transform 1 0 32844 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1644511149
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1644511149
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_381
timestamp 1644511149
transform 1 0 36156 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_401
timestamp 1644511149
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1644511149
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1644511149
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_421
timestamp 1644511149
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_433
timestamp 1644511149
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_445
timestamp 1644511149
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_457
timestamp 1644511149
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1644511149
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1644511149
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_477
timestamp 1644511149
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_489
timestamp 1644511149
transform 1 0 46092 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_512
timestamp 1644511149
transform 1 0 48208 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_9
timestamp 1644511149
transform 1 0 1932 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_13
timestamp 1644511149
transform 1 0 2300 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_25
timestamp 1644511149
transform 1 0 3404 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_37
timestamp 1644511149
transform 1 0 4508 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_49
timestamp 1644511149
transform 1 0 5612 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1644511149
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1644511149
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1644511149
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_93
timestamp 1644511149
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1644511149
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1644511149
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_113
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_125
timestamp 1644511149
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_137
timestamp 1644511149
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_149
timestamp 1644511149
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1644511149
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1644511149
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_169
timestamp 1644511149
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_181
timestamp 1644511149
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_193
timestamp 1644511149
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_205
timestamp 1644511149
transform 1 0 19964 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_214
timestamp 1644511149
transform 1 0 20792 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_222
timestamp 1644511149
transform 1 0 21528 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_225
timestamp 1644511149
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_237
timestamp 1644511149
transform 1 0 22908 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_241
timestamp 1644511149
transform 1 0 23276 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_258
timestamp 1644511149
transform 1 0 24840 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_69_272
timestamp 1644511149
transform 1 0 26128 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_281
timestamp 1644511149
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_293
timestamp 1644511149
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_305
timestamp 1644511149
transform 1 0 29164 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_311
timestamp 1644511149
transform 1 0 29716 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_321
timestamp 1644511149
transform 1 0 30636 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_332
timestamp 1644511149
transform 1 0 31648 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_342
timestamp 1644511149
transform 1 0 32568 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_362
timestamp 1644511149
transform 1 0 34408 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_374
timestamp 1644511149
transform 1 0 35512 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_386
timestamp 1644511149
transform 1 0 36616 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_69_393
timestamp 1644511149
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_405
timestamp 1644511149
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_417
timestamp 1644511149
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_429
timestamp 1644511149
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1644511149
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1644511149
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_449
timestamp 1644511149
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_461
timestamp 1644511149
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_473
timestamp 1644511149
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_485
timestamp 1644511149
transform 1 0 45724 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_493
timestamp 1644511149
transform 1 0 46460 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_498
timestamp 1644511149
transform 1 0 46920 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_69_508
timestamp 1644511149
transform 1 0 47840 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_3
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_11
timestamp 1644511149
transform 1 0 2116 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_23
timestamp 1644511149
transform 1 0 3220 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1644511149
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1644511149
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1644511149
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1644511149
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1644511149
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1644511149
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_97
timestamp 1644511149
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_109
timestamp 1644511149
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_121
timestamp 1644511149
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1644511149
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1644511149
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_153
timestamp 1644511149
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_165
timestamp 1644511149
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_177
timestamp 1644511149
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1644511149
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1644511149
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_197
timestamp 1644511149
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_209
timestamp 1644511149
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_221
timestamp 1644511149
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_233
timestamp 1644511149
transform 1 0 22540 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_239
timestamp 1644511149
transform 1 0 23092 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_244
timestamp 1644511149
transform 1 0 23552 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_253
timestamp 1644511149
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_265
timestamp 1644511149
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_277
timestamp 1644511149
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_289
timestamp 1644511149
transform 1 0 27692 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_297
timestamp 1644511149
transform 1 0 28428 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_304
timestamp 1644511149
transform 1 0 29072 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_309
timestamp 1644511149
transform 1 0 29532 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_316
timestamp 1644511149
transform 1 0 30176 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_328
timestamp 1644511149
transform 1 0 31280 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_341
timestamp 1644511149
transform 1 0 32476 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_354
timestamp 1644511149
transform 1 0 33672 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_362
timestamp 1644511149
transform 1 0 34408 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_365
timestamp 1644511149
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_377
timestamp 1644511149
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_389
timestamp 1644511149
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_401
timestamp 1644511149
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1644511149
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1644511149
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_421
timestamp 1644511149
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_433
timestamp 1644511149
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_445
timestamp 1644511149
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_457
timestamp 1644511149
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1644511149
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1644511149
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_477
timestamp 1644511149
transform 1 0 44988 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_483
timestamp 1644511149
transform 1 0 45540 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_487
timestamp 1644511149
transform 1 0 45908 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_512
timestamp 1644511149
transform 1 0 48208 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_3
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_11
timestamp 1644511149
transform 1 0 2116 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_18
timestamp 1644511149
transform 1 0 2760 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_30
timestamp 1644511149
transform 1 0 3864 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_42
timestamp 1644511149
transform 1 0 4968 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_54
timestamp 1644511149
transform 1 0 6072 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1644511149
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_93
timestamp 1644511149
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1644511149
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1644511149
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_125
timestamp 1644511149
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_137
timestamp 1644511149
transform 1 0 13708 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_145
timestamp 1644511149
transform 1 0 14444 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_164
timestamp 1644511149
transform 1 0 16192 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_169
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_181
timestamp 1644511149
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_193
timestamp 1644511149
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_205
timestamp 1644511149
transform 1 0 19964 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_71_219
timestamp 1644511149
transform 1 0 21252 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1644511149
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_230
timestamp 1644511149
transform 1 0 22264 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_242
timestamp 1644511149
transform 1 0 23368 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_251
timestamp 1644511149
transform 1 0 24196 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_263
timestamp 1644511149
transform 1 0 25300 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_275
timestamp 1644511149
transform 1 0 26404 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1644511149
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_281
timestamp 1644511149
transform 1 0 26956 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_71_297
timestamp 1644511149
transform 1 0 28428 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_307
timestamp 1644511149
transform 1 0 29348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_319
timestamp 1644511149
transform 1 0 30452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_331
timestamp 1644511149
transform 1 0 31556 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1644511149
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_337
timestamp 1644511149
transform 1 0 32108 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_355
timestamp 1644511149
transform 1 0 33764 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_367
timestamp 1644511149
transform 1 0 34868 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_379
timestamp 1644511149
transform 1 0 35972 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1644511149
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_393
timestamp 1644511149
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_405
timestamp 1644511149
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_417
timestamp 1644511149
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_429
timestamp 1644511149
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1644511149
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1644511149
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_449
timestamp 1644511149
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_461
timestamp 1644511149
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_473
timestamp 1644511149
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_485
timestamp 1644511149
transform 1 0 45724 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_493
timestamp 1644511149
transform 1 0 46460 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_71_498
timestamp 1644511149
transform 1 0 46920 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_71_505
timestamp 1644511149
transform 1 0 47564 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_512
timestamp 1644511149
transform 1 0 48208 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_24
timestamp 1644511149
transform 1 0 3312 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1644511149
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1644511149
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1644511149
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1644511149
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1644511149
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1644511149
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_97
timestamp 1644511149
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_109
timestamp 1644511149
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_121
timestamp 1644511149
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1644511149
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1644511149
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1644511149
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_153
timestamp 1644511149
transform 1 0 15180 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_178
timestamp 1644511149
transform 1 0 17480 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_190
timestamp 1644511149
transform 1 0 18584 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_72_197
timestamp 1644511149
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_209
timestamp 1644511149
transform 1 0 20332 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_227
timestamp 1644511149
transform 1 0 21988 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_231
timestamp 1644511149
transform 1 0 22356 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_248
timestamp 1644511149
transform 1 0 23920 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_261
timestamp 1644511149
transform 1 0 25116 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_269
timestamp 1644511149
transform 1 0 25852 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_286
timestamp 1644511149
transform 1 0 27416 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_290
timestamp 1644511149
transform 1 0 27784 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_299
timestamp 1644511149
transform 1 0 28612 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1644511149
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_325
timestamp 1644511149
transform 1 0 31004 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_337
timestamp 1644511149
transform 1 0 32108 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_349
timestamp 1644511149
transform 1 0 33212 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_361
timestamp 1644511149
transform 1 0 34316 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_365
timestamp 1644511149
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_377
timestamp 1644511149
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_389
timestamp 1644511149
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_401
timestamp 1644511149
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1644511149
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1644511149
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_421
timestamp 1644511149
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_433
timestamp 1644511149
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_445
timestamp 1644511149
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_457
timestamp 1644511149
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1644511149
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1644511149
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_477
timestamp 1644511149
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_489
timestamp 1644511149
transform 1 0 46092 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_512
timestamp 1644511149
transform 1 0 48208 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_3
timestamp 1644511149
transform 1 0 1380 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_7
timestamp 1644511149
transform 1 0 1748 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_11
timestamp 1644511149
transform 1 0 2116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_23
timestamp 1644511149
transform 1 0 3220 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_35
timestamp 1644511149
transform 1 0 4324 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_47
timestamp 1644511149
transform 1 0 5428 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1644511149
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1644511149
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_93
timestamp 1644511149
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1644511149
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1644511149
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1644511149
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1644511149
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_137
timestamp 1644511149
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_149
timestamp 1644511149
transform 1 0 14812 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_73_160
timestamp 1644511149
transform 1 0 15824 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_169
timestamp 1644511149
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_181
timestamp 1644511149
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_193
timestamp 1644511149
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_205
timestamp 1644511149
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1644511149
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1644511149
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_233
timestamp 1644511149
transform 1 0 22540 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_241
timestamp 1644511149
transform 1 0 23276 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_248
timestamp 1644511149
transform 1 0 23920 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_268
timestamp 1644511149
transform 1 0 25760 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_281
timestamp 1644511149
transform 1 0 26956 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_293
timestamp 1644511149
transform 1 0 28060 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_313
timestamp 1644511149
transform 1 0 29900 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_323
timestamp 1644511149
transform 1 0 30820 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1644511149
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_337
timestamp 1644511149
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_349
timestamp 1644511149
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_361
timestamp 1644511149
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_373
timestamp 1644511149
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1644511149
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1644511149
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_393
timestamp 1644511149
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_405
timestamp 1644511149
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_417
timestamp 1644511149
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_429
timestamp 1644511149
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1644511149
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1644511149
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_449
timestamp 1644511149
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_461
timestamp 1644511149
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_473
timestamp 1644511149
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_485
timestamp 1644511149
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1644511149
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1644511149
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_508
timestamp 1644511149
transform 1 0 47840 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1644511149
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1644511149
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1644511149
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1644511149
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1644511149
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_53
timestamp 1644511149
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_65
timestamp 1644511149
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1644511149
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1644511149
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_85
timestamp 1644511149
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_97
timestamp 1644511149
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_109
timestamp 1644511149
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_121
timestamp 1644511149
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1644511149
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1644511149
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1644511149
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_153
timestamp 1644511149
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_165
timestamp 1644511149
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_177
timestamp 1644511149
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1644511149
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1644511149
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_197
timestamp 1644511149
transform 1 0 19228 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_74_209
timestamp 1644511149
transform 1 0 20332 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_217
timestamp 1644511149
transform 1 0 21068 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_74_236
timestamp 1644511149
transform 1 0 22816 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_242
timestamp 1644511149
transform 1 0 23368 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_248
timestamp 1644511149
transform 1 0 23920 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_74_253
timestamp 1644511149
transform 1 0 24380 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_272
timestamp 1644511149
transform 1 0 26128 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_284
timestamp 1644511149
transform 1 0 27232 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_296
timestamp 1644511149
transform 1 0 28336 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_303
timestamp 1644511149
transform 1 0 28980 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1644511149
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_325
timestamp 1644511149
transform 1 0 31004 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_337
timestamp 1644511149
transform 1 0 32108 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_349
timestamp 1644511149
transform 1 0 33212 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_74_361
timestamp 1644511149
transform 1 0 34316 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_365
timestamp 1644511149
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_377
timestamp 1644511149
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_389
timestamp 1644511149
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_401
timestamp 1644511149
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1644511149
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1644511149
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_421
timestamp 1644511149
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_433
timestamp 1644511149
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_445
timestamp 1644511149
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_457
timestamp 1644511149
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1644511149
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1644511149
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_477
timestamp 1644511149
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_489
timestamp 1644511149
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_501
timestamp 1644511149
transform 1 0 47196 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_507
timestamp 1644511149
transform 1 0 47748 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_512
timestamp 1644511149
transform 1 0 48208 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_3
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_13
timestamp 1644511149
transform 1 0 2300 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_25
timestamp 1644511149
transform 1 0 3404 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_37
timestamp 1644511149
transform 1 0 4508 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_49
timestamp 1644511149
transform 1 0 5612 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1644511149
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1644511149
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1644511149
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_93
timestamp 1644511149
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1644511149
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1644511149
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_113
timestamp 1644511149
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_125
timestamp 1644511149
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_137
timestamp 1644511149
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_149
timestamp 1644511149
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1644511149
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1644511149
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_169
timestamp 1644511149
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_181
timestamp 1644511149
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_193
timestamp 1644511149
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_205
timestamp 1644511149
transform 1 0 19964 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_215
timestamp 1644511149
transform 1 0 20884 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1644511149
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_75_225
timestamp 1644511149
transform 1 0 21804 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_231
timestamp 1644511149
transform 1 0 22356 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_243
timestamp 1644511149
transform 1 0 23460 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_251
timestamp 1644511149
transform 1 0 24196 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_75_261
timestamp 1644511149
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1644511149
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1644511149
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_287
timestamp 1644511149
transform 1 0 27508 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_299
timestamp 1644511149
transform 1 0 28612 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_311
timestamp 1644511149
transform 1 0 29716 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_323
timestamp 1644511149
transform 1 0 30820 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1644511149
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_337
timestamp 1644511149
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_349
timestamp 1644511149
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_361
timestamp 1644511149
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_373
timestamp 1644511149
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1644511149
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1644511149
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_393
timestamp 1644511149
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_405
timestamp 1644511149
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_417
timestamp 1644511149
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_429
timestamp 1644511149
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1644511149
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1644511149
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_449
timestamp 1644511149
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_461
timestamp 1644511149
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_473
timestamp 1644511149
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_485
timestamp 1644511149
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_500
timestamp 1644511149
transform 1 0 47104 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_75_505
timestamp 1644511149
transform 1 0 47564 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_512
timestamp 1644511149
transform 1 0 48208 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_3
timestamp 1644511149
transform 1 0 1380 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_13
timestamp 1644511149
transform 1 0 2300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_25
timestamp 1644511149
transform 1 0 3404 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1644511149
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1644511149
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1644511149
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_65
timestamp 1644511149
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1644511149
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1644511149
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_85
timestamp 1644511149
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_97
timestamp 1644511149
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_109
timestamp 1644511149
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_121
timestamp 1644511149
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1644511149
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1644511149
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_141
timestamp 1644511149
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_153
timestamp 1644511149
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_165
timestamp 1644511149
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_177
timestamp 1644511149
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1644511149
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1644511149
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_197
timestamp 1644511149
transform 1 0 19228 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_205
timestamp 1644511149
transform 1 0 19964 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_212
timestamp 1644511149
transform 1 0 20608 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_224
timestamp 1644511149
transform 1 0 21712 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_236
timestamp 1644511149
transform 1 0 22816 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_76_248
timestamp 1644511149
transform 1 0 23920 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_262
timestamp 1644511149
transform 1 0 25208 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_274
timestamp 1644511149
transform 1 0 26312 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_286
timestamp 1644511149
transform 1 0 27416 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_298
timestamp 1644511149
transform 1 0 28520 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_306
timestamp 1644511149
transform 1 0 29256 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_76_309
timestamp 1644511149
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_321
timestamp 1644511149
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_333
timestamp 1644511149
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_345
timestamp 1644511149
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1644511149
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1644511149
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_365
timestamp 1644511149
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_377
timestamp 1644511149
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_389
timestamp 1644511149
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_401
timestamp 1644511149
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1644511149
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1644511149
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_421
timestamp 1644511149
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_433
timestamp 1644511149
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_445
timestamp 1644511149
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_457
timestamp 1644511149
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1644511149
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1644511149
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_477
timestamp 1644511149
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_489
timestamp 1644511149
transform 1 0 46092 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_512
timestamp 1644511149
transform 1 0 48208 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_3
timestamp 1644511149
transform 1 0 1380 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_9
timestamp 1644511149
transform 1 0 1932 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_31
timestamp 1644511149
transform 1 0 3956 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_43
timestamp 1644511149
transform 1 0 5060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1644511149
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1644511149
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1644511149
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1644511149
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_93
timestamp 1644511149
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1644511149
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1644511149
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_113
timestamp 1644511149
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_125
timestamp 1644511149
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_137
timestamp 1644511149
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_149
timestamp 1644511149
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1644511149
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1644511149
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_169
timestamp 1644511149
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_181
timestamp 1644511149
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_193
timestamp 1644511149
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_205
timestamp 1644511149
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1644511149
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1644511149
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_225
timestamp 1644511149
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_237
timestamp 1644511149
transform 1 0 22908 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_243
timestamp 1644511149
transform 1 0 23460 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_260
timestamp 1644511149
transform 1 0 25024 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_272
timestamp 1644511149
transform 1 0 26128 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_281
timestamp 1644511149
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_293
timestamp 1644511149
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_305
timestamp 1644511149
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_317
timestamp 1644511149
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1644511149
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1644511149
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_337
timestamp 1644511149
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_349
timestamp 1644511149
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_361
timestamp 1644511149
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_373
timestamp 1644511149
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1644511149
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1644511149
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_393
timestamp 1644511149
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_405
timestamp 1644511149
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_417
timestamp 1644511149
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_429
timestamp 1644511149
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1644511149
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1644511149
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_449
timestamp 1644511149
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_461
timestamp 1644511149
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_473
timestamp 1644511149
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_485
timestamp 1644511149
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_500
timestamp 1644511149
transform 1 0 47104 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_508
timestamp 1644511149
transform 1 0 47840 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_78_3
timestamp 1644511149
transform 1 0 1380 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_78_14
timestamp 1644511149
transform 1 0 2392 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_78_23
timestamp 1644511149
transform 1 0 3220 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1644511149
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1644511149
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_41
timestamp 1644511149
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_53
timestamp 1644511149
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_65
timestamp 1644511149
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1644511149
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1644511149
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_88
timestamp 1644511149
transform 1 0 9200 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_100
timestamp 1644511149
transform 1 0 10304 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_112
timestamp 1644511149
transform 1 0 11408 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_124
timestamp 1644511149
transform 1 0 12512 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_136
timestamp 1644511149
transform 1 0 13616 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1644511149
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_153
timestamp 1644511149
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_165
timestamp 1644511149
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_177
timestamp 1644511149
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1644511149
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1644511149
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_197
timestamp 1644511149
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_209
timestamp 1644511149
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_221
timestamp 1644511149
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_233
timestamp 1644511149
transform 1 0 22540 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_78_248
timestamp 1644511149
transform 1 0 23920 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_253
timestamp 1644511149
transform 1 0 24380 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_277
timestamp 1644511149
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_289
timestamp 1644511149
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1644511149
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1644511149
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_309
timestamp 1644511149
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_321
timestamp 1644511149
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_333
timestamp 1644511149
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_345
timestamp 1644511149
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1644511149
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1644511149
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_365
timestamp 1644511149
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_377
timestamp 1644511149
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_389
timestamp 1644511149
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_401
timestamp 1644511149
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1644511149
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1644511149
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_421
timestamp 1644511149
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_433
timestamp 1644511149
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_445
timestamp 1644511149
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_457
timestamp 1644511149
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1644511149
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1644511149
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_78_477
timestamp 1644511149
transform 1 0 44988 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_483
timestamp 1644511149
transform 1 0 45540 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_487
timestamp 1644511149
transform 1 0 45908 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_512
timestamp 1644511149
transform 1 0 48208 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_3
timestamp 1644511149
transform 1 0 1380 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_13
timestamp 1644511149
transform 1 0 2300 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_20
timestamp 1644511149
transform 1 0 2944 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_32
timestamp 1644511149
transform 1 0 4048 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_44
timestamp 1644511149
transform 1 0 5152 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1644511149
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_69
timestamp 1644511149
transform 1 0 7452 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_73
timestamp 1644511149
transform 1 0 7820 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_95
timestamp 1644511149
transform 1 0 9844 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_107
timestamp 1644511149
transform 1 0 10948 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1644511149
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_113
timestamp 1644511149
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_125
timestamp 1644511149
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_137
timestamp 1644511149
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_149
timestamp 1644511149
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1644511149
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1644511149
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_169
timestamp 1644511149
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_181
timestamp 1644511149
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_193
timestamp 1644511149
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_205
timestamp 1644511149
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1644511149
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1644511149
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_225
timestamp 1644511149
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_237
timestamp 1644511149
transform 1 0 22908 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_243
timestamp 1644511149
transform 1 0 23460 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_260
timestamp 1644511149
transform 1 0 25024 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_272
timestamp 1644511149
transform 1 0 26128 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_281
timestamp 1644511149
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_293
timestamp 1644511149
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_305
timestamp 1644511149
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_317
timestamp 1644511149
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1644511149
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1644511149
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_337
timestamp 1644511149
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_349
timestamp 1644511149
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_361
timestamp 1644511149
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_373
timestamp 1644511149
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1644511149
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1644511149
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_393
timestamp 1644511149
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_405
timestamp 1644511149
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_417
timestamp 1644511149
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_429
timestamp 1644511149
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1644511149
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1644511149
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_449
timestamp 1644511149
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_461
timestamp 1644511149
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_473
timestamp 1644511149
transform 1 0 44620 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_479
timestamp 1644511149
transform 1 0 45172 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_486
timestamp 1644511149
transform 1 0 45816 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_493
timestamp 1644511149
transform 1 0 46460 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_500
timestamp 1644511149
transform 1 0 47104 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_508
timestamp 1644511149
transform 1 0 47840 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_80_24
timestamp 1644511149
transform 1 0 3312 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_29
timestamp 1644511149
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_41
timestamp 1644511149
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_53
timestamp 1644511149
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_65
timestamp 1644511149
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1644511149
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1644511149
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_85
timestamp 1644511149
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_97
timestamp 1644511149
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_109
timestamp 1644511149
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_121
timestamp 1644511149
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1644511149
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1644511149
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_141
timestamp 1644511149
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_153
timestamp 1644511149
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_165
timestamp 1644511149
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_177
timestamp 1644511149
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1644511149
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1644511149
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_197
timestamp 1644511149
transform 1 0 19228 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_204
timestamp 1644511149
transform 1 0 19872 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_216
timestamp 1644511149
transform 1 0 20976 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_228
timestamp 1644511149
transform 1 0 22080 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_240
timestamp 1644511149
transform 1 0 23184 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_253
timestamp 1644511149
transform 1 0 24380 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_259
timestamp 1644511149
transform 1 0 24932 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_272
timestamp 1644511149
transform 1 0 26128 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_284
timestamp 1644511149
transform 1 0 27232 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_296
timestamp 1644511149
transform 1 0 28336 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_309
timestamp 1644511149
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_321
timestamp 1644511149
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_333
timestamp 1644511149
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_345
timestamp 1644511149
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1644511149
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1644511149
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_365
timestamp 1644511149
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_377
timestamp 1644511149
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_389
timestamp 1644511149
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_401
timestamp 1644511149
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_413
timestamp 1644511149
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1644511149
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_421
timestamp 1644511149
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_433
timestamp 1644511149
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_445
timestamp 1644511149
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_457
timestamp 1644511149
transform 1 0 43148 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_465
timestamp 1644511149
transform 1 0 43884 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_471
timestamp 1644511149
transform 1 0 44436 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1644511149
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_480
timestamp 1644511149
transform 1 0 45264 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_487
timestamp 1644511149
transform 1 0 45908 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_512
timestamp 1644511149
transform 1 0 48208 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_7
timestamp 1644511149
transform 1 0 1748 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_14
timestamp 1644511149
transform 1 0 2392 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_21
timestamp 1644511149
transform 1 0 3036 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_28
timestamp 1644511149
transform 1 0 3680 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_35
timestamp 1644511149
transform 1 0 4324 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_47
timestamp 1644511149
transform 1 0 5428 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1644511149
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1644511149
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_69
timestamp 1644511149
transform 1 0 7452 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_73
timestamp 1644511149
transform 1 0 7820 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_77
timestamp 1644511149
transform 1 0 8188 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_89
timestamp 1644511149
transform 1 0 9292 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_101
timestamp 1644511149
transform 1 0 10396 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_109
timestamp 1644511149
transform 1 0 11132 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_113
timestamp 1644511149
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_125
timestamp 1644511149
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_137
timestamp 1644511149
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_149
timestamp 1644511149
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1644511149
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1644511149
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_169
timestamp 1644511149
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_181
timestamp 1644511149
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_193
timestamp 1644511149
transform 1 0 18860 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_220
timestamp 1644511149
transform 1 0 21344 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_225
timestamp 1644511149
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_237
timestamp 1644511149
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_249
timestamp 1644511149
transform 1 0 24012 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_255
timestamp 1644511149
transform 1 0 24564 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_276
timestamp 1644511149
transform 1 0 26496 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_281
timestamp 1644511149
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_296
timestamp 1644511149
transform 1 0 28336 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_308
timestamp 1644511149
transform 1 0 29440 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_320
timestamp 1644511149
transform 1 0 30544 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_332
timestamp 1644511149
transform 1 0 31648 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_337
timestamp 1644511149
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_349
timestamp 1644511149
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_361
timestamp 1644511149
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_373
timestamp 1644511149
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1644511149
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1644511149
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_393
timestamp 1644511149
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_405
timestamp 1644511149
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_417
timestamp 1644511149
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_429
timestamp 1644511149
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1644511149
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1644511149
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_449
timestamp 1644511149
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_461
timestamp 1644511149
transform 1 0 43516 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_468
timestamp 1644511149
transform 1 0 44160 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_475
timestamp 1644511149
transform 1 0 44804 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_500
timestamp 1644511149
transform 1 0 47104 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_508
timestamp 1644511149
transform 1 0 47840 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_82_24
timestamp 1644511149
transform 1 0 3312 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_32
timestamp 1644511149
transform 1 0 4048 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_39
timestamp 1644511149
transform 1 0 4692 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_50
timestamp 1644511149
transform 1 0 5704 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_62
timestamp 1644511149
transform 1 0 6808 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_74
timestamp 1644511149
transform 1 0 7912 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_82
timestamp 1644511149
transform 1 0 8648 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_88
timestamp 1644511149
transform 1 0 9200 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_100
timestamp 1644511149
transform 1 0 10304 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_112
timestamp 1644511149
transform 1 0 11408 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_124
timestamp 1644511149
transform 1 0 12512 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_136
timestamp 1644511149
transform 1 0 13616 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_141
timestamp 1644511149
transform 1 0 14076 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_146
timestamp 1644511149
transform 1 0 14536 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_158
timestamp 1644511149
transform 1 0 15640 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_170
timestamp 1644511149
transform 1 0 16744 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_182
timestamp 1644511149
transform 1 0 17848 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_194
timestamp 1644511149
transform 1 0 18952 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_197
timestamp 1644511149
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_209
timestamp 1644511149
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_221
timestamp 1644511149
transform 1 0 21436 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_228
timestamp 1644511149
transform 1 0 22080 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_240
timestamp 1644511149
transform 1 0 23184 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_256
timestamp 1644511149
transform 1 0 24656 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_280
timestamp 1644511149
transform 1 0 26864 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_293
timestamp 1644511149
transform 1 0 28060 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_300
timestamp 1644511149
transform 1 0 28704 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_309
timestamp 1644511149
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_321
timestamp 1644511149
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_333
timestamp 1644511149
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_345
timestamp 1644511149
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 1644511149
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1644511149
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_365
timestamp 1644511149
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_377
timestamp 1644511149
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_389
timestamp 1644511149
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_401
timestamp 1644511149
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1644511149
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1644511149
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_421
timestamp 1644511149
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_433
timestamp 1644511149
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_445
timestamp 1644511149
transform 1 0 42044 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_82_456
timestamp 1644511149
transform 1 0 43056 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_465
timestamp 1644511149
transform 1 0 43884 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_472
timestamp 1644511149
transform 1 0 44528 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_477
timestamp 1644511149
transform 1 0 44988 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_482
timestamp 1644511149
transform 1 0 45448 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_490
timestamp 1644511149
transform 1 0 46184 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_512
timestamp 1644511149
transform 1 0 48208 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_6
timestamp 1644511149
transform 1 0 1656 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_16
timestamp 1644511149
transform 1 0 2576 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_83_23
timestamp 1644511149
transform 1 0 3220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_83_32
timestamp 1644511149
transform 1 0 4048 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_83_42
timestamp 1644511149
transform 1 0 4968 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_83_49
timestamp 1644511149
transform 1 0 5612 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1644511149
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_57
timestamp 1644511149
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_90
timestamp 1644511149
transform 1 0 9384 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_94
timestamp 1644511149
transform 1 0 9752 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_98
timestamp 1644511149
transform 1 0 10120 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_83_110
timestamp 1644511149
transform 1 0 11224 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_83_113
timestamp 1644511149
transform 1 0 11500 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_117
timestamp 1644511149
transform 1 0 11868 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_129
timestamp 1644511149
transform 1 0 12972 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_141
timestamp 1644511149
transform 1 0 14076 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_83_148
timestamp 1644511149
transform 1 0 14720 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_160
timestamp 1644511149
transform 1 0 15824 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_83_172
timestamp 1644511149
transform 1 0 16928 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_83_179
timestamp 1644511149
transform 1 0 17572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_191
timestamp 1644511149
transform 1 0 18676 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_199
timestamp 1644511149
transform 1 0 19412 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_83_204
timestamp 1644511149
transform 1 0 19872 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_83_216
timestamp 1644511149
transform 1 0 20976 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_220
timestamp 1644511149
transform 1 0 21344 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_246
timestamp 1644511149
transform 1 0 23736 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_83_253
timestamp 1644511149
transform 1 0 24380 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_259
timestamp 1644511149
transform 1 0 24932 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_276
timestamp 1644511149
transform 1 0 26496 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_83_284
timestamp 1644511149
transform 1 0 27232 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_292
timestamp 1644511149
transform 1 0 27968 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_314
timestamp 1644511149
transform 1 0 29992 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_83_321
timestamp 1644511149
transform 1 0 30636 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_83_333
timestamp 1644511149
transform 1 0 31740 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_83_340
timestamp 1644511149
transform 1 0 32384 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_83_351
timestamp 1644511149
transform 1 0 33396 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_376
timestamp 1644511149
transform 1 0 35696 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_83_383
timestamp 1644511149
transform 1 0 36340 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1644511149
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_393
timestamp 1644511149
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_405
timestamp 1644511149
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_83_417
timestamp 1644511149
transform 1 0 39468 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_421
timestamp 1644511149
transform 1 0 39836 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_425
timestamp 1644511149
transform 1 0 40204 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_429
timestamp 1644511149
transform 1 0 40572 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_433
timestamp 1644511149
transform 1 0 40940 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_437
timestamp 1644511149
transform 1 0 41308 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_444
timestamp 1644511149
transform 1 0 41952 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_83_449
timestamp 1644511149
transform 1 0 42412 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_83_454
timestamp 1644511149
transform 1 0 42872 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_460
timestamp 1644511149
transform 1 0 43424 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_464
timestamp 1644511149
transform 1 0 43792 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_489
timestamp 1644511149
transform 1 0 46092 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_493
timestamp 1644511149
transform 1 0 46460 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_500
timestamp 1644511149
transform 1 0 47104 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_505
timestamp 1644511149
transform 1 0 47564 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_512
timestamp 1644511149
transform 1 0 48208 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_24
timestamp 1644511149
transform 1 0 3312 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_29
timestamp 1644511149
transform 1 0 3772 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_84_37
timestamp 1644511149
transform 1 0 4508 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_45
timestamp 1644511149
transform 1 0 5244 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_67
timestamp 1644511149
transform 1 0 7268 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_84_74
timestamp 1644511149
transform 1 0 7912 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_82
timestamp 1644511149
transform 1 0 8648 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_84_85
timestamp 1644511149
transform 1 0 8924 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_89
timestamp 1644511149
transform 1 0 9292 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_114
timestamp 1644511149
transform 1 0 11592 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_84_121
timestamp 1644511149
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1644511149
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1644511149
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_141
timestamp 1644511149
transform 1 0 14076 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_166
timestamp 1644511149
transform 1 0 16376 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_191
timestamp 1644511149
transform 1 0 18676 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1644511149
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_197
timestamp 1644511149
transform 1 0 19228 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_84_226
timestamp 1644511149
transform 1 0 21896 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_240
timestamp 1644511149
transform 1 0 23184 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_247
timestamp 1644511149
transform 1 0 23828 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1644511149
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_253
timestamp 1644511149
transform 1 0 24380 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_257
timestamp 1644511149
transform 1 0 24748 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_264
timestamp 1644511149
transform 1 0 25392 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_289
timestamp 1644511149
transform 1 0 27692 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_296
timestamp 1644511149
transform 1 0 28336 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_300
timestamp 1644511149
transform 1 0 28704 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_304
timestamp 1644511149
transform 1 0 29072 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_84_309
timestamp 1644511149
transform 1 0 29532 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_84_318
timestamp 1644511149
transform 1 0 30360 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_325
timestamp 1644511149
transform 1 0 31004 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_84_350
timestamp 1644511149
transform 1 0 33304 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_84_359
timestamp 1644511149
transform 1 0 34132 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 1644511149
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_365
timestamp 1644511149
transform 1 0 34684 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_84_373
timestamp 1644511149
transform 1 0 35420 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_84_379
timestamp 1644511149
transform 1 0 35972 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_404
timestamp 1644511149
transform 1 0 38272 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_84_411
timestamp 1644511149
transform 1 0 38916 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1644511149
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_424
timestamp 1644511149
transform 1 0 40112 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_432
timestamp 1644511149
transform 1 0 40848 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_84_455
timestamp 1644511149
transform 1 0 42964 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_463
timestamp 1644511149
transform 1 0 43700 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1644511149
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1644511149
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_481
timestamp 1644511149
transform 1 0 45356 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_489
timestamp 1644511149
transform 1 0 46092 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_84_512
timestamp 1644511149
transform 1 0 48208 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_3
timestamp 1644511149
transform 1 0 1380 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_25
timestamp 1644511149
transform 1 0 3404 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_85_50
timestamp 1644511149
transform 1 0 5704 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_85_57
timestamp 1644511149
transform 1 0 6348 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_85_81
timestamp 1644511149
transform 1 0 8556 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_85_106
timestamp 1644511149
transform 1 0 10856 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_85_134
timestamp 1644511149
transform 1 0 13432 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_85_150
timestamp 1644511149
transform 1 0 14904 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_164
timestamp 1644511149
transform 1 0 16192 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_190
timestamp 1644511149
transform 1 0 18584 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_202
timestamp 1644511149
transform 1 0 19688 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_85_209
timestamp 1644511149
transform 1 0 20332 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_85_220
timestamp 1644511149
transform 1 0 21344 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_85_225
timestamp 1644511149
transform 1 0 21804 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_85_231
timestamp 1644511149
transform 1 0 22356 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_85_256
timestamp 1644511149
transform 1 0 24656 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_85_265
timestamp 1644511149
transform 1 0 25484 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_85_273
timestamp 1644511149
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1644511149
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_281
timestamp 1644511149
transform 1 0 26956 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_85_289
timestamp 1644511149
transform 1 0 27692 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_85_301
timestamp 1644511149
transform 1 0 28796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_85_326
timestamp 1644511149
transform 1 0 31096 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_85_334
timestamp 1644511149
transform 1 0 31832 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_85_358
timestamp 1644511149
transform 1 0 34040 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_85_366
timestamp 1644511149
transform 1 0 34776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_388
timestamp 1644511149
transform 1 0 36800 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_85_396
timestamp 1644511149
transform 1 0 37536 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_85_404
timestamp 1644511149
transform 1 0 38272 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_408
timestamp 1644511149
transform 1 0 38640 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_433
timestamp 1644511149
transform 1 0 40940 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_437
timestamp 1644511149
transform 1 0 41308 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_444
timestamp 1644511149
transform 1 0 41952 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_85_449
timestamp 1644511149
transform 1 0 42412 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_85_472
timestamp 1644511149
transform 1 0 44528 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_85_497
timestamp 1644511149
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1644511149
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_85_505
timestamp 1644511149
transform 1 0 47564 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_512
timestamp 1644511149
transform 1 0 48208 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_3
timestamp 1644511149
transform 1 0 1380 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_13
timestamp 1644511149
transform 1 0 2300 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_17
timestamp 1644511149
transform 1 0 2668 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_24
timestamp 1644511149
transform 1 0 3312 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_50
timestamp 1644511149
transform 1 0 5704 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_86_57
timestamp 1644511149
transform 1 0 6348 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_67
timestamp 1644511149
transform 1 0 7268 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_86_74
timestamp 1644511149
transform 1 0 7912 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_82
timestamp 1644511149
transform 1 0 8648 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_86_85
timestamp 1644511149
transform 1 0 8924 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_89
timestamp 1644511149
transform 1 0 9292 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_96
timestamp 1644511149
transform 1 0 9936 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_86_103
timestamp 1644511149
transform 1 0 10580 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_111
timestamp 1644511149
transform 1 0 11316 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_113
timestamp 1644511149
transform 1 0 11500 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_121
timestamp 1644511149
transform 1 0 12236 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_125
timestamp 1644511149
transform 1 0 12604 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_136
timestamp 1644511149
transform 1 0 13616 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_86_151
timestamp 1644511149
transform 1 0 14996 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_159
timestamp 1644511149
transform 1 0 15732 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_86_164
timestamp 1644511149
transform 1 0 16192 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_86_172
timestamp 1644511149
transform 1 0 16928 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_180
timestamp 1644511149
transform 1 0 17664 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_86_192
timestamp 1644511149
transform 1 0 18768 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_197
timestamp 1644511149
transform 1 0 19228 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_202
timestamp 1644511149
transform 1 0 19688 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_210
timestamp 1644511149
transform 1 0 20424 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_216
timestamp 1644511149
transform 1 0 20976 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_220
timestamp 1644511149
transform 1 0 21344 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_225
timestamp 1644511149
transform 1 0 21804 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_86_248
timestamp 1644511149
transform 1 0 23920 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_274
timestamp 1644511149
transform 1 0 26312 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_86_302
timestamp 1644511149
transform 1 0 28888 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_86_309
timestamp 1644511149
transform 1 0 29532 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_86_332
timestamp 1644511149
transform 1 0 31648 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_340
timestamp 1644511149
transform 1 0 32384 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_86_347
timestamp 1644511149
transform 1 0 33028 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_359
timestamp 1644511149
transform 1 0 34132 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1644511149
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_365
timestamp 1644511149
transform 1 0 34684 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_86_373
timestamp 1644511149
transform 1 0 35420 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_86_379
timestamp 1644511149
transform 1 0 35972 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_391
timestamp 1644511149
transform 1 0 37076 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_393
timestamp 1644511149
transform 1 0 37260 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_401
timestamp 1644511149
transform 1 0 37996 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_86_406
timestamp 1644511149
transform 1 0 38456 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_86_416
timestamp 1644511149
transform 1 0 39376 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_442
timestamp 1644511149
transform 1 0 41768 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_86_449
timestamp 1644511149
transform 1 0 42412 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_86_472
timestamp 1644511149
transform 1 0 44528 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_477
timestamp 1644511149
transform 1 0 44988 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_86_500
timestamp 1644511149
transform 1 0 47104 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_505
timestamp 1644511149
transform 1 0 47564 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_512
timestamp 1644511149
transform 1 0 48208 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 48852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 48852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 48852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 48852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 48852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 48852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 48852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 48852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 48852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 48852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 48852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 48852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 48852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 48852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 48852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 48852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 48852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 48852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 48852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 48852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 48852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 48852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 48852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 48852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 48852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 48852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 48852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 48852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 48852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 48852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 48852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 48852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 48852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 48852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 48852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 48852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 48852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 48852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 48852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 48852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 48852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 48852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 48852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 48852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 48852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 48852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 48852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 48852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 48852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 48852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 48852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 48852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 48852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 48852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 48852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 48852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 48852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 48852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 48852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 48852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 48852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 48852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 48852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 48852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 48852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 48852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 48852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 48852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 48852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 48852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 48852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 48852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 48852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 48852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 48852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 48852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1644511149
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1644511149
transform -1 0 48852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1644511149
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1644511149
transform -1 0 48852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1644511149
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1644511149
transform -1 0 48852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1644511149
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1644511149
transform -1 0 48852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1644511149
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1644511149
transform -1 0 48852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1644511149
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1644511149
transform -1 0 48852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1644511149
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1644511149
transform -1 0 48852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1644511149
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1644511149
transform -1 0 48852 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1644511149
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1644511149
transform -1 0 48852 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1644511149
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1644511149
transform -1 0 48852 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1644511149
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1644511149
transform -1 0 48852 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1644511149
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1644511149
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1644511149
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1644511149
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1644511149
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1644511149
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1644511149
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1644511149
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1644511149
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1644511149
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1644511149
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1644511149
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1644511149
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1644511149
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1644511149
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1644511149
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1644511149
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1644511149
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1644511149
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1644511149
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1644511149
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1644511149
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1644511149
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1644511149
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1644511149
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1644511149
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1644511149
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1644511149
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1644511149
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1644511149
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1644511149
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1644511149
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1644511149
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1644511149
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1644511149
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1644511149
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1644511149
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1644511149
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1644511149
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1644511149
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1644511149
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1644511149
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1644511149
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1644511149
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1644511149
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1644511149
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1644511149
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1644511149
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1644511149
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1644511149
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1644511149
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1644511149
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1644511149
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1644511149
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1644511149
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1644511149
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1644511149
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1644511149
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1644511149
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1644511149
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1644511149
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1644511149
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1644511149
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1644511149
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1644511149
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1644511149
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1644511149
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1644511149
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1644511149
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1644511149
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1644511149
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1644511149
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1644511149
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1644511149
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1644511149
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1644511149
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1644511149
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1644511149
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1644511149
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1644511149
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1644511149
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1644511149
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1644511149
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1644511149
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1644511149
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1644511149
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1644511149
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1644511149
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1644511149
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1644511149
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1644511149
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1644511149
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1644511149
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1644511149
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1644511149
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1644511149
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1644511149
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1644511149
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1644511149
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1644511149
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1644511149
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1644511149
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1644511149
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1644511149
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1644511149
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1644511149
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1644511149
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1644511149
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1644511149
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1644511149
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1644511149
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1644511149
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1644511149
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1644511149
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1644511149
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1644511149
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1644511149
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1644511149
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1644511149
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1644511149
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1644511149
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1644511149
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1644511149
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1644511149
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1644511149
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1644511149
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1644511149
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1644511149
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1644511149
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1644511149
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1644511149
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1644511149
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1644511149
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1644511149
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1644511149
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1644511149
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1644511149
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1644511149
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1644511149
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1644511149
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1644511149
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1644511149
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1644511149
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1644511149
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1644511149
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1644511149
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1644511149
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1644511149
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1644511149
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1644511149
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1644511149
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1644511149
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1644511149
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1644511149
transform 1 0 6256 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1644511149
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1644511149
transform 1 0 11408 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1644511149
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1644511149
transform 1 0 16560 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1644511149
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1644511149
transform 1 0 21712 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1644511149
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1644511149
transform 1 0 26864 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1644511149
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1644511149
transform 1 0 32016 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1644511149
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1644511149
transform 1 0 37168 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1644511149
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1644511149
transform 1 0 42320 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1644511149
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1644511149
transform 1 0 47472 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _0934_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26036 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0935_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22356 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0936_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19596 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0937_
timestamp 1644511149
transform 1 0 18216 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0938_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0939_
timestamp 1644511149
transform 1 0 17940 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0940_
timestamp 1644511149
transform 1 0 18308 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0941_
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0942_
timestamp 1644511149
transform 1 0 33488 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0943_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20148 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0944_
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0945_
timestamp 1644511149
transform 1 0 33304 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0946_
timestamp 1644511149
transform 1 0 33396 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0947_
timestamp 1644511149
transform 1 0 32844 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0948_
timestamp 1644511149
transform 1 0 33764 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0949_
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0950_
timestamp 1644511149
transform 1 0 18676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0951_
timestamp 1644511149
transform 1 0 36432 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0952_
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0953_
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0954_
timestamp 1644511149
transform 1 0 36616 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0955_
timestamp 1644511149
transform 1 0 16100 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0956_
timestamp 1644511149
transform 1 0 18124 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0957_
timestamp 1644511149
transform 1 0 10028 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0958_
timestamp 1644511149
transform 1 0 18492 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0959_
timestamp 1644511149
transform 1 0 12420 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0960_
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0961_
timestamp 1644511149
transform 1 0 9476 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0962_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0963_
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0964_
timestamp 1644511149
transform 1 0 4784 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0965_
timestamp 1644511149
transform 1 0 10488 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0966_
timestamp 1644511149
transform 1 0 4140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0967_
timestamp 1644511149
transform 1 0 24932 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _0968_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31556 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _0969_
timestamp 1644511149
transform 1 0 16652 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0970_
timestamp 1644511149
transform 1 0 26036 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1644511149
transform 1 0 35696 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0972_
timestamp 1644511149
transform 1 0 2852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0973_
timestamp 1644511149
transform 1 0 46644 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0974_
timestamp 1644511149
transform 1 0 31188 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  _0975_
timestamp 1644511149
transform 1 0 31096 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _0976_
timestamp 1644511149
transform 1 0 30728 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0977_
timestamp 1644511149
transform 1 0 9016 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0978_
timestamp 1644511149
transform 1 0 2116 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0979_
timestamp 1644511149
transform 1 0 2116 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0980_
timestamp 1644511149
transform 1 0 30912 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _0981_
timestamp 1644511149
transform 1 0 32476 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _0982_
timestamp 1644511149
transform 1 0 17296 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0983_
timestamp 1644511149
transform 1 0 11684 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0984_
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0985_
timestamp 1644511149
transform 1 0 45632 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0986_
timestamp 1644511149
transform 1 0 45172 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0987_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30544 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0988_
timestamp 1644511149
transform 1 0 39836 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0989_
timestamp 1644511149
transform 1 0 9844 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0990_
timestamp 1644511149
transform 1 0 7636 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0991_
timestamp 1644511149
transform 1 0 46736 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0992_
timestamp 1644511149
transform 1 0 7084 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0993_
timestamp 1644511149
transform 1 0 31556 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0994_
timestamp 1644511149
transform 1 0 31188 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0995_
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0996_
timestamp 1644511149
transform 1 0 37444 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0997_
timestamp 1644511149
transform 1 0 36708 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0998_
timestamp 1644511149
transform 1 0 38088 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _0999_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1000_
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1001_
timestamp 1644511149
transform 1 0 45632 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1002_
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1003_
timestamp 1644511149
transform 1 0 8924 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1004_
timestamp 1644511149
transform 1 0 13800 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1005_
timestamp 1644511149
transform 1 0 20056 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _1006_
timestamp 1644511149
transform 1 0 20056 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1007_
timestamp 1644511149
transform 1 0 26956 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1008_
timestamp 1644511149
transform 1 0 47564 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1009_
timestamp 1644511149
transform 1 0 42596 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1010_
timestamp 1644511149
transform 1 0 47564 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1011_
timestamp 1644511149
transform 1 0 2944 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1012_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20148 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1013_
timestamp 1644511149
transform 1 0 47564 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1014_
timestamp 1644511149
transform 1 0 20884 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1015_
timestamp 1644511149
transform 1 0 47564 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1016_
timestamp 1644511149
transform 1 0 7452 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1017_
timestamp 1644511149
transform 1 0 9200 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1018_
timestamp 1644511149
transform 1 0 20148 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1019_
timestamp 1644511149
transform 1 0 2760 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1020_
timestamp 1644511149
transform 1 0 13248 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1021_
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1022_
timestamp 1644511149
transform 1 0 20884 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1023_
timestamp 1644511149
transform 1 0 15180 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1024_
timestamp 1644511149
transform 1 0 19780 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1025_
timestamp 1644511149
transform 1 0 20792 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1026_
timestamp 1644511149
transform 1 0 19596 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1027_
timestamp 1644511149
transform 1 0 19596 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1028_
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1029_
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1030_
timestamp 1644511149
transform 1 0 20056 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1031_
timestamp 1644511149
transform 1 0 2024 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1032_
timestamp 1644511149
transform 1 0 11776 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1033_
timestamp 1644511149
transform 1 0 2668 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1034_
timestamp 1644511149
transform 1 0 2116 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1035_
timestamp 1644511149
transform 1 0 40296 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1036_
timestamp 1644511149
transform 1 0 30084 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _1037_
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1038_
timestamp 1644511149
transform 1 0 37812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1039_
timestamp 1644511149
transform 1 0 4600 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1040_
timestamp 1644511149
transform 1 0 36248 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1041_
timestamp 1644511149
transform 1 0 36340 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1042_
timestamp 1644511149
transform 1 0 38364 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1043_
timestamp 1644511149
transform 1 0 30544 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1044_
timestamp 1644511149
transform 1 0 15548 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1045_
timestamp 1644511149
transform 1 0 33028 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1046_
timestamp 1644511149
transform 1 0 12052 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1047_
timestamp 1644511149
transform 1 0 21804 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1048_
timestamp 1644511149
transform 1 0 33120 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1049_
timestamp 1644511149
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1050_
timestamp 1644511149
transform 1 0 14260 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1051_
timestamp 1644511149
transform 1 0 2760 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1052_
timestamp 1644511149
transform 1 0 2024 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1053_
timestamp 1644511149
transform 1 0 2024 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1054_
timestamp 1644511149
transform 1 0 46736 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _1055_
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1056_
timestamp 1644511149
transform 1 0 43884 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1057_
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1058_
timestamp 1644511149
transform 1 0 28428 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1059_
timestamp 1644511149
transform 1 0 4784 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1060_
timestamp 1644511149
transform 1 0 46644 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _1061_
timestamp 1644511149
transform 1 0 31740 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _1062_
timestamp 1644511149
transform 1 0 46092 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1063_
timestamp 1644511149
transform 1 0 47196 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1064_
timestamp 1644511149
transform 1 0 32108 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1065_
timestamp 1644511149
transform 1 0 41308 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1066_
timestamp 1644511149
transform 1 0 5336 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1067_
timestamp 1644511149
transform 1 0 23368 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  _1068_
timestamp 1644511149
transform 1 0 24748 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _1069_
timestamp 1644511149
transform 1 0 38640 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1070_
timestamp 1644511149
transform 1 0 19964 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1071_
timestamp 1644511149
transform 1 0 2208 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1072_
timestamp 1644511149
transform 1 0 30176 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1073_
timestamp 1644511149
transform 1 0 2944 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _1074_
timestamp 1644511149
transform 1 0 23552 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1075_
timestamp 1644511149
transform 1 0 23552 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1076_
timestamp 1644511149
transform 1 0 11960 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1077_
timestamp 1644511149
transform 1 0 2852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1078_
timestamp 1644511149
transform 1 0 23276 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1079_
timestamp 1644511149
transform 1 0 46736 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1080_
timestamp 1644511149
transform 1 0 22816 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1081_
timestamp 1644511149
transform 1 0 43516 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1082_
timestamp 1644511149
transform 1 0 47564 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1083_
timestamp 1644511149
transform 1 0 2852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1084_
timestamp 1644511149
transform 1 0 30084 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1085_
timestamp 1644511149
transform 1 0 46828 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1086_
timestamp 1644511149
transform 1 0 24380 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1087_
timestamp 1644511149
transform 1 0 44988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1088_
timestamp 1644511149
transform 1 0 47564 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1089_
timestamp 1644511149
transform 1 0 46828 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1090_
timestamp 1644511149
transform 1 0 8924 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1091_
timestamp 1644511149
transform 1 0 46828 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _1092_
timestamp 1644511149
transform 1 0 23552 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1093_
timestamp 1644511149
transform 1 0 47564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1094_
timestamp 1644511149
transform 1 0 2116 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1095_
timestamp 1644511149
transform 1 0 2484 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1096_
timestamp 1644511149
transform 1 0 36156 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1097_
timestamp 1644511149
transform 1 0 46828 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1098_
timestamp 1644511149
transform 1 0 24840 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  _1099_
timestamp 1644511149
transform 1 0 27232 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1100_
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1101_
timestamp 1644511149
transform 1 0 44252 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1102_
timestamp 1644511149
transform 1 0 2116 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1103_
timestamp 1644511149
transform 1 0 44528 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1104_
timestamp 1644511149
transform 1 0 24104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _1105_
timestamp 1644511149
transform 1 0 25024 0 1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _1106_
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1107_
timestamp 1644511149
transform 1 0 47564 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1108_
timestamp 1644511149
transform 1 0 1380 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1109_
timestamp 1644511149
transform 1 0 12328 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1110_
timestamp 1644511149
transform 1 0 46184 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1111_
timestamp 1644511149
transform 1 0 25024 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1112_
timestamp 1644511149
transform 1 0 2024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1113_
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1114_
timestamp 1644511149
transform 1 0 21068 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1115_
timestamp 1644511149
transform 1 0 2024 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1116_
timestamp 1644511149
transform 1 0 2024 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _1117_
timestamp 1644511149
transform 1 0 25024 0 -1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1118_
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1119_
timestamp 1644511149
transform 1 0 2852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1120_
timestamp 1644511149
transform 1 0 6072 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1121_
timestamp 1644511149
transform 1 0 36064 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1122_
timestamp 1644511149
transform 1 0 46644 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _1123_
timestamp 1644511149
transform 1 0 24656 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _1124_
timestamp 1644511149
transform 1 0 2116 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1125_
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1126_
timestamp 1644511149
transform 1 0 2116 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1127_
timestamp 1644511149
transform 1 0 5428 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1128_
timestamp 1644511149
transform 1 0 28796 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1129_
timestamp 1644511149
transform 1 0 14168 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1130_
timestamp 1644511149
transform 1 0 6808 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1131_
timestamp 1644511149
transform 1 0 15364 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1132_
timestamp 1644511149
transform 1 0 15732 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1133_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1134_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1135_
timestamp 1644511149
transform 1 0 12788 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1136_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16744 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1137_
timestamp 1644511149
transform 1 0 17480 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1138_
timestamp 1644511149
transform 1 0 17204 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1139_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16376 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _1140_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1141_
timestamp 1644511149
transform 1 0 21528 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1142_
timestamp 1644511149
transform 1 0 20700 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1143_
timestamp 1644511149
transform 1 0 15824 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1144_
timestamp 1644511149
transform 1 0 27140 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1145_
timestamp 1644511149
transform 1 0 28612 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1146_
timestamp 1644511149
transform 1 0 30820 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1147_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29072 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1148_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24196 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1149_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24840 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1150_
timestamp 1644511149
transform 1 0 30452 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1151_
timestamp 1644511149
transform 1 0 24472 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1152_
timestamp 1644511149
transform 1 0 25116 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1153_
timestamp 1644511149
transform 1 0 28612 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1154_
timestamp 1644511149
transform 1 0 28520 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1155_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27140 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1156_
timestamp 1644511149
transform 1 0 25576 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_1  _1157_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1158_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15364 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1159_
timestamp 1644511149
transform 1 0 15640 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1160_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1161_
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1162_
timestamp 1644511149
transform 1 0 15548 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1163_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26036 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1164_
timestamp 1644511149
transform 1 0 26680 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1165_
timestamp 1644511149
transform 1 0 27416 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1166_
timestamp 1644511149
transform 1 0 26680 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1167_
timestamp 1644511149
transform 1 0 17112 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1168_
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1169_
timestamp 1644511149
transform 1 0 20332 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1170_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19688 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1171_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21068 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1172_
timestamp 1644511149
transform 1 0 24656 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1173_
timestamp 1644511149
transform 1 0 24288 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1174_
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1175_
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1176_
timestamp 1644511149
transform 1 0 10120 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1177_
timestamp 1644511149
transform 1 0 10856 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1178_
timestamp 1644511149
transform 1 0 12420 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1179_
timestamp 1644511149
transform 1 0 9200 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1180_
timestamp 1644511149
transform 1 0 15272 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1181_
timestamp 1644511149
transform 1 0 16100 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1182_
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1183_
timestamp 1644511149
transform 1 0 13432 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1184_
timestamp 1644511149
transform 1 0 14720 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1185_
timestamp 1644511149
transform 1 0 7452 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1186_
timestamp 1644511149
transform 1 0 28336 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_2  _1187_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 47288 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1188_
timestamp 1644511149
transform 1 0 28612 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1189_
timestamp 1644511149
transform 1 0 28244 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1190_
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1191_
timestamp 1644511149
transform 1 0 30820 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1192_
timestamp 1644511149
transform 1 0 29440 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1193_
timestamp 1644511149
transform 1 0 31096 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1194_
timestamp 1644511149
transform 1 0 31188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1195_
timestamp 1644511149
transform 1 0 31004 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1196_
timestamp 1644511149
transform 1 0 26220 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1197_
timestamp 1644511149
transform 1 0 27416 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1198_
timestamp 1644511149
transform 1 0 27324 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1199_
timestamp 1644511149
transform 1 0 19596 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1200_
timestamp 1644511149
transform 1 0 26864 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1201_
timestamp 1644511149
transform 1 0 25484 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_4  _1202_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26128 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1203_
timestamp 1644511149
transform 1 0 18492 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1204_
timestamp 1644511149
transform 1 0 18308 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1205_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17848 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1206_
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1207_
timestamp 1644511149
transform 1 0 18216 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1208_
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1209_
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1210_
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1211_
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1212_
timestamp 1644511149
transform 1 0 18308 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1213_
timestamp 1644511149
transform 1 0 17204 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1214_
timestamp 1644511149
transform 1 0 18032 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1215_
timestamp 1644511149
transform 1 0 31648 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1216_
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1217_
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1218_
timestamp 1644511149
transform 1 0 30912 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1219_
timestamp 1644511149
transform 1 0 32660 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1220_
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1221_
timestamp 1644511149
transform 1 0 33028 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1222_
timestamp 1644511149
transform 1 0 32200 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1223_
timestamp 1644511149
transform 1 0 33580 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1224_
timestamp 1644511149
transform 1 0 31648 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1225_
timestamp 1644511149
transform 1 0 32476 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1226_
timestamp 1644511149
transform 1 0 31188 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1227_
timestamp 1644511149
transform 1 0 32384 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1228_
timestamp 1644511149
transform 1 0 31832 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1229_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1230_
timestamp 1644511149
transform 1 0 33212 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1231_
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1232_
timestamp 1644511149
transform 1 0 33028 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1233_
timestamp 1644511149
transform 1 0 31924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1234_
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1235_
timestamp 1644511149
transform 1 0 33120 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1236_
timestamp 1644511149
transform 1 0 36064 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1237_
timestamp 1644511149
transform 1 0 17664 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1238_
timestamp 1644511149
transform 1 0 33856 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1239_
timestamp 1644511149
transform 1 0 36064 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1240_
timestamp 1644511149
transform 1 0 34960 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1241_
timestamp 1644511149
transform 1 0 14168 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1242_
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1243_
timestamp 1644511149
transform 1 0 16836 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1244_
timestamp 1644511149
transform 1 0 16836 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1245_
timestamp 1644511149
transform 1 0 13524 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1246_
timestamp 1644511149
transform 1 0 14720 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1247_
timestamp 1644511149
transform 1 0 14536 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1248_
timestamp 1644511149
transform 1 0 15088 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1249_
timestamp 1644511149
transform 1 0 13156 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1250_
timestamp 1644511149
transform 1 0 15640 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1251_
timestamp 1644511149
transform 1 0 17296 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1252_
timestamp 1644511149
transform 1 0 18124 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1253_
timestamp 1644511149
transform 1 0 16192 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1254_
timestamp 1644511149
transform 1 0 14168 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1255_
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1256_
timestamp 1644511149
transform 1 0 12604 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1257_
timestamp 1644511149
transform 1 0 12328 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1258_
timestamp 1644511149
transform 1 0 9844 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1259_
timestamp 1644511149
transform 1 0 9200 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1260_
timestamp 1644511149
transform 1 0 9384 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1261_
timestamp 1644511149
transform 1 0 9384 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1262_
timestamp 1644511149
transform 1 0 10488 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1263_
timestamp 1644511149
transform 1 0 9016 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1264_
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1265_
timestamp 1644511149
transform 1 0 26680 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1266_
timestamp 1644511149
transform 1 0 22264 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1267_
timestamp 1644511149
transform 1 0 17112 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1268_
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1269_
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1270_
timestamp 1644511149
transform 1 0 11316 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1271_
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1272_
timestamp 1644511149
transform 1 0 20976 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1273_
timestamp 1644511149
transform 1 0 18768 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1274_
timestamp 1644511149
transform 1 0 22540 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1275_
timestamp 1644511149
transform 1 0 21528 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1276_
timestamp 1644511149
transform 1 0 16836 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and4_2  _1277_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25760 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1278_
timestamp 1644511149
transform 1 0 20608 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1279_
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1280_
timestamp 1644511149
transform 1 0 12880 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1281_
timestamp 1644511149
transform 1 0 14352 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1282_
timestamp 1644511149
transform 1 0 15456 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1283_
timestamp 1644511149
transform 1 0 17296 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1284_
timestamp 1644511149
transform 1 0 16744 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1285_
timestamp 1644511149
transform 1 0 17480 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1286_
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1287_
timestamp 1644511149
transform 1 0 12880 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1288_
timestamp 1644511149
transform 1 0 19780 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1289_
timestamp 1644511149
transform 1 0 20976 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1290_
timestamp 1644511149
transform 1 0 19504 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1291_
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1292_
timestamp 1644511149
transform 1 0 18032 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1293_
timestamp 1644511149
transform 1 0 17756 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1294_
timestamp 1644511149
transform 1 0 17848 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1295_
timestamp 1644511149
transform 1 0 16468 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1296_
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1297_
timestamp 1644511149
transform 1 0 20424 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1298_
timestamp 1644511149
transform 1 0 20700 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1299_
timestamp 1644511149
transform 1 0 20608 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1300_
timestamp 1644511149
transform 1 0 20516 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1301_
timestamp 1644511149
transform 1 0 20608 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1302_
timestamp 1644511149
transform 1 0 20240 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1303_
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1304_
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1305_
timestamp 1644511149
transform 1 0 20424 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1306_
timestamp 1644511149
transform 1 0 21896 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1307_
timestamp 1644511149
transform 1 0 22080 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1308_
timestamp 1644511149
transform 1 0 20332 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1309_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20424 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1310_
timestamp 1644511149
transform 1 0 20056 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1311_
timestamp 1644511149
transform 1 0 20608 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1312_
timestamp 1644511149
transform 1 0 22632 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1313_
timestamp 1644511149
transform 1 0 22632 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1314_
timestamp 1644511149
transform 1 0 22724 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1315_
timestamp 1644511149
transform 1 0 21804 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1316_
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1317_
timestamp 1644511149
transform 1 0 20332 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1318_
timestamp 1644511149
transform 1 0 22172 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1319_
timestamp 1644511149
transform 1 0 34960 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1320_
timestamp 1644511149
transform 1 0 35144 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1321_
timestamp 1644511149
transform 1 0 36156 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1322_
timestamp 1644511149
transform 1 0 36248 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1323_
timestamp 1644511149
transform 1 0 34960 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1324_
timestamp 1644511149
transform 1 0 35052 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1325_
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1326_
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1327_
timestamp 1644511149
transform 1 0 20516 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1328_
timestamp 1644511149
transform 1 0 21620 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1329_
timestamp 1644511149
transform 1 0 19688 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1330_
timestamp 1644511149
transform 1 0 20700 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1331_
timestamp 1644511149
transform 1 0 19596 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1332_
timestamp 1644511149
transform 1 0 20792 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1333_
timestamp 1644511149
transform 1 0 19688 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1334_
timestamp 1644511149
transform 1 0 19504 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1335_
timestamp 1644511149
transform 1 0 18952 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1336_
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1337_
timestamp 1644511149
transform 1 0 27232 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1338_
timestamp 1644511149
transform 1 0 27232 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1339_
timestamp 1644511149
transform 1 0 22448 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1340_
timestamp 1644511149
transform 1 0 47564 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1341_
timestamp 1644511149
transform 1 0 28428 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1342_
timestamp 1644511149
transform 1 0 29348 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1343_
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1344_
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1345_
timestamp 1644511149
transform 1 0 29624 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1346_
timestamp 1644511149
transform 1 0 30820 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1347_
timestamp 1644511149
transform 1 0 29532 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1348_
timestamp 1644511149
transform 1 0 28520 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1349_
timestamp 1644511149
transform 1 0 30084 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1350_
timestamp 1644511149
transform 1 0 31004 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_2  _1351_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25116 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1352_
timestamp 1644511149
transform 1 0 27692 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1353_
timestamp 1644511149
transform 1 0 28060 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1354_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27416 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1355_
timestamp 1644511149
transform 1 0 28704 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1356_
timestamp 1644511149
transform 1 0 25852 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1357_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23276 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1358_
timestamp 1644511149
transform 1 0 23460 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1359_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24472 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1360_
timestamp 1644511149
transform 1 0 23092 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1361_
timestamp 1644511149
transform 1 0 23460 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1362_
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1363_
timestamp 1644511149
transform 1 0 27692 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1364_
timestamp 1644511149
transform 1 0 23368 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1365_
timestamp 1644511149
transform 1 0 24104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1366_
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _1367_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25484 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1368_
timestamp 1644511149
transform 1 0 23092 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1369_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23000 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1370_
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1371_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23184 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1372_
timestamp 1644511149
transform 1 0 24656 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1373_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1374_
timestamp 1644511149
transform 1 0 25300 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1375_
timestamp 1644511149
transform 1 0 26680 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1376_
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1377_
timestamp 1644511149
transform 1 0 27692 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1378_
timestamp 1644511149
transform 1 0 25668 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1379_
timestamp 1644511149
transform 1 0 25576 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1380_
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1381_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25852 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1382_
timestamp 1644511149
transform 1 0 26036 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1383_
timestamp 1644511149
transform 1 0 26864 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1384_
timestamp 1644511149
transform 1 0 28152 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1385_
timestamp 1644511149
transform 1 0 27232 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1386_
timestamp 1644511149
transform 1 0 28152 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1387_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27968 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1388_
timestamp 1644511149
transform 1 0 29348 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1389_
timestamp 1644511149
transform 1 0 27876 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1390_
timestamp 1644511149
transform 1 0 28704 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1391_
timestamp 1644511149
transform 1 0 28520 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1392_
timestamp 1644511149
transform 1 0 27784 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1393_
timestamp 1644511149
transform 1 0 26956 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1394_
timestamp 1644511149
transform 1 0 29900 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1395_
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1396_
timestamp 1644511149
transform 1 0 27600 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1397_
timestamp 1644511149
transform 1 0 27416 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1398_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28244 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1399_
timestamp 1644511149
transform 1 0 28244 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1400_
timestamp 1644511149
transform 1 0 29072 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1401_
timestamp 1644511149
transform 1 0 29808 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1402_
timestamp 1644511149
transform 1 0 28888 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1403_
timestamp 1644511149
transform 1 0 27600 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1404_
timestamp 1644511149
transform 1 0 27508 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1405_
timestamp 1644511149
transform 1 0 28428 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1406_
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1407_
timestamp 1644511149
transform 1 0 28888 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1408_
timestamp 1644511149
transform 1 0 28612 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1409_
timestamp 1644511149
transform 1 0 26956 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1410_
timestamp 1644511149
transform 1 0 30728 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1411_
timestamp 1644511149
transform 1 0 29256 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1412_
timestamp 1644511149
transform 1 0 28244 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1413_
timestamp 1644511149
transform 1 0 27232 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1414_
timestamp 1644511149
transform 1 0 27692 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1415_
timestamp 1644511149
transform 1 0 28980 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1416_
timestamp 1644511149
transform 1 0 27508 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1417_
timestamp 1644511149
transform 1 0 26128 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1418_
timestamp 1644511149
transform 1 0 27508 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1419_
timestamp 1644511149
transform 1 0 26864 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1420_
timestamp 1644511149
transform 1 0 26680 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1421_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25852 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1422_
timestamp 1644511149
transform 1 0 25484 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1423_
timestamp 1644511149
transform 1 0 27692 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1424_
timestamp 1644511149
transform 1 0 27232 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1425_
timestamp 1644511149
transform 1 0 25484 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1426_
timestamp 1644511149
transform 1 0 26680 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1427_
timestamp 1644511149
transform 1 0 28888 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1428_
timestamp 1644511149
transform 1 0 25668 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1429_
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1430_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26220 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1431_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27048 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1432_
timestamp 1644511149
transform 1 0 28152 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1433_
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1434_
timestamp 1644511149
transform 1 0 24288 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o31ai_1  _1435_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25484 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1436_
timestamp 1644511149
transform 1 0 24748 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1437_
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1438_
timestamp 1644511149
transform 1 0 23184 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1439_
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1440_
timestamp 1644511149
transform 1 0 23276 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1441_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23552 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1442_
timestamp 1644511149
transform 1 0 22356 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1443_
timestamp 1644511149
transform 1 0 27416 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1444_
timestamp 1644511149
transform 1 0 27324 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1445_
timestamp 1644511149
transform 1 0 28520 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1446_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27784 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1447_
timestamp 1644511149
transform 1 0 27416 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1448_
timestamp 1644511149
transform 1 0 25668 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1449_
timestamp 1644511149
transform 1 0 25392 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1450_
timestamp 1644511149
transform 1 0 24932 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1451_
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1452_
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1453_
timestamp 1644511149
transform 1 0 24012 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1454_
timestamp 1644511149
transform 1 0 24288 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _1455_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14168 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1456_
timestamp 1644511149
transform 1 0 10672 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1457_
timestamp 1644511149
transform 1 0 10120 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1458_
timestamp 1644511149
transform 1 0 9292 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1459_
timestamp 1644511149
transform 1 0 8372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1460_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9936 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1461_
timestamp 1644511149
transform 1 0 9844 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1462_
timestamp 1644511149
transform 1 0 14260 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1463_
timestamp 1644511149
transform 1 0 14168 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1464_
timestamp 1644511149
transform 1 0 13248 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1465_
timestamp 1644511149
transform 1 0 13616 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1466_
timestamp 1644511149
transform 1 0 15180 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1467_
timestamp 1644511149
transform 1 0 15364 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1468_
timestamp 1644511149
transform 1 0 14720 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1469_
timestamp 1644511149
transform 1 0 15272 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1470_
timestamp 1644511149
transform 1 0 14720 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1471_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1472_
timestamp 1644511149
transform 1 0 11684 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _1473_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14444 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1474_
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1475_
timestamp 1644511149
transform 1 0 15548 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _1476_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1477_
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1478_
timestamp 1644511149
transform 1 0 9936 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22oi_1  _1479_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1480_
timestamp 1644511149
transform 1 0 10212 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1481_
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1482_
timestamp 1644511149
transform 1 0 12696 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1483_
timestamp 1644511149
transform 1 0 14904 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1484_
timestamp 1644511149
transform 1 0 14168 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1485_
timestamp 1644511149
transform 1 0 14260 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1486_
timestamp 1644511149
transform 1 0 12696 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1487_
timestamp 1644511149
transform 1 0 11868 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1488_
timestamp 1644511149
transform 1 0 12972 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1489_
timestamp 1644511149
transform 1 0 13800 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1490_
timestamp 1644511149
transform 1 0 14628 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1491_
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1492_
timestamp 1644511149
transform 1 0 13708 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _1493_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12696 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1494_
timestamp 1644511149
transform 1 0 11960 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1495_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11592 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1496_
timestamp 1644511149
transform 1 0 11316 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1497_
timestamp 1644511149
transform 1 0 11500 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1498_
timestamp 1644511149
transform 1 0 12144 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1499_
timestamp 1644511149
transform 1 0 11684 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1500_
timestamp 1644511149
transform 1 0 12420 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1501_
timestamp 1644511149
transform 1 0 11224 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1502_
timestamp 1644511149
transform 1 0 10672 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1503_
timestamp 1644511149
transform 1 0 9936 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1504_
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1505_
timestamp 1644511149
transform 1 0 9476 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1506_
timestamp 1644511149
transform 1 0 10304 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1507_
timestamp 1644511149
transform 1 0 9108 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1508_
timestamp 1644511149
transform 1 0 9108 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1509_
timestamp 1644511149
transform 1 0 10488 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1510_
timestamp 1644511149
transform 1 0 8372 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1511_
timestamp 1644511149
transform 1 0 8280 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1512_
timestamp 1644511149
transform 1 0 7728 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1513_
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1514_
timestamp 1644511149
transform 1 0 9384 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1515_
timestamp 1644511149
transform 1 0 7820 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1516_
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1517_
timestamp 1644511149
transform 1 0 17572 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1518_
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1519_
timestamp 1644511149
transform 1 0 25484 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1520_
timestamp 1644511149
transform 1 0 18308 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1521_
timestamp 1644511149
transform 1 0 26128 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1522_
timestamp 1644511149
transform 1 0 26680 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1523_
timestamp 1644511149
transform 1 0 26036 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1524_
timestamp 1644511149
transform 1 0 24656 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1525_
timestamp 1644511149
transform 1 0 24748 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1526_
timestamp 1644511149
transform 1 0 27508 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1527_
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1528_
timestamp 1644511149
transform 1 0 28428 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1529_
timestamp 1644511149
transform 1 0 27324 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1530_
timestamp 1644511149
transform 1 0 32660 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1531_
timestamp 1644511149
transform 1 0 28244 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1532_
timestamp 1644511149
transform 1 0 27968 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1533_
timestamp 1644511149
transform 1 0 27232 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1534_
timestamp 1644511149
transform 1 0 29808 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1535_
timestamp 1644511149
transform 1 0 29808 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1536_
timestamp 1644511149
transform 1 0 29440 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1537_
timestamp 1644511149
transform 1 0 30728 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1538_
timestamp 1644511149
transform 1 0 31464 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1539_
timestamp 1644511149
transform 1 0 31188 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1540_
timestamp 1644511149
transform 1 0 30912 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1541_
timestamp 1644511149
transform 1 0 24380 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1542_
timestamp 1644511149
transform 1 0 26128 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1543_
timestamp 1644511149
transform 1 0 33396 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1544_
timestamp 1644511149
transform 1 0 32568 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1545_
timestamp 1644511149
transform 1 0 32476 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1546_
timestamp 1644511149
transform 1 0 27232 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1547_
timestamp 1644511149
transform 1 0 33396 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1548_
timestamp 1644511149
transform 1 0 32016 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1549_
timestamp 1644511149
transform 1 0 32476 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1550_
timestamp 1644511149
transform 1 0 28612 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1551_
timestamp 1644511149
transform 1 0 32844 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1552_
timestamp 1644511149
transform 1 0 32200 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1553_
timestamp 1644511149
transform 1 0 32292 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1554_
timestamp 1644511149
transform 1 0 27600 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1555_
timestamp 1644511149
transform 1 0 26772 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1556_
timestamp 1644511149
transform 1 0 28612 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1557_
timestamp 1644511149
transform 1 0 25760 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1558_
timestamp 1644511149
transform 1 0 30268 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1559_
timestamp 1644511149
transform 1 0 30636 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1560_
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1561_
timestamp 1644511149
transform 1 0 26128 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1562_
timestamp 1644511149
transform 1 0 28520 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1563_
timestamp 1644511149
transform 1 0 28152 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1564_
timestamp 1644511149
transform 1 0 27048 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1565_
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1566_
timestamp 1644511149
transform 1 0 27416 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1567_
timestamp 1644511149
transform 1 0 27968 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1568_
timestamp 1644511149
transform 1 0 26864 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1569_
timestamp 1644511149
transform 1 0 30452 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1570_
timestamp 1644511149
transform 1 0 29900 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1571_
timestamp 1644511149
transform 1 0 29624 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1572_
timestamp 1644511149
transform 1 0 29348 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1573_
timestamp 1644511149
transform 1 0 32200 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1574_
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1575_
timestamp 1644511149
transform 1 0 29164 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1576_
timestamp 1644511149
transform 1 0 31096 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1577_
timestamp 1644511149
transform 1 0 33396 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1578_
timestamp 1644511149
transform 1 0 33028 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1579_
timestamp 1644511149
transform 1 0 31924 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1580_
timestamp 1644511149
transform 1 0 26128 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1581_
timestamp 1644511149
transform 1 0 32752 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1582_
timestamp 1644511149
transform 1 0 31556 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1583_
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1584_
timestamp 1644511149
transform 1 0 26588 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1585_
timestamp 1644511149
transform 1 0 29808 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1586_
timestamp 1644511149
transform 1 0 28980 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1587_
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1588_
timestamp 1644511149
transform 1 0 28244 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1589_
timestamp 1644511149
transform 1 0 30360 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1590_
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1591_
timestamp 1644511149
transform 1 0 28888 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1592_
timestamp 1644511149
transform 1 0 27048 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1593_
timestamp 1644511149
transform 1 0 25852 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1594_
timestamp 1644511149
transform 1 0 31004 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1595_
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1596_
timestamp 1644511149
transform 1 0 26772 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1597_
timestamp 1644511149
transform 1 0 27968 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1598_
timestamp 1644511149
transform 1 0 25668 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1599_
timestamp 1644511149
transform 1 0 28520 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1600_
timestamp 1644511149
transform 1 0 29164 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1601_
timestamp 1644511149
transform 1 0 28796 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1602_
timestamp 1644511149
transform 1 0 28336 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1603_
timestamp 1644511149
transform 1 0 23184 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1604_
timestamp 1644511149
transform 1 0 29808 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1605_
timestamp 1644511149
transform 1 0 29716 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1606_
timestamp 1644511149
transform 1 0 30360 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1607_
timestamp 1644511149
transform 1 0 31648 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1608_
timestamp 1644511149
transform 1 0 32108 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1609_
timestamp 1644511149
transform 1 0 32108 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1610_
timestamp 1644511149
transform 1 0 32844 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1611_
timestamp 1644511149
transform 1 0 31188 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1612_
timestamp 1644511149
transform 1 0 23092 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1613_
timestamp 1644511149
transform 1 0 24012 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1614_
timestamp 1644511149
transform 1 0 33212 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  _1615_
timestamp 1644511149
transform 1 0 30912 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1616_
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1617_
timestamp 1644511149
transform 1 0 32844 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1618_
timestamp 1644511149
transform 1 0 33120 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1619_
timestamp 1644511149
transform 1 0 25484 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1620_
timestamp 1644511149
transform 1 0 32200 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1621_
timestamp 1644511149
transform 1 0 32384 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1622_
timestamp 1644511149
transform 1 0 28704 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1623_
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1624_
timestamp 1644511149
transform 1 0 25392 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1625_
timestamp 1644511149
transform 1 0 27692 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1626_
timestamp 1644511149
transform 1 0 25668 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1627_
timestamp 1644511149
transform 1 0 28428 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1628_
timestamp 1644511149
transform 1 0 23184 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1629_
timestamp 1644511149
transform 1 0 27324 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1630_
timestamp 1644511149
transform 1 0 30268 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1631_
timestamp 1644511149
transform 1 0 27876 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1632_
timestamp 1644511149
transform 1 0 21436 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1633_
timestamp 1644511149
transform 1 0 22540 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1634_
timestamp 1644511149
transform 1 0 26956 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1635_
timestamp 1644511149
transform 1 0 26496 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1636_
timestamp 1644511149
transform 1 0 28796 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1637_
timestamp 1644511149
transform 1 0 27692 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1638_
timestamp 1644511149
transform 1 0 23736 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1639_
timestamp 1644511149
transform 1 0 22632 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1640_
timestamp 1644511149
transform 1 0 23000 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1641_
timestamp 1644511149
transform 1 0 23000 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1642_
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1643_
timestamp 1644511149
transform 1 0 19320 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1644_
timestamp 1644511149
transform 1 0 22908 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1645_
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1646_
timestamp 1644511149
transform 1 0 21344 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1647_
timestamp 1644511149
transform 1 0 23644 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1648_
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1649_
timestamp 1644511149
transform 1 0 24564 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1650_
timestamp 1644511149
transform 1 0 24472 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1651_
timestamp 1644511149
transform 1 0 20700 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1652_
timestamp 1644511149
transform 1 0 20332 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1653_
timestamp 1644511149
transform 1 0 20332 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1654_
timestamp 1644511149
transform 1 0 23000 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1655_
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1656_
timestamp 1644511149
transform 1 0 18676 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1657_
timestamp 1644511149
transform 1 0 21344 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1658_
timestamp 1644511149
transform 1 0 20608 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1659_
timestamp 1644511149
transform 1 0 22172 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1660_
timestamp 1644511149
transform 1 0 18308 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1661_
timestamp 1644511149
transform 1 0 18768 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1662_
timestamp 1644511149
transform 1 0 23000 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1663_
timestamp 1644511149
transform 1 0 23184 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1664_
timestamp 1644511149
transform 1 0 22172 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1665_
timestamp 1644511149
transform 1 0 22080 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1666_
timestamp 1644511149
transform 1 0 19872 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1667_
timestamp 1644511149
transform 1 0 23000 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1668_
timestamp 1644511149
transform 1 0 18032 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1669_
timestamp 1644511149
transform 1 0 19044 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1670_
timestamp 1644511149
transform 1 0 24012 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1671_
timestamp 1644511149
transform 1 0 23828 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1672_
timestamp 1644511149
transform 1 0 21620 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1673_
timestamp 1644511149
transform 1 0 23460 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1674_
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1675_
timestamp 1644511149
transform 1 0 20884 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1676_
timestamp 1644511149
transform 1 0 21436 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1677_
timestamp 1644511149
transform 1 0 19780 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1678_
timestamp 1644511149
transform 1 0 18676 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1679_
timestamp 1644511149
transform 1 0 20424 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1680_
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1681_
timestamp 1644511149
transform 1 0 21252 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1682_
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1683_
timestamp 1644511149
transform 1 0 23644 0 -1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1684_
timestamp 1644511149
transform 1 0 22632 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1685_
timestamp 1644511149
transform 1 0 22448 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1686_
timestamp 1644511149
transform 1 0 20884 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1687_
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1688_
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1689_
timestamp 1644511149
transform 1 0 20424 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1690_
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1691_
timestamp 1644511149
transform 1 0 19688 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1692_
timestamp 1644511149
transform 1 0 18584 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1693_
timestamp 1644511149
transform 1 0 20332 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1694_
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1695_
timestamp 1644511149
transform 1 0 19872 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1696_
timestamp 1644511149
transform 1 0 22908 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1697_
timestamp 1644511149
transform 1 0 33396 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1698_
timestamp 1644511149
transform 1 0 34224 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1699_
timestamp 1644511149
transform 1 0 22540 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1700_
timestamp 1644511149
transform 1 0 37260 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1701_
timestamp 1644511149
transform 1 0 35972 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1702_
timestamp 1644511149
transform 1 0 35604 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1703_
timestamp 1644511149
transform 1 0 35788 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1704_
timestamp 1644511149
transform 1 0 35420 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1705_
timestamp 1644511149
transform 1 0 36064 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1706_
timestamp 1644511149
transform 1 0 24472 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1707_
timestamp 1644511149
transform 1 0 22816 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1708_
timestamp 1644511149
transform 1 0 23184 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1709_
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1710_
timestamp 1644511149
transform 1 0 22080 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1711_
timestamp 1644511149
transform 1 0 21712 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1712_
timestamp 1644511149
transform 1 0 21896 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1713_
timestamp 1644511149
transform 1 0 21804 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1714_
timestamp 1644511149
transform 1 0 23460 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1715_
timestamp 1644511149
transform 1 0 24380 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1716_
timestamp 1644511149
transform 1 0 23460 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1717_
timestamp 1644511149
transform 1 0 24380 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1718_
timestamp 1644511149
transform 1 0 21804 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1719_
timestamp 1644511149
transform 1 0 20608 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1720_
timestamp 1644511149
transform 1 0 20516 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1721_
timestamp 1644511149
transform 1 0 32016 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1722_
timestamp 1644511149
transform 1 0 20976 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1723_
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1724_
timestamp 1644511149
transform 1 0 25300 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1725_
timestamp 1644511149
transform 1 0 29900 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1726_
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1727_
timestamp 1644511149
transform 1 0 28336 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1728_
timestamp 1644511149
transform 1 0 33948 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1729_
timestamp 1644511149
transform 1 0 32568 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1730_
timestamp 1644511149
transform 1 0 29624 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1731_
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1732_
timestamp 1644511149
transform 1 0 33304 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1733_
timestamp 1644511149
transform 1 0 34868 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1734_
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1735_
timestamp 1644511149
transform 1 0 35512 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1736_
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1737_
timestamp 1644511149
transform 1 0 35512 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1738_
timestamp 1644511149
transform 1 0 34408 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1739_
timestamp 1644511149
transform 1 0 35696 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1740_
timestamp 1644511149
transform 1 0 33488 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1741_
timestamp 1644511149
transform 1 0 16284 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1742_
timestamp 1644511149
transform 1 0 15640 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1743_
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1744_
timestamp 1644511149
transform 1 0 15456 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1745_
timestamp 1644511149
transform 1 0 17204 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1746_
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1747_
timestamp 1644511149
transform 1 0 17940 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1748_
timestamp 1644511149
transform 1 0 17388 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1749_
timestamp 1644511149
transform 1 0 17940 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1750_
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1751_
timestamp 1644511149
transform 1 0 18860 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1752_
timestamp 1644511149
transform 1 0 17848 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1753_
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1754_
timestamp 1644511149
transform 1 0 11776 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1755_
timestamp 1644511149
transform 1 0 10396 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1756_
timestamp 1644511149
transform 1 0 10212 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1757_
timestamp 1644511149
transform 1 0 9568 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1758_
timestamp 1644511149
transform 1 0 10396 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1759_
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _1760_
timestamp 1644511149
transform 1 0 15272 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1761_
timestamp 1644511149
transform 1 0 14628 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1762_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14720 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1763_
timestamp 1644511149
transform 1 0 19504 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1764_
timestamp 1644511149
transform 1 0 23368 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1765_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1766_
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1767_
timestamp 1644511149
transform 1 0 19320 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1768_
timestamp 1644511149
transform 1 0 18492 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1769_
timestamp 1644511149
transform 1 0 17020 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1770_
timestamp 1644511149
transform 1 0 17112 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1771_
timestamp 1644511149
transform 1 0 31188 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1772_
timestamp 1644511149
transform 1 0 32384 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1773_
timestamp 1644511149
transform 1 0 32384 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1774_
timestamp 1644511149
transform 1 0 32568 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1775_
timestamp 1644511149
transform 1 0 32384 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1776_
timestamp 1644511149
transform 1 0 31924 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1777_
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1778_
timestamp 1644511149
transform 1 0 34224 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1779_
timestamp 1644511149
transform 1 0 34776 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1780_
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1781_
timestamp 1644511149
transform 1 0 17020 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1782_
timestamp 1644511149
transform 1 0 14536 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1783_
timestamp 1644511149
transform 1 0 12328 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1784_
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1785_
timestamp 1644511149
transform 1 0 12328 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1786_
timestamp 1644511149
transform 1 0 8004 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1787_
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1788_
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1789_
timestamp 1644511149
transform 1 0 10304 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1790_
timestamp 1644511149
transform 1 0 10764 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1791_
timestamp 1644511149
transform 1 0 17112 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1792_
timestamp 1644511149
transform 1 0 12972 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1793_
timestamp 1644511149
transform 1 0 15180 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1794_
timestamp 1644511149
transform 1 0 16836 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1795_
timestamp 1644511149
transform 1 0 13064 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1796_
timestamp 1644511149
transform 1 0 18216 0 -1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1797_
timestamp 1644511149
transform 1 0 17296 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1798_
timestamp 1644511149
transform 1 0 16008 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1799_
timestamp 1644511149
transform 1 0 20424 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1800_
timestamp 1644511149
transform 1 0 22264 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1801_
timestamp 1644511149
transform 1 0 20240 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1802_
timestamp 1644511149
transform 1 0 22448 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1803_
timestamp 1644511149
transform 1 0 19596 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1804_
timestamp 1644511149
transform 1 0 20240 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1805_
timestamp 1644511149
transform 1 0 23368 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1806_
timestamp 1644511149
transform 1 0 20976 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1807_
timestamp 1644511149
transform 1 0 35144 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1808_
timestamp 1644511149
transform 1 0 35052 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1809_
timestamp 1644511149
transform 1 0 34960 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1810_
timestamp 1644511149
transform 1 0 20792 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1811_
timestamp 1644511149
transform 1 0 19872 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1812_
timestamp 1644511149
transform 1 0 19872 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1813_
timestamp 1644511149
transform 1 0 20332 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1814_
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1815_
timestamp 1644511149
transform 1 0 22632 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1816_
timestamp 1644511149
transform 1 0 6808 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1817_
timestamp 1644511149
transform 1 0 22448 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1818_
timestamp 1644511149
transform 1 0 23460 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1819_
timestamp 1644511149
transform 1 0 23000 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1820_
timestamp 1644511149
transform 1 0 25208 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1821_
timestamp 1644511149
transform 1 0 27416 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1822_
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1823_
timestamp 1644511149
transform 1 0 29992 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1824_
timestamp 1644511149
transform 1 0 30452 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1825_
timestamp 1644511149
transform 1 0 29900 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1826_
timestamp 1644511149
transform 1 0 29992 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1827_
timestamp 1644511149
transform 1 0 29808 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1828_
timestamp 1644511149
transform 1 0 24932 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1829_
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1830_
timestamp 1644511149
transform 1 0 29348 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1831_
timestamp 1644511149
transform 1 0 22448 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1832_
timestamp 1644511149
transform 1 0 22816 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1833_
timestamp 1644511149
transform 1 0 26680 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1834_
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1835_
timestamp 1644511149
transform 1 0 13340 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1836_
timestamp 1644511149
transform 1 0 22448 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1837_
timestamp 1644511149
transform 1 0 14260 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1838_
timestamp 1644511149
transform 1 0 14168 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1839_
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1840_
timestamp 1644511149
transform 1 0 11960 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1841_
timestamp 1644511149
transform 1 0 7728 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1842_
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1843_
timestamp 1644511149
transform 1 0 6992 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1844_
timestamp 1644511149
transform 1 0 7820 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1845_
timestamp 1644511149
transform 1 0 24840 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1846_
timestamp 1644511149
transform 1 0 27876 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1847_
timestamp 1644511149
transform 1 0 27692 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1848_
timestamp 1644511149
transform 1 0 30176 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1849_
timestamp 1644511149
transform 1 0 32476 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1850_
timestamp 1644511149
transform 1 0 33672 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1851_
timestamp 1644511149
transform 1 0 33580 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1852_
timestamp 1644511149
transform 1 0 33028 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1853_
timestamp 1644511149
transform 1 0 26312 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1854_
timestamp 1644511149
transform 1 0 29716 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1855_
timestamp 1644511149
transform 1 0 27508 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1856_
timestamp 1644511149
transform 1 0 27048 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1857_
timestamp 1644511149
transform 1 0 29992 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1858_
timestamp 1644511149
transform 1 0 33028 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1859_
timestamp 1644511149
transform 1 0 34868 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1860_
timestamp 1644511149
transform 1 0 32384 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1861_
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1862_
timestamp 1644511149
transform 1 0 29992 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1863_
timestamp 1644511149
transform 1 0 26680 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1864_
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1865_
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1866_
timestamp 1644511149
transform 1 0 30268 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1867_
timestamp 1644511149
transform 1 0 32292 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1868_
timestamp 1644511149
transform 1 0 32936 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1869_
timestamp 1644511149
transform 1 0 33764 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1870_
timestamp 1644511149
transform 1 0 32384 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1871_
timestamp 1644511149
transform 1 0 25852 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1872_
timestamp 1644511149
transform 1 0 25024 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1873_
timestamp 1644511149
transform 1 0 28428 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1874_
timestamp 1644511149
transform 1 0 29532 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1875_
timestamp 1644511149
transform 1 0 25944 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1876_
timestamp 1644511149
transform 1 0 29532 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1877_
timestamp 1644511149
transform 1 0 22448 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1878_
timestamp 1644511149
transform 1 0 21988 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1879_
timestamp 1644511149
transform 1 0 21804 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1880_
timestamp 1644511149
transform 1 0 24472 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1881_
timestamp 1644511149
transform 1 0 24656 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1882_
timestamp 1644511149
transform 1 0 19964 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1883_
timestamp 1644511149
transform 1 0 19044 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1884_
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1885_
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1886_
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1887_
timestamp 1644511149
transform 1 0 23644 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1888_
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1889_
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1890_
timestamp 1644511149
transform 1 0 23920 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1891_
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1892_
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1893_
timestamp 1644511149
transform 1 0 18584 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1894_
timestamp 1644511149
transform 1 0 21896 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1895_
timestamp 1644511149
transform 1 0 23828 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1896_
timestamp 1644511149
transform 1 0 18584 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1897_
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1898_
timestamp 1644511149
transform 1 0 19872 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1899_
timestamp 1644511149
transform 1 0 34684 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1900_
timestamp 1644511149
transform 1 0 36524 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1901_
timestamp 1644511149
transform 1 0 35604 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1902_
timestamp 1644511149
transform 1 0 36248 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1903_
timestamp 1644511149
transform 1 0 23368 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1904_
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1905_
timestamp 1644511149
transform 1 0 21344 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1906_
timestamp 1644511149
transform 1 0 24656 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1907_
timestamp 1644511149
transform 1 0 24288 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1908_
timestamp 1644511149
transform 1 0 20516 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1909_
timestamp 1644511149
transform 1 0 23460 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1910_
timestamp 1644511149
transform 1 0 29348 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1911_
timestamp 1644511149
transform 1 0 32752 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1912_
timestamp 1644511149
transform 1 0 32660 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1913_
timestamp 1644511149
transform 1 0 35144 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1914_
timestamp 1644511149
transform 1 0 35328 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1915_
timestamp 1644511149
transform 1 0 34960 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1916_
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1917_
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1918_
timestamp 1644511149
transform 1 0 16744 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1919_
timestamp 1644511149
transform 1 0 18492 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1920_
timestamp 1644511149
transform 1 0 18124 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1921_
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1922_
timestamp 1644511149
transform 1 0 11776 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1923_
timestamp 1644511149
transform 1 0 8464 0 -1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1924_
timestamp 1644511149
transform 1 0 9476 0 -1 31552
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1925_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14168 0 -1 34816
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1926_
timestamp 1644511149
transform 1 0 14628 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1927_
timestamp 1644511149
transform 1 0 15548 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1928_
timestamp 1644511149
transform 1 0 15364 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1929__200 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 40480 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1930__201
timestamp 1644511149
transform 1 0 32108 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1931__202
timestamp 1644511149
transform 1 0 9016 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1932__203
timestamp 1644511149
transform 1 0 2668 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1933__96
timestamp 1644511149
transform 1 0 3404 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1934__97
timestamp 1644511149
transform 1 0 25208 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1935__98
timestamp 1644511149
transform 1 0 16652 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1936__99
timestamp 1644511149
transform 1 0 25852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1937__100
timestamp 1644511149
transform 1 0 37260 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1938__101
timestamp 1644511149
transform 1 0 2024 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1939__102
timestamp 1644511149
transform 1 0 47564 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1940__103
timestamp 1644511149
transform 1 0 1472 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1941__104
timestamp 1644511149
transform 1 0 1840 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1942__105
timestamp 1644511149
transform 1 0 1472 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1943__106
timestamp 1644511149
transform 1 0 31280 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1944__107
timestamp 1644511149
transform 1 0 15916 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1945__108
timestamp 1644511149
transform 1 0 2760 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1946__109
timestamp 1644511149
transform 1 0 32752 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1947__110
timestamp 1644511149
transform 1 0 4416 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1948__111
timestamp 1644511149
transform 1 0 46828 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1949__112
timestamp 1644511149
transform 1 0 23460 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1950__113
timestamp 1644511149
transform 1 0 11592 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1951__114
timestamp 1644511149
transform 1 0 29808 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1952__115
timestamp 1644511149
transform 1 0 20240 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1953__116
timestamp 1644511149
transform 1 0 40756 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1954__117
timestamp 1644511149
transform 1 0 46828 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1955__118
timestamp 1644511149
transform 1 0 3772 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1956__119
timestamp 1644511149
transform 1 0 41032 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1957__120
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1958__121
timestamp 1644511149
transform 1 0 1840 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1959__122
timestamp 1644511149
transform 1 0 18032 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1960__123
timestamp 1644511149
transform 1 0 20056 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1961__124
timestamp 1644511149
transform 1 0 15272 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1962__125
timestamp 1644511149
transform 1 0 28796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1963__126
timestamp 1644511149
transform 1 0 2116 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1964__127
timestamp 1644511149
transform 1 0 47472 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1965__128
timestamp 1644511149
transform 1 0 30360 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1966__129
timestamp 1644511149
transform 1 0 2024 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1967__130
timestamp 1644511149
transform 1 0 22080 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1968__131
timestamp 1644511149
transform 1 0 4048 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1969__132
timestamp 1644511149
transform 1 0 38364 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1970__133
timestamp 1644511149
transform 1 0 3772 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1971__134
timestamp 1644511149
transform 1 0 47564 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1972__135
timestamp 1644511149
transform 1 0 38640 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1973__136
timestamp 1644511149
transform 1 0 45632 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1974__137
timestamp 1644511149
transform 1 0 3404 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1975__138
timestamp 1644511149
transform 1 0 35696 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1976__139
timestamp 1644511149
transform 1 0 12236 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1977__140
timestamp 1644511149
transform 1 0 46184 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1978__141
timestamp 1644511149
transform 1 0 44988 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1979__142
timestamp 1644511149
transform 1 0 39560 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1980__143
timestamp 1644511149
transform 1 0 9660 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1981__144
timestamp 1644511149
transform 1 0 7636 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1982__145
timestamp 1644511149
transform 1 0 47564 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1983__146
timestamp 1644511149
transform 1 0 33856 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1984__147
timestamp 1644511149
transform 1 0 14444 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1985__148
timestamp 1644511149
transform 1 0 2668 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1986__149
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1987__150
timestamp 1644511149
transform 1 0 2668 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1988__151
timestamp 1644511149
transform 1 0 46828 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1989__152
timestamp 1644511149
transform 1 0 44068 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1990__153
timestamp 1644511149
transform 1 0 2760 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1991__154
timestamp 1644511149
transform 1 0 28060 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1992__155
timestamp 1644511149
transform 1 0 45540 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1993__156
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1994__157
timestamp 1644511149
transform 1 0 47840 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1995__158
timestamp 1644511149
transform 1 0 10304 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1996__159
timestamp 1644511149
transform 1 0 12880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1997__160
timestamp 1644511149
transform 1 0 28060 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1998__161
timestamp 1644511149
transform 1 0 43608 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1999__162
timestamp 1644511149
transform 1 0 6716 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2000__163
timestamp 1644511149
transform 1 0 42780 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2001__164
timestamp 1644511149
transform 1 0 4416 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2002__165
timestamp 1644511149
transform 1 0 47564 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2003__166
timestamp 1644511149
transform 1 0 2116 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2004__167
timestamp 1644511149
transform 1 0 47564 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2005__168
timestamp 1644511149
transform 1 0 20700 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2006__169
timestamp 1644511149
transform 1 0 47564 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2007__170
timestamp 1644511149
transform 1 0 43884 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2008__171
timestamp 1644511149
transform 1 0 47472 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2009__172
timestamp 1644511149
transform 1 0 46828 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2010__173
timestamp 1644511149
transform 1 0 44712 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2011__174
timestamp 1644511149
transform 1 0 6440 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2012__175
timestamp 1644511149
transform 1 0 45632 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2013__176
timestamp 1644511149
transform 1 0 7912 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2014__177
timestamp 1644511149
transform 1 0 46828 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2015__178
timestamp 1644511149
transform 1 0 46828 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2016__179
timestamp 1644511149
transform 1 0 1840 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2017__180
timestamp 1644511149
transform 1 0 1840 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2018__181
timestamp 1644511149
transform 1 0 36340 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2019__182
timestamp 1644511149
transform 1 0 45632 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2020__183
timestamp 1644511149
transform 1 0 2760 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2021__184
timestamp 1644511149
transform 1 0 44160 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2022__185
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2023__186
timestamp 1644511149
transform 1 0 41676 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2024__187
timestamp 1644511149
transform 1 0 24380 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2025__188
timestamp 1644511149
transform 1 0 1840 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2026__189
timestamp 1644511149
transform 1 0 47472 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2027__190
timestamp 1644511149
transform 1 0 4048 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2028__191
timestamp 1644511149
transform 1 0 10948 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2029__192
timestamp 1644511149
transform 1 0 44896 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2030__193
timestamp 1644511149
transform 1 0 1840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2031__194
timestamp 1644511149
transform 1 0 32752 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2032__195
timestamp 1644511149
transform 1 0 21068 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2033__196
timestamp 1644511149
transform 1 0 2668 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2034__197
timestamp 1644511149
transform 1 0 2668 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2035__198
timestamp 1644511149
transform 1 0 39376 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2036__199
timestamp 1644511149
transform 1 0 2024 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2037_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7268 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2038_
timestamp 1644511149
transform 1 0 16008 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2039_
timestamp 1644511149
transform 1 0 25668 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2040_
timestamp 1644511149
transform 1 0 20056 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2041_
timestamp 1644511149
transform 1 0 17572 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2042_
timestamp 1644511149
transform 1 0 18124 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2043_
timestamp 1644511149
transform 1 0 31648 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2044_
timestamp 1644511149
transform 1 0 33580 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2045_
timestamp 1644511149
transform 1 0 32844 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2046_
timestamp 1644511149
transform 1 0 33488 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2047_
timestamp 1644511149
transform 1 0 33120 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2048_
timestamp 1644511149
transform 1 0 33672 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2049_
timestamp 1644511149
transform 1 0 32568 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2050_
timestamp 1644511149
transform 1 0 36340 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2051_
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2052_
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2053_
timestamp 1644511149
transform 1 0 37260 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2054_
timestamp 1644511149
transform 1 0 15548 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2055_
timestamp 1644511149
transform 1 0 9936 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2056_
timestamp 1644511149
transform 1 0 17756 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2057_
timestamp 1644511149
transform 1 0 12420 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2058_
timestamp 1644511149
transform 1 0 8740 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2059_
timestamp 1644511149
transform 1 0 9200 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2060_
timestamp 1644511149
transform 1 0 8096 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2061_
timestamp 1644511149
transform 1 0 4692 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2062_
timestamp 1644511149
transform 1 0 11500 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2063_
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2064_
timestamp 1644511149
transform 1 0 25760 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2065_
timestamp 1644511149
transform 1 0 16652 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2066_
timestamp 1644511149
transform 1 0 25760 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2067_
timestamp 1644511149
transform 1 0 36340 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2068_
timestamp 1644511149
transform 1 0 2024 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2069_
timestamp 1644511149
transform 1 0 46276 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_2  _2070_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6624 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_8  _2071_
timestamp 1644511149
transform 1 0 14076 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2072_
timestamp 1644511149
transform 1 0 29164 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2073_
timestamp 1644511149
transform 1 0 5336 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2074_
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2075_
timestamp 1644511149
transform 1 0 40020 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2076_
timestamp 1644511149
transform 1 0 32108 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2077_
timestamp 1644511149
transform 1 0 8924 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2078_
timestamp 1644511149
transform 1 0 1748 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2079_
timestamp 1644511149
transform 1 0 1748 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2080_
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2081_
timestamp 1644511149
transform 1 0 31188 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2082_
timestamp 1644511149
transform 1 0 16744 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2083_
timestamp 1644511149
transform 1 0 2024 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2084_
timestamp 1644511149
transform 1 0 31372 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2085_
timestamp 1644511149
transform 1 0 3956 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2086_
timestamp 1644511149
transform 1 0 46276 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2087_
timestamp 1644511149
transform 1 0 23368 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2088_
timestamp 1644511149
transform 1 0 11500 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2089_
timestamp 1644511149
transform 1 0 29716 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2090_
timestamp 1644511149
transform 1 0 20056 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2091_
timestamp 1644511149
transform 1 0 41400 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2092_
timestamp 1644511149
transform 1 0 46276 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2093_
timestamp 1644511149
transform 1 0 3772 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2094_
timestamp 1644511149
transform 1 0 41032 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2095_
timestamp 1644511149
transform 1 0 1748 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2096_
timestamp 1644511149
transform 1 0 1748 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2097_
timestamp 1644511149
transform 1 0 17940 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2098_
timestamp 1644511149
transform 1 0 19964 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2099_
timestamp 1644511149
transform 1 0 14904 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2100_
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2101_
timestamp 1644511149
transform 1 0 1932 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2102_
timestamp 1644511149
transform 1 0 46276 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2103_
timestamp 1644511149
transform 1 0 29716 0 1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2104_
timestamp 1644511149
transform 1 0 2024 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2105_
timestamp 1644511149
transform 1 0 22724 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2106_
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2107_
timestamp 1644511149
transform 1 0 39008 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2108_
timestamp 1644511149
transform 1 0 3772 0 1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2109_
timestamp 1644511149
transform 1 0 46276 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2110_
timestamp 1644511149
transform 1 0 38640 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2111_
timestamp 1644511149
transform 1 0 46276 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2112_
timestamp 1644511149
transform 1 0 1380 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2113_
timestamp 1644511149
transform 1 0 11684 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2114_
timestamp 1644511149
transform 1 0 18308 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2115_
timestamp 1644511149
transform 1 0 19412 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2116_
timestamp 1644511149
transform 1 0 20148 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2117_
timestamp 1644511149
transform 1 0 20792 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2118_
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2119_
timestamp 1644511149
transform 1 0 9108 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2120_
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2121_
timestamp 1644511149
transform 1 0 34868 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2122_
timestamp 1644511149
transform 1 0 12236 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2123_
timestamp 1644511149
transform 1 0 46276 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2124_
timestamp 1644511149
transform 1 0 44896 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2125_
timestamp 1644511149
transform 1 0 39836 0 1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2126_
timestamp 1644511149
transform 1 0 9660 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2127_
timestamp 1644511149
transform 1 0 6624 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2128_
timestamp 1644511149
transform 1 0 46276 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2129_
timestamp 1644511149
transform 1 0 6532 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2130_
timestamp 1644511149
transform 1 0 30360 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2131_
timestamp 1644511149
transform 1 0 36984 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2132_
timestamp 1644511149
transform 1 0 37444 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2133_
timestamp 1644511149
transform 1 0 37352 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2134_
timestamp 1644511149
transform 1 0 37352 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2135_
timestamp 1644511149
transform 1 0 36892 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2136_
timestamp 1644511149
transform 1 0 36064 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2137_
timestamp 1644511149
transform 1 0 36156 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2138_
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2139_
timestamp 1644511149
transform 1 0 15548 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2140_
timestamp 1644511149
transform 1 0 33396 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2141_
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2142_
timestamp 1644511149
transform 1 0 21804 0 -1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2143_
timestamp 1644511149
transform 1 0 33764 0 -1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2144_
timestamp 1644511149
transform 1 0 14444 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2145_
timestamp 1644511149
transform 1 0 1380 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2146_
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2147_
timestamp 1644511149
transform 1 0 1748 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2148_
timestamp 1644511149
transform 1 0 46276 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2149_
timestamp 1644511149
transform 1 0 43976 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2150_
timestamp 1644511149
transform 1 0 2116 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2151_
timestamp 1644511149
transform 1 0 28060 0 -1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2152_
timestamp 1644511149
transform 1 0 46276 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2153_
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2154_
timestamp 1644511149
transform 1 0 46276 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2155_
timestamp 1644511149
transform 1 0 7452 0 -1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2156_
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2157_
timestamp 1644511149
transform 1 0 26956 0 1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2158_
timestamp 1644511149
transform 1 0 46276 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2159_
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2160_
timestamp 1644511149
transform 1 0 42596 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2161_
timestamp 1644511149
transform 1 0 1472 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2162_
timestamp 1644511149
transform 1 0 46276 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2163_
timestamp 1644511149
transform 1 0 2024 0 -1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2164_
timestamp 1644511149
transform 1 0 46276 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2165_
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2166_
timestamp 1644511149
transform 1 0 46276 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2167_
timestamp 1644511149
transform 1 0 45172 0 1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2168_
timestamp 1644511149
transform 1 0 46276 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2169_
timestamp 1644511149
transform 1 0 46276 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2170_
timestamp 1644511149
transform 1 0 44988 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2171_
timestamp 1644511149
transform 1 0 6440 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2172_
timestamp 1644511149
transform 1 0 46276 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2173_
timestamp 1644511149
transform 1 0 7912 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2174_
timestamp 1644511149
transform 1 0 46276 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2175_
timestamp 1644511149
transform 1 0 46276 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2176_
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2177_
timestamp 1644511149
transform 1 0 1380 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2178_
timestamp 1644511149
transform 1 0 36248 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2179_
timestamp 1644511149
transform 1 0 46276 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2180_
timestamp 1644511149
transform 1 0 1748 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2181_
timestamp 1644511149
transform 1 0 44160 0 -1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2182_
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2183_
timestamp 1644511149
transform 1 0 42596 0 1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2184_
timestamp 1644511149
transform 1 0 24380 0 1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2185_
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2186_
timestamp 1644511149
transform 1 0 46276 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2187_
timestamp 1644511149
transform 1 0 1380 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2188_
timestamp 1644511149
transform 1 0 11592 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2189_
timestamp 1644511149
transform 1 0 45172 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2190_
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2191_
timestamp 1644511149
transform 1 0 32200 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2192_
timestamp 1644511149
transform 1 0 21988 0 1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2193_
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2194_
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2195_
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2196_
timestamp 1644511149
transform 1 0 2024 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i
timestamp 1644511149
transform 1 0 22080 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 22632 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 23552 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 18400 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 30084 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 20700 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 28428 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 18400 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 17848 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 28244 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_4_0_wb_clk_i
timestamp 1644511149
transform 1 0 18308 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_5_0_wb_clk_i
timestamp 1644511149
transform 1 0 19688 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_6_0_wb_clk_i
timestamp 1644511149
transform 1 0 30452 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_7_0_wb_clk_i
timestamp 1644511149
transform 1 0 30636 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 19780 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 15732 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 19596 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_4_0_wb_clk_i
timestamp 1644511149
transform 1 0 25852 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_5_0_wb_clk_i
timestamp 1644511149
transform 1 0 28888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_6_0_wb_clk_i
timestamp 1644511149
transform 1 0 30176 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_7_0_wb_clk_i
timestamp 1644511149
transform 1 0 32384 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_8_0_wb_clk_i
timestamp 1644511149
transform 1 0 17572 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_9_0_wb_clk_i
timestamp 1644511149
transform 1 0 19964 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_10_0_wb_clk_i
timestamp 1644511149
transform 1 0 17664 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_11_0_wb_clk_i
timestamp 1644511149
transform 1 0 20424 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_12_0_wb_clk_i
timestamp 1644511149
transform 1 0 29348 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_13_0_wb_clk_i
timestamp 1644511149
transform 1 0 31464 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_14_0_wb_clk_i
timestamp 1644511149
transform 1 0 28060 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_15_0_wb_clk_i
timestamp 1644511149
transform 1 0 31372 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input1
timestamp 1644511149
transform 1 0 47656 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input2
timestamp 1644511149
transform 1 0 1748 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp 1644511149
transform 1 0 14076 0 1 48960
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1644511149
transform 1 0 22632 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1644511149
transform 1 0 1748 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input6
timestamp 1644511149
transform 1 0 47656 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input7
timestamp 1644511149
transform 1 0 47840 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1644511149
transform 1 0 22264 0 1 47872
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1644511149
transform 1 0 12696 0 1 48960
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1644511149
transform 1 0 17848 0 1 48960
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input11
timestamp 1644511149
transform 1 0 27140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input12
timestamp 1644511149
transform 1 0 32936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input13
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input14
timestamp 1644511149
transform 1 0 10212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input15
timestamp 1644511149
transform 1 0 1748 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1644511149
transform 1 0 15272 0 -1 48960
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 1644511149
transform 1 0 47840 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1644511149
transform 1 0 47288 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp 1644511149
transform 1 0 46184 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1644511149
transform 1 0 47932 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1644511149
transform 1 0 21068 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1644511149
transform 1 0 1748 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1644511149
transform 1 0 4140 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1644511149
transform 1 0 47840 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1644511149
transform 1 0 1748 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input26
timestamp 1644511149
transform 1 0 47656 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1644511149
transform 1 0 13984 0 -1 48960
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1644511149
transform 1 0 47840 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1644511149
transform 1 0 47840 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input30
timestamp 1644511149
transform 1 0 1380 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input31
timestamp 1644511149
transform 1 0 4600 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1644511149
transform 1 0 20056 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1644511149
transform 1 0 1748 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input34
timestamp 1644511149
transform 1 0 39008 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1644511149
transform 1 0 27324 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input36
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input37
timestamp 1644511149
transform 1 0 38088 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input38
timestamp 1644511149
transform 1 0 20056 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input40
timestamp 1644511149
transform 1 0 6716 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1644511149
transform 1 0 47840 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input42
timestamp 1644511149
transform 1 0 1748 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1644511149
transform 1 0 27876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input44
timestamp 1644511149
transform 1 0 1748 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1644511149
transform 1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input46
timestamp 1644511149
transform 1 0 43240 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input47
timestamp 1644511149
transform 1 0 44988 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1644511149
transform 1 0 1748 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1644511149
transform 1 0 25208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1644511149
transform 1 0 36156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input51
timestamp 1644511149
transform 1 0 47840 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input52
timestamp 1644511149
transform 1 0 19320 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input53
timestamp 1644511149
transform 1 0 25944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input54
timestamp 1644511149
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1644511149
transform 1 0 28428 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1644511149
transform 1 0 47932 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1644511149
transform 1 0 47840 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input58
timestamp 1644511149
transform 1 0 17480 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input59
timestamp 1644511149
transform 1 0 47656 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1644511149
transform 1 0 47840 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input61
timestamp 1644511149
transform 1 0 35052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input62
timestamp 1644511149
transform 1 0 47656 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1644511149
transform 1 0 33856 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input64
timestamp 1644511149
transform 1 0 14536 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input65
timestamp 1644511149
transform 1 0 1748 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input66
timestamp 1644511149
transform 1 0 46276 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1644511149
transform 1 0 47840 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1644511149
transform 1 0 25852 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input69
timestamp 1644511149
transform 1 0 47840 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input70
timestamp 1644511149
transform 1 0 1748 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input71
timestamp 1644511149
transform 1 0 2760 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input72
timestamp 1644511149
transform 1 0 2024 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp 1644511149
transform 1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1644511149
transform 1 0 9936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input75
timestamp 1644511149
transform 1 0 47840 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input76
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input77
timestamp 1644511149
transform 1 0 41400 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input78
timestamp 1644511149
transform 1 0 47656 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input79
timestamp 1644511149
transform 1 0 11868 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input80
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input81
timestamp 1644511149
transform 1 0 47840 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input82
timestamp 1644511149
transform 1 0 46552 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input83
timestamp 1644511149
transform 1 0 1748 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input84
timestamp 1644511149
transform 1 0 47840 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input85
timestamp 1644511149
transform 1 0 1748 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input86
timestamp 1644511149
transform 1 0 38456 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input87
timestamp 1644511149
transform 1 0 47840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input88
timestamp 1644511149
transform 1 0 8648 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input90
timestamp 1644511149
transform 1 0 47840 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input91
timestamp 1644511149
transform 1 0 43884 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input92
timestamp 1644511149
transform 1 0 47840 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input93
timestamp 1644511149
transform 1 0 47840 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input94
timestamp 1644511149
transform 1 0 1748 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input95
timestamp 1644511149
transform 1 0 47840 0 1 25024
box -38 -48 406 592
<< labels >>
rlabel metal3 s 49200 31968 50000 32088 6 active
port 0 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 25134 51200 25190 52000 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 49200 15648 50000 15768 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 21270 51200 21326 52000 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 49200 2048 50000 2168 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 io_in[18]
port 10 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 49200 18368 50000 18488 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 0 30608 800 30728 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 49200 21088 50000 21208 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 49200 32648 50000 32768 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 49200 23128 50000 23248 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 2594 51200 2650 52000 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 46386 51200 46442 52000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 9034 51200 9090 52000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 31574 51200 31630 52000 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 49200 47608 50000 47728 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 49200 20408 50000 20528 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 35438 51200 35494 52000 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 49200 2728 50000 2848 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 3882 51200 3938 52000 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 io_oeb[0]
port 39 nsew signal bidirectional
rlabel metal3 s 49200 24488 50000 24608 6 io_oeb[10]
port 40 nsew signal bidirectional
rlabel metal2 s 45098 0 45154 800 6 io_oeb[11]
port 41 nsew signal bidirectional
rlabel metal2 s 5814 0 5870 800 6 io_oeb[12]
port 42 nsew signal bidirectional
rlabel metal2 s 48318 0 48374 800 6 io_oeb[13]
port 43 nsew signal bidirectional
rlabel metal2 s 7746 51200 7802 52000 6 io_oeb[14]
port 44 nsew signal bidirectional
rlabel metal3 s 49200 43528 50000 43648 6 io_oeb[15]
port 45 nsew signal bidirectional
rlabel metal3 s 49200 4768 50000 4888 6 io_oeb[16]
port 46 nsew signal bidirectional
rlabel metal3 s 0 6808 800 6928 6 io_oeb[17]
port 47 nsew signal bidirectional
rlabel metal3 s 0 41488 800 41608 6 io_oeb[18]
port 48 nsew signal bidirectional
rlabel metal2 s 36726 0 36782 800 6 io_oeb[19]
port 49 nsew signal bidirectional
rlabel metal2 s 43166 51200 43222 52000 6 io_oeb[1]
port 50 nsew signal bidirectional
rlabel metal3 s 49200 46928 50000 47048 6 io_oeb[20]
port 51 nsew signal bidirectional
rlabel metal3 s 0 9528 800 9648 6 io_oeb[21]
port 52 nsew signal bidirectional
rlabel metal2 s 45098 51200 45154 52000 6 io_oeb[22]
port 53 nsew signal bidirectional
rlabel metal3 s 0 26528 800 26648 6 io_oeb[23]
port 54 nsew signal bidirectional
rlabel metal3 s 49200 51688 50000 51808 6 io_oeb[24]
port 55 nsew signal bidirectional
rlabel metal2 s 24490 51200 24546 52000 6 io_oeb[25]
port 56 nsew signal bidirectional
rlabel metal3 s 0 23128 800 23248 6 io_oeb[26]
port 57 nsew signal bidirectional
rlabel metal3 s 49200 28568 50000 28688 6 io_oeb[27]
port 58 nsew signal bidirectional
rlabel metal2 s 1306 51200 1362 52000 6 io_oeb[28]
port 59 nsew signal bidirectional
rlabel metal2 s 12254 0 12310 800 6 io_oeb[29]
port 60 nsew signal bidirectional
rlabel metal3 s 0 51688 800 51808 6 io_oeb[2]
port 61 nsew signal bidirectional
rlabel metal2 s 49606 51200 49662 52000 6 io_oeb[30]
port 62 nsew signal bidirectional
rlabel metal3 s 0 3408 800 3528 6 io_oeb[31]
port 63 nsew signal bidirectional
rlabel metal2 s 33506 0 33562 800 6 io_oeb[32]
port 64 nsew signal bidirectional
rlabel metal2 s 22558 51200 22614 52000 6 io_oeb[33]
port 65 nsew signal bidirectional
rlabel metal3 s 0 17688 800 17808 6 io_oeb[34]
port 66 nsew signal bidirectional
rlabel metal3 s 0 13608 800 13728 6 io_oeb[35]
port 67 nsew signal bidirectional
rlabel metal2 s 39946 0 40002 800 6 io_oeb[36]
port 68 nsew signal bidirectional
rlabel metal3 s 0 39448 800 39568 6 io_oeb[37]
port 69 nsew signal bidirectional
rlabel metal3 s 49200 45568 50000 45688 6 io_oeb[3]
port 70 nsew signal bidirectional
rlabel metal3 s 0 44888 800 45008 6 io_oeb[4]
port 71 nsew signal bidirectional
rlabel metal3 s 49200 36728 50000 36848 6 io_oeb[5]
port 72 nsew signal bidirectional
rlabel metal2 s 21270 0 21326 800 6 io_oeb[6]
port 73 nsew signal bidirectional
rlabel metal3 s 49200 17008 50000 17128 6 io_oeb[7]
port 74 nsew signal bidirectional
rlabel metal3 s 49200 49648 50000 49768 6 io_oeb[8]
port 75 nsew signal bidirectional
rlabel metal3 s 49200 16328 50000 16448 6 io_oeb[9]
port 76 nsew signal bidirectional
rlabel metal2 s 36082 51200 36138 52000 6 io_out[0]
port 77 nsew signal bidirectional
rlabel metal3 s 49200 44208 50000 44328 6 io_out[10]
port 78 nsew signal bidirectional
rlabel metal3 s 49200 9528 50000 9648 6 io_out[11]
port 79 nsew signal bidirectional
rlabel metal2 s 48962 0 49018 800 6 io_out[12]
port 80 nsew signal bidirectional
rlabel metal2 s 47030 0 47086 800 6 io_out[13]
port 81 nsew signal bidirectional
rlabel metal3 s 49200 12248 50000 12368 6 io_out[14]
port 82 nsew signal bidirectional
rlabel metal2 s 37370 0 37426 800 6 io_out[15]
port 83 nsew signal bidirectional
rlabel metal2 s 37370 51200 37426 52000 6 io_out[16]
port 84 nsew signal bidirectional
rlabel metal2 s 38658 51200 38714 52000 6 io_out[17]
port 85 nsew signal bidirectional
rlabel metal2 s 15474 51200 15530 52000 6 io_out[18]
port 86 nsew signal bidirectional
rlabel metal3 s 49200 3408 50000 3528 6 io_out[19]
port 87 nsew signal bidirectional
rlabel metal2 s 12898 0 12954 800 6 io_out[1]
port 88 nsew signal bidirectional
rlabel metal2 s 11610 0 11666 800 6 io_out[20]
port 89 nsew signal bidirectional
rlabel metal3 s 0 48288 800 48408 6 io_out[21]
port 90 nsew signal bidirectional
rlabel metal2 s 34794 51200 34850 52000 6 io_out[22]
port 91 nsew signal bidirectional
rlabel metal2 s 14830 51200 14886 52000 6 io_out[23]
port 92 nsew signal bidirectional
rlabel metal3 s 0 46248 800 46368 6 io_out[24]
port 93 nsew signal bidirectional
rlabel metal3 s 0 34008 800 34128 6 io_out[25]
port 94 nsew signal bidirectional
rlabel metal3 s 0 27208 800 27328 6 io_out[26]
port 95 nsew signal bidirectional
rlabel metal3 s 49200 7488 50000 7608 6 io_out[27]
port 96 nsew signal bidirectional
rlabel metal2 s 44454 0 44510 800 6 io_out[28]
port 97 nsew signal bidirectional
rlabel metal3 s 0 5448 800 5568 6 io_out[29]
port 98 nsew signal bidirectional
rlabel metal3 s 49200 35368 50000 35488 6 io_out[2]
port 99 nsew signal bidirectional
rlabel metal2 s 28354 51200 28410 52000 6 io_out[30]
port 100 nsew signal bidirectional
rlabel metal3 s 49200 46248 50000 46368 6 io_out[31]
port 101 nsew signal bidirectional
rlabel metal2 s 42522 0 42578 800 6 io_out[32]
port 102 nsew signal bidirectional
rlabel metal3 s 49200 10888 50000 11008 6 io_out[33]
port 103 nsew signal bidirectional
rlabel metal3 s 0 51008 800 51128 6 io_out[34]
port 104 nsew signal bidirectional
rlabel metal2 s 13542 0 13598 800 6 io_out[35]
port 105 nsew signal bidirectional
rlabel metal2 s 27066 51200 27122 52000 6 io_out[36]
port 106 nsew signal bidirectional
rlabel metal2 s 48318 51200 48374 52000 6 io_out[37]
port 107 nsew signal bidirectional
rlabel metal2 s 45742 51200 45798 52000 6 io_out[3]
port 108 nsew signal bidirectional
rlabel metal2 s 39946 51200 40002 52000 6 io_out[4]
port 109 nsew signal bidirectional
rlabel metal2 s 10322 51200 10378 52000 6 io_out[5]
port 110 nsew signal bidirectional
rlabel metal2 s 7102 51200 7158 52000 6 io_out[6]
port 111 nsew signal bidirectional
rlabel metal3 s 49200 34008 50000 34128 6 io_out[7]
port 112 nsew signal bidirectional
rlabel metal2 s 2594 0 2650 800 6 io_out[8]
port 113 nsew signal bidirectional
rlabel metal2 s 8390 51200 8446 52000 6 io_out[9]
port 114 nsew signal bidirectional
rlabel metal3 s 0 8168 800 8288 6 rambus_wb_ack_i
port 115 nsew signal input
rlabel metal3 s 49200 40128 50000 40248 6 rambus_wb_adr_o[0]
port 116 nsew signal bidirectional
rlabel metal3 s 0 46928 800 47048 6 rambus_wb_adr_o[1]
port 117 nsew signal bidirectional
rlabel metal2 s 10966 51200 11022 52000 6 rambus_wb_adr_o[2]
port 118 nsew signal bidirectional
rlabel metal3 s 49200 6128 50000 6248 6 rambus_wb_adr_o[3]
port 119 nsew signal bidirectional
rlabel metal3 s 49200 51008 50000 51128 6 rambus_wb_adr_o[4]
port 120 nsew signal bidirectional
rlabel metal3 s 49200 17688 50000 17808 6 rambus_wb_adr_o[5]
port 121 nsew signal bidirectional
rlabel metal3 s 49200 6808 50000 6928 6 rambus_wb_adr_o[6]
port 122 nsew signal bidirectional
rlabel metal3 s 49200 29248 50000 29368 6 rambus_wb_adr_o[7]
port 123 nsew signal bidirectional
rlabel metal2 s 9034 0 9090 800 6 rambus_wb_adr_o[8]
port 124 nsew signal bidirectional
rlabel metal3 s 0 2048 800 2168 6 rambus_wb_adr_o[9]
port 125 nsew signal bidirectional
rlabel metal3 s 0 18368 800 18488 6 rambus_wb_clk_o
port 126 nsew signal bidirectional
rlabel metal2 s 5170 51200 5226 52000 6 rambus_wb_cyc_o
port 127 nsew signal bidirectional
rlabel metal2 s 13542 51200 13598 52000 6 rambus_wb_dat_i[0]
port 128 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 rambus_wb_dat_i[10]
port 129 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 rambus_wb_dat_i[11]
port 130 nsew signal input
rlabel metal3 s 49200 688 50000 808 6 rambus_wb_dat_i[12]
port 131 nsew signal input
rlabel metal3 s 49200 13608 50000 13728 6 rambus_wb_dat_i[13]
port 132 nsew signal input
rlabel metal2 s 21914 51200 21970 52000 6 rambus_wb_dat_i[14]
port 133 nsew signal input
rlabel metal2 s 12898 51200 12954 52000 6 rambus_wb_dat_i[15]
port 134 nsew signal input
rlabel metal2 s 18050 51200 18106 52000 6 rambus_wb_dat_i[16]
port 135 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 rambus_wb_dat_i[17]
port 136 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 rambus_wb_dat_i[18]
port 137 nsew signal input
rlabel metal3 s 0 34688 800 34808 6 rambus_wb_dat_i[19]
port 138 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 rambus_wb_dat_i[1]
port 139 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 rambus_wb_dat_i[20]
port 140 nsew signal input
rlabel metal2 s 16118 51200 16174 52000 6 rambus_wb_dat_i[21]
port 141 nsew signal input
rlabel metal3 s 49200 8168 50000 8288 6 rambus_wb_dat_i[22]
port 142 nsew signal input
rlabel metal3 s 49200 31288 50000 31408 6 rambus_wb_dat_i[23]
port 143 nsew signal input
rlabel metal3 s 49200 33328 50000 33448 6 rambus_wb_dat_i[24]
port 144 nsew signal input
rlabel metal3 s 49200 38768 50000 38888 6 rambus_wb_dat_i[25]
port 145 nsew signal input
rlabel metal2 s 23846 51200 23902 52000 6 rambus_wb_dat_i[26]
port 146 nsew signal input
rlabel metal3 s 0 36728 800 36848 6 rambus_wb_dat_i[27]
port 147 nsew signal input
rlabel metal2 s 18 51200 74 52000 6 rambus_wb_dat_i[28]
port 148 nsew signal input
rlabel metal3 s 49200 42168 50000 42288 6 rambus_wb_dat_i[29]
port 149 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 rambus_wb_dat_i[2]
port 150 nsew signal input
rlabel metal3 s 49200 10208 50000 10328 6 rambus_wb_dat_i[30]
port 151 nsew signal input
rlabel metal2 s 14186 51200 14242 52000 6 rambus_wb_dat_i[31]
port 152 nsew signal input
rlabel metal3 s 49200 29928 50000 30048 6 rambus_wb_dat_i[3]
port 153 nsew signal input
rlabel metal3 s 49200 23808 50000 23928 6 rambus_wb_dat_i[4]
port 154 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 rambus_wb_dat_i[5]
port 155 nsew signal input
rlabel metal2 s 4526 51200 4582 52000 6 rambus_wb_dat_i[6]
port 156 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 rambus_wb_dat_i[7]
port 157 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 rambus_wb_dat_i[8]
port 158 nsew signal input
rlabel metal2 s 40590 51200 40646 52000 6 rambus_wb_dat_i[9]
port 159 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 rambus_wb_dat_o[0]
port 160 nsew signal bidirectional
rlabel metal2 s 30286 0 30342 800 6 rambus_wb_dat_o[10]
port 161 nsew signal bidirectional
rlabel metal2 s 20626 0 20682 800 6 rambus_wb_dat_o[11]
port 162 nsew signal bidirectional
rlabel metal2 s 41878 0 41934 800 6 rambus_wb_dat_o[12]
port 163 nsew signal bidirectional
rlabel metal3 s 49200 34688 50000 34808 6 rambus_wb_dat_o[13]
port 164 nsew signal bidirectional
rlabel metal3 s 0 50328 800 50448 6 rambus_wb_dat_o[14]
port 165 nsew signal bidirectional
rlabel metal2 s 42522 51200 42578 52000 6 rambus_wb_dat_o[15]
port 166 nsew signal bidirectional
rlabel metal2 s 1306 0 1362 800 6 rambus_wb_dat_o[16]
port 167 nsew signal bidirectional
rlabel metal3 s 0 29928 800 30048 6 rambus_wb_dat_o[17]
port 168 nsew signal bidirectional
rlabel metal2 s 18050 0 18106 800 6 rambus_wb_dat_o[18]
port 169 nsew signal bidirectional
rlabel metal2 s 20626 51200 20682 52000 6 rambus_wb_dat_o[19]
port 170 nsew signal bidirectional
rlabel metal3 s 0 10208 800 10328 6 rambus_wb_dat_o[1]
port 171 nsew signal bidirectional
rlabel metal2 s 15474 0 15530 800 6 rambus_wb_dat_o[20]
port 172 nsew signal bidirectional
rlabel metal2 s 30930 0 30986 800 6 rambus_wb_dat_o[21]
port 173 nsew signal bidirectional
rlabel metal3 s 0 31968 800 32088 6 rambus_wb_dat_o[22]
port 174 nsew signal bidirectional
rlabel metal3 s 49200 19728 50000 19848 6 rambus_wb_dat_o[23]
port 175 nsew signal bidirectional
rlabel metal2 s 30930 51200 30986 52000 6 rambus_wb_dat_o[24]
port 176 nsew signal bidirectional
rlabel metal3 s 0 16328 800 16448 6 rambus_wb_dat_o[25]
port 177 nsew signal bidirectional
rlabel metal2 s 23202 51200 23258 52000 6 rambus_wb_dat_o[26]
port 178 nsew signal bidirectional
rlabel metal3 s 0 28568 800 28688 6 rambus_wb_dat_o[27]
port 179 nsew signal bidirectional
rlabel metal3 s 49200 50328 50000 50448 6 rambus_wb_dat_o[28]
port 180 nsew signal bidirectional
rlabel metal3 s 0 48968 800 49088 6 rambus_wb_dat_o[29]
port 181 nsew signal bidirectional
rlabel metal2 s 31574 0 31630 800 6 rambus_wb_dat_o[2]
port 182 nsew signal bidirectional
rlabel metal3 s 49200 41488 50000 41608 6 rambus_wb_dat_o[30]
port 183 nsew signal bidirectional
rlabel metal2 s 46386 0 46442 800 6 rambus_wb_dat_o[31]
port 184 nsew signal bidirectional
rlabel metal2 s 17406 51200 17462 52000 6 rambus_wb_dat_o[3]
port 185 nsew signal bidirectional
rlabel metal3 s 0 32648 800 32768 6 rambus_wb_dat_o[4]
port 186 nsew signal bidirectional
rlabel metal2 s 32218 51200 32274 52000 6 rambus_wb_dat_o[5]
port 187 nsew signal bidirectional
rlabel metal2 s 5170 0 5226 800 6 rambus_wb_dat_o[6]
port 188 nsew signal bidirectional
rlabel metal3 s 49200 14288 50000 14408 6 rambus_wb_dat_o[7]
port 189 nsew signal bidirectional
rlabel metal2 s 23846 0 23902 800 6 rambus_wb_dat_o[8]
port 190 nsew signal bidirectional
rlabel metal2 s 12254 51200 12310 52000 6 rambus_wb_dat_o[9]
port 191 nsew signal bidirectional
rlabel metal3 s 0 8848 800 8968 6 rambus_wb_rst_o
port 192 nsew signal bidirectional
rlabel metal2 s 41234 0 41290 800 6 rambus_wb_sel_o[0]
port 193 nsew signal bidirectional
rlabel metal2 s 32862 51200 32918 52000 6 rambus_wb_sel_o[1]
port 194 nsew signal bidirectional
rlabel metal2 s 9678 51200 9734 52000 6 rambus_wb_sel_o[2]
port 195 nsew signal bidirectional
rlabel metal3 s 0 33328 800 33448 6 rambus_wb_sel_o[3]
port 196 nsew signal bidirectional
rlabel metal2 s 29642 51200 29698 52000 6 rambus_wb_stb_o
port 197 nsew signal bidirectional
rlabel metal3 s 0 4768 800 4888 6 rambus_wb_we_o
port 198 nsew signal bidirectional
rlabel metal4 s 4208 2128 4528 49552 6 vccd1
port 199 nsew power input
rlabel metal4 s 34928 2128 35248 49552 6 vccd1
port 199 nsew power input
rlabel metal4 s 19568 2128 19888 49552 6 vssd1
port 200 nsew ground input
rlabel metal3 s 49200 1368 50000 1488 6 wb_clk_i
port 201 nsew signal input
rlabel metal2 s 26422 51200 26478 52000 6 wb_rst_i
port 202 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 wbs_ack_o
port 203 nsew signal bidirectional
rlabel metal3 s 0 31288 800 31408 6 wbs_adr_i[0]
port 204 nsew signal input
rlabel metal2 s 38014 51200 38070 52000 6 wbs_adr_i[10]
port 205 nsew signal input
rlabel metal2 s 19982 51200 20038 52000 6 wbs_adr_i[11]
port 206 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 wbs_adr_i[12]
port 207 nsew signal input
rlabel metal2 s 6458 51200 6514 52000 6 wbs_adr_i[13]
port 208 nsew signal input
rlabel metal3 s 49200 27888 50000 28008 6 wbs_adr_i[14]
port 209 nsew signal input
rlabel metal3 s 0 688 800 808 6 wbs_adr_i[15]
port 210 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 wbs_adr_i[16]
port 211 nsew signal input
rlabel metal3 s 0 44208 800 44328 6 wbs_adr_i[17]
port 212 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 wbs_adr_i[18]
port 213 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 wbs_adr_i[19]
port 214 nsew signal input
rlabel metal2 s 44454 51200 44510 52000 6 wbs_adr_i[1]
port 215 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 wbs_adr_i[20]
port 216 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 wbs_adr_i[21]
port 217 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wbs_adr_i[22]
port 218 nsew signal input
rlabel metal3 s 49200 5448 50000 5568 6 wbs_adr_i[23]
port 219 nsew signal input
rlabel metal2 s 19338 51200 19394 52000 6 wbs_adr_i[24]
port 220 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_adr_i[25]
port 221 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_adr_i[26]
port 222 nsew signal input
rlabel metal2 s 28998 51200 29054 52000 6 wbs_adr_i[27]
port 223 nsew signal input
rlabel metal3 s 49200 22448 50000 22568 6 wbs_adr_i[28]
port 224 nsew signal input
rlabel metal3 s 49200 40808 50000 40928 6 wbs_adr_i[29]
port 225 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_adr_i[2]
port 226 nsew signal input
rlabel metal2 s 48962 51200 49018 52000 6 wbs_adr_i[30]
port 227 nsew signal input
rlabel metal3 s 49200 14968 50000 15088 6 wbs_adr_i[31]
port 228 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 wbs_adr_i[3]
port 229 nsew signal input
rlabel metal2 s 47674 51200 47730 52000 6 wbs_adr_i[4]
port 230 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 wbs_adr_i[5]
port 231 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 wbs_adr_i[6]
port 232 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 wbs_adr_i[7]
port 233 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 wbs_adr_i[8]
port 234 nsew signal input
rlabel metal3 s 49200 8848 50000 8968 6 wbs_adr_i[9]
port 235 nsew signal input
rlabel metal2 s 25778 51200 25834 52000 6 wbs_cyc_i
port 236 nsew signal input
rlabel metal3 s 49200 38088 50000 38208 6 wbs_dat_i[0]
port 237 nsew signal input
rlabel metal2 s 662 51200 718 52000 6 wbs_dat_i[10]
port 238 nsew signal input
rlabel metal2 s 3238 51200 3294 52000 6 wbs_dat_i[11]
port 239 nsew signal input
rlabel metal2 s 1950 51200 2006 52000 6 wbs_dat_i[12]
port 240 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wbs_dat_i[13]
port 241 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 wbs_dat_i[14]
port 242 nsew signal input
rlabel metal3 s 49200 21768 50000 21888 6 wbs_dat_i[15]
port 243 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 wbs_dat_i[16]
port 244 nsew signal input
rlabel metal2 s 41878 51200 41934 52000 6 wbs_dat_i[17]
port 245 nsew signal input
rlabel metal3 s 49200 48968 50000 49088 6 wbs_dat_i[18]
port 246 nsew signal input
rlabel metal2 s 11610 51200 11666 52000 6 wbs_dat_i[19]
port 247 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_dat_i[1]
port 248 nsew signal input
rlabel metal3 s 49200 25848 50000 25968 6 wbs_dat_i[20]
port 249 nsew signal input
rlabel metal3 s 49200 48288 50000 48408 6 wbs_dat_i[21]
port 250 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 wbs_dat_i[22]
port 251 nsew signal input
rlabel metal3 s 49200 36048 50000 36168 6 wbs_dat_i[23]
port 252 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 wbs_dat_i[24]
port 253 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 wbs_dat_i[25]
port 254 nsew signal input
rlabel metal2 s 47030 51200 47086 52000 6 wbs_dat_i[26]
port 255 nsew signal input
rlabel metal2 s 18694 51200 18750 52000 6 wbs_dat_i[27]
port 256 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_i[28]
port 257 nsew signal input
rlabel metal3 s 49200 27208 50000 27328 6 wbs_dat_i[29]
port 258 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 wbs_dat_i[2]
port 259 nsew signal input
rlabel metal3 s 49200 11568 50000 11688 6 wbs_dat_i[30]
port 260 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 wbs_dat_i[31]
port 261 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 wbs_dat_i[3]
port 262 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_dat_i[4]
port 263 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 wbs_dat_i[5]
port 264 nsew signal input
rlabel metal3 s 49200 19048 50000 19168 6 wbs_dat_i[6]
port 265 nsew signal input
rlabel metal2 s 43810 51200 43866 52000 6 wbs_dat_i[7]
port 266 nsew signal input
rlabel metal3 s 49200 42848 50000 42968 6 wbs_dat_i[8]
port 267 nsew signal input
rlabel metal3 s 49200 8 50000 128 6 wbs_dat_i[9]
port 268 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_o[0]
port 269 nsew signal bidirectional
rlabel metal3 s 49200 26528 50000 26648 6 wbs_dat_o[10]
port 270 nsew signal bidirectional
rlabel metal2 s 662 0 718 800 6 wbs_dat_o[11]
port 271 nsew signal bidirectional
rlabel metal3 s 49200 44888 50000 45008 6 wbs_dat_o[12]
port 272 nsew signal bidirectional
rlabel metal2 s 41234 51200 41290 52000 6 wbs_dat_o[13]
port 273 nsew signal bidirectional
rlabel metal3 s 49200 4088 50000 4208 6 wbs_dat_o[14]
port 274 nsew signal bidirectional
rlabel metal2 s 39302 51200 39358 52000 6 wbs_dat_o[15]
port 275 nsew signal bidirectional
rlabel metal3 s 0 19728 800 19848 6 wbs_dat_o[16]
port 276 nsew signal bidirectional
rlabel metal3 s 0 21768 800 21888 6 wbs_dat_o[17]
port 277 nsew signal bidirectional
rlabel metal2 s 32218 0 32274 800 6 wbs_dat_o[18]
port 278 nsew signal bidirectional
rlabel metal2 s 18 0 74 800 6 wbs_dat_o[19]
port 279 nsew signal bidirectional
rlabel metal2 s 38014 0 38070 800 6 wbs_dat_o[1]
port 280 nsew signal bidirectional
rlabel metal3 s 0 29248 800 29368 6 wbs_dat_o[20]
port 281 nsew signal bidirectional
rlabel metal3 s 0 4088 800 4208 6 wbs_dat_o[21]
port 282 nsew signal bidirectional
rlabel metal3 s 0 12928 800 13048 6 wbs_dat_o[22]
port 283 nsew signal bidirectional
rlabel metal3 s 0 21088 800 21208 6 wbs_dat_o[23]
port 284 nsew signal bidirectional
rlabel metal2 s 10322 0 10378 800 6 wbs_dat_o[24]
port 285 nsew signal bidirectional
rlabel metal2 s 3238 0 3294 800 6 wbs_dat_o[25]
port 286 nsew signal bidirectional
rlabel metal2 s 27710 51200 27766 52000 6 wbs_dat_o[26]
port 287 nsew signal bidirectional
rlabel metal2 s 16762 51200 16818 52000 6 wbs_dat_o[27]
port 288 nsew signal bidirectional
rlabel metal2 s 26422 0 26478 800 6 wbs_dat_o[28]
port 289 nsew signal bidirectional
rlabel metal2 s 36726 51200 36782 52000 6 wbs_dat_o[29]
port 290 nsew signal bidirectional
rlabel metal3 s 49200 12928 50000 13048 6 wbs_dat_o[2]
port 291 nsew signal bidirectional
rlabel metal3 s 0 36048 800 36168 6 wbs_dat_o[30]
port 292 nsew signal bidirectional
rlabel metal3 s 49200 39448 50000 39568 6 wbs_dat_o[31]
port 293 nsew signal bidirectional
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_o[3]
port 294 nsew signal bidirectional
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_o[4]
port 295 nsew signal bidirectional
rlabel metal3 s 0 6128 800 6248 6 wbs_dat_o[5]
port 296 nsew signal bidirectional
rlabel metal3 s 49200 37408 50000 37528 6 wbs_dat_o[6]
port 297 nsew signal bidirectional
rlabel metal2 s 29642 0 29698 800 6 wbs_dat_o[7]
port 298 nsew signal bidirectional
rlabel metal2 s 34150 51200 34206 52000 6 wbs_dat_o[8]
port 299 nsew signal bidirectional
rlabel metal2 s 33506 51200 33562 52000 6 wbs_dat_o[9]
port 300 nsew signal bidirectional
rlabel metal3 s 0 49648 800 49768 6 wbs_sel_i[0]
port 301 nsew signal input
rlabel metal2 s 5814 51200 5870 52000 6 wbs_sel_i[1]
port 302 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 wbs_sel_i[2]
port 303 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 wbs_sel_i[3]
port 304 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 wbs_stb_i
port 305 nsew signal input
rlabel metal3 s 49200 25168 50000 25288 6 wbs_we_i
port 306 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 50000 52000
<< end >>
