magic
tech sky130A
magscale 1 2
timestamp 1647555614
<< viali >>
rect 29009 49317 29043 49351
rect 14289 49249 14323 49283
rect 14565 49249 14599 49283
rect 17877 49249 17911 49283
rect 18153 49249 18187 49283
rect 22017 49249 22051 49283
rect 22569 49249 22603 49283
rect 24869 49249 24903 49283
rect 29745 49249 29779 49283
rect 30941 49249 30975 49283
rect 40693 49249 40727 49283
rect 42809 49249 42843 49283
rect 44465 49249 44499 49283
rect 46857 49249 46891 49283
rect 1869 49181 1903 49215
rect 4261 49181 4295 49215
rect 5089 49181 5123 49215
rect 6837 49181 6871 49215
rect 7665 49181 7699 49215
rect 10333 49181 10367 49215
rect 10977 49181 11011 49215
rect 11989 49181 12023 49215
rect 13277 49181 13311 49215
rect 16129 49181 16163 49215
rect 17141 49181 17175 49215
rect 17325 49181 17359 49215
rect 19441 49181 19475 49215
rect 20085 49181 20119 49215
rect 21005 49181 21039 49215
rect 24409 49181 24443 49215
rect 27445 49181 27479 49215
rect 27629 49181 27663 49215
rect 28273 49181 28307 49215
rect 28825 49181 28859 49215
rect 33609 49181 33643 49215
rect 35817 49181 35851 49215
rect 36461 49181 36495 49215
rect 38209 49181 38243 49215
rect 40969 49181 41003 49215
rect 42625 49181 42659 49215
rect 45201 49181 45235 49215
rect 47777 49181 47811 49215
rect 2789 49113 2823 49147
rect 2973 49113 3007 49147
rect 4629 49113 4663 49147
rect 19625 49113 19659 49147
rect 22201 49113 22235 49147
rect 24593 49113 24627 49147
rect 29929 49113 29963 49147
rect 45385 49113 45419 49147
rect 1961 49045 1995 49079
rect 5273 49045 5307 49079
rect 6929 49045 6963 49079
rect 8953 49045 8987 49079
rect 12081 49045 12115 49079
rect 13461 49045 13495 49079
rect 20269 49045 20303 49079
rect 32137 49045 32171 49079
rect 38301 49045 38335 49079
rect 47869 49045 47903 49079
rect 47869 48841 47903 48875
rect 22017 48773 22051 48807
rect 25973 48773 26007 48807
rect 47777 48773 47811 48807
rect 1409 48705 1443 48739
rect 4353 48705 4387 48739
rect 8953 48705 8987 48739
rect 11529 48705 11563 48739
rect 19257 48705 19291 48739
rect 27353 48705 27387 48739
rect 29653 48705 29687 48739
rect 32137 48705 32171 48739
rect 34897 48705 34931 48739
rect 2053 48637 2087 48671
rect 2237 48637 2271 48671
rect 2881 48637 2915 48671
rect 6377 48637 6411 48671
rect 6561 48637 6595 48671
rect 7205 48637 7239 48671
rect 9137 48637 9171 48671
rect 9689 48637 9723 48671
rect 11713 48637 11747 48671
rect 12449 48637 12483 48671
rect 14197 48637 14231 48671
rect 14381 48637 14415 48671
rect 15209 48637 15243 48671
rect 16957 48637 16991 48671
rect 17141 48637 17175 48671
rect 17417 48637 17451 48671
rect 19441 48637 19475 48671
rect 19717 48637 19751 48671
rect 22661 48637 22695 48671
rect 22845 48637 22879 48671
rect 23489 48637 23523 48671
rect 27537 48637 27571 48671
rect 28825 48637 28859 48671
rect 29837 48637 29871 48671
rect 30113 48637 30147 48671
rect 32321 48637 32355 48671
rect 33149 48637 33183 48671
rect 35081 48637 35115 48671
rect 36093 48637 36127 48671
rect 39129 48637 39163 48671
rect 39589 48637 39623 48671
rect 39773 48637 39807 48671
rect 40049 48637 40083 48671
rect 42441 48637 42475 48671
rect 42625 48637 42659 48671
rect 42901 48637 42935 48671
rect 45201 48637 45235 48671
rect 45385 48637 45419 48671
rect 45753 48637 45787 48671
rect 5273 48569 5307 48603
rect 25421 48569 25455 48603
rect 1501 48501 1535 48535
rect 4537 48501 4571 48535
rect 22109 48501 22143 48535
rect 26065 48501 26099 48535
rect 9413 48297 9447 48331
rect 14565 48297 14599 48331
rect 39957 48297 39991 48331
rect 7573 48229 7607 48263
rect 16129 48229 16163 48263
rect 19349 48229 19383 48263
rect 22661 48229 22695 48263
rect 24501 48229 24535 48263
rect 25237 48229 25271 48263
rect 28733 48229 28767 48263
rect 29837 48229 29871 48263
rect 41153 48229 41187 48263
rect 1593 48161 1627 48195
rect 3893 48161 3927 48195
rect 4905 48161 4939 48195
rect 10517 48161 10551 48195
rect 11069 48161 11103 48195
rect 16589 48161 16623 48195
rect 17417 48161 17451 48195
rect 20269 48161 20303 48195
rect 20729 48161 20763 48195
rect 27077 48161 27111 48195
rect 32229 48161 32263 48195
rect 35541 48161 35575 48195
rect 36737 48161 36771 48195
rect 43177 48161 43211 48195
rect 46765 48161 46799 48195
rect 1409 48093 1443 48127
rect 3801 48093 3835 48127
rect 4445 48093 4479 48127
rect 6929 48093 6963 48127
rect 9321 48093 9355 48127
rect 12909 48093 12943 48127
rect 14473 48093 14507 48127
rect 19257 48093 19291 48127
rect 22569 48093 22603 48127
rect 23397 48093 23431 48127
rect 24409 48093 24443 48127
rect 25881 48093 25915 48127
rect 26341 48093 26375 48127
rect 28641 48093 28675 48127
rect 29745 48093 29779 48127
rect 30389 48093 30423 48127
rect 31033 48093 31067 48127
rect 33333 48093 33367 48127
rect 34897 48093 34931 48127
rect 39865 48093 39899 48127
rect 41061 48093 41095 48127
rect 41797 48093 41831 48127
rect 42625 48093 42659 48127
rect 45017 48093 45051 48127
rect 46305 48093 46339 48127
rect 3249 48025 3283 48059
rect 4629 48025 4663 48059
rect 10701 48025 10735 48059
rect 13093 48025 13127 48059
rect 16773 48025 16807 48059
rect 20453 48025 20487 48059
rect 26525 48025 26559 48059
rect 30481 48025 30515 48059
rect 31217 48025 31251 48059
rect 34989 48025 35023 48059
rect 35725 48025 35759 48059
rect 42809 48025 42843 48059
rect 46489 48025 46523 48059
rect 33425 47957 33459 47991
rect 41889 47957 41923 47991
rect 45201 47957 45235 47991
rect 5365 47753 5399 47787
rect 6561 47753 6595 47787
rect 11621 47753 11655 47787
rect 12265 47753 12299 47787
rect 16037 47753 16071 47787
rect 19165 47753 19199 47787
rect 20177 47753 20211 47787
rect 27077 47753 27111 47787
rect 30113 47753 30147 47787
rect 32229 47753 32263 47787
rect 35909 47753 35943 47787
rect 41797 47753 41831 47787
rect 46305 47753 46339 47787
rect 2145 47685 2179 47719
rect 21925 47685 21959 47719
rect 33517 47685 33551 47719
rect 42717 47685 42751 47719
rect 43453 47685 43487 47719
rect 45109 47685 45143 47719
rect 47777 47685 47811 47719
rect 1961 47617 1995 47651
rect 4721 47617 4755 47651
rect 5273 47617 5307 47651
rect 6469 47617 6503 47651
rect 7113 47617 7147 47651
rect 11529 47617 11563 47651
rect 12173 47617 12207 47651
rect 14381 47617 14415 47651
rect 15945 47617 15979 47651
rect 16773 47617 16807 47651
rect 19073 47617 19107 47651
rect 20085 47617 20119 47651
rect 21833 47617 21867 47651
rect 22661 47617 22695 47651
rect 24133 47617 24167 47651
rect 26985 47617 27019 47651
rect 27721 47617 27755 47651
rect 30021 47617 30055 47651
rect 31309 47617 31343 47651
rect 32137 47617 32171 47651
rect 33333 47617 33367 47651
rect 35817 47617 35851 47651
rect 41705 47617 41739 47651
rect 42625 47617 42659 47651
rect 45569 47617 45603 47651
rect 46213 47617 46247 47651
rect 46857 47617 46891 47651
rect 3065 47549 3099 47583
rect 7297 47549 7331 47583
rect 7757 47549 7791 47583
rect 16957 47549 16991 47583
rect 17233 47549 17267 47583
rect 27905 47549 27939 47583
rect 28365 47549 28399 47583
rect 34713 47549 34747 47583
rect 43269 47549 43303 47583
rect 47961 47481 47995 47515
rect 23949 47413 23983 47447
rect 45661 47413 45695 47447
rect 46949 47413 46983 47447
rect 2513 47209 2547 47243
rect 3985 47209 4019 47243
rect 7665 47209 7699 47243
rect 16957 47209 16991 47243
rect 42349 47209 42383 47243
rect 43453 47209 43487 47243
rect 30665 47141 30699 47175
rect 44097 47141 44131 47175
rect 45201 47073 45235 47107
rect 45569 47073 45603 47107
rect 1409 47005 1443 47039
rect 2421 47005 2455 47039
rect 3249 47005 3283 47039
rect 7573 47005 7607 47039
rect 16865 47005 16899 47039
rect 19257 47005 19291 47039
rect 28089 47005 28123 47039
rect 28181 47005 28215 47039
rect 43913 47005 43947 47039
rect 45017 47005 45051 47039
rect 47961 47005 47995 47039
rect 20085 46937 20119 46971
rect 48145 46937 48179 46971
rect 1593 46869 1627 46903
rect 44649 46665 44683 46699
rect 47685 46665 47719 46699
rect 3801 46597 3835 46631
rect 18245 46597 18279 46631
rect 1961 46529 1995 46563
rect 17969 46529 18003 46563
rect 19073 46529 19107 46563
rect 42809 46529 42843 46563
rect 44097 46529 44131 46563
rect 44557 46529 44591 46563
rect 47041 46529 47075 46563
rect 47593 46529 47627 46563
rect 2145 46461 2179 46495
rect 20085 46461 20119 46495
rect 43453 46461 43487 46495
rect 45201 46461 45235 46495
rect 45385 46461 45419 46495
rect 2513 46121 2547 46155
rect 18613 46121 18647 46155
rect 44465 46121 44499 46155
rect 45201 46121 45235 46155
rect 46305 45985 46339 46019
rect 48145 45985 48179 46019
rect 1409 45917 1443 45951
rect 2421 45917 2455 45951
rect 3249 45917 3283 45951
rect 3985 45917 4019 45951
rect 13277 45917 13311 45951
rect 18429 45917 18463 45951
rect 19257 45917 19291 45951
rect 45109 45917 45143 45951
rect 20085 45849 20119 45883
rect 46489 45849 46523 45883
rect 1593 45781 1627 45815
rect 13369 45781 13403 45815
rect 13093 45509 13127 45543
rect 47685 45509 47719 45543
rect 2053 45441 2087 45475
rect 2697 45441 2731 45475
rect 18981 45441 19015 45475
rect 44833 45441 44867 45475
rect 45477 45441 45511 45475
rect 46397 45441 46431 45475
rect 46857 45441 46891 45475
rect 47593 45441 47627 45475
rect 2881 45373 2915 45407
rect 4077 45373 4111 45407
rect 12909 45373 12943 45407
rect 13829 45373 13863 45407
rect 19349 45373 19383 45407
rect 1593 45237 1627 45271
rect 2145 45237 2179 45271
rect 46949 45237 46983 45271
rect 3893 45033 3927 45067
rect 13185 45033 13219 45067
rect 1409 44897 1443 44931
rect 2789 44897 2823 44931
rect 46489 44897 46523 44931
rect 48145 44897 48179 44931
rect 3801 44829 3835 44863
rect 45201 44829 45235 44863
rect 45845 44829 45879 44863
rect 46305 44829 46339 44863
rect 1593 44761 1627 44795
rect 2053 44421 2087 44455
rect 45385 44421 45419 44455
rect 1869 44353 1903 44387
rect 45201 44353 45235 44387
rect 47777 44353 47811 44387
rect 2881 44285 2915 44319
rect 46857 44285 46891 44319
rect 2789 43945 2823 43979
rect 1869 43741 1903 43775
rect 2697 43741 2731 43775
rect 45845 43741 45879 43775
rect 46305 43741 46339 43775
rect 46489 43673 46523 43707
rect 48145 43673 48179 43707
rect 1961 43605 1995 43639
rect 46949 43401 46983 43435
rect 1869 43333 1903 43367
rect 46857 43265 46891 43299
rect 47869 43265 47903 43299
rect 2145 43061 2179 43095
rect 48053 43061 48087 43095
rect 47317 42721 47351 42755
rect 47225 42653 47259 42687
rect 47961 42585 47995 42619
rect 48053 42517 48087 42551
rect 46765 42177 46799 42211
rect 2053 41973 2087 42007
rect 46857 41973 46891 42007
rect 47777 41973 47811 42007
rect 1409 41633 1443 41667
rect 1869 41633 1903 41667
rect 46305 41633 46339 41667
rect 46489 41633 46523 41667
rect 1593 41497 1627 41531
rect 48145 41497 48179 41531
rect 2605 41225 2639 41259
rect 1869 41089 1903 41123
rect 2513 41089 2547 41123
rect 46489 41089 46523 41123
rect 46213 41021 46247 41055
rect 2053 40953 2087 40987
rect 47777 40885 47811 40919
rect 46305 40545 46339 40579
rect 1409 40477 1443 40511
rect 22661 40477 22695 40511
rect 22753 40477 22787 40511
rect 22845 40477 22879 40511
rect 23029 40477 23063 40511
rect 46489 40409 46523 40443
rect 48145 40409 48179 40443
rect 1593 40341 1627 40375
rect 22385 40341 22419 40375
rect 21189 40137 21223 40171
rect 23213 40137 23247 40171
rect 22100 40069 22134 40103
rect 21005 40001 21039 40035
rect 21281 40001 21315 40035
rect 23929 40001 23963 40035
rect 47593 40001 47627 40035
rect 47685 40001 47719 40035
rect 21833 39933 21867 39967
rect 23673 39933 23707 39967
rect 20821 39797 20855 39831
rect 25053 39797 25087 39831
rect 23121 39593 23155 39627
rect 20453 39457 20487 39491
rect 2237 39389 2271 39423
rect 17417 39389 17451 39423
rect 18337 39389 18371 39423
rect 23397 39389 23431 39423
rect 23486 39389 23520 39423
rect 23581 39389 23615 39423
rect 23765 39389 23799 39423
rect 24409 39389 24443 39423
rect 26893 39389 26927 39423
rect 47685 39389 47719 39423
rect 20720 39321 20754 39355
rect 24654 39321 24688 39355
rect 27138 39321 27172 39355
rect 17601 39253 17635 39287
rect 18429 39253 18463 39287
rect 21833 39253 21867 39287
rect 25789 39253 25823 39287
rect 28273 39253 28307 39287
rect 20453 39049 20487 39083
rect 22661 39049 22695 39083
rect 23213 39049 23247 39083
rect 26985 39049 27019 39083
rect 48053 39049 48087 39083
rect 2053 38913 2087 38947
rect 17233 38913 17267 38947
rect 18613 38913 18647 38947
rect 20729 38913 20763 38947
rect 20821 38913 20855 38947
rect 20913 38913 20947 38947
rect 21097 38913 21131 38947
rect 22477 38913 22511 38947
rect 22753 38913 22787 38947
rect 23469 38913 23503 38947
rect 23581 38913 23615 38947
rect 23673 38913 23707 38947
rect 23857 38913 23891 38947
rect 25053 38913 25087 38947
rect 25309 38913 25343 38947
rect 27261 38913 27295 38947
rect 27353 38913 27387 38947
rect 27445 38913 27479 38947
rect 27629 38913 27663 38947
rect 30389 38913 30423 38947
rect 30573 38913 30607 38947
rect 47961 38913 47995 38947
rect 2237 38845 2271 38879
rect 3065 38845 3099 38879
rect 18889 38845 18923 38879
rect 22293 38845 22327 38879
rect 17509 38709 17543 38743
rect 19993 38709 20027 38743
rect 26433 38709 26467 38743
rect 30757 38709 30791 38743
rect 2973 38505 3007 38539
rect 21833 38505 21867 38539
rect 22385 38505 22419 38539
rect 23305 38437 23339 38471
rect 24777 38437 24811 38471
rect 18153 38369 18187 38403
rect 19441 38369 19475 38403
rect 46305 38369 46339 38403
rect 48145 38369 48179 38403
rect 2881 38301 2915 38335
rect 15669 38301 15703 38335
rect 16313 38301 16347 38335
rect 19257 38301 19291 38335
rect 21097 38301 21131 38335
rect 22569 38301 22603 38335
rect 22753 38301 22787 38335
rect 22845 38301 22879 38335
rect 23489 38301 23523 38335
rect 23765 38301 23799 38335
rect 25053 38301 25087 38335
rect 25145 38301 25179 38335
rect 25237 38301 25271 38335
rect 25421 38301 25455 38335
rect 29561 38301 29595 38335
rect 31677 38301 31711 38335
rect 31766 38301 31800 38335
rect 31861 38301 31895 38335
rect 32045 38301 32079 38335
rect 15761 38233 15795 38267
rect 16497 38233 16531 38267
rect 21741 38233 21775 38267
rect 29806 38233 29840 38267
rect 31401 38233 31435 38267
rect 46489 38233 46523 38267
rect 23673 38165 23707 38199
rect 30941 38165 30975 38199
rect 19717 37893 19751 37927
rect 27905 37893 27939 37927
rect 30665 37893 30699 37927
rect 1869 37825 1903 37859
rect 8953 37825 8987 37859
rect 15669 37825 15703 37859
rect 17233 37825 17267 37859
rect 18613 37825 18647 37859
rect 20453 37825 20487 37859
rect 22089 37825 22123 37859
rect 22182 37825 22216 37859
rect 22293 37825 22327 37859
rect 22477 37825 22511 37859
rect 23029 37825 23063 37859
rect 23213 37825 23247 37859
rect 25421 37825 25455 37859
rect 25605 37825 25639 37859
rect 28181 37825 28215 37859
rect 28270 37825 28304 37859
rect 28365 37825 28399 37859
rect 28549 37825 28583 37859
rect 29377 37825 29411 37859
rect 30941 37825 30975 37859
rect 31033 37825 31067 37859
rect 31125 37825 31159 37859
rect 31309 37825 31343 37859
rect 32393 37825 32427 37859
rect 47869 37825 47903 37859
rect 15853 37757 15887 37791
rect 17417 37757 17451 37791
rect 20729 37757 20763 37791
rect 29469 37757 29503 37791
rect 29653 37757 29687 37791
rect 32137 37757 32171 37791
rect 2053 37689 2087 37723
rect 9045 37621 9079 37655
rect 21833 37621 21867 37655
rect 23397 37621 23431 37655
rect 25789 37621 25823 37655
rect 29009 37621 29043 37655
rect 33517 37621 33551 37655
rect 48053 37621 48087 37655
rect 23121 37417 23155 37451
rect 25053 37417 25087 37451
rect 29009 37417 29043 37451
rect 32873 37349 32907 37383
rect 1409 37281 1443 37315
rect 9137 37281 9171 37315
rect 9413 37281 9447 37315
rect 15577 37281 15611 37315
rect 23581 37281 23615 37315
rect 23765 37281 23799 37315
rect 30757 37281 30791 37315
rect 1685 37213 1719 37247
rect 8953 37213 8987 37247
rect 15117 37213 15151 37247
rect 17417 37213 17451 37247
rect 19257 37213 19291 37247
rect 21097 37213 21131 37247
rect 21364 37213 21398 37247
rect 24869 37213 24903 37247
rect 25973 37213 26007 37247
rect 26065 37213 26099 37247
rect 26157 37213 26191 37247
rect 26341 37213 26375 37247
rect 26801 37213 26835 37247
rect 28641 37213 28675 37247
rect 30665 37213 30699 37247
rect 31493 37213 31527 37247
rect 31749 37213 31783 37247
rect 47133 37213 47167 37247
rect 47961 37213 47995 37247
rect 15301 37145 15335 37179
rect 18245 37145 18279 37179
rect 20361 37145 20395 37179
rect 24685 37145 24719 37179
rect 25697 37145 25731 37179
rect 27046 37145 27080 37179
rect 28825 37145 28859 37179
rect 30573 37145 30607 37179
rect 22477 37077 22511 37111
rect 23489 37077 23523 37111
rect 28181 37077 28215 37111
rect 30205 37077 30239 37111
rect 47225 37077 47259 37111
rect 9597 36873 9631 36907
rect 15577 36873 15611 36907
rect 21833 36873 21867 36907
rect 24685 36873 24719 36907
rect 26249 36873 26283 36907
rect 29561 36873 29595 36907
rect 31125 36873 31159 36907
rect 13369 36805 13403 36839
rect 19349 36805 19383 36839
rect 30757 36805 30791 36839
rect 8217 36737 8251 36771
rect 8484 36737 8518 36771
rect 11529 36737 11563 36771
rect 14464 36737 14498 36771
rect 17233 36737 17267 36771
rect 18613 36737 18647 36771
rect 20729 36737 20763 36771
rect 22017 36737 22051 36771
rect 22201 36737 22235 36771
rect 22293 36737 22327 36771
rect 22753 36737 22787 36771
rect 23020 36737 23054 36771
rect 25053 36737 25087 36771
rect 25881 36737 25915 36771
rect 26065 36737 26099 36771
rect 27241 36737 27275 36771
rect 29929 36737 29963 36771
rect 30941 36737 30975 36771
rect 11713 36669 11747 36703
rect 14197 36669 14231 36703
rect 17417 36669 17451 36703
rect 20453 36669 20487 36703
rect 25145 36669 25179 36703
rect 25329 36669 25363 36703
rect 26985 36669 27019 36703
rect 30021 36669 30055 36703
rect 30205 36669 30239 36703
rect 2329 36533 2363 36567
rect 24133 36533 24167 36567
rect 28365 36533 28399 36567
rect 47777 36533 47811 36567
rect 11529 36329 11563 36363
rect 16497 36329 16531 36363
rect 18613 36329 18647 36363
rect 25145 36329 25179 36363
rect 26341 36329 26375 36363
rect 24685 36261 24719 36295
rect 20085 36193 20119 36227
rect 22661 36193 22695 36227
rect 25697 36193 25731 36227
rect 46305 36193 46339 36227
rect 46489 36193 46523 36227
rect 48145 36193 48179 36227
rect 2973 36125 3007 36159
rect 11437 36125 11471 36159
rect 15117 36125 15151 36159
rect 17233 36125 17267 36159
rect 17325 36125 17359 36159
rect 17417 36125 17451 36159
rect 17601 36125 17635 36159
rect 19257 36125 19291 36159
rect 22385 36125 22419 36159
rect 25513 36125 25547 36159
rect 25605 36125 25639 36159
rect 26571 36125 26605 36159
rect 26709 36125 26743 36159
rect 26801 36125 26835 36159
rect 26985 36125 27019 36159
rect 27721 36125 27755 36159
rect 31125 36125 31159 36159
rect 31217 36125 31251 36159
rect 31330 36125 31364 36159
rect 31493 36125 31527 36159
rect 15384 36057 15418 36091
rect 18337 36057 18371 36091
rect 20269 36057 20303 36091
rect 21925 36057 21959 36091
rect 24501 36057 24535 36091
rect 27537 36057 27571 36091
rect 3065 35989 3099 36023
rect 16957 35989 16991 36023
rect 19441 35989 19475 36023
rect 30849 35989 30883 36023
rect 9045 35785 9079 35819
rect 15209 35785 15243 35819
rect 18245 35785 18279 35819
rect 21925 35785 21959 35819
rect 22937 35785 22971 35819
rect 25053 35785 25087 35819
rect 28365 35785 28399 35819
rect 29101 35785 29135 35819
rect 30481 35785 30515 35819
rect 30849 35785 30883 35819
rect 2237 35717 2271 35751
rect 15945 35717 15979 35751
rect 17110 35717 17144 35751
rect 19993 35717 20027 35751
rect 29653 35717 29687 35751
rect 30021 35717 30055 35751
rect 32382 35717 32416 35751
rect 2053 35649 2087 35683
rect 9229 35649 9263 35683
rect 15117 35649 15151 35683
rect 15761 35649 15795 35683
rect 19257 35649 19291 35683
rect 20867 35649 20901 35683
rect 21005 35649 21039 35683
rect 21118 35649 21152 35683
rect 21281 35649 21315 35683
rect 21833 35649 21867 35683
rect 23167 35649 23201 35683
rect 23305 35649 23339 35683
rect 23397 35649 23431 35683
rect 23581 35649 23615 35683
rect 24041 35649 24075 35683
rect 24317 35649 24351 35683
rect 25421 35649 25455 35683
rect 26249 35649 26283 35683
rect 26341 35649 26375 35683
rect 28273 35649 28307 35683
rect 29009 35649 29043 35683
rect 29837 35649 29871 35683
rect 46857 35649 46891 35683
rect 47869 35649 47903 35683
rect 2789 35581 2823 35615
rect 16865 35581 16899 35615
rect 24225 35581 24259 35615
rect 25513 35581 25547 35615
rect 25697 35581 25731 35615
rect 30941 35581 30975 35615
rect 31033 35581 31067 35615
rect 32137 35581 32171 35615
rect 16129 35445 16163 35479
rect 20637 35445 20671 35479
rect 24041 35445 24075 35479
rect 24501 35445 24535 35479
rect 33517 35445 33551 35479
rect 46949 35445 46983 35479
rect 48053 35445 48087 35479
rect 1961 35241 1995 35275
rect 15853 35241 15887 35275
rect 17509 35241 17543 35275
rect 27629 35173 27663 35207
rect 28089 35173 28123 35207
rect 29009 35173 29043 35207
rect 31217 35173 31251 35207
rect 18337 35105 18371 35139
rect 20085 35105 20119 35139
rect 22569 35105 22603 35139
rect 30389 35105 30423 35139
rect 12173 35037 12207 35071
rect 16129 35037 16163 35071
rect 16221 35037 16255 35071
rect 16313 35037 16347 35071
rect 16497 35037 16531 35071
rect 17141 35037 17175 35071
rect 17325 35037 17359 35071
rect 18061 35037 18095 35071
rect 19257 35037 19291 35071
rect 20352 35037 20386 35071
rect 22017 35037 22051 35071
rect 23397 35037 23431 35071
rect 26617 35037 26651 35071
rect 28273 35037 28307 35071
rect 28825 35037 28859 35071
rect 31861 35037 31895 35071
rect 31953 35037 31987 35071
rect 32045 35037 32079 35071
rect 32229 35037 32263 35071
rect 32781 35037 32815 35071
rect 45845 35037 45879 35071
rect 46305 35037 46339 35071
rect 1869 34969 1903 35003
rect 12418 34969 12452 35003
rect 24869 34969 24903 35003
rect 25053 34969 25087 35003
rect 25605 34969 25639 35003
rect 27261 34969 27295 35003
rect 27445 34969 27479 35003
rect 30297 34969 30331 35003
rect 31585 34969 31619 35003
rect 33048 34969 33082 35003
rect 46489 34969 46523 35003
rect 48145 34969 48179 35003
rect 13553 34901 13587 34935
rect 19441 34901 19475 34935
rect 21465 34901 21499 34935
rect 23213 34901 23247 34935
rect 25697 34901 25731 34935
rect 26709 34901 26743 34935
rect 29837 34901 29871 34935
rect 30205 34901 30239 34935
rect 34161 34901 34195 34935
rect 12173 34697 12207 34731
rect 14749 34697 14783 34731
rect 21833 34697 21867 34731
rect 27445 34697 27479 34731
rect 27813 34697 27847 34731
rect 47685 34697 47719 34731
rect 15853 34629 15887 34663
rect 18153 34629 18187 34663
rect 27905 34629 27939 34663
rect 29469 34629 29503 34663
rect 30389 34629 30423 34663
rect 30573 34629 30607 34663
rect 2053 34561 2087 34595
rect 12449 34561 12483 34595
rect 12541 34561 12575 34595
rect 12633 34561 12667 34595
rect 12817 34561 12851 34595
rect 13645 34561 13679 34595
rect 13829 34561 13863 34595
rect 14473 34561 14507 34595
rect 14657 34561 14691 34595
rect 16911 34561 16945 34595
rect 17046 34561 17080 34595
rect 17141 34561 17175 34595
rect 17325 34561 17359 34595
rect 17969 34561 18003 34595
rect 19441 34561 19475 34595
rect 20821 34561 20855 34595
rect 21189 34561 21223 34595
rect 22017 34561 22051 34595
rect 22201 34561 22235 34595
rect 22293 34561 22327 34595
rect 23397 34561 23431 34595
rect 24225 34561 24259 34595
rect 24409 34561 24443 34595
rect 25053 34561 25087 34595
rect 25145 34561 25179 34595
rect 25973 34561 26007 34595
rect 26249 34561 26283 34595
rect 29745 34561 29779 34595
rect 45201 34561 45235 34595
rect 47593 34561 47627 34595
rect 2697 34493 2731 34527
rect 13737 34493 13771 34527
rect 16037 34493 16071 34527
rect 20085 34493 20119 34527
rect 23489 34493 23523 34527
rect 23673 34493 23707 34527
rect 26157 34493 26191 34527
rect 28089 34493 28123 34527
rect 29653 34493 29687 34527
rect 45385 34493 45419 34527
rect 46857 34493 46891 34527
rect 24593 34425 24627 34459
rect 1593 34357 1627 34391
rect 2145 34357 2179 34391
rect 16681 34357 16715 34391
rect 23029 34357 23063 34391
rect 24317 34357 24351 34391
rect 25053 34357 25087 34391
rect 25421 34357 25455 34391
rect 26157 34357 26191 34391
rect 26433 34357 26467 34391
rect 29469 34357 29503 34391
rect 29929 34357 29963 34391
rect 30757 34357 30791 34391
rect 14105 34153 14139 34187
rect 14565 34153 14599 34187
rect 24777 34153 24811 34187
rect 25053 34153 25087 34187
rect 26617 34153 26651 34187
rect 27077 34085 27111 34119
rect 1409 34017 1443 34051
rect 1593 34017 1627 34051
rect 2789 34017 2823 34051
rect 9597 34017 9631 34051
rect 10333 34017 10367 34051
rect 12725 34017 12759 34051
rect 13001 34017 13035 34051
rect 14197 34017 14231 34051
rect 15485 34017 15519 34051
rect 17049 34017 17083 34051
rect 17325 34017 17359 34051
rect 19441 34017 19475 34051
rect 25973 34017 26007 34051
rect 26801 34017 26835 34051
rect 28457 34017 28491 34051
rect 30205 34017 30239 34051
rect 35817 34017 35851 34051
rect 37657 34017 37691 34051
rect 46305 34017 46339 34051
rect 46489 34017 46523 34051
rect 48145 34017 48179 34051
rect 9505 33949 9539 33983
rect 14105 33949 14139 33983
rect 14381 33949 14415 33983
rect 15209 33949 15243 33983
rect 19717 33949 19751 33983
rect 22753 33949 22787 33983
rect 24777 33949 24811 33983
rect 24869 33949 24903 33983
rect 25513 33949 25547 33983
rect 25881 33949 25915 33983
rect 26617 33949 26651 33983
rect 26893 33949 26927 33983
rect 28273 33949 28307 33983
rect 30757 33949 30791 33983
rect 10578 33881 10612 33915
rect 22937 33881 22971 33915
rect 24593 33881 24627 33915
rect 28365 33881 28399 33915
rect 30021 33881 30055 33915
rect 36001 33881 36035 33915
rect 9873 33813 9907 33847
rect 11713 33813 11747 33847
rect 18613 33813 18647 33847
rect 23121 33813 23155 33847
rect 25605 33813 25639 33847
rect 27905 33813 27939 33847
rect 30849 33813 30883 33847
rect 10333 33609 10367 33643
rect 11989 33609 12023 33643
rect 13001 33609 13035 33643
rect 17509 33609 17543 33643
rect 29745 33609 29779 33643
rect 33885 33609 33919 33643
rect 35909 33609 35943 33643
rect 46949 33609 46983 33643
rect 11897 33541 11931 33575
rect 18981 33541 19015 33575
rect 22201 33541 22235 33575
rect 26249 33541 26283 33575
rect 27537 33541 27571 33575
rect 1869 33473 1903 33507
rect 8401 33473 8435 33507
rect 8668 33473 8702 33507
rect 10563 33473 10597 33507
rect 10701 33473 10735 33507
rect 10798 33473 10832 33507
rect 10977 33473 11011 33507
rect 11805 33473 11839 33507
rect 12725 33473 12759 33507
rect 13645 33473 13679 33507
rect 14289 33473 14323 33507
rect 14556 33473 14590 33507
rect 17141 33473 17175 33507
rect 17325 33473 17359 33507
rect 19165 33473 19199 33507
rect 19901 33473 19935 33507
rect 20168 33473 20202 33507
rect 22017 33473 22051 33507
rect 22293 33473 22327 33507
rect 23673 33473 23707 33507
rect 27721 33473 27755 33507
rect 28365 33473 28399 33507
rect 28621 33473 28655 33507
rect 30665 33473 30699 33507
rect 30757 33473 30791 33507
rect 30849 33473 30883 33507
rect 31033 33473 31067 33507
rect 32772 33473 32806 33507
rect 35817 33473 35851 33507
rect 46857 33473 46891 33507
rect 47961 33473 47995 33507
rect 2053 33405 2087 33439
rect 2789 33405 2823 33439
rect 12173 33405 12207 33439
rect 12265 33405 12299 33439
rect 13001 33405 13035 33439
rect 13461 33405 13495 33439
rect 32505 33405 32539 33439
rect 11529 33337 11563 33371
rect 21281 33337 21315 33371
rect 23857 33337 23891 33371
rect 26433 33337 26467 33371
rect 27905 33337 27939 33371
rect 9781 33269 9815 33303
rect 12817 33269 12851 33303
rect 13829 33269 13863 33303
rect 15669 33269 15703 33303
rect 21833 33269 21867 33303
rect 30389 33269 30423 33303
rect 48053 33269 48087 33303
rect 2789 33065 2823 33099
rect 10333 33065 10367 33099
rect 11253 33065 11287 33099
rect 13461 33065 13495 33099
rect 20453 33065 20487 33099
rect 27813 33065 27847 33099
rect 33057 33065 33091 33099
rect 47685 33065 47719 33099
rect 26249 32997 26283 33031
rect 12265 32929 12299 32963
rect 27169 32929 27203 32963
rect 30297 32929 30331 32963
rect 31217 32929 31251 32963
rect 2237 32861 2271 32895
rect 2697 32861 2731 32895
rect 10241 32861 10275 32895
rect 10425 32861 10459 32895
rect 10885 32861 10919 32895
rect 11989 32861 12023 32895
rect 14473 32861 14507 32895
rect 14933 32861 14967 32895
rect 18521 32861 18555 32895
rect 19257 32861 19291 32895
rect 20709 32861 20743 32895
rect 20802 32861 20836 32895
rect 20913 32858 20947 32892
rect 21097 32861 21131 32895
rect 22201 32861 22235 32895
rect 26433 32861 26467 32895
rect 28043 32861 28077 32895
rect 28181 32861 28215 32895
rect 28278 32861 28312 32895
rect 28457 32861 28491 32895
rect 30113 32861 30147 32895
rect 31473 32861 31507 32895
rect 33333 32861 33367 32895
rect 33425 32861 33459 32895
rect 33517 32861 33551 32895
rect 33701 32861 33735 32895
rect 11069 32793 11103 32827
rect 13369 32793 13403 32827
rect 22446 32793 22480 32827
rect 26985 32793 27019 32827
rect 15301 32725 15335 32759
rect 18613 32725 18647 32759
rect 19349 32725 19383 32759
rect 23581 32725 23615 32759
rect 29745 32725 29779 32759
rect 30205 32725 30239 32759
rect 32597 32725 32631 32759
rect 13185 32521 13219 32555
rect 14473 32521 14507 32555
rect 18981 32521 19015 32555
rect 23397 32521 23431 32555
rect 25421 32521 25455 32555
rect 27997 32521 28031 32555
rect 31309 32521 31343 32555
rect 18889 32453 18923 32487
rect 25513 32453 25547 32487
rect 27169 32453 27203 32487
rect 30941 32453 30975 32487
rect 2053 32385 2087 32419
rect 10379 32385 10413 32419
rect 10517 32385 10551 32419
rect 10614 32385 10648 32419
rect 10793 32385 10827 32419
rect 12081 32385 12115 32419
rect 12265 32385 12299 32419
rect 13093 32385 13127 32419
rect 13277 32385 13311 32419
rect 13737 32385 13771 32419
rect 13925 32385 13959 32419
rect 14013 32385 14047 32419
rect 14289 32385 14323 32419
rect 14933 32385 14967 32419
rect 15117 32385 15151 32419
rect 16957 32385 16991 32419
rect 17224 32385 17258 32419
rect 19901 32385 19935 32419
rect 22017 32385 22051 32419
rect 22284 32385 22318 32419
rect 24225 32385 24259 32419
rect 27353 32385 27387 32419
rect 28365 32385 28399 32419
rect 30113 32385 30147 32419
rect 31125 32385 31159 32419
rect 32689 32385 32723 32419
rect 32945 32385 32979 32419
rect 47685 32385 47719 32419
rect 2237 32317 2271 32351
rect 2881 32317 2915 32351
rect 14105 32317 14139 32351
rect 24317 32317 24351 32351
rect 24501 32317 24535 32351
rect 25605 32317 25639 32351
rect 28457 32317 28491 32351
rect 28641 32317 28675 32351
rect 30205 32317 30239 32351
rect 30297 32317 30331 32351
rect 47869 32317 47903 32351
rect 10149 32181 10183 32215
rect 12173 32181 12207 32215
rect 15301 32181 15335 32215
rect 18337 32181 18371 32215
rect 20085 32181 20119 32215
rect 23857 32181 23891 32215
rect 25053 32181 25087 32215
rect 27537 32181 27571 32215
rect 29745 32181 29779 32215
rect 34069 32181 34103 32215
rect 2973 31977 3007 32011
rect 9689 31977 9723 32011
rect 15853 31977 15887 32011
rect 22017 31977 22051 32011
rect 23121 31977 23155 32011
rect 26801 31977 26835 32011
rect 30021 31977 30055 32011
rect 31309 31977 31343 32011
rect 31769 31977 31803 32011
rect 11529 31909 11563 31943
rect 18337 31909 18371 31943
rect 30481 31909 30515 31943
rect 32965 31909 32999 31943
rect 12265 31841 12299 31875
rect 13461 31841 13495 31875
rect 16957 31841 16991 31875
rect 19257 31841 19291 31875
rect 19441 31841 19475 31875
rect 30205 31841 30239 31875
rect 33517 31841 33551 31875
rect 37841 31841 37875 31875
rect 1869 31773 1903 31807
rect 2053 31773 2087 31807
rect 2881 31773 2915 31807
rect 9689 31773 9723 31807
rect 9873 31773 9907 31807
rect 10609 31773 10643 31807
rect 10698 31767 10732 31801
rect 10793 31773 10827 31807
rect 10977 31773 11011 31807
rect 11805 31773 11839 31807
rect 12541 31773 12575 31807
rect 12633 31773 12667 31807
rect 12725 31773 12759 31807
rect 12909 31773 12943 31807
rect 13369 31773 13403 31807
rect 13553 31773 13587 31807
rect 16129 31773 16163 31807
rect 16221 31773 16255 31807
rect 16313 31773 16347 31807
rect 16497 31773 16531 31807
rect 21097 31773 21131 31807
rect 22293 31773 22327 31807
rect 22385 31773 22419 31807
rect 22477 31773 22511 31807
rect 22661 31773 22695 31807
rect 23397 31773 23431 31807
rect 23489 31773 23523 31807
rect 23581 31773 23615 31807
rect 23765 31773 23799 31807
rect 24501 31773 24535 31807
rect 25421 31773 25455 31807
rect 28273 31773 28307 31807
rect 28365 31773 28399 31807
rect 28457 31773 28491 31807
rect 28641 31773 28675 31807
rect 30021 31773 30055 31807
rect 30297 31773 30331 31807
rect 30941 31773 30975 31807
rect 31125 31773 31159 31807
rect 31999 31773 32033 31807
rect 32137 31773 32171 31807
rect 32234 31773 32268 31807
rect 32413 31773 32447 31807
rect 33425 31773 33459 31807
rect 36001 31773 36035 31807
rect 47961 31773 47995 31807
rect 11529 31705 11563 31739
rect 17202 31705 17236 31739
rect 24685 31705 24719 31739
rect 25666 31705 25700 31739
rect 36185 31705 36219 31739
rect 10333 31637 10367 31671
rect 11713 31637 11747 31671
rect 24869 31637 24903 31671
rect 27997 31637 28031 31671
rect 33333 31637 33367 31671
rect 48053 31637 48087 31671
rect 13461 31433 13495 31467
rect 14473 31433 14507 31467
rect 23489 31433 23523 31467
rect 25329 31433 25363 31467
rect 28089 31433 28123 31467
rect 30849 31433 30883 31467
rect 36093 31433 36127 31467
rect 9220 31365 9254 31399
rect 10885 31365 10919 31399
rect 16681 31365 16715 31399
rect 17785 31365 17819 31399
rect 17969 31365 18003 31399
rect 18889 31365 18923 31399
rect 23121 31365 23155 31399
rect 24593 31365 24627 31399
rect 28733 31365 28767 31399
rect 29653 31365 29687 31399
rect 7113 31297 7147 31331
rect 7380 31297 7414 31331
rect 10793 31297 10827 31331
rect 10977 31297 11011 31331
rect 11989 31297 12023 31331
rect 12173 31297 12207 31331
rect 13369 31297 13403 31331
rect 14013 31297 14047 31331
rect 14289 31297 14323 31331
rect 14933 31297 14967 31331
rect 15117 31297 15151 31331
rect 15209 31297 15243 31331
rect 16911 31297 16945 31331
rect 17049 31297 17083 31331
rect 17141 31297 17175 31331
rect 17325 31297 17359 31331
rect 21097 31297 21131 31331
rect 21833 31297 21867 31331
rect 23305 31297 23339 31331
rect 24501 31297 24535 31331
rect 25585 31297 25619 31331
rect 25678 31297 25712 31331
rect 25794 31297 25828 31331
rect 25973 31297 26007 31331
rect 27997 31297 28031 31331
rect 29469 31297 29503 31331
rect 30481 31297 30515 31331
rect 30665 31297 30699 31331
rect 32137 31297 32171 31331
rect 32321 31297 32355 31331
rect 36001 31297 36035 31331
rect 1961 31229 1995 31263
rect 2145 31229 2179 31263
rect 3065 31229 3099 31263
rect 8953 31229 8987 31263
rect 14105 31229 14139 31263
rect 18153 31229 18187 31263
rect 18705 31229 18739 31263
rect 20545 31229 20579 31263
rect 22109 31229 22143 31263
rect 24777 31229 24811 31263
rect 14933 31161 14967 31195
rect 8493 31093 8527 31127
rect 10333 31093 10367 31127
rect 12357 31093 12391 31127
rect 14289 31093 14323 31127
rect 21189 31093 21223 31127
rect 24133 31093 24167 31127
rect 28825 31093 28859 31127
rect 32505 31093 32539 31127
rect 2237 30889 2271 30923
rect 2881 30889 2915 30923
rect 10425 30889 10459 30923
rect 10609 30889 10643 30923
rect 13001 30889 13035 30923
rect 14289 30889 14323 30923
rect 16497 30889 16531 30923
rect 26801 30889 26835 30923
rect 30481 30889 30515 30923
rect 36093 30889 36127 30923
rect 15301 30821 15335 30855
rect 17509 30821 17543 30855
rect 18245 30753 18279 30787
rect 21189 30753 21223 30787
rect 22937 30753 22971 30787
rect 2789 30685 2823 30719
rect 11069 30685 11103 30719
rect 11345 30685 11379 30719
rect 12633 30685 12667 30719
rect 12817 30685 12851 30719
rect 13093 30685 13127 30719
rect 14197 30685 14231 30719
rect 15117 30685 15151 30719
rect 16681 30685 16715 30719
rect 17141 30685 17175 30719
rect 18061 30685 18095 30719
rect 19717 30685 19751 30719
rect 20913 30685 20947 30719
rect 22661 30685 22695 30719
rect 24409 30685 24443 30719
rect 25421 30685 25455 30719
rect 27537 30685 27571 30719
rect 28273 30685 28307 30719
rect 31125 30685 31159 30719
rect 31217 30685 31251 30719
rect 31309 30685 31343 30719
rect 31493 30685 31527 30719
rect 31953 30685 31987 30719
rect 34713 30685 34747 30719
rect 10241 30617 10275 30651
rect 12725 30617 12759 30651
rect 17325 30617 17359 30651
rect 24593 30617 24627 30651
rect 25666 30617 25700 30651
rect 30849 30617 30883 30651
rect 32198 30617 32232 30651
rect 34958 30617 34992 30651
rect 10451 30549 10485 30583
rect 12357 30549 12391 30583
rect 19809 30549 19843 30583
rect 24777 30549 24811 30583
rect 27629 30549 27663 30583
rect 28365 30549 28399 30583
rect 33333 30549 33367 30583
rect 11805 30345 11839 30379
rect 13369 30345 13403 30379
rect 14381 30345 14415 30379
rect 21189 30345 21223 30379
rect 24869 30345 24903 30379
rect 32137 30345 32171 30379
rect 10609 30277 10643 30311
rect 11621 30277 11655 30311
rect 12173 30277 12207 30311
rect 13277 30277 13311 30311
rect 26065 30277 26099 30311
rect 28794 30277 28828 30311
rect 30481 30277 30515 30311
rect 32597 30277 32631 30311
rect 34897 30277 34931 30311
rect 10517 30209 10551 30243
rect 10701 30209 10735 30243
rect 11897 30209 11931 30243
rect 11989 30209 12023 30243
rect 14381 30209 14415 30243
rect 15209 30209 15243 30243
rect 17417 30209 17451 30243
rect 19717 30209 19751 30243
rect 19901 30209 19935 30243
rect 20269 30209 20303 30243
rect 21005 30209 21039 30243
rect 21833 30209 21867 30243
rect 22937 30209 22971 30243
rect 23949 30209 23983 30243
rect 24041 30209 24075 30243
rect 24133 30209 24167 30243
rect 24317 30209 24351 30243
rect 25145 30209 25179 30243
rect 25237 30209 25271 30243
rect 25329 30209 25363 30243
rect 25513 30209 25547 30243
rect 27721 30209 27755 30243
rect 27826 30209 27860 30243
rect 27926 30215 27960 30249
rect 28089 30209 28123 30243
rect 32505 30209 32539 30243
rect 33885 30209 33919 30243
rect 33977 30209 34011 30243
rect 34069 30209 34103 30243
rect 34253 30209 34287 30243
rect 35081 30209 35115 30243
rect 1961 30141 1995 30175
rect 2145 30141 2179 30175
rect 2881 30141 2915 30175
rect 14197 30141 14231 30175
rect 14749 30141 14783 30175
rect 17141 30141 17175 30175
rect 19993 30141 20027 30175
rect 20085 30141 20119 30175
rect 26249 30141 26283 30175
rect 28549 30141 28583 30175
rect 32781 30141 32815 30175
rect 35265 30141 35299 30175
rect 22017 30073 22051 30107
rect 29929 30073 29963 30107
rect 15301 30005 15335 30039
rect 20453 30005 20487 30039
rect 23121 30005 23155 30039
rect 23673 30005 23707 30039
rect 27445 30005 27479 30039
rect 30573 30005 30607 30039
rect 33609 30005 33643 30039
rect 2237 29801 2271 29835
rect 2881 29801 2915 29835
rect 15301 29801 15335 29835
rect 15853 29801 15887 29835
rect 19349 29801 19383 29835
rect 21557 29801 21591 29835
rect 22661 29801 22695 29835
rect 23397 29801 23431 29835
rect 25789 29801 25823 29835
rect 26893 29801 26927 29835
rect 27813 29801 27847 29835
rect 8401 29665 8435 29699
rect 13001 29665 13035 29699
rect 14657 29665 14691 29699
rect 17417 29665 17451 29699
rect 20453 29665 20487 29699
rect 30021 29665 30055 29699
rect 30205 29665 30239 29699
rect 47593 29665 47627 29699
rect 2789 29597 2823 29631
rect 8033 29597 8067 29631
rect 10885 29597 10919 29631
rect 12725 29597 12759 29631
rect 14933 29597 14967 29631
rect 15025 29597 15059 29631
rect 15393 29597 15427 29631
rect 16037 29597 16071 29631
rect 16129 29597 16163 29631
rect 17141 29597 17175 29631
rect 17233 29597 17267 29631
rect 18153 29597 18187 29631
rect 18245 29597 18279 29631
rect 18337 29597 18371 29631
rect 18521 29597 18555 29631
rect 19257 29597 19291 29631
rect 20177 29597 20211 29631
rect 22385 29597 22419 29631
rect 22477 29597 22511 29631
rect 23581 29597 23615 29631
rect 23857 29597 23891 29631
rect 24409 29597 24443 29631
rect 27629 29597 27663 29631
rect 28825 29597 28859 29631
rect 31861 29597 31895 29631
rect 31953 29597 31987 29631
rect 32045 29597 32079 29631
rect 32229 29597 32263 29631
rect 35061 29597 35095 29631
rect 35173 29597 35207 29631
rect 35265 29597 35299 29631
rect 35443 29597 35477 29631
rect 47317 29597 47351 29631
rect 8217 29529 8251 29563
rect 8953 29529 8987 29563
rect 9137 29529 9171 29563
rect 11152 29529 11186 29563
rect 15853 29529 15887 29563
rect 24654 29529 24688 29563
rect 26801 29529 26835 29563
rect 27445 29529 27479 29563
rect 29009 29529 29043 29563
rect 9321 29461 9355 29495
rect 12265 29461 12299 29495
rect 15117 29461 15151 29495
rect 17417 29461 17451 29495
rect 17877 29461 17911 29495
rect 23765 29461 23799 29495
rect 29561 29461 29595 29495
rect 29929 29461 29963 29495
rect 31585 29461 31619 29495
rect 34805 29461 34839 29495
rect 17233 29257 17267 29291
rect 20453 29257 20487 29291
rect 23213 29257 23247 29291
rect 25789 29257 25823 29291
rect 29561 29257 29595 29291
rect 31309 29257 31343 29291
rect 33149 29257 33183 29291
rect 34713 29257 34747 29291
rect 36553 29257 36587 29291
rect 15853 29189 15887 29223
rect 18674 29189 18708 29223
rect 23949 29189 23983 29223
rect 27537 29189 27571 29223
rect 31217 29189 31251 29223
rect 34345 29189 34379 29223
rect 35418 29189 35452 29223
rect 7205 29121 7239 29155
rect 7472 29121 7506 29155
rect 9275 29121 9309 29155
rect 9413 29121 9447 29155
rect 9505 29121 9539 29155
rect 9689 29121 9723 29155
rect 12541 29121 12575 29155
rect 13001 29121 13035 29155
rect 13185 29121 13219 29155
rect 13829 29121 13863 29155
rect 14096 29121 14130 29155
rect 15669 29121 15703 29155
rect 15945 29121 15979 29155
rect 17693 29121 17727 29155
rect 20361 29121 20395 29155
rect 20545 29121 20579 29155
rect 21833 29121 21867 29155
rect 22109 29121 22143 29155
rect 23397 29121 23431 29155
rect 24133 29121 24167 29155
rect 25605 29121 25639 29155
rect 28437 29121 28471 29155
rect 33057 29121 33091 29155
rect 34529 29121 34563 29155
rect 35173 29121 35207 29155
rect 46305 29121 46339 29155
rect 47593 29121 47627 29155
rect 9045 29053 9079 29087
rect 17417 29053 17451 29087
rect 18429 29053 18463 29087
rect 22201 29053 22235 29087
rect 28181 29053 28215 29087
rect 31401 29053 31435 29087
rect 33333 29053 33367 29087
rect 8585 28985 8619 29019
rect 12357 28985 12391 29019
rect 15669 28985 15703 29019
rect 17601 28985 17635 29019
rect 19809 28985 19843 29019
rect 27721 28985 27755 29019
rect 32689 28985 32723 29019
rect 47685 28985 47719 29019
rect 2053 28917 2087 28951
rect 13093 28917 13127 28951
rect 15209 28917 15243 28951
rect 30849 28917 30883 28951
rect 46397 28917 46431 28951
rect 14197 28713 14231 28747
rect 31401 28713 31435 28747
rect 33241 28713 33275 28747
rect 18705 28645 18739 28679
rect 20177 28645 20211 28679
rect 1409 28577 1443 28611
rect 2789 28577 2823 28611
rect 7021 28577 7055 28611
rect 27077 28577 27111 28611
rect 34713 28577 34747 28611
rect 36645 28577 36679 28611
rect 46305 28577 46339 28611
rect 46489 28577 46523 28611
rect 48145 28577 48179 28611
rect 9229 28509 9263 28543
rect 9318 28509 9352 28543
rect 9413 28509 9447 28543
rect 9597 28509 9631 28543
rect 10149 28509 10183 28543
rect 14381 28509 14415 28543
rect 14657 28509 14691 28543
rect 15761 28509 15795 28543
rect 16037 28509 16071 28543
rect 16497 28509 16531 28543
rect 20361 28509 20395 28543
rect 20453 28509 20487 28543
rect 23029 28509 23063 28543
rect 25697 28509 25731 28543
rect 26985 28509 27019 28543
rect 27997 28509 28031 28543
rect 28089 28509 28123 28543
rect 28181 28509 28215 28543
rect 28365 28509 28399 28543
rect 30389 28509 30423 28543
rect 30573 28509 30607 28543
rect 31861 28509 31895 28543
rect 33701 28509 33735 28543
rect 34989 28509 35023 28543
rect 36001 28509 36035 28543
rect 1593 28441 1627 28475
rect 7288 28441 7322 28475
rect 8953 28441 8987 28475
rect 14565 28441 14599 28475
rect 15577 28441 15611 28475
rect 16742 28441 16776 28475
rect 18337 28441 18371 28475
rect 18521 28441 18555 28475
rect 20177 28441 20211 28475
rect 25881 28441 25915 28475
rect 26893 28441 26927 28475
rect 31033 28441 31067 28475
rect 31217 28441 31251 28475
rect 32106 28441 32140 28475
rect 33885 28441 33919 28475
rect 36093 28441 36127 28475
rect 36829 28441 36863 28475
rect 38485 28441 38519 28475
rect 8401 28373 8435 28407
rect 10241 28373 10275 28407
rect 15945 28373 15979 28407
rect 17877 28373 17911 28407
rect 23121 28373 23155 28407
rect 26065 28373 26099 28407
rect 26525 28373 26559 28407
rect 27721 28373 27755 28407
rect 34069 28373 34103 28407
rect 2145 28169 2179 28203
rect 12541 28169 12575 28203
rect 16773 28169 16807 28203
rect 17509 28169 17543 28203
rect 48053 28169 48087 28203
rect 9413 28101 9447 28135
rect 18429 28101 18463 28135
rect 20168 28101 20202 28135
rect 23213 28101 23247 28135
rect 27252 28101 27286 28135
rect 2053 28033 2087 28067
rect 9589 28023 9623 28057
rect 9681 28033 9715 28067
rect 9873 28033 9907 28067
rect 9965 28033 9999 28067
rect 11713 28033 11747 28067
rect 12725 28033 12759 28067
rect 13001 28033 13035 28067
rect 15577 28033 15611 28067
rect 16681 28033 16715 28067
rect 17325 28033 17359 28067
rect 18613 28033 18647 28067
rect 19901 28033 19935 28067
rect 26065 28033 26099 28067
rect 26154 28033 26188 28067
rect 26254 28033 26288 28067
rect 26433 28033 26467 28067
rect 29377 28033 29411 28067
rect 29466 28033 29500 28067
rect 29561 28033 29595 28067
rect 29745 28033 29779 28067
rect 32853 28033 32887 28067
rect 35265 28033 35299 28067
rect 35357 28033 35391 28067
rect 35449 28033 35483 28067
rect 35633 28033 35667 28067
rect 47869 28033 47903 28067
rect 11621 27965 11655 27999
rect 15301 27965 15335 27999
rect 17693 27965 17727 27999
rect 23029 27965 23063 27999
rect 23489 27965 23523 27999
rect 26985 27965 27019 27999
rect 32597 27965 32631 27999
rect 12081 27897 12115 27931
rect 12817 27897 12851 27931
rect 12909 27897 12943 27931
rect 33977 27897 34011 27931
rect 17693 27829 17727 27863
rect 21281 27829 21315 27863
rect 25789 27829 25823 27863
rect 28365 27829 28399 27863
rect 29101 27829 29135 27863
rect 34989 27829 35023 27863
rect 47041 27829 47075 27863
rect 20545 27625 20579 27659
rect 27353 27625 27387 27659
rect 28181 27625 28215 27659
rect 29009 27625 29043 27659
rect 32045 27625 32079 27659
rect 33517 27625 33551 27659
rect 35449 27625 35483 27659
rect 10149 27557 10183 27591
rect 11161 27557 11195 27591
rect 17601 27557 17635 27591
rect 20729 27557 20763 27591
rect 24501 27557 24535 27591
rect 37289 27557 37323 27591
rect 1869 27489 1903 27523
rect 9965 27489 9999 27523
rect 10701 27489 10735 27523
rect 12173 27489 12207 27523
rect 24685 27489 24719 27523
rect 46305 27489 46339 27523
rect 48145 27489 48179 27523
rect 1409 27421 1443 27455
rect 9873 27421 9907 27455
rect 10793 27421 10827 27455
rect 12440 27421 12474 27455
rect 14841 27421 14875 27455
rect 17417 27421 17451 27455
rect 20269 27421 20303 27455
rect 22477 27421 22511 27455
rect 24409 27421 24443 27455
rect 25973 27421 26007 27455
rect 28641 27421 28675 27455
rect 29561 27421 29595 27455
rect 29817 27421 29851 27455
rect 32301 27421 32335 27455
rect 32410 27415 32444 27449
rect 32526 27421 32560 27455
rect 32689 27421 32723 27455
rect 35265 27421 35299 27455
rect 35909 27421 35943 27455
rect 36165 27421 36199 27455
rect 1593 27353 1627 27387
rect 9505 27353 9539 27387
rect 15108 27353 15142 27387
rect 22744 27353 22778 27387
rect 26240 27353 26274 27387
rect 27813 27353 27847 27387
rect 27997 27353 28031 27387
rect 28825 27353 28859 27387
rect 33149 27353 33183 27387
rect 33333 27353 33367 27387
rect 35081 27353 35115 27387
rect 46489 27353 46523 27387
rect 13553 27285 13587 27319
rect 16221 27285 16255 27319
rect 23857 27285 23891 27319
rect 24685 27285 24719 27319
rect 30941 27285 30975 27319
rect 2145 27081 2179 27115
rect 9597 27081 9631 27115
rect 22937 27081 22971 27115
rect 10793 27013 10827 27047
rect 14197 27013 14231 27047
rect 15117 27013 15151 27047
rect 2053 26945 2087 26979
rect 2881 26945 2915 26979
rect 8677 26945 8711 26979
rect 8861 26945 8895 26979
rect 9045 26945 9079 26979
rect 9873 26945 9907 26979
rect 9978 26951 10012 26985
rect 10078 26945 10112 26979
rect 10241 26945 10275 26979
rect 10701 26945 10735 26979
rect 10885 26945 10919 26979
rect 14841 26945 14875 26979
rect 23213 26945 23247 26979
rect 23305 26945 23339 26979
rect 23397 26945 23431 26979
rect 23581 26945 23615 26979
rect 27077 26945 27111 26979
rect 32689 26945 32723 26979
rect 32781 26945 32815 26979
rect 32873 26945 32907 26979
rect 33057 26945 33091 26979
rect 33977 26945 34011 26979
rect 34069 26945 34103 26979
rect 34161 26945 34195 26979
rect 34345 26945 34379 26979
rect 35081 26945 35115 26979
rect 35173 26945 35207 26979
rect 35265 26945 35299 26979
rect 35449 26945 35483 26979
rect 35909 26945 35943 26979
rect 36093 26945 36127 26979
rect 8953 26877 8987 26911
rect 15117 26877 15151 26911
rect 27261 26877 27295 26911
rect 28089 26877 28123 26911
rect 29745 26877 29779 26911
rect 29929 26877 29963 26911
rect 31585 26877 31619 26911
rect 36277 26877 36311 26911
rect 1593 26741 1627 26775
rect 9137 26741 9171 26775
rect 14289 26741 14323 26775
rect 14933 26741 14967 26775
rect 32413 26741 32447 26775
rect 33701 26741 33735 26775
rect 34805 26741 34839 26775
rect 6193 26537 6227 26571
rect 9781 26537 9815 26571
rect 21557 26537 21591 26571
rect 27169 26537 27203 26571
rect 29929 26537 29963 26571
rect 34161 26537 34195 26571
rect 38945 26537 38979 26571
rect 6653 26469 6687 26503
rect 10609 26469 10643 26503
rect 12081 26469 12115 26503
rect 14105 26469 14139 26503
rect 36737 26469 36771 26503
rect 1409 26401 1443 26435
rect 2789 26401 2823 26435
rect 6285 26401 6319 26435
rect 31861 26401 31895 26435
rect 32137 26401 32171 26435
rect 6469 26333 6503 26367
rect 9395 26333 9429 26367
rect 9495 26333 9529 26367
rect 9597 26333 9631 26367
rect 10425 26333 10459 26367
rect 12357 26333 12391 26367
rect 14105 26333 14139 26367
rect 14381 26333 14415 26367
rect 14841 26333 14875 26367
rect 15301 26333 15335 26367
rect 17831 26333 17865 26367
rect 17966 26327 18000 26361
rect 18082 26333 18116 26367
rect 18245 26333 18279 26367
rect 19533 26333 19567 26367
rect 20177 26333 20211 26367
rect 27077 26333 27111 26367
rect 29837 26333 29871 26367
rect 30757 26333 30791 26367
rect 33793 26333 33827 26367
rect 35357 26333 35391 26367
rect 35613 26333 35647 26367
rect 38117 26333 38151 26367
rect 38761 26333 38795 26367
rect 1593 26265 1627 26299
rect 5917 26265 5951 26299
rect 6193 26265 6227 26299
rect 10241 26265 10275 26299
rect 12081 26265 12115 26299
rect 19349 26265 19383 26299
rect 20422 26265 20456 26299
rect 31125 26265 31159 26299
rect 33977 26265 34011 26299
rect 47961 26265 47995 26299
rect 48145 26265 48179 26299
rect 12265 26197 12299 26231
rect 14289 26197 14323 26231
rect 15117 26197 15151 26231
rect 15209 26197 15243 26231
rect 17601 26197 17635 26231
rect 19717 26197 19751 26231
rect 38209 26197 38243 26231
rect 2237 25993 2271 26027
rect 12633 25993 12667 26027
rect 18429 25993 18463 26027
rect 20085 25993 20119 26027
rect 23397 25993 23431 26027
rect 33701 25993 33735 26027
rect 35633 25993 35667 26027
rect 22937 25925 22971 25959
rect 24777 25925 24811 25959
rect 31309 25925 31343 25959
rect 38301 25925 38335 25959
rect 46949 25925 46983 25959
rect 1593 25857 1627 25891
rect 2145 25857 2179 25891
rect 10241 25857 10275 25891
rect 12173 25857 12207 25891
rect 12449 25857 12483 25891
rect 13737 25857 13771 25891
rect 14565 25857 14599 25891
rect 14841 25857 14875 25891
rect 16948 25857 16982 25891
rect 19073 25857 19107 25891
rect 19165 25857 19199 25891
rect 19257 25857 19291 25891
rect 19441 25857 19475 25891
rect 20315 25857 20349 25891
rect 20453 25857 20487 25891
rect 20545 25857 20579 25891
rect 20729 25857 20763 25891
rect 23213 25857 23247 25891
rect 23857 25857 23891 25891
rect 24133 25857 24167 25891
rect 24961 25857 24995 25891
rect 25053 25857 25087 25891
rect 26157 25857 26191 25891
rect 26341 25857 26375 25891
rect 29929 25857 29963 25891
rect 30941 25857 30975 25891
rect 32577 25857 32611 25891
rect 34253 25857 34287 25891
rect 34520 25857 34554 25891
rect 38117 25857 38151 25891
rect 46857 25857 46891 25891
rect 6837 25789 6871 25823
rect 7021 25789 7055 25823
rect 8677 25789 8711 25823
rect 9965 25789 9999 25823
rect 12265 25789 12299 25823
rect 13645 25789 13679 25823
rect 14657 25789 14691 25823
rect 16681 25789 16715 25823
rect 23121 25789 23155 25823
rect 23949 25789 23983 25823
rect 30113 25789 30147 25823
rect 32321 25789 32355 25823
rect 39957 25789 39991 25823
rect 1409 25721 1443 25755
rect 14105 25721 14139 25755
rect 15025 25721 15059 25755
rect 24317 25721 24351 25755
rect 26157 25721 26191 25755
rect 12173 25653 12207 25687
rect 14565 25653 14599 25687
rect 18061 25653 18095 25687
rect 18797 25653 18831 25687
rect 22569 25653 22603 25687
rect 22937 25653 22971 25687
rect 23765 25653 23799 25687
rect 24133 25653 24167 25687
rect 24777 25653 24811 25687
rect 25237 25653 25271 25687
rect 47777 25653 47811 25687
rect 7021 25449 7055 25483
rect 9229 25449 9263 25483
rect 9965 25449 9999 25483
rect 10149 25449 10183 25483
rect 11069 25449 11103 25483
rect 12357 25449 12391 25483
rect 12541 25449 12575 25483
rect 14289 25449 14323 25483
rect 14473 25449 14507 25483
rect 21465 25449 21499 25483
rect 22201 25449 22235 25483
rect 23581 25449 23615 25483
rect 23765 25449 23799 25483
rect 37657 25449 37691 25483
rect 38117 25449 38151 25483
rect 9321 25313 9355 25347
rect 10701 25313 10735 25347
rect 25237 25313 25271 25347
rect 38117 25313 38151 25347
rect 46305 25313 46339 25347
rect 6929 25245 6963 25279
rect 9045 25245 9079 25279
rect 9137 25245 9171 25279
rect 9781 25245 9815 25279
rect 9965 25245 9999 25279
rect 10793 25245 10827 25279
rect 13001 25245 13035 25279
rect 17233 25245 17267 25279
rect 20085 25245 20119 25279
rect 22017 25245 22051 25279
rect 24409 25245 24443 25279
rect 25145 25245 25179 25279
rect 25329 25245 25363 25279
rect 31125 25245 31159 25279
rect 32689 25245 32723 25279
rect 38025 25245 38059 25279
rect 38301 25245 38335 25279
rect 12173 25177 12207 25211
rect 12373 25177 12407 25211
rect 14105 25177 14139 25211
rect 14321 25177 14355 25211
rect 17500 25177 17534 25211
rect 19257 25177 19291 25211
rect 19441 25177 19475 25211
rect 20330 25177 20364 25211
rect 23397 25177 23431 25211
rect 31953 25177 31987 25211
rect 46489 25177 46523 25211
rect 48145 25177 48179 25211
rect 13093 25109 13127 25143
rect 18613 25109 18647 25143
rect 19625 25109 19659 25143
rect 23581 25109 23615 25143
rect 24593 25109 24627 25143
rect 32781 25109 32815 25143
rect 38485 25109 38519 25143
rect 14105 24905 14139 24939
rect 18429 24905 18463 24939
rect 20085 24905 20119 24939
rect 23857 24905 23891 24939
rect 24777 24905 24811 24939
rect 24961 24905 24995 24939
rect 18245 24837 18279 24871
rect 24593 24837 24627 24871
rect 31493 24837 31527 24871
rect 37473 24837 37507 24871
rect 7665 24769 7699 24803
rect 8309 24769 8343 24803
rect 13829 24769 13863 24803
rect 17233 24769 17267 24803
rect 17417 24769 17451 24803
rect 17601 24769 17635 24803
rect 18061 24769 18095 24803
rect 20361 24769 20395 24803
rect 20453 24769 20487 24803
rect 20545 24769 20579 24803
rect 20729 24769 20763 24803
rect 22063 24769 22097 24803
rect 22201 24772 22235 24806
rect 22293 24769 22327 24803
rect 22477 24769 22511 24803
rect 23765 24769 23799 24803
rect 23949 24769 23983 24803
rect 24685 24769 24719 24803
rect 25513 24769 25547 24803
rect 27261 24769 27295 24803
rect 27353 24769 27387 24803
rect 27445 24769 27479 24803
rect 27629 24769 27663 24803
rect 29423 24769 29457 24803
rect 29542 24769 29576 24803
rect 29674 24772 29708 24806
rect 29837 24769 29871 24803
rect 30849 24769 30883 24803
rect 31309 24769 31343 24803
rect 32597 24769 32631 24803
rect 33609 24769 33643 24803
rect 36553 24769 36587 24803
rect 36645 24769 36679 24803
rect 39129 24769 39163 24803
rect 47961 24769 47995 24803
rect 8493 24701 8527 24735
rect 8769 24701 8803 24735
rect 11529 24701 11563 24735
rect 11713 24701 11747 24735
rect 13369 24701 13403 24735
rect 14105 24701 14139 24735
rect 33793 24701 33827 24735
rect 35449 24701 35483 24735
rect 37289 24701 37323 24735
rect 7757 24633 7791 24667
rect 24409 24633 24443 24667
rect 25605 24633 25639 24667
rect 48145 24633 48179 24667
rect 13921 24565 13955 24599
rect 21833 24565 21867 24599
rect 26985 24565 27019 24599
rect 29193 24565 29227 24599
rect 32689 24565 32723 24599
rect 1593 24361 1627 24395
rect 10425 24361 10459 24395
rect 12449 24361 12483 24395
rect 13277 24361 13311 24395
rect 13461 24361 13495 24395
rect 14105 24361 14139 24395
rect 22661 24361 22695 24395
rect 34805 24361 34839 24395
rect 29009 24293 29043 24327
rect 3801 24225 3835 24259
rect 10149 24225 10183 24259
rect 13093 24225 13127 24259
rect 18153 24225 18187 24259
rect 20269 24225 20303 24259
rect 26801 24225 26835 24259
rect 32505 24225 32539 24259
rect 37289 24225 37323 24259
rect 47593 24225 47627 24259
rect 1409 24157 1443 24191
rect 3065 24157 3099 24191
rect 10057 24157 10091 24191
rect 12357 24157 12391 24191
rect 12541 24157 12575 24191
rect 13277 24157 13311 24191
rect 14105 24157 14139 24191
rect 14289 24157 14323 24191
rect 17877 24157 17911 24191
rect 19901 24157 19935 24191
rect 20085 24157 20119 24191
rect 24593 24157 24627 24191
rect 24685 24157 24719 24191
rect 25145 24157 25179 24191
rect 25973 24157 26007 24191
rect 26065 24157 26099 24191
rect 26157 24157 26191 24191
rect 26341 24157 26375 24191
rect 29561 24157 29595 24191
rect 29828 24157 29862 24191
rect 32321 24157 32355 24191
rect 34713 24157 34747 24191
rect 47317 24157 47351 24191
rect 3157 24089 3191 24123
rect 3985 24089 4019 24123
rect 5641 24089 5675 24123
rect 13001 24089 13035 24123
rect 21373 24089 21407 24123
rect 25053 24089 25087 24123
rect 25697 24089 25731 24123
rect 27046 24089 27080 24123
rect 28641 24089 28675 24123
rect 28825 24089 28859 24123
rect 34161 24089 34195 24123
rect 37473 24089 37507 24123
rect 39129 24089 39163 24123
rect 14473 24021 14507 24055
rect 28181 24021 28215 24055
rect 30941 24021 30975 24055
rect 19349 23817 19383 23851
rect 31125 23817 31159 23851
rect 37473 23817 37507 23851
rect 17233 23749 17267 23783
rect 29101 23749 29135 23783
rect 7849 23681 7883 23715
rect 8116 23681 8150 23715
rect 13185 23681 13219 23715
rect 13921 23681 13955 23715
rect 14657 23681 14691 23715
rect 19533 23681 19567 23715
rect 23397 23681 23431 23715
rect 23673 23681 23707 23715
rect 24409 23681 24443 23715
rect 24685 23681 24719 23715
rect 25605 23681 25639 23715
rect 26985 23681 27019 23715
rect 27241 23681 27275 23715
rect 28917 23681 28951 23715
rect 30001 23681 30035 23715
rect 37381 23681 37415 23715
rect 18061 23613 18095 23647
rect 18337 23613 18371 23647
rect 23489 23613 23523 23647
rect 24501 23613 24535 23647
rect 25329 23613 25363 23647
rect 29745 23613 29779 23647
rect 33241 23613 33275 23647
rect 33425 23613 33459 23647
rect 35081 23613 35115 23647
rect 17417 23545 17451 23579
rect 2053 23477 2087 23511
rect 9229 23477 9263 23511
rect 13277 23477 13311 23511
rect 14013 23477 14047 23511
rect 14749 23477 14783 23511
rect 23397 23477 23431 23511
rect 23857 23477 23891 23511
rect 24685 23477 24719 23511
rect 24869 23477 24903 23511
rect 28365 23477 28399 23511
rect 29285 23477 29319 23511
rect 23765 23273 23799 23307
rect 27537 23273 27571 23307
rect 29561 23273 29595 23307
rect 33241 23273 33275 23307
rect 47869 23273 47903 23307
rect 8953 23205 8987 23239
rect 15485 23205 15519 23239
rect 17325 23205 17359 23239
rect 22201 23205 22235 23239
rect 1409 23137 1443 23171
rect 2789 23137 2823 23171
rect 13093 23137 13127 23171
rect 20821 23137 20855 23171
rect 25881 23137 25915 23171
rect 47409 23137 47443 23171
rect 8217 23069 8251 23103
rect 9229 23069 9263 23103
rect 9334 23066 9368 23100
rect 9434 23063 9468 23097
rect 9609 23069 9643 23103
rect 11851 23069 11885 23103
rect 11989 23069 12023 23103
rect 12081 23069 12115 23103
rect 12265 23069 12299 23103
rect 12725 23069 12759 23103
rect 14105 23069 14139 23103
rect 15945 23069 15979 23103
rect 18061 23069 18095 23103
rect 18153 23069 18187 23103
rect 18245 23069 18279 23103
rect 18429 23069 18463 23103
rect 19449 23069 19483 23103
rect 21088 23069 21122 23103
rect 22753 23069 22787 23103
rect 23489 23069 23523 23103
rect 24685 23069 24719 23103
rect 25605 23069 25639 23103
rect 27353 23069 27387 23103
rect 28595 23069 28629 23103
rect 28733 23069 28767 23103
rect 28825 23066 28859 23100
rect 29009 23069 29043 23103
rect 29817 23069 29851 23103
rect 29929 23069 29963 23103
rect 30021 23069 30055 23103
rect 30205 23069 30239 23103
rect 33149 23069 33183 23103
rect 47501 23069 47535 23103
rect 47869 23069 47903 23103
rect 1593 23001 1627 23035
rect 8033 23001 8067 23035
rect 8401 23001 8435 23035
rect 12909 23001 12943 23035
rect 14350 23001 14384 23035
rect 16190 23001 16224 23035
rect 24961 23001 24995 23035
rect 27169 23001 27203 23035
rect 11621 22933 11655 22967
rect 17785 22933 17819 22967
rect 19257 22933 19291 22967
rect 22845 22933 22879 22967
rect 28365 22933 28399 22967
rect 48053 22933 48087 22967
rect 1593 22729 1627 22763
rect 2329 22729 2363 22763
rect 14197 22729 14231 22763
rect 15485 22729 15519 22763
rect 27353 22729 27387 22763
rect 28825 22729 28859 22763
rect 47961 22729 47995 22763
rect 9045 22661 9079 22695
rect 11774 22661 11808 22695
rect 13553 22661 13587 22695
rect 22078 22661 22112 22695
rect 32382 22661 32416 22695
rect 1409 22593 1443 22627
rect 2237 22593 2271 22627
rect 7205 22593 7239 22627
rect 7472 22593 7506 22627
rect 9229 22593 9263 22627
rect 11529 22593 11563 22627
rect 13369 22593 13403 22627
rect 14473 22593 14507 22627
rect 14565 22593 14599 22627
rect 14657 22593 14691 22627
rect 14841 22593 14875 22627
rect 15209 22593 15243 22627
rect 15761 22593 15795 22627
rect 15853 22593 15887 22627
rect 15945 22593 15979 22627
rect 16129 22593 16163 22627
rect 16865 22593 16899 22627
rect 17509 22593 17543 22627
rect 17776 22593 17810 22627
rect 19349 22593 19383 22627
rect 19605 22593 19639 22627
rect 21833 22593 21867 22627
rect 24133 22593 24167 22627
rect 24317 22593 24351 22627
rect 24409 22593 24443 22627
rect 25053 22593 25087 22627
rect 25329 22593 25363 22627
rect 26157 22593 26191 22627
rect 26985 22593 27019 22627
rect 27169 22593 27203 22627
rect 28457 22593 28491 22627
rect 28641 22593 28675 22627
rect 29285 22593 29319 22627
rect 29541 22593 29575 22627
rect 32137 22593 32171 22627
rect 48145 22593 48179 22627
rect 10057 22525 10091 22559
rect 10333 22525 10367 22559
rect 13737 22525 13771 22559
rect 25237 22525 25271 22559
rect 24593 22457 24627 22491
rect 25973 22457 26007 22491
rect 33517 22457 33551 22491
rect 8585 22389 8619 22423
rect 9413 22389 9447 22423
rect 12909 22389 12943 22423
rect 16957 22389 16991 22423
rect 18889 22389 18923 22423
rect 20729 22389 20763 22423
rect 23213 22389 23247 22423
rect 24225 22389 24259 22423
rect 25329 22389 25363 22423
rect 25513 22389 25547 22423
rect 30665 22389 30699 22423
rect 13001 22185 13035 22219
rect 15945 22185 15979 22219
rect 16589 22185 16623 22219
rect 18337 22185 18371 22219
rect 20821 22185 20855 22219
rect 30389 22185 30423 22219
rect 33793 22185 33827 22219
rect 6469 22049 6503 22083
rect 8953 22049 8987 22083
rect 11621 22049 11655 22083
rect 19257 22049 19291 22083
rect 22017 22049 22051 22083
rect 48145 22049 48179 22083
rect 9229 21981 9263 22015
rect 9318 21975 9352 22009
rect 9434 21981 9468 22015
rect 9597 21981 9631 22015
rect 16497 21981 16531 22015
rect 19533 21981 19567 22015
rect 19625 21981 19659 22015
rect 19717 21981 19751 22015
rect 19901 21981 19935 22015
rect 21005 21981 21039 22015
rect 24685 21981 24719 22015
rect 30619 21981 30653 22015
rect 30738 21981 30772 22015
rect 30854 21981 30888 22015
rect 31033 21981 31067 22015
rect 31769 21981 31803 22015
rect 31858 21981 31892 22015
rect 31953 21975 31987 22009
rect 32137 21981 32171 22015
rect 32597 21981 32631 22015
rect 33425 21981 33459 22015
rect 33609 21981 33643 22015
rect 34713 21981 34747 22015
rect 36553 21981 36587 22015
rect 6653 21913 6687 21947
rect 8309 21913 8343 21947
rect 10425 21913 10459 21947
rect 11866 21913 11900 21947
rect 15577 21913 15611 21947
rect 15761 21913 15795 21947
rect 17969 21913 18003 21947
rect 18153 21913 18187 21947
rect 21833 21913 21867 21947
rect 24409 21913 24443 21947
rect 32781 21913 32815 21947
rect 34897 21913 34931 21947
rect 47961 21913 47995 21947
rect 10517 21845 10551 21879
rect 21465 21845 21499 21879
rect 21925 21845 21959 21879
rect 24507 21845 24541 21879
rect 24593 21845 24627 21879
rect 31493 21845 31527 21879
rect 32965 21845 32999 21879
rect 6745 21641 6779 21675
rect 11621 21641 11655 21675
rect 18981 21641 19015 21675
rect 24041 21641 24075 21675
rect 33885 21641 33919 21675
rect 12725 21573 12759 21607
rect 14013 21573 14047 21607
rect 17785 21573 17819 21607
rect 18613 21573 18647 21607
rect 22753 21573 22787 21607
rect 24133 21573 24167 21607
rect 32750 21573 32784 21607
rect 6653 21505 6687 21539
rect 9505 21505 9539 21539
rect 9594 21508 9628 21542
rect 9689 21505 9723 21539
rect 9873 21505 9907 21539
rect 11851 21505 11885 21539
rect 12002 21511 12036 21545
rect 12102 21505 12136 21539
rect 12265 21505 12299 21539
rect 12909 21505 12943 21539
rect 17969 21505 18003 21539
rect 18797 21505 18831 21539
rect 22661 21505 22695 21539
rect 24961 21505 24995 21539
rect 25228 21505 25262 21539
rect 31217 21505 31251 21539
rect 31309 21505 31343 21539
rect 31401 21505 31435 21539
rect 31585 21505 31619 21539
rect 13093 21437 13127 21471
rect 13829 21437 13863 21471
rect 14289 21437 14323 21471
rect 22937 21437 22971 21471
rect 24225 21437 24259 21471
rect 32505 21437 32539 21471
rect 34529 21437 34563 21471
rect 34713 21437 34747 21471
rect 36369 21437 36403 21471
rect 9229 21301 9263 21335
rect 18153 21301 18187 21335
rect 22293 21301 22327 21335
rect 23673 21301 23707 21335
rect 26341 21301 26375 21335
rect 30941 21301 30975 21335
rect 11161 21097 11195 21131
rect 21741 21097 21775 21131
rect 23121 21097 23155 21131
rect 25421 21097 25455 21131
rect 32229 21097 32263 21131
rect 34805 21097 34839 21131
rect 18429 21029 18463 21063
rect 22753 21029 22787 21063
rect 17049 20961 17083 20995
rect 21281 20961 21315 20995
rect 22201 20961 22235 20995
rect 24961 20961 24995 20995
rect 25053 20961 25087 20995
rect 26157 20961 26191 20995
rect 30481 20961 30515 20995
rect 30757 20961 30791 20995
rect 6653 20893 6687 20927
rect 8033 20893 8067 20927
rect 8953 20893 8987 20927
rect 9220 20893 9254 20927
rect 10793 20893 10827 20927
rect 14197 20893 14231 20927
rect 21005 20893 21039 20927
rect 21097 20893 21131 20927
rect 21925 20893 21959 20927
rect 22017 20893 22051 20927
rect 22293 20893 22327 20927
rect 22937 20893 22971 20927
rect 23213 20893 23247 20927
rect 23857 20893 23891 20927
rect 24685 20893 24719 20927
rect 24869 20893 24903 20927
rect 25237 20893 25271 20927
rect 25881 20893 25915 20927
rect 25973 20893 26007 20927
rect 26617 20893 26651 20927
rect 26801 20893 26835 20927
rect 27629 20893 27663 20927
rect 32689 20893 32723 20927
rect 32945 20893 32979 20927
rect 34713 20893 34747 20927
rect 8217 20825 8251 20859
rect 10977 20825 11011 20859
rect 14442 20825 14476 20859
rect 17294 20825 17328 20859
rect 21281 20825 21315 20859
rect 27874 20825 27908 20859
rect 31861 20825 31895 20859
rect 32045 20825 32079 20859
rect 6745 20757 6779 20791
rect 8401 20757 8435 20791
rect 10333 20757 10367 20791
rect 15577 20757 15611 20791
rect 23673 20757 23707 20791
rect 26157 20757 26191 20791
rect 26709 20757 26743 20791
rect 29009 20757 29043 20791
rect 34069 20757 34103 20791
rect 13921 20553 13955 20587
rect 16865 20553 16899 20587
rect 23489 20553 23523 20587
rect 34437 20553 34471 20587
rect 5733 20485 5767 20519
rect 6561 20485 6595 20519
rect 10517 20485 10551 20519
rect 19441 20485 19475 20519
rect 22201 20485 22235 20519
rect 22385 20485 22419 20519
rect 27905 20485 27939 20519
rect 5641 20417 5675 20451
rect 8677 20417 8711 20451
rect 8944 20417 8978 20451
rect 10701 20417 10735 20451
rect 13277 20417 13311 20451
rect 14177 20417 14211 20451
rect 14289 20417 14323 20451
rect 14402 20417 14436 20451
rect 14565 20417 14599 20451
rect 15945 20417 15979 20451
rect 16129 20417 16163 20451
rect 17141 20417 17175 20451
rect 17233 20417 17267 20451
rect 17325 20417 17359 20451
rect 17509 20417 17543 20451
rect 18245 20417 18279 20451
rect 18337 20417 18371 20451
rect 18429 20417 18463 20451
rect 18613 20417 18647 20451
rect 19073 20417 19107 20451
rect 19257 20417 19291 20451
rect 20177 20417 20211 20451
rect 20913 20417 20947 20451
rect 21097 20417 21131 20451
rect 23305 20417 23339 20451
rect 24317 20417 24351 20451
rect 25145 20417 25179 20451
rect 25973 20417 26007 20451
rect 27813 20417 27847 20451
rect 28825 20417 28859 20451
rect 30849 20417 30883 20451
rect 32137 20417 32171 20451
rect 32321 20417 32355 20451
rect 34345 20417 34379 20451
rect 6377 20349 6411 20383
rect 8033 20349 8067 20383
rect 16037 20349 16071 20383
rect 20453 20349 20487 20383
rect 27997 20349 28031 20383
rect 29101 20349 29135 20383
rect 20269 20281 20303 20315
rect 22569 20281 22603 20315
rect 25421 20281 25455 20315
rect 30665 20281 30699 20315
rect 10057 20213 10091 20247
rect 10885 20213 10919 20247
rect 13369 20213 13403 20247
rect 17969 20213 18003 20247
rect 20361 20213 20395 20247
rect 21005 20213 21039 20247
rect 21281 20213 21315 20247
rect 24501 20213 24535 20247
rect 26157 20213 26191 20247
rect 27445 20213 27479 20247
rect 28641 20213 28675 20247
rect 29009 20213 29043 20247
rect 32505 20213 32539 20247
rect 47777 20213 47811 20247
rect 8953 20009 8987 20043
rect 18705 20009 18739 20043
rect 27721 20009 27755 20043
rect 21097 19941 21131 19975
rect 23581 19941 23615 19975
rect 6469 19873 6503 19907
rect 6653 19873 6687 19907
rect 6929 19873 6963 19907
rect 10149 19873 10183 19907
rect 21649 19873 21683 19907
rect 22569 19873 22603 19907
rect 22753 19873 22787 19907
rect 24777 19873 24811 19907
rect 46305 19873 46339 19907
rect 9183 19805 9217 19839
rect 9321 19805 9355 19839
rect 9413 19802 9447 19836
rect 9597 19805 9631 19839
rect 10425 19805 10459 19839
rect 14289 19805 14323 19839
rect 17325 19805 17359 19839
rect 17592 19805 17626 19839
rect 19257 19805 19291 19839
rect 22477 19805 22511 19839
rect 22661 19805 22695 19839
rect 23397 19805 23431 19839
rect 25053 19805 25087 19839
rect 26433 19805 26467 19839
rect 26709 19805 26743 19839
rect 27169 19805 27203 19839
rect 27537 19805 27571 19839
rect 30297 19805 30331 19839
rect 31815 19805 31849 19839
rect 31953 19805 31987 19839
rect 32045 19805 32079 19839
rect 32229 19805 32263 19839
rect 32965 19805 32999 19839
rect 33057 19805 33091 19839
rect 33149 19805 33183 19839
rect 33333 19805 33367 19839
rect 48145 19805 48179 19839
rect 14105 19737 14139 19771
rect 19524 19737 19558 19771
rect 21557 19737 21591 19771
rect 26249 19737 26283 19771
rect 27353 19737 27387 19771
rect 27445 19737 27479 19771
rect 46489 19737 46523 19771
rect 14473 19669 14507 19703
rect 20637 19669 20671 19703
rect 21465 19669 21499 19703
rect 22293 19669 22327 19703
rect 26617 19669 26651 19703
rect 30527 19669 30561 19703
rect 31585 19669 31619 19703
rect 32689 19669 32723 19703
rect 15945 19465 15979 19499
rect 17693 19465 17727 19499
rect 20269 19465 20303 19499
rect 23397 19465 23431 19499
rect 27905 19465 27939 19499
rect 30021 19465 30055 19499
rect 33517 19465 33551 19499
rect 46949 19465 46983 19499
rect 12541 19397 12575 19431
rect 14197 19397 14231 19431
rect 15853 19397 15887 19431
rect 17601 19397 17635 19431
rect 21925 19397 21959 19431
rect 23949 19397 23983 19431
rect 26065 19397 26099 19431
rect 31217 19397 31251 19431
rect 31585 19397 31619 19431
rect 32404 19397 32438 19431
rect 2145 19329 2179 19363
rect 9404 19329 9438 19363
rect 14933 19329 14967 19363
rect 15025 19329 15059 19363
rect 15117 19329 15151 19363
rect 15301 19329 15335 19363
rect 16681 19329 16715 19363
rect 20637 19329 20671 19363
rect 20729 19329 20763 19363
rect 22201 19329 22235 19363
rect 23121 19329 23155 19363
rect 23213 19329 23247 19363
rect 24869 19329 24903 19363
rect 26249 19329 26283 19363
rect 27813 19329 27847 19363
rect 28641 19329 28675 19363
rect 28908 19329 28942 19363
rect 31401 19329 31435 19363
rect 32137 19329 32171 19363
rect 46857 19329 46891 19363
rect 47961 19329 47995 19363
rect 9137 19261 9171 19295
rect 12357 19261 12391 19295
rect 16773 19261 16807 19295
rect 20913 19261 20947 19295
rect 22017 19261 22051 19295
rect 23397 19261 23431 19295
rect 24593 19261 24627 19295
rect 27997 19261 28031 19295
rect 10517 19193 10551 19227
rect 24133 19193 24167 19227
rect 1685 19125 1719 19159
rect 2237 19125 2271 19159
rect 14657 19125 14691 19159
rect 21925 19125 21959 19159
rect 22385 19125 22419 19159
rect 26433 19125 26467 19159
rect 27445 19125 27479 19159
rect 48053 19125 48087 19159
rect 9597 18921 9631 18955
rect 12633 18921 12667 18955
rect 20407 18921 20441 18955
rect 21189 18921 21223 18955
rect 25421 18921 25455 18955
rect 26249 18921 26283 18955
rect 27077 18921 27111 18955
rect 27537 18921 27571 18955
rect 28825 18921 28859 18955
rect 26433 18853 26467 18887
rect 1409 18785 1443 18819
rect 1593 18785 1627 18819
rect 2789 18785 2823 18819
rect 20545 18785 20579 18819
rect 21281 18785 21315 18819
rect 26157 18785 26191 18819
rect 28365 18785 28399 18819
rect 28457 18785 28491 18819
rect 9827 18717 9861 18751
rect 9965 18717 9999 18751
rect 10057 18714 10091 18748
rect 10241 18717 10275 18751
rect 11253 18717 11287 18751
rect 13277 18717 13311 18751
rect 14335 18717 14369 18751
rect 14473 18717 14507 18751
rect 14565 18717 14599 18751
rect 14749 18717 14783 18751
rect 15669 18717 15703 18751
rect 17509 18717 17543 18751
rect 17693 18717 17727 18751
rect 20269 18717 20303 18751
rect 20729 18717 20763 18751
rect 21465 18717 21499 18751
rect 22109 18717 22143 18751
rect 23397 18717 23431 18751
rect 23489 18717 23523 18751
rect 24409 18717 24443 18751
rect 24777 18717 24811 18751
rect 25237 18717 25271 18751
rect 25973 18717 26007 18751
rect 26249 18717 26283 18751
rect 26985 18717 27019 18751
rect 27353 18717 27387 18751
rect 28089 18717 28123 18751
rect 28273 18717 28307 18751
rect 28641 18717 28675 18751
rect 30849 18717 30883 18751
rect 31116 18717 31150 18751
rect 11520 18649 11554 18683
rect 13093 18649 13127 18683
rect 13461 18649 13495 18683
rect 15936 18649 15970 18683
rect 21189 18649 21223 18683
rect 22201 18649 22235 18683
rect 23673 18649 23707 18683
rect 24593 18649 24627 18683
rect 14105 18581 14139 18615
rect 17049 18581 17083 18615
rect 17693 18581 17727 18615
rect 20729 18581 20763 18615
rect 21649 18581 21683 18615
rect 32229 18581 32263 18615
rect 14197 18377 14231 18411
rect 16681 18377 16715 18411
rect 17785 18377 17819 18411
rect 20545 18377 20579 18411
rect 25789 18377 25823 18411
rect 27813 18377 27847 18411
rect 15761 18309 15795 18343
rect 15945 18309 15979 18343
rect 17049 18309 17083 18343
rect 17601 18309 17635 18343
rect 21005 18309 21039 18343
rect 23305 18309 23339 18343
rect 25697 18309 25731 18343
rect 28641 18309 28675 18343
rect 12817 18241 12851 18275
rect 13084 18241 13118 18275
rect 14913 18241 14947 18275
rect 15025 18241 15059 18275
rect 15117 18241 15151 18275
rect 15301 18241 15335 18275
rect 16865 18241 16899 18275
rect 17141 18241 17175 18275
rect 17877 18241 17911 18275
rect 18613 18241 18647 18275
rect 20913 18241 20947 18275
rect 22109 18241 22143 18275
rect 23121 18241 23155 18275
rect 24133 18241 24167 18275
rect 24961 18241 24995 18275
rect 27261 18241 27295 18275
rect 28917 18241 28951 18275
rect 1777 18173 1811 18207
rect 1961 18173 1995 18207
rect 2789 18173 2823 18207
rect 16129 18173 16163 18207
rect 21189 18173 21223 18207
rect 22017 18173 22051 18207
rect 22201 18173 22235 18207
rect 22293 18173 22327 18207
rect 27537 18173 27571 18207
rect 28825 18173 28859 18207
rect 32873 18173 32907 18207
rect 33057 18173 33091 18207
rect 34529 18173 34563 18207
rect 25145 18105 25179 18139
rect 29101 18105 29135 18139
rect 4261 18037 4295 18071
rect 14657 18037 14691 18071
rect 17601 18037 17635 18071
rect 18705 18037 18739 18071
rect 21833 18037 21867 18071
rect 23489 18037 23523 18071
rect 23949 18037 23983 18071
rect 27629 18037 27663 18071
rect 28733 18037 28767 18071
rect 2145 17833 2179 17867
rect 16037 17833 16071 17867
rect 19441 17833 19475 17867
rect 21189 17833 21223 17867
rect 23397 17833 23431 17867
rect 24593 17833 24627 17867
rect 25329 17833 25363 17867
rect 26801 17833 26835 17867
rect 27997 17833 28031 17867
rect 34805 17833 34839 17867
rect 8309 17765 8343 17799
rect 16773 17765 16807 17799
rect 18613 17765 18647 17799
rect 27169 17765 27203 17799
rect 7757 17697 7791 17731
rect 11345 17697 11379 17731
rect 12725 17697 12759 17731
rect 27629 17697 27663 17731
rect 28733 17697 28767 17731
rect 31401 17697 31435 17731
rect 33057 17697 33091 17731
rect 1593 17629 1627 17663
rect 2053 17629 2087 17663
rect 2697 17629 2731 17663
rect 9873 17629 9907 17663
rect 13001 17629 13035 17663
rect 14657 17629 14691 17663
rect 17233 17629 17267 17663
rect 17500 17629 17534 17663
rect 19349 17629 19383 17663
rect 21373 17629 21407 17663
rect 21649 17629 21683 17663
rect 22109 17629 22143 17663
rect 23213 17629 23247 17663
rect 23397 17629 23431 17663
rect 23489 17629 23523 17663
rect 25237 17629 25271 17663
rect 26801 17629 26835 17663
rect 26985 17629 27019 17663
rect 27813 17629 27847 17663
rect 30757 17629 30791 17663
rect 33701 17629 33735 17663
rect 34713 17629 34747 17663
rect 47685 17629 47719 17663
rect 7849 17561 7883 17595
rect 10057 17561 10091 17595
rect 14924 17561 14958 17595
rect 16589 17561 16623 17595
rect 24409 17561 24443 17595
rect 26157 17561 26191 17595
rect 28549 17561 28583 17595
rect 30849 17561 30883 17595
rect 31585 17561 31619 17595
rect 2789 17493 2823 17527
rect 21557 17493 21591 17527
rect 22293 17493 22327 17527
rect 23673 17493 23707 17527
rect 24609 17493 24643 17527
rect 24777 17493 24811 17527
rect 26249 17493 26283 17527
rect 33793 17493 33827 17527
rect 8861 17289 8895 17323
rect 10057 17289 10091 17323
rect 20913 17289 20947 17323
rect 22293 17289 22327 17323
rect 24133 17289 24167 17323
rect 24961 17289 24995 17323
rect 25605 17289 25639 17323
rect 27445 17289 27479 17323
rect 1961 17221 1995 17255
rect 22937 17221 22971 17255
rect 24501 17221 24535 17255
rect 27905 17221 27939 17255
rect 28089 17221 28123 17255
rect 28273 17221 28307 17255
rect 33517 17221 33551 17255
rect 1777 17153 1811 17187
rect 8769 17153 8803 17187
rect 9965 17153 9999 17187
rect 10609 17153 10643 17187
rect 10793 17153 10827 17187
rect 11851 17153 11885 17187
rect 11989 17153 12023 17187
rect 12081 17153 12115 17187
rect 12265 17153 12299 17187
rect 12725 17153 12759 17187
rect 14289 17153 14323 17187
rect 15557 17153 15591 17187
rect 15669 17153 15703 17187
rect 15782 17153 15816 17187
rect 15945 17153 15979 17187
rect 17877 17153 17911 17187
rect 18705 17153 18739 17187
rect 19800 17153 19834 17187
rect 22201 17153 22235 17187
rect 22385 17153 22419 17187
rect 23121 17153 23155 17187
rect 23213 17153 23247 17187
rect 23857 17153 23891 17187
rect 24777 17153 24811 17187
rect 25513 17153 25547 17187
rect 27077 17153 27111 17187
rect 27261 17153 27295 17187
rect 29092 17153 29126 17187
rect 47593 17153 47627 17187
rect 2789 17085 2823 17119
rect 10977 17085 11011 17119
rect 14013 17085 14047 17119
rect 19533 17085 19567 17119
rect 24593 17085 24627 17119
rect 28825 17085 28859 17119
rect 33333 17085 33367 17119
rect 33793 17085 33827 17119
rect 23397 17017 23431 17051
rect 11621 16949 11655 16983
rect 12955 16949 12989 16983
rect 15301 16949 15335 16983
rect 17969 16949 18003 16983
rect 18889 16949 18923 16983
rect 23213 16949 23247 16983
rect 23673 16949 23707 16983
rect 24685 16949 24719 16983
rect 30205 16949 30239 16983
rect 47685 16949 47719 16983
rect 1961 16745 1995 16779
rect 18429 16745 18463 16779
rect 19993 16745 20027 16779
rect 20545 16745 20579 16779
rect 30297 16745 30331 16779
rect 17417 16677 17451 16711
rect 27629 16677 27663 16711
rect 11437 16609 11471 16643
rect 14381 16609 14415 16643
rect 24409 16609 24443 16643
rect 27169 16609 27203 16643
rect 28549 16609 28583 16643
rect 28641 16609 28675 16643
rect 29929 16609 29963 16643
rect 46305 16609 46339 16643
rect 48145 16609 48179 16643
rect 1869 16541 1903 16575
rect 10793 16541 10827 16575
rect 11704 16541 11738 16575
rect 14648 16541 14682 16575
rect 18337 16541 18371 16575
rect 20729 16541 20763 16575
rect 20913 16541 20947 16575
rect 21005 16541 21039 16575
rect 21557 16541 21591 16575
rect 24665 16541 24699 16575
rect 27261 16541 27295 16575
rect 28457 16541 28491 16575
rect 29561 16541 29595 16575
rect 29745 16541 29779 16575
rect 29837 16541 29871 16575
rect 30113 16541 30147 16575
rect 31769 16541 31803 16575
rect 17233 16473 17267 16507
rect 19717 16473 19751 16507
rect 31585 16473 31619 16507
rect 46489 16473 46523 16507
rect 10885 16405 10919 16439
rect 12817 16405 12851 16439
rect 15761 16405 15795 16439
rect 21649 16405 21683 16439
rect 25789 16405 25823 16439
rect 28089 16405 28123 16439
rect 31953 16405 31987 16439
rect 14841 16201 14875 16235
rect 27445 16201 27479 16235
rect 29653 16201 29687 16235
rect 11713 16133 11747 16167
rect 14473 16133 14507 16167
rect 16037 16133 16071 16167
rect 16865 16133 16899 16167
rect 30297 16133 30331 16167
rect 11529 16065 11563 16099
rect 14657 16065 14691 16099
rect 15945 16065 15979 16099
rect 16681 16065 16715 16099
rect 18981 16065 19015 16099
rect 20913 16065 20947 16099
rect 25145 16065 25179 16099
rect 28641 16065 28675 16099
rect 29561 16065 29595 16099
rect 31217 16065 31251 16099
rect 31309 16065 31343 16099
rect 31401 16065 31435 16099
rect 31585 16065 31619 16099
rect 32137 16065 32171 16099
rect 32393 16065 32427 16099
rect 11989 15997 12023 16031
rect 18521 15997 18555 16031
rect 19533 15997 19567 16031
rect 26985 15997 27019 16031
rect 28733 15997 28767 16031
rect 28825 15997 28859 16031
rect 21097 15929 21131 15963
rect 27261 15929 27295 15963
rect 25329 15861 25363 15895
rect 28273 15861 28307 15895
rect 30389 15861 30423 15895
rect 30941 15861 30975 15895
rect 33517 15861 33551 15895
rect 47777 15861 47811 15895
rect 21005 15657 21039 15691
rect 22569 15657 22603 15691
rect 25145 15657 25179 15691
rect 26801 15657 26835 15691
rect 27445 15657 27479 15691
rect 32873 15589 32907 15623
rect 18061 15521 18095 15555
rect 28641 15521 28675 15555
rect 46305 15521 46339 15555
rect 46489 15521 46523 15555
rect 48145 15521 48179 15555
rect 17877 15453 17911 15487
rect 19717 15453 19751 15487
rect 20729 15453 20763 15487
rect 20821 15453 20855 15487
rect 21097 15453 21131 15487
rect 25053 15453 25087 15487
rect 26617 15453 26651 15487
rect 26893 15453 26927 15487
rect 27353 15453 27387 15487
rect 27445 15453 27479 15487
rect 28273 15453 28307 15487
rect 28457 15453 28491 15487
rect 28549 15453 28583 15487
rect 28825 15453 28859 15487
rect 29561 15453 29595 15487
rect 31493 15453 31527 15487
rect 31760 15453 31794 15487
rect 22385 15385 22419 15419
rect 26433 15385 26467 15419
rect 29009 15385 29043 15419
rect 29806 15385 29840 15419
rect 19809 15317 19843 15351
rect 20545 15317 20579 15351
rect 22585 15317 22619 15351
rect 22753 15317 22787 15351
rect 27721 15317 27755 15351
rect 30941 15317 30975 15351
rect 20269 15113 20303 15147
rect 21189 15113 21223 15147
rect 22201 15113 22235 15147
rect 22753 15113 22787 15147
rect 30941 15113 30975 15147
rect 46857 15113 46891 15147
rect 17693 15045 17727 15079
rect 19165 15045 19199 15079
rect 20177 15045 20211 15079
rect 21833 15045 21867 15079
rect 24041 15045 24075 15079
rect 32321 15045 32355 15079
rect 18337 14977 18371 15011
rect 21097 14977 21131 15011
rect 21281 14977 21315 15011
rect 22017 14977 22051 15011
rect 22661 14977 22695 15011
rect 22845 14977 22879 15011
rect 23581 14977 23615 15011
rect 23673 14977 23707 15011
rect 25145 14977 25179 15011
rect 27353 14977 27387 15011
rect 27629 14977 27663 15011
rect 31217 14977 31251 15011
rect 31309 14977 31343 15011
rect 31401 14977 31435 15011
rect 31585 14977 31619 15011
rect 32137 14977 32171 15011
rect 47041 14977 47075 15011
rect 47593 14977 47627 15011
rect 20453 14909 20487 14943
rect 23949 14909 23983 14943
rect 32505 14909 32539 14943
rect 17877 14841 17911 14875
rect 19809 14773 19843 14807
rect 23397 14773 23431 14807
rect 25329 14773 25363 14807
rect 27169 14773 27203 14807
rect 27537 14773 27571 14807
rect 47685 14773 47719 14807
rect 20085 14569 20119 14603
rect 21005 14569 21039 14603
rect 24593 14569 24627 14603
rect 25329 14569 25363 14603
rect 28181 14569 28215 14603
rect 23397 14501 23431 14535
rect 24501 14501 24535 14535
rect 26341 14501 26375 14535
rect 21649 14433 21683 14467
rect 22753 14433 22787 14467
rect 24685 14433 24719 14467
rect 46489 14433 46523 14467
rect 17141 14365 17175 14399
rect 19441 14365 19475 14399
rect 20269 14365 20303 14399
rect 20545 14365 20579 14399
rect 23682 14365 23716 14399
rect 24409 14365 24443 14399
rect 26157 14365 26191 14399
rect 27169 14365 27203 14399
rect 27537 14365 27571 14399
rect 28181 14365 28215 14399
rect 28365 14365 28399 14399
rect 31493 14365 31527 14399
rect 46305 14365 46339 14399
rect 17969 14297 18003 14331
rect 20453 14297 20487 14331
rect 21373 14297 21407 14331
rect 22661 14297 22695 14331
rect 23397 14297 23431 14331
rect 25237 14297 25271 14331
rect 27353 14297 27387 14331
rect 27445 14297 27479 14331
rect 48145 14297 48179 14331
rect 17325 14229 17359 14263
rect 18061 14229 18095 14263
rect 19257 14229 19291 14263
rect 21465 14229 21499 14263
rect 22201 14229 22235 14263
rect 22569 14229 22603 14263
rect 23581 14229 23615 14263
rect 27721 14229 27755 14263
rect 31585 14229 31619 14263
rect 24593 14025 24627 14059
rect 26985 14025 27019 14059
rect 29377 14025 29411 14059
rect 18512 13957 18546 13991
rect 20637 13957 20671 13991
rect 20729 13957 20763 13991
rect 32413 13957 32447 13991
rect 2053 13889 2087 13923
rect 17417 13889 17451 13923
rect 17509 13889 17543 13923
rect 17693 13889 17727 13923
rect 17785 13889 17819 13923
rect 20361 13889 20395 13923
rect 20509 13889 20543 13923
rect 20867 13889 20901 13923
rect 22201 13889 22235 13923
rect 23213 13889 23247 13923
rect 23480 13889 23514 13923
rect 27169 13889 27203 13923
rect 27261 13889 27295 13923
rect 27445 13889 27479 13923
rect 27537 13889 27571 13923
rect 27997 13889 28031 13923
rect 28253 13889 28287 13923
rect 31033 13889 31067 13923
rect 31125 13889 31159 13923
rect 31217 13889 31251 13923
rect 31401 13889 31435 13923
rect 34069 13889 34103 13923
rect 47869 13889 47903 13923
rect 18245 13821 18279 13855
rect 22293 13821 22327 13855
rect 22477 13821 22511 13855
rect 32229 13821 32263 13855
rect 19625 13753 19659 13787
rect 48053 13753 48087 13787
rect 2145 13685 2179 13719
rect 2881 13685 2915 13719
rect 17233 13685 17267 13719
rect 21005 13685 21039 13719
rect 21833 13685 21867 13719
rect 30757 13685 30791 13719
rect 20637 13481 20671 13515
rect 22293 13481 22327 13515
rect 23489 13481 23523 13515
rect 26341 13481 26375 13515
rect 26801 13481 26835 13515
rect 32505 13481 32539 13515
rect 47685 13481 47719 13515
rect 21465 13413 21499 13447
rect 1409 13345 1443 13379
rect 1593 13345 1627 13379
rect 2789 13345 2823 13379
rect 14565 13345 14599 13379
rect 21557 13345 21591 13379
rect 22293 13345 22327 13379
rect 26525 13345 26559 13379
rect 28181 13345 28215 13379
rect 31125 13345 31159 13379
rect 14105 13277 14139 13311
rect 16865 13277 16899 13311
rect 19257 13277 19291 13311
rect 19524 13277 19558 13311
rect 21281 13277 21315 13311
rect 21373 13277 21407 13311
rect 22477 13277 22511 13311
rect 26617 13277 26651 13311
rect 28089 13277 28123 13311
rect 30665 13277 30699 13311
rect 31381 13277 31415 13311
rect 14289 13209 14323 13243
rect 17132 13209 17166 13243
rect 22017 13209 22051 13243
rect 23121 13209 23155 13243
rect 23305 13209 23339 13243
rect 26341 13209 26375 13243
rect 27997 13209 28031 13243
rect 18245 13141 18279 13175
rect 22661 13141 22695 13175
rect 27629 13141 27663 13175
rect 30481 13141 30515 13175
rect 14013 12937 14047 12971
rect 18153 12937 18187 12971
rect 21189 12937 21223 12971
rect 22477 12937 22511 12971
rect 26433 12937 26467 12971
rect 27353 12937 27387 12971
rect 28917 12937 28951 12971
rect 32505 12937 32539 12971
rect 21097 12869 21131 12903
rect 24225 12869 24259 12903
rect 24409 12869 24443 12903
rect 25973 12869 26007 12903
rect 27813 12869 27847 12903
rect 28549 12869 28583 12903
rect 32137 12869 32171 12903
rect 32321 12869 32355 12903
rect 1685 12801 1719 12835
rect 9781 12801 9815 12835
rect 13921 12801 13955 12835
rect 17877 12801 17911 12835
rect 17969 12801 18003 12835
rect 22017 12801 22051 12835
rect 22293 12801 22327 12835
rect 24501 12801 24535 12835
rect 25145 12801 25179 12835
rect 26249 12801 26283 12835
rect 27721 12801 27755 12835
rect 28733 12801 28767 12835
rect 30573 12801 30607 12835
rect 1409 12733 1443 12767
rect 10057 12733 10091 12767
rect 22109 12733 22143 12767
rect 25237 12733 25271 12767
rect 26157 12733 26191 12767
rect 27905 12733 27939 12767
rect 30297 12733 30331 12767
rect 22201 12597 22235 12631
rect 24225 12597 24259 12631
rect 25329 12597 25363 12631
rect 25513 12597 25547 12631
rect 25973 12597 26007 12631
rect 23765 12393 23799 12427
rect 25145 12393 25179 12427
rect 25789 12393 25823 12427
rect 18613 12325 18647 12359
rect 21833 12257 21867 12291
rect 23673 12257 23707 12291
rect 23853 12257 23887 12291
rect 24777 12257 24811 12291
rect 25973 12257 26007 12291
rect 27537 12257 27571 12291
rect 11621 12189 11655 12223
rect 18429 12189 18463 12223
rect 19717 12189 19751 12223
rect 21557 12189 21591 12223
rect 21741 12189 21775 12223
rect 21925 12189 21959 12223
rect 22109 12189 22143 12223
rect 23581 12189 23615 12223
rect 24961 12189 24995 12223
rect 25237 12189 25271 12223
rect 25697 12189 25731 12223
rect 27169 12189 27203 12223
rect 27353 12189 27387 12223
rect 27445 12189 27479 12223
rect 27721 12189 27755 12223
rect 28457 12189 28491 12223
rect 30113 12189 30147 12223
rect 30389 12189 30423 12223
rect 31677 12189 31711 12223
rect 31769 12189 31803 12223
rect 31861 12189 31895 12223
rect 32045 12189 32079 12223
rect 28641 12121 28675 12155
rect 11713 12053 11747 12087
rect 19809 12053 19843 12087
rect 22293 12053 22327 12087
rect 26249 12053 26283 12087
rect 27905 12053 27939 12087
rect 31401 12053 31435 12087
rect 18429 11849 18463 11883
rect 23489 11849 23523 11883
rect 24041 11849 24075 11883
rect 25513 11849 25547 11883
rect 27169 11849 27203 11883
rect 31493 11849 31527 11883
rect 22293 11781 22327 11815
rect 25881 11781 25915 11815
rect 26985 11781 27019 11815
rect 39129 11781 39163 11815
rect 18797 11713 18831 11747
rect 20177 11713 20211 11747
rect 20361 11713 20395 11747
rect 22201 11713 22235 11747
rect 23029 11713 23063 11747
rect 24409 11713 24443 11747
rect 24501 11713 24535 11747
rect 25973 11713 26007 11747
rect 27261 11713 27295 11747
rect 27988 11713 28022 11747
rect 30297 11713 30331 11747
rect 30389 11713 30423 11747
rect 30481 11713 30515 11747
rect 30665 11713 30699 11747
rect 31125 11713 31159 11747
rect 31309 11713 31343 11747
rect 37289 11713 37323 11747
rect 19073 11645 19107 11679
rect 22385 11645 22419 11679
rect 24593 11645 24627 11679
rect 26065 11645 26099 11679
rect 27721 11645 27755 11679
rect 37473 11645 37507 11679
rect 21833 11577 21867 11611
rect 20545 11509 20579 11543
rect 23305 11509 23339 11543
rect 26985 11509 27019 11543
rect 29101 11509 29135 11543
rect 30021 11509 30055 11543
rect 18705 11305 18739 11339
rect 22569 11305 22603 11339
rect 25789 11305 25823 11339
rect 28825 11305 28859 11339
rect 30021 11305 30055 11339
rect 37381 11305 37415 11339
rect 2053 11169 2087 11203
rect 11529 11169 11563 11203
rect 11713 11169 11747 11203
rect 13093 11169 13127 11203
rect 19257 11169 19291 11203
rect 26525 11169 26559 11203
rect 28273 11169 28307 11203
rect 2513 11101 2547 11135
rect 17325 11101 17359 11135
rect 19533 11101 19567 11135
rect 21189 11101 21223 11135
rect 24409 11101 24443 11135
rect 26249 11101 26283 11135
rect 26433 11101 26467 11135
rect 26617 11101 26651 11135
rect 26801 11101 26835 11135
rect 28733 11101 28767 11135
rect 28917 11101 28951 11135
rect 30481 11101 30515 11135
rect 30748 11101 30782 11135
rect 37289 11101 37323 11135
rect 47133 11101 47167 11135
rect 47961 11101 47995 11135
rect 1869 11033 1903 11067
rect 17592 11033 17626 11067
rect 21456 11033 21490 11067
rect 24676 11033 24710 11067
rect 28089 11033 28123 11067
rect 29653 11033 29687 11067
rect 29837 11033 29871 11067
rect 2605 10965 2639 10999
rect 26985 10965 27019 10999
rect 31861 10965 31895 10999
rect 47225 10965 47259 10999
rect 18797 10761 18831 10795
rect 21281 10761 21315 10795
rect 24685 10761 24719 10795
rect 25329 10761 25363 10795
rect 1961 10693 1995 10727
rect 18153 10693 18187 10727
rect 18337 10693 18371 10727
rect 25237 10693 25271 10727
rect 30012 10693 30046 10727
rect 17969 10625 18003 10659
rect 19073 10625 19107 10659
rect 19165 10625 19199 10659
rect 19257 10625 19291 10659
rect 19441 10625 19475 10659
rect 19901 10625 19935 10659
rect 20168 10625 20202 10659
rect 23949 10625 23983 10659
rect 24133 10625 24167 10659
rect 24225 10625 24259 10659
rect 24501 10625 24535 10659
rect 47777 10625 47811 10659
rect 1777 10557 1811 10591
rect 2973 10557 3007 10591
rect 24317 10557 24351 10591
rect 29745 10557 29779 10591
rect 31125 10421 31159 10455
rect 47869 10421 47903 10455
rect 1593 10217 1627 10251
rect 20085 10217 20119 10251
rect 27169 10217 27203 10251
rect 25789 10081 25823 10115
rect 46305 10081 46339 10115
rect 46489 10081 46523 10115
rect 48145 10081 48179 10115
rect 2237 10013 2271 10047
rect 2697 10013 2731 10047
rect 20341 10013 20375 10047
rect 20434 10013 20468 10047
rect 20550 10010 20584 10044
rect 20729 10013 20763 10047
rect 26056 10013 26090 10047
rect 19257 9945 19291 9979
rect 19441 9945 19475 9979
rect 2789 9877 2823 9911
rect 19625 9877 19659 9911
rect 2145 9605 2179 9639
rect 24409 9605 24443 9639
rect 1961 9537 1995 9571
rect 17325 9537 17359 9571
rect 17592 9537 17626 9571
rect 19441 9537 19475 9571
rect 19533 9537 19567 9571
rect 19625 9537 19659 9571
rect 19809 9537 19843 9571
rect 23029 9537 23063 9571
rect 27077 9537 27111 9571
rect 27261 9537 27295 9571
rect 28161 9537 28195 9571
rect 29929 9537 29963 9571
rect 30573 9537 30607 9571
rect 2881 9469 2915 9503
rect 23305 9469 23339 9503
rect 27905 9469 27939 9503
rect 19165 9401 19199 9435
rect 18705 9333 18739 9367
rect 24501 9333 24535 9367
rect 27445 9333 27479 9367
rect 29285 9333 29319 9367
rect 30021 9333 30055 9367
rect 30665 9333 30699 9367
rect 27261 9129 27295 9163
rect 19257 8993 19291 9027
rect 22845 8993 22879 9027
rect 30021 8993 30055 9027
rect 30297 8993 30331 9027
rect 21281 8925 21315 8959
rect 23121 8925 23155 8959
rect 24731 8925 24765 8959
rect 24866 8925 24900 8959
rect 24961 8925 24995 8959
rect 25145 8925 25179 8959
rect 26433 8925 26467 8959
rect 27491 8925 27525 8959
rect 27626 8925 27660 8959
rect 27721 8925 27755 8959
rect 27905 8925 27939 8959
rect 29837 8925 29871 8959
rect 19524 8857 19558 8891
rect 21097 8857 21131 8891
rect 22017 8857 22051 8891
rect 22201 8857 22235 8891
rect 26617 8857 26651 8891
rect 47961 8857 47995 8891
rect 20637 8789 20671 8823
rect 21465 8789 21499 8823
rect 22385 8789 22419 8823
rect 24501 8789 24535 8823
rect 26801 8789 26835 8823
rect 48053 8789 48087 8823
rect 47869 8585 47903 8619
rect 22017 8517 22051 8551
rect 23112 8517 23146 8551
rect 29929 8517 29963 8551
rect 1869 8449 1903 8483
rect 17969 8449 18003 8483
rect 20591 8449 20625 8483
rect 20710 8449 20744 8483
rect 20821 8449 20855 8483
rect 21005 8449 21039 8483
rect 21833 8449 21867 8483
rect 22845 8449 22879 8483
rect 24869 8449 24903 8483
rect 25125 8449 25159 8483
rect 26985 8449 27019 8483
rect 27252 8449 27286 8483
rect 29745 8449 29779 8483
rect 47777 8449 47811 8483
rect 18153 8381 18187 8415
rect 19349 8381 19383 8415
rect 31217 8381 31251 8415
rect 2145 8313 2179 8347
rect 22201 8313 22235 8347
rect 24225 8313 24259 8347
rect 26249 8313 26283 8347
rect 20361 8245 20395 8279
rect 28365 8245 28399 8279
rect 18521 8041 18555 8075
rect 22937 8041 22971 8075
rect 25881 8041 25915 8075
rect 26617 8041 26651 8075
rect 19257 7905 19291 7939
rect 20729 7905 20763 7939
rect 1409 7837 1443 7871
rect 18429 7837 18463 7871
rect 21557 7837 21591 7871
rect 21813 7837 21847 7871
rect 24639 7837 24673 7871
rect 24758 7837 24792 7871
rect 24874 7837 24908 7871
rect 25053 7837 25087 7871
rect 25513 7837 25547 7871
rect 26893 7837 26927 7871
rect 26985 7837 27019 7871
rect 27082 7837 27116 7871
rect 27261 7837 27295 7871
rect 46305 7837 46339 7871
rect 19441 7769 19475 7803
rect 23397 7769 23431 7803
rect 23581 7769 23615 7803
rect 23765 7769 23799 7803
rect 25697 7769 25731 7803
rect 46489 7769 46523 7803
rect 48145 7769 48179 7803
rect 1593 7701 1627 7735
rect 24409 7701 24443 7735
rect 18889 7497 18923 7531
rect 19441 7497 19475 7531
rect 24133 7497 24167 7531
rect 46765 7497 46799 7531
rect 23020 7429 23054 7463
rect 36645 7429 36679 7463
rect 37473 7429 37507 7463
rect 18797 7361 18831 7395
rect 19717 7361 19751 7395
rect 19809 7361 19843 7395
rect 19901 7361 19935 7395
rect 20085 7361 20119 7395
rect 22753 7361 22787 7395
rect 36553 7361 36587 7395
rect 37289 7361 37323 7395
rect 46673 7361 46707 7395
rect 47777 7361 47811 7395
rect 38025 7293 38059 7327
rect 2053 7157 2087 7191
rect 1409 6817 1443 6851
rect 2789 6817 2823 6851
rect 45845 6817 45879 6851
rect 22891 6749 22925 6783
rect 23010 6749 23044 6783
rect 23110 6749 23144 6783
rect 23305 6749 23339 6783
rect 1593 6681 1627 6715
rect 46029 6681 46063 6715
rect 47685 6681 47719 6715
rect 22661 6613 22695 6647
rect 2237 6409 2271 6443
rect 45937 6409 45971 6443
rect 2145 6273 2179 6307
rect 45845 6273 45879 6307
rect 47777 6069 47811 6103
rect 24685 5865 24719 5899
rect 25053 5865 25087 5899
rect 25513 5865 25547 5899
rect 46305 5729 46339 5763
rect 1777 5661 1811 5695
rect 2237 5661 2271 5695
rect 2973 5661 3007 5695
rect 25237 5661 25271 5695
rect 25329 5661 25363 5695
rect 25053 5593 25087 5627
rect 46489 5593 46523 5627
rect 48145 5593 48179 5627
rect 2329 5525 2363 5559
rect 3065 5525 3099 5559
rect 46949 5321 46983 5355
rect 2329 5253 2363 5287
rect 31493 5253 31527 5287
rect 32413 5253 32447 5287
rect 47961 5253 47995 5287
rect 2145 5185 2179 5219
rect 31401 5185 31435 5219
rect 46857 5185 46891 5219
rect 2789 5117 2823 5151
rect 32229 5117 32263 5151
rect 34069 5117 34103 5151
rect 48145 5049 48179 5083
rect 1685 4981 1719 5015
rect 1409 4641 1443 4675
rect 1593 4641 1627 4675
rect 2789 4641 2823 4675
rect 45201 4573 45235 4607
rect 45845 4573 45879 4607
rect 46305 4573 46339 4607
rect 46489 4505 46523 4539
rect 48145 4505 48179 4539
rect 2053 4097 2087 4131
rect 2697 4097 2731 4131
rect 4905 4097 4939 4131
rect 6745 4097 6779 4131
rect 7481 4097 7515 4131
rect 11897 4097 11931 4131
rect 12633 4097 12667 4131
rect 30757 4097 30791 4131
rect 32137 4097 32171 4131
rect 36185 4097 36219 4131
rect 38025 4097 38059 4131
rect 41705 4097 41739 4131
rect 45845 4097 45879 4131
rect 46857 4097 46891 4131
rect 46949 4097 46983 4131
rect 47869 4097 47903 4131
rect 38761 4029 38795 4063
rect 38945 4029 38979 4063
rect 39773 4029 39807 4063
rect 42441 4029 42475 4063
rect 42625 4029 42659 4063
rect 42901 4029 42935 4063
rect 32965 3961 32999 3995
rect 38117 3961 38151 3995
rect 41797 3961 41831 3995
rect 1593 3893 1627 3927
rect 2145 3893 2179 3927
rect 2789 3893 2823 3927
rect 3525 3893 3559 3927
rect 4445 3893 4479 3927
rect 4997 3893 5031 3927
rect 6837 3893 6871 3927
rect 7573 3893 7607 3927
rect 11989 3893 12023 3927
rect 12725 3893 12759 3927
rect 20177 3893 20211 3927
rect 29561 3893 29595 3927
rect 30205 3893 30239 3927
rect 30849 3893 30883 3927
rect 32229 3893 32263 3927
rect 36277 3893 36311 3927
rect 41245 3893 41279 3927
rect 45385 3893 45419 3927
rect 45937 3893 45971 3927
rect 48053 3893 48087 3927
rect 38945 3689 38979 3723
rect 1409 3553 1443 3587
rect 1593 3553 1627 3587
rect 1869 3553 1903 3587
rect 4445 3553 4479 3587
rect 5181 3553 5215 3587
rect 17233 3553 17267 3587
rect 19993 3553 20027 3587
rect 20637 3553 20671 3587
rect 31309 3553 31343 3587
rect 31585 3553 31619 3587
rect 36553 3553 36587 3587
rect 36829 3553 36863 3587
rect 41521 3553 41555 3587
rect 41981 3553 42015 3587
rect 46029 3553 46063 3587
rect 46213 3553 46247 3587
rect 46489 3553 46523 3587
rect 3801 3485 3835 3519
rect 8125 3485 8159 3519
rect 11805 3485 11839 3519
rect 12449 3485 12483 3519
rect 14565 3485 14599 3519
rect 15025 3485 15059 3519
rect 17693 3485 17727 3519
rect 23121 3485 23155 3519
rect 23581 3485 23615 3519
rect 25329 3485 25363 3519
rect 25973 3485 26007 3519
rect 27813 3485 27847 3519
rect 28733 3485 28767 3519
rect 29745 3485 29779 3519
rect 30665 3485 30699 3519
rect 31125 3485 31159 3519
rect 36369 3485 36403 3519
rect 39865 3485 39899 3519
rect 40877 3485 40911 3519
rect 43821 3485 43855 3519
rect 45017 3485 45051 3519
rect 4629 3417 4663 3451
rect 7297 3417 7331 3451
rect 7481 3417 7515 3451
rect 20177 3417 20211 3451
rect 25421 3417 25455 3451
rect 26157 3417 26191 3451
rect 40969 3417 41003 3451
rect 41705 3417 41739 3451
rect 3893 3349 3927 3383
rect 15117 3349 15151 3383
rect 17785 3349 17819 3383
rect 23673 3349 23707 3383
rect 28825 3349 28859 3383
rect 29837 3349 29871 3383
rect 39957 3349 39991 3383
rect 43913 3349 43947 3383
rect 45109 3349 45143 3383
rect 1961 3145 1995 3179
rect 20361 3145 20395 3179
rect 1869 3077 1903 3111
rect 3525 3077 3559 3111
rect 6837 3077 6871 3111
rect 12173 3077 12207 3111
rect 14473 3077 14507 3111
rect 17509 3077 17543 3111
rect 23397 3077 23431 3111
rect 29929 3077 29963 3111
rect 32321 3077 32355 3111
rect 40141 3077 40175 3111
rect 44189 3077 44223 3111
rect 2513 3009 2547 3043
rect 6653 3009 6687 3043
rect 8953 3009 8987 3043
rect 11989 3009 12023 3043
rect 14289 3009 14323 3043
rect 17325 3009 17359 3043
rect 20269 3009 20303 3043
rect 23213 3009 23247 3043
rect 26249 3009 26283 3043
rect 29745 3009 29779 3043
rect 32137 3009 32171 3043
rect 36553 3009 36587 3043
rect 42625 3009 42659 3043
rect 46397 3009 46431 3043
rect 46581 3009 46615 3043
rect 47869 3009 47903 3043
rect 3341 2941 3375 2975
rect 3801 2941 3835 2975
rect 7113 2941 7147 2975
rect 12909 2941 12943 2975
rect 15485 2941 15519 2975
rect 18061 2941 18095 2975
rect 23857 2941 23891 2975
rect 30297 2941 30331 2975
rect 33517 2941 33551 2975
rect 39957 2941 39991 2975
rect 41153 2941 41187 2975
rect 44005 2941 44039 2975
rect 44465 2941 44499 2975
rect 48053 2873 48087 2907
rect 2697 2805 2731 2839
rect 5825 2805 5859 2839
rect 9137 2805 9171 2839
rect 3985 2601 4019 2635
rect 10425 2601 10459 2635
rect 17785 2533 17819 2567
rect 23397 2533 23431 2567
rect 25881 2533 25915 2567
rect 35081 2533 35115 2567
rect 47961 2533 47995 2567
rect 1409 2465 1443 2499
rect 1869 2465 1903 2499
rect 6377 2465 6411 2499
rect 6561 2465 6595 2499
rect 6929 2465 6963 2499
rect 9229 2465 9263 2499
rect 11529 2465 11563 2499
rect 12265 2465 12299 2499
rect 14749 2465 14783 2499
rect 24869 2465 24903 2499
rect 28089 2465 28123 2499
rect 29561 2465 29595 2499
rect 29745 2465 29779 2499
rect 30941 2465 30975 2499
rect 38761 2465 38795 2499
rect 39957 2465 39991 2499
rect 44281 2465 44315 2499
rect 45017 2465 45051 2499
rect 45201 2465 45235 2499
rect 45569 2465 45603 2499
rect 4629 2397 4663 2431
rect 8953 2397 8987 2431
rect 20085 2397 20119 2431
rect 22661 2397 22695 2431
rect 23581 2397 23615 2431
rect 24593 2397 24627 2431
rect 26065 2397 26099 2431
rect 27077 2397 27111 2431
rect 27813 2397 27847 2431
rect 32965 2397 32999 2431
rect 34897 2397 34931 2431
rect 36369 2397 36403 2431
rect 38485 2397 38519 2431
rect 1593 2329 1627 2363
rect 10333 2329 10367 2363
rect 11713 2329 11747 2363
rect 14565 2329 14599 2363
rect 17601 2329 17635 2363
rect 33977 2329 34011 2363
rect 43361 2329 43395 2363
rect 47777 2329 47811 2363
rect 4813 2261 4847 2295
rect 20269 2261 20303 2295
rect 22845 2261 22879 2295
rect 27261 2261 27295 2295
rect 33149 2261 33183 2295
rect 34069 2261 34103 2295
rect 36185 2261 36219 2295
rect 43453 2261 43487 2295
<< metal1 >>
rect 1104 49530 48852 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 48852 49530
rect 1104 49456 48852 49478
rect 20438 49416 20444 49428
rect 14568 49388 20444 49416
rect 14182 49240 14188 49292
rect 14240 49280 14246 49292
rect 14568 49289 14596 49388
rect 20438 49376 20444 49388
rect 20496 49376 20502 49428
rect 24210 49348 24216 49360
rect 18156 49320 24216 49348
rect 14277 49283 14335 49289
rect 14277 49280 14289 49283
rect 14240 49252 14289 49280
rect 14240 49240 14246 49252
rect 14277 49249 14289 49252
rect 14323 49249 14335 49283
rect 14277 49243 14335 49249
rect 14553 49283 14611 49289
rect 14553 49249 14565 49283
rect 14599 49249 14611 49283
rect 14553 49243 14611 49249
rect 17865 49283 17923 49289
rect 17865 49249 17877 49283
rect 17911 49280 17923 49283
rect 18046 49280 18052 49292
rect 17911 49252 18052 49280
rect 17911 49249 17923 49252
rect 17865 49243 17923 49249
rect 18046 49240 18052 49252
rect 18104 49240 18110 49292
rect 18156 49289 18184 49320
rect 24210 49308 24216 49320
rect 24268 49308 24274 49360
rect 28997 49351 29055 49357
rect 28997 49317 29009 49351
rect 29043 49348 29055 49351
rect 29086 49348 29092 49360
rect 29043 49320 29092 49348
rect 29043 49317 29055 49320
rect 28997 49311 29055 49317
rect 29086 49308 29092 49320
rect 29144 49308 29150 49360
rect 46198 49348 46204 49360
rect 42812 49320 46204 49348
rect 18141 49283 18199 49289
rect 18141 49249 18153 49283
rect 18187 49249 18199 49283
rect 21358 49280 21364 49292
rect 18141 49243 18199 49249
rect 19260 49252 21364 49280
rect 658 49172 664 49224
rect 716 49212 722 49224
rect 1857 49215 1915 49221
rect 1857 49212 1869 49215
rect 716 49184 1869 49212
rect 716 49172 722 49184
rect 1857 49181 1869 49184
rect 1903 49181 1915 49215
rect 1857 49175 1915 49181
rect 3602 49172 3608 49224
rect 3660 49212 3666 49224
rect 4249 49215 4307 49221
rect 4249 49212 4261 49215
rect 3660 49184 4261 49212
rect 3660 49172 3666 49184
rect 4249 49181 4261 49184
rect 4295 49181 4307 49215
rect 4249 49175 4307 49181
rect 4890 49172 4896 49224
rect 4948 49212 4954 49224
rect 5077 49215 5135 49221
rect 5077 49212 5089 49215
rect 4948 49184 5089 49212
rect 4948 49172 4954 49184
rect 5077 49181 5089 49184
rect 5123 49181 5135 49215
rect 5077 49175 5135 49181
rect 6454 49172 6460 49224
rect 6512 49212 6518 49224
rect 6825 49215 6883 49221
rect 6825 49212 6837 49215
rect 6512 49184 6837 49212
rect 6512 49172 6518 49184
rect 6825 49181 6837 49184
rect 6871 49181 6883 49215
rect 6825 49175 6883 49181
rect 7098 49172 7104 49224
rect 7156 49212 7162 49224
rect 7653 49215 7711 49221
rect 7653 49212 7665 49215
rect 7156 49184 7665 49212
rect 7156 49172 7162 49184
rect 7653 49181 7665 49184
rect 7699 49181 7711 49215
rect 10318 49212 10324 49224
rect 10279 49184 10324 49212
rect 7653 49175 7711 49181
rect 10318 49172 10324 49184
rect 10376 49172 10382 49224
rect 10965 49215 11023 49221
rect 10965 49181 10977 49215
rect 11011 49212 11023 49215
rect 11514 49212 11520 49224
rect 11011 49184 11520 49212
rect 11011 49181 11023 49184
rect 10965 49175 11023 49181
rect 11514 49172 11520 49184
rect 11572 49172 11578 49224
rect 11606 49172 11612 49224
rect 11664 49212 11670 49224
rect 11977 49215 12035 49221
rect 11977 49212 11989 49215
rect 11664 49184 11989 49212
rect 11664 49172 11670 49184
rect 11977 49181 11989 49184
rect 12023 49181 12035 49215
rect 13262 49212 13268 49224
rect 13223 49184 13268 49212
rect 11977 49175 12035 49181
rect 13262 49172 13268 49184
rect 13320 49172 13326 49224
rect 16117 49215 16175 49221
rect 16117 49181 16129 49215
rect 16163 49212 16175 49215
rect 16574 49212 16580 49224
rect 16163 49184 16580 49212
rect 16163 49181 16175 49184
rect 16117 49175 16175 49181
rect 16574 49172 16580 49184
rect 16632 49172 16638 49224
rect 16666 49172 16672 49224
rect 16724 49212 16730 49224
rect 17129 49215 17187 49221
rect 17129 49212 17141 49215
rect 16724 49184 17141 49212
rect 16724 49172 16730 49184
rect 17129 49181 17141 49184
rect 17175 49181 17187 49215
rect 17129 49175 17187 49181
rect 17313 49215 17371 49221
rect 17313 49181 17325 49215
rect 17359 49212 17371 49215
rect 19260 49212 19288 49252
rect 21358 49240 21364 49252
rect 21416 49240 21422 49292
rect 22005 49283 22063 49289
rect 22005 49249 22017 49283
rect 22051 49280 22063 49283
rect 22370 49280 22376 49292
rect 22051 49252 22376 49280
rect 22051 49249 22063 49252
rect 22005 49243 22063 49249
rect 22370 49240 22376 49252
rect 22428 49240 22434 49292
rect 22554 49280 22560 49292
rect 22515 49252 22560 49280
rect 22554 49240 22560 49252
rect 22612 49240 22618 49292
rect 24762 49240 24768 49292
rect 24820 49280 24826 49292
rect 24857 49283 24915 49289
rect 24857 49280 24869 49283
rect 24820 49252 24869 49280
rect 24820 49240 24826 49252
rect 24857 49249 24869 49252
rect 24903 49249 24915 49283
rect 24857 49243 24915 49249
rect 29733 49283 29791 49289
rect 29733 49249 29745 49283
rect 29779 49280 29791 49283
rect 30650 49280 30656 49292
rect 29779 49252 30656 49280
rect 29779 49249 29791 49252
rect 29733 49243 29791 49249
rect 30650 49240 30656 49252
rect 30708 49240 30714 49292
rect 30926 49280 30932 49292
rect 30887 49252 30932 49280
rect 30926 49240 30932 49252
rect 30984 49240 30990 49292
rect 40678 49280 40684 49292
rect 40639 49252 40684 49280
rect 40678 49240 40684 49252
rect 40736 49240 40742 49292
rect 42812 49289 42840 49320
rect 46198 49308 46204 49320
rect 46256 49308 46262 49360
rect 42797 49283 42855 49289
rect 42797 49249 42809 49283
rect 42843 49249 42855 49283
rect 42797 49243 42855 49249
rect 44453 49283 44511 49289
rect 44453 49249 44465 49283
rect 44499 49280 44511 49283
rect 46658 49280 46664 49292
rect 44499 49252 46664 49280
rect 44499 49249 44511 49252
rect 44453 49243 44511 49249
rect 46658 49240 46664 49252
rect 46716 49240 46722 49292
rect 46842 49280 46848 49292
rect 46803 49252 46848 49280
rect 46842 49240 46848 49252
rect 46900 49240 46906 49292
rect 19426 49212 19432 49224
rect 17359 49184 19288 49212
rect 19387 49184 19432 49212
rect 17359 49181 17371 49184
rect 17313 49175 17371 49181
rect 19426 49172 19432 49184
rect 19484 49172 19490 49224
rect 20070 49212 20076 49224
rect 20031 49184 20076 49212
rect 20070 49172 20076 49184
rect 20128 49172 20134 49224
rect 20990 49212 20996 49224
rect 20951 49184 20996 49212
rect 20990 49172 20996 49184
rect 21048 49172 21054 49224
rect 24397 49215 24455 49221
rect 24397 49181 24409 49215
rect 24443 49181 24455 49215
rect 24397 49175 24455 49181
rect 2774 49144 2780 49156
rect 2735 49116 2780 49144
rect 2774 49104 2780 49116
rect 2832 49104 2838 49156
rect 2958 49144 2964 49156
rect 2919 49116 2964 49144
rect 2958 49104 2964 49116
rect 3016 49104 3022 49156
rect 4617 49147 4675 49153
rect 4617 49113 4629 49147
rect 4663 49144 4675 49147
rect 4706 49144 4712 49156
rect 4663 49116 4712 49144
rect 4663 49113 4675 49116
rect 4617 49107 4675 49113
rect 4706 49104 4712 49116
rect 4764 49104 4770 49156
rect 19613 49147 19671 49153
rect 19613 49113 19625 49147
rect 19659 49144 19671 49147
rect 21082 49144 21088 49156
rect 19659 49116 21088 49144
rect 19659 49113 19671 49116
rect 19613 49107 19671 49113
rect 21082 49104 21088 49116
rect 21140 49104 21146 49156
rect 22186 49144 22192 49156
rect 22147 49116 22192 49144
rect 22186 49104 22192 49116
rect 22244 49104 22250 49156
rect 1762 49036 1768 49088
rect 1820 49076 1826 49088
rect 1949 49079 2007 49085
rect 1949 49076 1961 49079
rect 1820 49048 1961 49076
rect 1820 49036 1826 49048
rect 1949 49045 1961 49048
rect 1995 49045 2007 49079
rect 5258 49076 5264 49088
rect 5219 49048 5264 49076
rect 1949 49039 2007 49045
rect 5258 49036 5264 49048
rect 5316 49036 5322 49088
rect 6454 49036 6460 49088
rect 6512 49076 6518 49088
rect 6917 49079 6975 49085
rect 6917 49076 6929 49079
rect 6512 49048 6929 49076
rect 6512 49036 6518 49048
rect 6917 49045 6929 49048
rect 6963 49045 6975 49079
rect 8938 49076 8944 49088
rect 8899 49048 8944 49076
rect 6917 49039 6975 49045
rect 8938 49036 8944 49048
rect 8996 49036 9002 49088
rect 11882 49036 11888 49088
rect 11940 49076 11946 49088
rect 12069 49079 12127 49085
rect 12069 49076 12081 49079
rect 11940 49048 12081 49076
rect 11940 49036 11946 49048
rect 12069 49045 12081 49048
rect 12115 49045 12127 49079
rect 13446 49076 13452 49088
rect 13407 49048 13452 49076
rect 12069 49039 12127 49045
rect 13446 49036 13452 49048
rect 13504 49036 13510 49088
rect 20257 49079 20315 49085
rect 20257 49045 20269 49079
rect 20303 49076 20315 49079
rect 20530 49076 20536 49088
rect 20303 49048 20536 49076
rect 20303 49045 20315 49048
rect 20257 49039 20315 49045
rect 20530 49036 20536 49048
rect 20588 49036 20594 49088
rect 24412 49076 24440 49175
rect 26418 49172 26424 49224
rect 26476 49212 26482 49224
rect 27433 49215 27491 49221
rect 27433 49212 27445 49215
rect 26476 49184 27445 49212
rect 26476 49172 26482 49184
rect 27433 49181 27445 49184
rect 27479 49181 27491 49215
rect 27433 49175 27491 49181
rect 27617 49215 27675 49221
rect 27617 49181 27629 49215
rect 27663 49212 27675 49215
rect 27982 49212 27988 49224
rect 27663 49184 27988 49212
rect 27663 49181 27675 49184
rect 27617 49175 27675 49181
rect 27982 49172 27988 49184
rect 28040 49172 28046 49224
rect 28261 49215 28319 49221
rect 28261 49181 28273 49215
rect 28307 49181 28319 49215
rect 28261 49175 28319 49181
rect 28813 49215 28871 49221
rect 28813 49181 28825 49215
rect 28859 49212 28871 49215
rect 28994 49212 29000 49224
rect 28859 49184 29000 49212
rect 28859 49181 28871 49184
rect 28813 49175 28871 49181
rect 24578 49144 24584 49156
rect 24539 49116 24584 49144
rect 24578 49104 24584 49116
rect 24636 49104 24642 49156
rect 27338 49104 27344 49156
rect 27396 49144 27402 49156
rect 28276 49144 28304 49175
rect 28994 49172 29000 49184
rect 29052 49172 29058 49224
rect 33318 49172 33324 49224
rect 33376 49212 33382 49224
rect 33597 49215 33655 49221
rect 33597 49212 33609 49215
rect 33376 49184 33609 49212
rect 33376 49172 33382 49184
rect 33597 49181 33609 49184
rect 33643 49181 33655 49215
rect 35802 49212 35808 49224
rect 35763 49184 35808 49212
rect 33597 49175 33655 49181
rect 35802 49172 35808 49184
rect 35860 49172 35866 49224
rect 36449 49215 36507 49221
rect 36449 49181 36461 49215
rect 36495 49181 36507 49215
rect 38194 49212 38200 49224
rect 38155 49184 38200 49212
rect 36449 49175 36507 49181
rect 29914 49144 29920 49156
rect 27396 49116 28304 49144
rect 29875 49116 29920 49144
rect 27396 49104 27402 49116
rect 29914 49104 29920 49116
rect 29972 49104 29978 49156
rect 30024 49116 32444 49144
rect 25222 49076 25228 49088
rect 24412 49048 25228 49076
rect 25222 49036 25228 49048
rect 25280 49036 25286 49088
rect 25314 49036 25320 49088
rect 25372 49076 25378 49088
rect 26602 49076 26608 49088
rect 25372 49048 26608 49076
rect 25372 49036 25378 49048
rect 26602 49036 26608 49048
rect 26660 49076 26666 49088
rect 27522 49076 27528 49088
rect 26660 49048 27528 49076
rect 26660 49036 26666 49048
rect 27522 49036 27528 49048
rect 27580 49036 27586 49088
rect 29638 49036 29644 49088
rect 29696 49076 29702 49088
rect 30024 49076 30052 49116
rect 32122 49076 32128 49088
rect 29696 49048 30052 49076
rect 32083 49048 32128 49076
rect 29696 49036 29702 49048
rect 32122 49036 32128 49048
rect 32180 49036 32186 49088
rect 32416 49076 32444 49116
rect 34882 49104 34888 49156
rect 34940 49144 34946 49156
rect 36464 49144 36492 49175
rect 38194 49172 38200 49184
rect 38252 49172 38258 49224
rect 39298 49172 39304 49224
rect 39356 49212 39362 49224
rect 40957 49215 41015 49221
rect 40957 49212 40969 49215
rect 39356 49184 40969 49212
rect 39356 49172 39362 49184
rect 40957 49181 40969 49184
rect 41003 49181 41015 49215
rect 40957 49175 41015 49181
rect 42334 49172 42340 49224
rect 42392 49212 42398 49224
rect 42613 49215 42671 49221
rect 42613 49212 42625 49215
rect 42392 49184 42625 49212
rect 42392 49172 42398 49184
rect 42613 49181 42625 49184
rect 42659 49181 42671 49215
rect 42613 49175 42671 49181
rect 44082 49172 44088 49224
rect 44140 49212 44146 49224
rect 45189 49215 45247 49221
rect 45189 49212 45201 49215
rect 44140 49184 45201 49212
rect 44140 49172 44146 49184
rect 45189 49181 45201 49184
rect 45235 49181 45247 49215
rect 47762 49212 47768 49224
rect 47723 49184 47768 49212
rect 45189 49175 45247 49181
rect 47762 49172 47768 49184
rect 47820 49172 47826 49224
rect 34940 49116 36492 49144
rect 37936 49116 38424 49144
rect 34940 49104 34946 49116
rect 37936 49076 37964 49116
rect 32416 49048 37964 49076
rect 38010 49036 38016 49088
rect 38068 49076 38074 49088
rect 38289 49079 38347 49085
rect 38289 49076 38301 49079
rect 38068 49048 38301 49076
rect 38068 49036 38074 49048
rect 38289 49045 38301 49048
rect 38335 49045 38347 49079
rect 38396 49076 38424 49116
rect 44634 49104 44640 49156
rect 44692 49144 44698 49156
rect 45373 49147 45431 49153
rect 45373 49144 45385 49147
rect 44692 49116 45385 49144
rect 44692 49104 44698 49116
rect 45373 49113 45385 49116
rect 45419 49113 45431 49147
rect 45373 49107 45431 49113
rect 47857 49079 47915 49085
rect 47857 49076 47869 49079
rect 38396 49048 47869 49076
rect 38289 49039 38347 49045
rect 47857 49045 47869 49048
rect 47903 49045 47915 49079
rect 47857 49039 47915 49045
rect 1104 48986 48852 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 48852 48986
rect 1104 48912 48852 48934
rect 25314 48872 25320 48884
rect 19260 48844 25320 48872
rect 1946 48764 1952 48816
rect 2004 48804 2010 48816
rect 2004 48776 4384 48804
rect 2004 48764 2010 48776
rect 1397 48739 1455 48745
rect 1397 48705 1409 48739
rect 1443 48736 1455 48739
rect 1670 48736 1676 48748
rect 1443 48708 1676 48736
rect 1443 48705 1455 48708
rect 1397 48699 1455 48705
rect 1670 48696 1676 48708
rect 1728 48696 1734 48748
rect 4356 48745 4384 48776
rect 4341 48739 4399 48745
rect 4341 48705 4353 48739
rect 4387 48705 4399 48739
rect 8938 48736 8944 48748
rect 8899 48708 8944 48736
rect 4341 48699 4399 48705
rect 8938 48696 8944 48708
rect 8996 48696 9002 48748
rect 11514 48736 11520 48748
rect 11475 48708 11520 48736
rect 11514 48696 11520 48708
rect 11572 48696 11578 48748
rect 19260 48745 19288 48844
rect 25314 48832 25320 48844
rect 25372 48832 25378 48884
rect 39666 48832 39672 48884
rect 39724 48872 39730 48884
rect 47857 48875 47915 48881
rect 47857 48872 47869 48875
rect 39724 48844 47869 48872
rect 39724 48832 39730 48844
rect 47857 48841 47869 48844
rect 47903 48841 47915 48875
rect 47857 48835 47915 48841
rect 22002 48804 22008 48816
rect 21963 48776 22008 48804
rect 22002 48764 22008 48776
rect 22060 48764 22066 48816
rect 25958 48804 25964 48816
rect 25919 48776 25964 48804
rect 25958 48764 25964 48776
rect 26016 48764 26022 48816
rect 27522 48764 27528 48816
rect 27580 48804 27586 48816
rect 47762 48804 47768 48816
rect 27580 48776 29684 48804
rect 47723 48776 47768 48804
rect 27580 48764 27586 48776
rect 19245 48739 19303 48745
rect 19245 48705 19257 48739
rect 19291 48705 19303 48739
rect 27338 48736 27344 48748
rect 27299 48708 27344 48736
rect 19245 48699 19303 48705
rect 27338 48696 27344 48708
rect 27396 48696 27402 48748
rect 29656 48745 29684 48776
rect 47762 48764 47768 48776
rect 47820 48764 47826 48816
rect 29641 48739 29699 48745
rect 29641 48705 29653 48739
rect 29687 48705 29699 48739
rect 32122 48736 32128 48748
rect 32083 48708 32128 48736
rect 29641 48699 29699 48705
rect 32122 48696 32128 48708
rect 32180 48696 32186 48748
rect 34882 48736 34888 48748
rect 34843 48708 34888 48736
rect 34882 48696 34888 48708
rect 34940 48696 34946 48748
rect 2041 48671 2099 48677
rect 2041 48637 2053 48671
rect 2087 48637 2099 48671
rect 2222 48668 2228 48680
rect 2183 48640 2228 48668
rect 2041 48631 2099 48637
rect 2056 48600 2084 48631
rect 2222 48628 2228 48640
rect 2280 48628 2286 48680
rect 2866 48668 2872 48680
rect 2827 48640 2872 48668
rect 2866 48628 2872 48640
rect 2924 48628 2930 48680
rect 6365 48671 6423 48677
rect 6365 48637 6377 48671
rect 6411 48637 6423 48671
rect 6546 48668 6552 48680
rect 6507 48640 6552 48668
rect 6365 48631 6423 48637
rect 5261 48603 5319 48609
rect 5261 48600 5273 48603
rect 2056 48572 5273 48600
rect 5261 48569 5273 48572
rect 5307 48569 5319 48603
rect 6380 48600 6408 48631
rect 6546 48628 6552 48640
rect 6604 48628 6610 48680
rect 7190 48668 7196 48680
rect 7151 48640 7196 48668
rect 7190 48628 7196 48640
rect 7248 48628 7254 48680
rect 9122 48668 9128 48680
rect 9083 48640 9128 48668
rect 9122 48628 9128 48640
rect 9180 48628 9186 48680
rect 9674 48668 9680 48680
rect 9635 48640 9680 48668
rect 9674 48628 9680 48640
rect 9732 48628 9738 48680
rect 11698 48668 11704 48680
rect 11659 48640 11704 48668
rect 11698 48628 11704 48640
rect 11756 48628 11762 48680
rect 12434 48628 12440 48680
rect 12492 48668 12498 48680
rect 14182 48668 14188 48680
rect 12492 48640 12537 48668
rect 14143 48640 14188 48668
rect 12492 48628 12498 48640
rect 14182 48628 14188 48640
rect 14240 48628 14246 48680
rect 14366 48668 14372 48680
rect 14327 48640 14372 48668
rect 14366 48628 14372 48640
rect 14424 48628 14430 48680
rect 15194 48668 15200 48680
rect 15155 48640 15200 48668
rect 15194 48628 15200 48640
rect 15252 48628 15258 48680
rect 16942 48668 16948 48680
rect 16903 48640 16948 48668
rect 16942 48628 16948 48640
rect 17000 48628 17006 48680
rect 17129 48671 17187 48677
rect 17129 48637 17141 48671
rect 17175 48637 17187 48671
rect 17129 48631 17187 48637
rect 7558 48600 7564 48612
rect 6380 48572 7564 48600
rect 5261 48563 5319 48569
rect 7558 48560 7564 48572
rect 7616 48560 7622 48612
rect 17144 48600 17172 48631
rect 17218 48628 17224 48680
rect 17276 48668 17282 48680
rect 17405 48671 17463 48677
rect 17405 48668 17417 48671
rect 17276 48640 17417 48668
rect 17276 48628 17282 48640
rect 17405 48637 17417 48640
rect 17451 48637 17463 48671
rect 19426 48668 19432 48680
rect 19387 48640 19432 48668
rect 17405 48631 17463 48637
rect 19426 48628 19432 48640
rect 19484 48628 19490 48680
rect 19705 48671 19763 48677
rect 19705 48637 19717 48671
rect 19751 48637 19763 48671
rect 22646 48668 22652 48680
rect 22607 48640 22652 48668
rect 19705 48631 19763 48637
rect 19334 48600 19340 48612
rect 17144 48572 19340 48600
rect 19334 48560 19340 48572
rect 19392 48560 19398 48612
rect 1489 48535 1547 48541
rect 1489 48501 1501 48535
rect 1535 48532 1547 48535
rect 2130 48532 2136 48544
rect 1535 48504 2136 48532
rect 1535 48501 1547 48504
rect 1489 48495 1547 48501
rect 2130 48492 2136 48504
rect 2188 48492 2194 48544
rect 4525 48535 4583 48541
rect 4525 48501 4537 48535
rect 4571 48532 4583 48535
rect 4614 48532 4620 48544
rect 4571 48504 4620 48532
rect 4571 48501 4583 48504
rect 4525 48495 4583 48501
rect 4614 48492 4620 48504
rect 4672 48492 4678 48544
rect 9030 48492 9036 48544
rect 9088 48532 9094 48544
rect 15102 48532 15108 48544
rect 9088 48504 15108 48532
rect 9088 48492 9094 48504
rect 15102 48492 15108 48504
rect 15160 48492 15166 48544
rect 17954 48492 17960 48544
rect 18012 48532 18018 48544
rect 19720 48532 19748 48631
rect 22646 48628 22652 48640
rect 22704 48628 22710 48680
rect 22830 48668 22836 48680
rect 22791 48640 22836 48668
rect 22830 48628 22836 48640
rect 22888 48628 22894 48680
rect 23474 48668 23480 48680
rect 23435 48640 23480 48668
rect 23474 48628 23480 48640
rect 23532 48628 23538 48680
rect 27525 48671 27583 48677
rect 27525 48637 27537 48671
rect 27571 48668 27583 48671
rect 28718 48668 28724 48680
rect 27571 48640 28724 48668
rect 27571 48637 27583 48640
rect 27525 48631 27583 48637
rect 28718 48628 28724 48640
rect 28776 48628 28782 48680
rect 28813 48671 28871 48677
rect 28813 48637 28825 48671
rect 28859 48637 28871 48671
rect 29822 48668 29828 48680
rect 29783 48640 29828 48668
rect 28813 48631 28871 48637
rect 25409 48603 25467 48609
rect 25409 48569 25421 48603
rect 25455 48600 25467 48603
rect 27614 48600 27620 48612
rect 25455 48572 27620 48600
rect 25455 48569 25467 48572
rect 25409 48563 25467 48569
rect 27614 48560 27620 48572
rect 27672 48560 27678 48612
rect 27706 48560 27712 48612
rect 27764 48600 27770 48612
rect 28828 48600 28856 48631
rect 29822 48628 29828 48640
rect 29880 48628 29886 48680
rect 30006 48628 30012 48680
rect 30064 48668 30070 48680
rect 30101 48671 30159 48677
rect 30101 48668 30113 48671
rect 30064 48640 30113 48668
rect 30064 48628 30070 48640
rect 30101 48637 30113 48640
rect 30147 48637 30159 48671
rect 32306 48668 32312 48680
rect 32267 48640 32312 48668
rect 30101 48631 30159 48637
rect 32306 48628 32312 48640
rect 32364 48628 32370 48680
rect 33134 48668 33140 48680
rect 33095 48640 33140 48668
rect 33134 48628 33140 48640
rect 33192 48628 33198 48680
rect 35069 48671 35127 48677
rect 35069 48637 35081 48671
rect 35115 48668 35127 48671
rect 35894 48668 35900 48680
rect 35115 48640 35900 48668
rect 35115 48637 35127 48640
rect 35069 48631 35127 48637
rect 35894 48628 35900 48640
rect 35952 48628 35958 48680
rect 36078 48668 36084 48680
rect 36039 48640 36084 48668
rect 36078 48628 36084 48640
rect 36136 48628 36142 48680
rect 39117 48671 39175 48677
rect 39117 48637 39129 48671
rect 39163 48668 39175 48671
rect 39577 48671 39635 48677
rect 39577 48668 39589 48671
rect 39163 48640 39589 48668
rect 39163 48637 39175 48640
rect 39117 48631 39175 48637
rect 39577 48637 39589 48640
rect 39623 48637 39635 48671
rect 39758 48668 39764 48680
rect 39719 48640 39764 48668
rect 39577 48631 39635 48637
rect 39758 48628 39764 48640
rect 39816 48628 39822 48680
rect 40034 48668 40040 48680
rect 39995 48640 40040 48668
rect 40034 48628 40040 48640
rect 40092 48628 40098 48680
rect 42426 48668 42432 48680
rect 42387 48640 42432 48668
rect 42426 48628 42432 48640
rect 42484 48628 42490 48680
rect 42610 48668 42616 48680
rect 42571 48640 42616 48668
rect 42610 48628 42616 48640
rect 42668 48628 42674 48680
rect 42794 48628 42800 48680
rect 42852 48668 42858 48680
rect 42889 48671 42947 48677
rect 42889 48668 42901 48671
rect 42852 48640 42901 48668
rect 42852 48628 42858 48640
rect 42889 48637 42901 48640
rect 42935 48637 42947 48671
rect 42889 48631 42947 48637
rect 45189 48671 45247 48677
rect 45189 48637 45201 48671
rect 45235 48637 45247 48671
rect 45370 48668 45376 48680
rect 45331 48640 45376 48668
rect 45189 48631 45247 48637
rect 27764 48572 28856 48600
rect 27764 48560 27770 48572
rect 33410 48560 33416 48612
rect 33468 48600 33474 48612
rect 33870 48600 33876 48612
rect 33468 48572 33876 48600
rect 33468 48560 33474 48572
rect 33870 48560 33876 48572
rect 33928 48560 33934 48612
rect 45204 48600 45232 48631
rect 45370 48628 45376 48640
rect 45428 48628 45434 48680
rect 45738 48668 45744 48680
rect 45699 48640 45744 48668
rect 45738 48628 45744 48640
rect 45796 48628 45802 48680
rect 45462 48600 45468 48612
rect 45204 48572 45468 48600
rect 45462 48560 45468 48572
rect 45520 48560 45526 48612
rect 22094 48532 22100 48544
rect 18012 48504 19748 48532
rect 22055 48504 22100 48532
rect 18012 48492 18018 48504
rect 22094 48492 22100 48504
rect 22152 48492 22158 48544
rect 24946 48492 24952 48544
rect 25004 48532 25010 48544
rect 26053 48535 26111 48541
rect 26053 48532 26065 48535
rect 25004 48504 26065 48532
rect 25004 48492 25010 48504
rect 26053 48501 26065 48504
rect 26099 48501 26111 48535
rect 26053 48495 26111 48501
rect 1104 48442 48852 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 48852 48442
rect 1104 48368 48852 48390
rect 3418 48288 3424 48340
rect 3476 48328 3482 48340
rect 9030 48328 9036 48340
rect 3476 48300 9036 48328
rect 3476 48288 3482 48300
rect 9030 48288 9036 48300
rect 9088 48288 9094 48340
rect 9122 48288 9128 48340
rect 9180 48328 9186 48340
rect 9401 48331 9459 48337
rect 9401 48328 9413 48331
rect 9180 48300 9413 48328
rect 9180 48288 9186 48300
rect 9401 48297 9413 48300
rect 9447 48297 9459 48331
rect 9401 48291 9459 48297
rect 14366 48288 14372 48340
rect 14424 48328 14430 48340
rect 14553 48331 14611 48337
rect 14553 48328 14565 48331
rect 14424 48300 14565 48328
rect 14424 48288 14430 48300
rect 14553 48297 14565 48300
rect 14599 48297 14611 48331
rect 14553 48291 14611 48297
rect 16206 48288 16212 48340
rect 16264 48328 16270 48340
rect 39666 48328 39672 48340
rect 16264 48300 39672 48328
rect 16264 48288 16270 48300
rect 39666 48288 39672 48300
rect 39724 48288 39730 48340
rect 39758 48288 39764 48340
rect 39816 48328 39822 48340
rect 39945 48331 40003 48337
rect 39945 48328 39957 48331
rect 39816 48300 39957 48328
rect 39816 48288 39822 48300
rect 39945 48297 39957 48300
rect 39991 48297 40003 48331
rect 39945 48291 40003 48297
rect 14 48220 20 48272
rect 72 48260 78 48272
rect 2774 48260 2780 48272
rect 72 48232 2780 48260
rect 72 48220 78 48232
rect 2774 48220 2780 48232
rect 2832 48220 2838 48272
rect 7558 48260 7564 48272
rect 7519 48232 7564 48260
rect 7558 48220 7564 48232
rect 7616 48220 7622 48272
rect 16117 48263 16175 48269
rect 9324 48232 15976 48260
rect 1581 48195 1639 48201
rect 1581 48161 1593 48195
rect 1627 48192 1639 48195
rect 3881 48195 3939 48201
rect 3881 48192 3893 48195
rect 1627 48164 3893 48192
rect 1627 48161 1639 48164
rect 1581 48155 1639 48161
rect 3881 48161 3893 48164
rect 3927 48161 3939 48195
rect 3881 48155 3939 48161
rect 4062 48152 4068 48204
rect 4120 48192 4126 48204
rect 4893 48195 4951 48201
rect 4893 48192 4905 48195
rect 4120 48164 4905 48192
rect 4120 48152 4126 48164
rect 4893 48161 4905 48164
rect 4939 48161 4951 48195
rect 4893 48155 4951 48161
rect 1397 48127 1455 48133
rect 1397 48093 1409 48127
rect 1443 48093 1455 48127
rect 1397 48087 1455 48093
rect 1412 48056 1440 48087
rect 3602 48084 3608 48136
rect 3660 48124 3666 48136
rect 3789 48127 3847 48133
rect 3789 48124 3801 48127
rect 3660 48096 3801 48124
rect 3660 48084 3666 48096
rect 3789 48093 3801 48096
rect 3835 48093 3847 48127
rect 4430 48124 4436 48136
rect 4391 48096 4436 48124
rect 3789 48087 3847 48093
rect 4430 48084 4436 48096
rect 4488 48084 4494 48136
rect 9324 48133 9352 48232
rect 10318 48152 10324 48204
rect 10376 48192 10382 48204
rect 10505 48195 10563 48201
rect 10505 48192 10517 48195
rect 10376 48164 10517 48192
rect 10376 48152 10382 48164
rect 10505 48161 10517 48164
rect 10551 48161 10563 48195
rect 10505 48155 10563 48161
rect 10686 48152 10692 48204
rect 10744 48192 10750 48204
rect 11057 48195 11115 48201
rect 11057 48192 11069 48195
rect 10744 48164 11069 48192
rect 10744 48152 10750 48164
rect 11057 48161 11069 48164
rect 11103 48161 11115 48195
rect 11057 48155 11115 48161
rect 6917 48127 6975 48133
rect 6917 48093 6929 48127
rect 6963 48093 6975 48127
rect 6917 48087 6975 48093
rect 9309 48127 9367 48133
rect 9309 48093 9321 48127
rect 9355 48093 9367 48127
rect 12894 48124 12900 48136
rect 12855 48096 12900 48124
rect 9309 48087 9367 48093
rect 3142 48056 3148 48068
rect 1412 48028 3148 48056
rect 3142 48016 3148 48028
rect 3200 48016 3206 48068
rect 3234 48016 3240 48068
rect 3292 48056 3298 48068
rect 4617 48059 4675 48065
rect 3292 48028 3337 48056
rect 3292 48016 3298 48028
rect 4617 48025 4629 48059
rect 4663 48056 4675 48059
rect 5350 48056 5356 48068
rect 4663 48028 5356 48056
rect 4663 48025 4675 48028
rect 4617 48019 4675 48025
rect 5350 48016 5356 48028
rect 5408 48016 5414 48068
rect 1946 47948 1952 48000
rect 2004 47988 2010 48000
rect 6932 47988 6960 48087
rect 12894 48084 12900 48096
rect 12952 48084 12958 48136
rect 14458 48124 14464 48136
rect 14419 48096 14464 48124
rect 14458 48084 14464 48096
rect 14516 48084 14522 48136
rect 10689 48059 10747 48065
rect 10689 48025 10701 48059
rect 10735 48056 10747 48059
rect 11606 48056 11612 48068
rect 10735 48028 11612 48056
rect 10735 48025 10747 48028
rect 10689 48019 10747 48025
rect 11606 48016 11612 48028
rect 11664 48016 11670 48068
rect 13081 48059 13139 48065
rect 13081 48025 13093 48059
rect 13127 48056 13139 48059
rect 13722 48056 13728 48068
rect 13127 48028 13728 48056
rect 13127 48025 13139 48028
rect 13081 48019 13139 48025
rect 13722 48016 13728 48028
rect 13780 48016 13786 48068
rect 2004 47960 6960 47988
rect 2004 47948 2010 47960
rect 10962 47948 10968 48000
rect 11020 47988 11026 48000
rect 13354 47988 13360 48000
rect 11020 47960 13360 47988
rect 11020 47948 11026 47960
rect 13354 47948 13360 47960
rect 13412 47948 13418 48000
rect 15948 47988 15976 48232
rect 16117 48229 16129 48263
rect 16163 48260 16175 48263
rect 16942 48260 16948 48272
rect 16163 48232 16948 48260
rect 16163 48229 16175 48232
rect 16117 48223 16175 48229
rect 16942 48220 16948 48232
rect 17000 48220 17006 48272
rect 19334 48260 19340 48272
rect 19295 48232 19340 48260
rect 19334 48220 19340 48232
rect 19392 48220 19398 48272
rect 20990 48260 20996 48272
rect 20272 48232 20996 48260
rect 16574 48192 16580 48204
rect 16535 48164 16580 48192
rect 16574 48152 16580 48164
rect 16632 48152 16638 48204
rect 17402 48192 17408 48204
rect 17363 48164 17408 48192
rect 17402 48152 17408 48164
rect 17460 48152 17466 48204
rect 20272 48201 20300 48232
rect 20990 48220 20996 48232
rect 21048 48220 21054 48272
rect 22649 48263 22707 48269
rect 22649 48229 22661 48263
rect 22695 48260 22707 48263
rect 22830 48260 22836 48272
rect 22695 48232 22836 48260
rect 22695 48229 22707 48232
rect 22649 48223 22707 48229
rect 22830 48220 22836 48232
rect 22888 48220 22894 48272
rect 24489 48263 24547 48269
rect 24489 48229 24501 48263
rect 24535 48260 24547 48263
rect 24578 48260 24584 48272
rect 24535 48232 24584 48260
rect 24535 48229 24547 48232
rect 24489 48223 24547 48229
rect 24578 48220 24584 48232
rect 24636 48220 24642 48272
rect 25222 48260 25228 48272
rect 25183 48232 25228 48260
rect 25222 48220 25228 48232
rect 25280 48220 25286 48272
rect 25332 48232 28672 48260
rect 20257 48195 20315 48201
rect 20257 48161 20269 48195
rect 20303 48161 20315 48195
rect 20257 48155 20315 48161
rect 20622 48152 20628 48204
rect 20680 48192 20686 48204
rect 20717 48195 20775 48201
rect 20717 48192 20729 48195
rect 20680 48164 20729 48192
rect 20680 48152 20686 48164
rect 20717 48161 20729 48164
rect 20763 48161 20775 48195
rect 25332 48192 25360 48232
rect 27062 48192 27068 48204
rect 20717 48155 20775 48161
rect 22066 48164 25360 48192
rect 27023 48164 27068 48192
rect 19245 48127 19303 48133
rect 19245 48093 19257 48127
rect 19291 48124 19303 48127
rect 20070 48124 20076 48136
rect 19291 48096 20076 48124
rect 19291 48093 19303 48096
rect 19245 48087 19303 48093
rect 20070 48084 20076 48096
rect 20128 48084 20134 48136
rect 16022 48016 16028 48068
rect 16080 48056 16086 48068
rect 16761 48059 16819 48065
rect 16761 48056 16773 48059
rect 16080 48028 16773 48056
rect 16080 48016 16086 48028
rect 16761 48025 16773 48028
rect 16807 48025 16819 48059
rect 16761 48019 16819 48025
rect 20162 48016 20168 48068
rect 20220 48056 20226 48068
rect 20441 48059 20499 48065
rect 20441 48056 20453 48059
rect 20220 48028 20453 48056
rect 20220 48016 20226 48028
rect 20441 48025 20453 48028
rect 20487 48025 20499 48059
rect 20441 48019 20499 48025
rect 20254 47988 20260 48000
rect 15948 47960 20260 47988
rect 20254 47948 20260 47960
rect 20312 47948 20318 48000
rect 20346 47948 20352 48000
rect 20404 47988 20410 48000
rect 22066 47988 22094 48164
rect 27062 48152 27068 48164
rect 27120 48152 27126 48204
rect 22557 48127 22615 48133
rect 22557 48093 22569 48127
rect 22603 48093 22615 48127
rect 22557 48087 22615 48093
rect 22572 48056 22600 48087
rect 22646 48084 22652 48136
rect 22704 48124 22710 48136
rect 23385 48127 23443 48133
rect 23385 48124 23397 48127
rect 22704 48096 23397 48124
rect 22704 48084 22710 48096
rect 23385 48093 23397 48096
rect 23431 48093 23443 48127
rect 24394 48124 24400 48136
rect 24355 48096 24400 48124
rect 23385 48087 23443 48093
rect 24394 48084 24400 48096
rect 24452 48084 24458 48136
rect 28644 48133 28672 48232
rect 28718 48220 28724 48272
rect 28776 48260 28782 48272
rect 29825 48263 29883 48269
rect 28776 48232 28821 48260
rect 28776 48220 28782 48232
rect 29825 48229 29837 48263
rect 29871 48260 29883 48263
rect 29914 48260 29920 48272
rect 29871 48232 29920 48260
rect 29871 48229 29883 48232
rect 29825 48223 29883 48229
rect 29914 48220 29920 48232
rect 29972 48220 29978 48272
rect 41141 48263 41199 48269
rect 32416 48232 40724 48260
rect 32214 48192 32220 48204
rect 32175 48164 32220 48192
rect 32214 48152 32220 48164
rect 32272 48152 32278 48204
rect 25869 48127 25927 48133
rect 25869 48093 25881 48127
rect 25915 48124 25927 48127
rect 26329 48127 26387 48133
rect 26329 48124 26341 48127
rect 25915 48096 26341 48124
rect 25915 48093 25927 48096
rect 25869 48087 25927 48093
rect 26329 48093 26341 48096
rect 26375 48093 26387 48127
rect 26329 48087 26387 48093
rect 28629 48127 28687 48133
rect 28629 48093 28641 48127
rect 28675 48093 28687 48127
rect 29730 48124 29736 48136
rect 29691 48096 29736 48124
rect 28629 48087 28687 48093
rect 29730 48084 29736 48096
rect 29788 48124 29794 48136
rect 30377 48127 30435 48133
rect 30377 48124 30389 48127
rect 29788 48096 30389 48124
rect 29788 48084 29794 48096
rect 30377 48093 30389 48096
rect 30423 48093 30435 48127
rect 31018 48124 31024 48136
rect 30979 48096 31024 48124
rect 30377 48087 30435 48093
rect 31018 48084 31024 48096
rect 31076 48084 31082 48136
rect 22922 48056 22928 48068
rect 22572 48028 22928 48056
rect 22922 48016 22928 48028
rect 22980 48016 22986 48068
rect 26513 48059 26571 48065
rect 26513 48025 26525 48059
rect 26559 48056 26571 48059
rect 27062 48056 27068 48068
rect 26559 48028 27068 48056
rect 26559 48025 26571 48028
rect 26513 48019 26571 48025
rect 27062 48016 27068 48028
rect 27120 48016 27126 48068
rect 30469 48059 30527 48065
rect 30469 48025 30481 48059
rect 30515 48056 30527 48059
rect 31205 48059 31263 48065
rect 31205 48056 31217 48059
rect 30515 48028 31217 48056
rect 30515 48025 30527 48028
rect 30469 48019 30527 48025
rect 31205 48025 31217 48028
rect 31251 48025 31263 48059
rect 31205 48019 31263 48025
rect 20404 47960 22094 47988
rect 20404 47948 20410 47960
rect 24394 47948 24400 48000
rect 24452 47988 24458 48000
rect 32416 47988 32444 48232
rect 35529 48195 35587 48201
rect 35529 48161 35541 48195
rect 35575 48192 35587 48195
rect 35802 48192 35808 48204
rect 35575 48164 35808 48192
rect 35575 48161 35587 48164
rect 35529 48155 35587 48161
rect 35802 48152 35808 48164
rect 35860 48152 35866 48204
rect 36722 48192 36728 48204
rect 36683 48164 36728 48192
rect 36722 48152 36728 48164
rect 36780 48152 36786 48204
rect 40696 48192 40724 48232
rect 41141 48229 41153 48263
rect 41187 48260 41199 48263
rect 42610 48260 42616 48272
rect 41187 48232 42616 48260
rect 41187 48229 41199 48232
rect 41141 48223 41199 48229
rect 42610 48220 42616 48232
rect 42668 48220 42674 48272
rect 47026 48220 47032 48272
rect 47084 48260 47090 48272
rect 49602 48260 49608 48272
rect 47084 48232 49608 48260
rect 47084 48220 47090 48232
rect 49602 48220 49608 48232
rect 49660 48220 49666 48272
rect 42518 48192 42524 48204
rect 40696 48164 42524 48192
rect 42518 48152 42524 48164
rect 42576 48152 42582 48204
rect 42794 48192 42800 48204
rect 42628 48164 42800 48192
rect 32490 48084 32496 48136
rect 32548 48124 32554 48136
rect 33321 48127 33379 48133
rect 33321 48124 33333 48127
rect 32548 48096 33333 48124
rect 32548 48084 32554 48096
rect 33321 48093 33333 48096
rect 33367 48093 33379 48127
rect 33321 48087 33379 48093
rect 34790 48084 34796 48136
rect 34848 48124 34854 48136
rect 34885 48127 34943 48133
rect 34885 48124 34897 48127
rect 34848 48096 34897 48124
rect 34848 48084 34854 48096
rect 34885 48093 34897 48096
rect 34931 48093 34943 48127
rect 34885 48087 34943 48093
rect 39853 48127 39911 48133
rect 39853 48093 39865 48127
rect 39899 48093 39911 48127
rect 41046 48124 41052 48136
rect 41007 48096 41052 48124
rect 39853 48087 39911 48093
rect 34977 48059 35035 48065
rect 34977 48025 34989 48059
rect 35023 48056 35035 48059
rect 35713 48059 35771 48065
rect 35713 48056 35725 48059
rect 35023 48028 35725 48056
rect 35023 48025 35035 48028
rect 34977 48019 35035 48025
rect 35713 48025 35725 48028
rect 35759 48025 35771 48059
rect 39868 48056 39896 48087
rect 41046 48084 41052 48096
rect 41104 48084 41110 48136
rect 41782 48124 41788 48136
rect 41743 48096 41788 48124
rect 41782 48084 41788 48096
rect 41840 48084 41846 48136
rect 42628 48133 42656 48164
rect 42794 48152 42800 48164
rect 42852 48152 42858 48204
rect 43162 48192 43168 48204
rect 43123 48164 43168 48192
rect 43162 48152 43168 48164
rect 43220 48152 43226 48204
rect 46750 48192 46756 48204
rect 46711 48164 46756 48192
rect 46750 48152 46756 48164
rect 46808 48152 46814 48204
rect 42613 48127 42671 48133
rect 42613 48093 42625 48127
rect 42659 48093 42671 48127
rect 42613 48087 42671 48093
rect 44726 48084 44732 48136
rect 44784 48124 44790 48136
rect 45005 48127 45063 48133
rect 45005 48124 45017 48127
rect 44784 48096 45017 48124
rect 44784 48084 44790 48096
rect 45005 48093 45017 48096
rect 45051 48093 45063 48127
rect 46290 48124 46296 48136
rect 46251 48096 46296 48124
rect 45005 48087 45063 48093
rect 46290 48084 46296 48096
rect 46348 48084 46354 48136
rect 39868 48028 42012 48056
rect 35713 48019 35771 48025
rect 24452 47960 32444 47988
rect 33413 47991 33471 47997
rect 24452 47948 24458 47960
rect 33413 47957 33425 47991
rect 33459 47988 33471 47991
rect 33502 47988 33508 48000
rect 33459 47960 33508 47988
rect 33459 47957 33471 47960
rect 33413 47951 33471 47957
rect 33502 47948 33508 47960
rect 33560 47948 33566 48000
rect 41874 47988 41880 48000
rect 41835 47960 41880 47988
rect 41874 47948 41880 47960
rect 41932 47948 41938 48000
rect 41984 47988 42012 48028
rect 42058 48016 42064 48068
rect 42116 48056 42122 48068
rect 42797 48059 42855 48065
rect 42797 48056 42809 48059
rect 42116 48028 42809 48056
rect 42116 48016 42122 48028
rect 42797 48025 42809 48028
rect 42843 48025 42855 48059
rect 42797 48019 42855 48025
rect 46477 48059 46535 48065
rect 46477 48025 46489 48059
rect 46523 48056 46535 48059
rect 47670 48056 47676 48068
rect 46523 48028 47676 48056
rect 46523 48025 46535 48028
rect 46477 48019 46535 48025
rect 47670 48016 47676 48028
rect 47728 48016 47734 48068
rect 44174 47988 44180 48000
rect 41984 47960 44180 47988
rect 44174 47948 44180 47960
rect 44232 47948 44238 48000
rect 45094 47948 45100 48000
rect 45152 47988 45158 48000
rect 45189 47991 45247 47997
rect 45189 47988 45201 47991
rect 45152 47960 45201 47988
rect 45152 47948 45158 47960
rect 45189 47957 45201 47960
rect 45235 47957 45247 47991
rect 45189 47951 45247 47957
rect 1104 47898 48852 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 48852 47898
rect 1104 47824 48852 47846
rect 1302 47744 1308 47796
rect 1360 47784 1366 47796
rect 3234 47784 3240 47796
rect 1360 47756 3240 47784
rect 1360 47744 1366 47756
rect 3234 47744 3240 47756
rect 3292 47744 3298 47796
rect 5350 47784 5356 47796
rect 5311 47756 5356 47784
rect 5350 47744 5356 47756
rect 5408 47744 5414 47796
rect 6546 47784 6552 47796
rect 6507 47756 6552 47784
rect 6546 47744 6552 47756
rect 6604 47744 6610 47796
rect 11606 47784 11612 47796
rect 11567 47756 11612 47784
rect 11606 47744 11612 47756
rect 11664 47744 11670 47796
rect 11698 47744 11704 47796
rect 11756 47784 11762 47796
rect 12253 47787 12311 47793
rect 12253 47784 12265 47787
rect 11756 47756 12265 47784
rect 11756 47744 11762 47756
rect 12253 47753 12265 47756
rect 12299 47753 12311 47787
rect 16022 47784 16028 47796
rect 15983 47756 16028 47784
rect 12253 47747 12311 47753
rect 16022 47744 16028 47756
rect 16080 47744 16086 47796
rect 17954 47784 17960 47796
rect 16684 47756 17960 47784
rect 2130 47716 2136 47728
rect 2091 47688 2136 47716
rect 2130 47676 2136 47688
rect 2188 47676 2194 47728
rect 5166 47676 5172 47728
rect 5224 47716 5230 47728
rect 16684 47716 16712 47756
rect 17954 47744 17960 47756
rect 18012 47744 18018 47796
rect 19153 47787 19211 47793
rect 19153 47753 19165 47787
rect 19199 47784 19211 47787
rect 19426 47784 19432 47796
rect 19199 47756 19432 47784
rect 19199 47753 19211 47756
rect 19153 47747 19211 47753
rect 19426 47744 19432 47756
rect 19484 47744 19490 47796
rect 20162 47784 20168 47796
rect 20123 47756 20168 47784
rect 20162 47744 20168 47756
rect 20220 47744 20226 47796
rect 20254 47744 20260 47796
rect 20312 47784 20318 47796
rect 27062 47784 27068 47796
rect 20312 47756 26234 47784
rect 27023 47756 27068 47784
rect 20312 47744 20318 47756
rect 18414 47716 18420 47728
rect 5224 47688 16712 47716
rect 16776 47688 18420 47716
rect 5224 47676 5230 47688
rect 1946 47648 1952 47660
rect 1907 47620 1952 47648
rect 1946 47608 1952 47620
rect 2004 47608 2010 47660
rect 4430 47608 4436 47660
rect 4488 47648 4494 47660
rect 4709 47651 4767 47657
rect 4709 47648 4721 47651
rect 4488 47620 4721 47648
rect 4488 47608 4494 47620
rect 4709 47617 4721 47620
rect 4755 47617 4767 47651
rect 4709 47611 4767 47617
rect 5261 47651 5319 47657
rect 5261 47617 5273 47651
rect 5307 47617 5319 47651
rect 5261 47611 5319 47617
rect 6457 47651 6515 47657
rect 6457 47617 6469 47651
rect 6503 47648 6515 47651
rect 6914 47648 6920 47660
rect 6503 47620 6920 47648
rect 6503 47617 6515 47620
rect 6457 47611 6515 47617
rect 3050 47580 3056 47592
rect 3011 47552 3056 47580
rect 3050 47540 3056 47552
rect 3108 47540 3114 47592
rect 5276 47444 5304 47611
rect 6914 47608 6920 47620
rect 6972 47608 6978 47660
rect 7098 47648 7104 47660
rect 7059 47620 7104 47648
rect 7098 47608 7104 47620
rect 7156 47608 7162 47660
rect 11514 47648 11520 47660
rect 11475 47620 11520 47648
rect 11514 47608 11520 47620
rect 11572 47608 11578 47660
rect 12066 47608 12072 47660
rect 12124 47648 12130 47660
rect 12161 47651 12219 47657
rect 12161 47648 12173 47651
rect 12124 47620 12173 47648
rect 12124 47608 12130 47620
rect 12161 47617 12173 47620
rect 12207 47617 12219 47651
rect 12161 47611 12219 47617
rect 14182 47608 14188 47660
rect 14240 47648 14246 47660
rect 14369 47651 14427 47657
rect 14369 47648 14381 47651
rect 14240 47620 14381 47648
rect 14240 47608 14246 47620
rect 14369 47617 14381 47620
rect 14415 47617 14427 47651
rect 14369 47611 14427 47617
rect 15562 47608 15568 47660
rect 15620 47648 15626 47660
rect 16776 47657 16804 47688
rect 18414 47676 18420 47688
rect 18472 47676 18478 47728
rect 21913 47719 21971 47725
rect 21913 47685 21925 47719
rect 21959 47716 21971 47719
rect 22186 47716 22192 47728
rect 21959 47688 22192 47716
rect 21959 47685 21971 47688
rect 21913 47679 21971 47685
rect 22186 47676 22192 47688
rect 22244 47676 22250 47728
rect 26206 47716 26234 47756
rect 27062 47744 27068 47756
rect 27120 47744 27126 47796
rect 29822 47744 29828 47796
rect 29880 47784 29886 47796
rect 30101 47787 30159 47793
rect 30101 47784 30113 47787
rect 29880 47756 30113 47784
rect 29880 47744 29886 47756
rect 30101 47753 30113 47756
rect 30147 47753 30159 47787
rect 30101 47747 30159 47753
rect 32217 47787 32275 47793
rect 32217 47753 32229 47787
rect 32263 47784 32275 47787
rect 32306 47784 32312 47796
rect 32263 47756 32312 47784
rect 32263 47753 32275 47756
rect 32217 47747 32275 47753
rect 32306 47744 32312 47756
rect 32364 47744 32370 47796
rect 35894 47744 35900 47796
rect 35952 47784 35958 47796
rect 41785 47787 41843 47793
rect 35952 47756 35997 47784
rect 35952 47744 35958 47756
rect 41785 47753 41797 47787
rect 41831 47784 41843 47787
rect 42058 47784 42064 47796
rect 41831 47756 42064 47784
rect 41831 47753 41843 47756
rect 41785 47747 41843 47753
rect 42058 47744 42064 47756
rect 42116 47744 42122 47796
rect 42518 47744 42524 47796
rect 42576 47784 42582 47796
rect 42576 47756 44680 47784
rect 42576 47744 42582 47756
rect 31846 47716 31852 47728
rect 26206 47688 31852 47716
rect 31846 47676 31852 47688
rect 31904 47716 31910 47728
rect 33502 47716 33508 47728
rect 31904 47688 32168 47716
rect 33463 47688 33508 47716
rect 31904 47676 31910 47688
rect 15933 47651 15991 47657
rect 15933 47648 15945 47651
rect 15620 47620 15945 47648
rect 15620 47608 15626 47620
rect 15933 47617 15945 47620
rect 15979 47617 15991 47651
rect 15933 47611 15991 47617
rect 16761 47651 16819 47657
rect 16761 47617 16773 47651
rect 16807 47617 16819 47651
rect 19058 47648 19064 47660
rect 19019 47620 19064 47648
rect 16761 47611 16819 47617
rect 19058 47608 19064 47620
rect 19116 47608 19122 47660
rect 19334 47608 19340 47660
rect 19392 47648 19398 47660
rect 20073 47651 20131 47657
rect 20073 47648 20085 47651
rect 19392 47620 20085 47648
rect 19392 47608 19398 47620
rect 20073 47617 20085 47620
rect 20119 47617 20131 47651
rect 20073 47611 20131 47617
rect 21726 47608 21732 47660
rect 21784 47648 21790 47660
rect 21821 47651 21879 47657
rect 21821 47648 21833 47651
rect 21784 47620 21833 47648
rect 21784 47608 21790 47620
rect 21821 47617 21833 47620
rect 21867 47617 21879 47651
rect 21821 47611 21879 47617
rect 22370 47608 22376 47660
rect 22428 47648 22434 47660
rect 22649 47651 22707 47657
rect 22649 47648 22661 47651
rect 22428 47620 22661 47648
rect 22428 47608 22434 47620
rect 22649 47617 22661 47620
rect 22695 47617 22707 47651
rect 24118 47648 24124 47660
rect 24079 47620 24124 47648
rect 22649 47611 22707 47617
rect 24118 47608 24124 47620
rect 24176 47608 24182 47660
rect 26973 47651 27031 47657
rect 26973 47617 26985 47651
rect 27019 47617 27031 47651
rect 26973 47611 27031 47617
rect 7285 47583 7343 47589
rect 7285 47549 7297 47583
rect 7331 47580 7343 47583
rect 7650 47580 7656 47592
rect 7331 47552 7656 47580
rect 7331 47549 7343 47552
rect 7285 47543 7343 47549
rect 7650 47540 7656 47552
rect 7708 47540 7714 47592
rect 7742 47540 7748 47592
rect 7800 47580 7806 47592
rect 16942 47580 16948 47592
rect 7800 47552 7845 47580
rect 16903 47552 16948 47580
rect 7800 47540 7806 47552
rect 16942 47540 16948 47552
rect 17000 47540 17006 47592
rect 17221 47583 17279 47589
rect 17221 47549 17233 47583
rect 17267 47549 17279 47583
rect 17221 47543 17279 47549
rect 15102 47472 15108 47524
rect 15160 47512 15166 47524
rect 17236 47512 17264 47543
rect 26988 47524 27016 47611
rect 27614 47608 27620 47660
rect 27672 47648 27678 47660
rect 27709 47651 27767 47657
rect 27709 47648 27721 47651
rect 27672 47620 27721 47648
rect 27672 47608 27678 47620
rect 27709 47617 27721 47620
rect 27755 47617 27767 47651
rect 30006 47648 30012 47660
rect 29967 47620 30012 47648
rect 27709 47611 27767 47617
rect 30006 47608 30012 47620
rect 30064 47608 30070 47660
rect 31018 47608 31024 47660
rect 31076 47648 31082 47660
rect 32140 47657 32168 47688
rect 33502 47676 33508 47688
rect 33560 47676 33566 47728
rect 42705 47719 42763 47725
rect 42705 47685 42717 47719
rect 42751 47716 42763 47719
rect 43441 47719 43499 47725
rect 43441 47716 43453 47719
rect 42751 47688 43453 47716
rect 42751 47685 42763 47688
rect 42705 47679 42763 47685
rect 43441 47685 43453 47688
rect 43487 47685 43499 47719
rect 43441 47679 43499 47685
rect 31297 47651 31355 47657
rect 31297 47648 31309 47651
rect 31076 47620 31309 47648
rect 31076 47608 31082 47620
rect 31297 47617 31309 47620
rect 31343 47617 31355 47651
rect 31297 47611 31355 47617
rect 32125 47651 32183 47657
rect 32125 47617 32137 47651
rect 32171 47617 32183 47651
rect 33318 47648 33324 47660
rect 33279 47620 33324 47648
rect 32125 47611 32183 47617
rect 33318 47608 33324 47620
rect 33376 47608 33382 47660
rect 35805 47651 35863 47657
rect 35805 47617 35817 47651
rect 35851 47617 35863 47651
rect 41690 47648 41696 47660
rect 41651 47620 41696 47648
rect 35805 47611 35863 47617
rect 27893 47583 27951 47589
rect 27893 47549 27905 47583
rect 27939 47580 27951 47583
rect 28166 47580 28172 47592
rect 27939 47552 28172 47580
rect 27939 47549 27951 47552
rect 27893 47543 27951 47549
rect 28166 47540 28172 47552
rect 28224 47540 28230 47592
rect 28350 47580 28356 47592
rect 28311 47552 28356 47580
rect 28350 47540 28356 47552
rect 28408 47540 28414 47592
rect 29822 47540 29828 47592
rect 29880 47580 29886 47592
rect 32490 47580 32496 47592
rect 29880 47552 32496 47580
rect 29880 47540 29886 47552
rect 32490 47540 32496 47552
rect 32548 47540 32554 47592
rect 34698 47580 34704 47592
rect 34659 47552 34704 47580
rect 34698 47540 34704 47552
rect 34756 47540 34762 47592
rect 26970 47512 26976 47524
rect 15160 47484 17264 47512
rect 26883 47484 26976 47512
rect 15160 47472 15166 47484
rect 26970 47472 26976 47484
rect 27028 47512 27034 47524
rect 30742 47512 30748 47524
rect 27028 47484 30748 47512
rect 27028 47472 27034 47484
rect 30742 47472 30748 47484
rect 30800 47472 30806 47524
rect 13262 47444 13268 47456
rect 5276 47416 13268 47444
rect 13262 47404 13268 47416
rect 13320 47404 13326 47456
rect 19058 47404 19064 47456
rect 19116 47444 19122 47456
rect 20070 47444 20076 47456
rect 19116 47416 20076 47444
rect 19116 47404 19122 47416
rect 20070 47404 20076 47416
rect 20128 47404 20134 47456
rect 23934 47444 23940 47456
rect 23895 47416 23940 47444
rect 23934 47404 23940 47416
rect 23992 47404 23998 47456
rect 34514 47404 34520 47456
rect 34572 47444 34578 47456
rect 35820 47444 35848 47611
rect 41690 47608 41696 47620
rect 41748 47648 41754 47660
rect 42613 47651 42671 47657
rect 42613 47648 42625 47651
rect 41748 47620 42625 47648
rect 41748 47608 41754 47620
rect 42613 47617 42625 47620
rect 42659 47617 42671 47651
rect 44652 47648 44680 47756
rect 46198 47744 46204 47796
rect 46256 47784 46262 47796
rect 46293 47787 46351 47793
rect 46293 47784 46305 47787
rect 46256 47756 46305 47784
rect 46256 47744 46262 47756
rect 46293 47753 46305 47756
rect 46339 47753 46351 47787
rect 48314 47784 48320 47796
rect 46293 47747 46351 47753
rect 47596 47756 48320 47784
rect 45097 47719 45155 47725
rect 45097 47685 45109 47719
rect 45143 47716 45155 47719
rect 47596 47716 47624 47756
rect 48314 47744 48320 47756
rect 48372 47744 48378 47796
rect 47762 47716 47768 47728
rect 45143 47688 47624 47716
rect 47723 47688 47768 47716
rect 45143 47685 45155 47688
rect 45097 47679 45155 47685
rect 47762 47676 47768 47688
rect 47820 47676 47826 47728
rect 45557 47651 45615 47657
rect 45557 47648 45569 47651
rect 44652 47620 45569 47648
rect 42613 47611 42671 47617
rect 45557 47617 45569 47620
rect 45603 47648 45615 47651
rect 46201 47651 46259 47657
rect 46201 47648 46213 47651
rect 45603 47620 46213 47648
rect 45603 47617 45615 47620
rect 45557 47611 45615 47617
rect 46201 47617 46213 47620
rect 46247 47617 46259 47651
rect 46201 47611 46259 47617
rect 46845 47651 46903 47657
rect 46845 47617 46857 47651
rect 46891 47617 46903 47651
rect 46845 47611 46903 47617
rect 43257 47583 43315 47589
rect 43257 47549 43269 47583
rect 43303 47580 43315 47583
rect 43438 47580 43444 47592
rect 43303 47552 43444 47580
rect 43303 47549 43315 47552
rect 43257 47543 43315 47549
rect 43438 47540 43444 47552
rect 43496 47540 43502 47592
rect 46014 47540 46020 47592
rect 46072 47580 46078 47592
rect 46860 47580 46888 47611
rect 46072 47552 46888 47580
rect 46072 47540 46078 47552
rect 40678 47472 40684 47524
rect 40736 47512 40742 47524
rect 47949 47515 48007 47521
rect 47949 47512 47961 47515
rect 40736 47484 47961 47512
rect 40736 47472 40742 47484
rect 47949 47481 47961 47484
rect 47995 47481 48007 47515
rect 47949 47475 48007 47481
rect 44542 47444 44548 47456
rect 34572 47416 44548 47444
rect 34572 47404 34578 47416
rect 44542 47404 44548 47416
rect 44600 47404 44606 47456
rect 45186 47404 45192 47456
rect 45244 47444 45250 47456
rect 45649 47447 45707 47453
rect 45649 47444 45661 47447
rect 45244 47416 45661 47444
rect 45244 47404 45250 47416
rect 45649 47413 45661 47416
rect 45695 47413 45707 47447
rect 45649 47407 45707 47413
rect 46382 47404 46388 47456
rect 46440 47444 46446 47456
rect 46937 47447 46995 47453
rect 46937 47444 46949 47447
rect 46440 47416 46949 47444
rect 46440 47404 46446 47416
rect 46937 47413 46949 47416
rect 46983 47413 46995 47447
rect 46937 47407 46995 47413
rect 1104 47354 48852 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 48852 47354
rect 1104 47280 48852 47302
rect 2222 47200 2228 47252
rect 2280 47240 2286 47252
rect 2501 47243 2559 47249
rect 2501 47240 2513 47243
rect 2280 47212 2513 47240
rect 2280 47200 2286 47212
rect 2501 47209 2513 47212
rect 2547 47209 2559 47243
rect 2501 47203 2559 47209
rect 3142 47200 3148 47252
rect 3200 47240 3206 47252
rect 3973 47243 4031 47249
rect 3973 47240 3985 47243
rect 3200 47212 3985 47240
rect 3200 47200 3206 47212
rect 3973 47209 3985 47212
rect 4019 47209 4031 47243
rect 7650 47240 7656 47252
rect 7611 47212 7656 47240
rect 3973 47203 4031 47209
rect 7650 47200 7656 47212
rect 7708 47200 7714 47252
rect 16942 47240 16948 47252
rect 16903 47212 16948 47240
rect 16942 47200 16948 47212
rect 17000 47200 17006 47252
rect 18046 47200 18052 47252
rect 18104 47240 18110 47252
rect 40678 47240 40684 47252
rect 18104 47212 40684 47240
rect 18104 47200 18110 47212
rect 40678 47200 40684 47212
rect 40736 47200 40742 47252
rect 42337 47243 42395 47249
rect 42337 47209 42349 47243
rect 42383 47240 42395 47243
rect 42426 47240 42432 47252
rect 42383 47212 42432 47240
rect 42383 47209 42395 47212
rect 42337 47203 42395 47209
rect 42426 47200 42432 47212
rect 42484 47200 42490 47252
rect 43438 47240 43444 47252
rect 43399 47212 43444 47240
rect 43438 47200 43444 47212
rect 43496 47200 43502 47252
rect 6914 47132 6920 47184
rect 6972 47172 6978 47184
rect 17862 47172 17868 47184
rect 6972 47144 17868 47172
rect 6972 47132 6978 47144
rect 17862 47132 17868 47144
rect 17920 47132 17926 47184
rect 18230 47132 18236 47184
rect 18288 47172 18294 47184
rect 26970 47172 26976 47184
rect 18288 47144 26976 47172
rect 18288 47132 18294 47144
rect 26970 47132 26976 47144
rect 27028 47132 27034 47184
rect 29822 47172 29828 47184
rect 27816 47144 29828 47172
rect 14458 47064 14464 47116
rect 14516 47104 14522 47116
rect 27816 47104 27844 47144
rect 29822 47132 29828 47144
rect 29880 47132 29886 47184
rect 30650 47172 30656 47184
rect 30611 47144 30656 47172
rect 30650 47132 30656 47144
rect 30708 47132 30714 47184
rect 30742 47132 30748 47184
rect 30800 47172 30806 47184
rect 41690 47172 41696 47184
rect 30800 47144 41696 47172
rect 30800 47132 30806 47144
rect 41690 47132 41696 47144
rect 41748 47132 41754 47184
rect 43990 47132 43996 47184
rect 44048 47172 44054 47184
rect 44085 47175 44143 47181
rect 44085 47172 44097 47175
rect 44048 47144 44097 47172
rect 44048 47132 44054 47144
rect 44085 47141 44097 47144
rect 44131 47141 44143 47175
rect 44085 47135 44143 47141
rect 30006 47104 30012 47116
rect 14516 47076 27844 47104
rect 27908 47076 30012 47104
rect 14516 47064 14522 47076
rect 1394 47036 1400 47048
rect 1355 47008 1400 47036
rect 1394 46996 1400 47008
rect 1452 46996 1458 47048
rect 2406 47036 2412 47048
rect 2367 47008 2412 47036
rect 2406 46996 2412 47008
rect 2464 46996 2470 47048
rect 2774 46996 2780 47048
rect 2832 47036 2838 47048
rect 3237 47039 3295 47045
rect 3237 47036 3249 47039
rect 2832 47008 3249 47036
rect 2832 46996 2838 47008
rect 3237 47005 3249 47008
rect 3283 47005 3295 47039
rect 3237 46999 3295 47005
rect 7561 47039 7619 47045
rect 7561 47005 7573 47039
rect 7607 47036 7619 47039
rect 7926 47036 7932 47048
rect 7607 47008 7932 47036
rect 7607 47005 7619 47008
rect 7561 46999 7619 47005
rect 7926 46996 7932 47008
rect 7984 46996 7990 47048
rect 16868 47045 16896 47076
rect 16853 47039 16911 47045
rect 16853 47005 16865 47039
rect 16899 47005 16911 47039
rect 19242 47036 19248 47048
rect 19203 47008 19248 47036
rect 16853 46999 16911 47005
rect 19242 46996 19248 47008
rect 19300 46996 19306 47048
rect 20088 47036 20300 47038
rect 27908 47036 27936 47076
rect 30006 47064 30012 47076
rect 30064 47104 30070 47116
rect 39850 47104 39856 47116
rect 30064 47076 39856 47104
rect 30064 47064 30070 47076
rect 39850 47064 39856 47076
rect 39908 47064 39914 47116
rect 45186 47104 45192 47116
rect 45147 47076 45192 47104
rect 45186 47064 45192 47076
rect 45244 47064 45250 47116
rect 45278 47064 45284 47116
rect 45336 47104 45342 47116
rect 45557 47107 45615 47113
rect 45557 47104 45569 47107
rect 45336 47076 45569 47104
rect 45336 47064 45342 47076
rect 45557 47073 45569 47076
rect 45603 47073 45615 47107
rect 45557 47067 45615 47073
rect 28074 47036 28080 47048
rect 20088 47010 27936 47036
rect 20088 46980 20116 47010
rect 20272 47008 27936 47010
rect 28035 47008 28080 47036
rect 28074 46996 28080 47008
rect 28132 46996 28138 47048
rect 28166 46996 28172 47048
rect 28224 47036 28230 47048
rect 43898 47036 43904 47048
rect 28224 47008 28269 47036
rect 43859 47008 43904 47036
rect 28224 46996 28230 47008
rect 43898 46996 43904 47008
rect 43956 46996 43962 47048
rect 45002 47036 45008 47048
rect 44963 47008 45008 47036
rect 45002 46996 45008 47008
rect 45060 46996 45066 47048
rect 47949 47039 48007 47045
rect 47949 47005 47961 47039
rect 47995 47036 48007 47039
rect 48958 47036 48964 47048
rect 47995 47008 48964 47036
rect 47995 47005 48007 47008
rect 47949 46999 48007 47005
rect 48958 46996 48964 47008
rect 49016 46996 49022 47048
rect 1596 46940 19932 46968
rect 1596 46909 1624 46940
rect 1581 46903 1639 46909
rect 1581 46869 1593 46903
rect 1627 46869 1639 46903
rect 19904 46900 19932 46940
rect 20070 46928 20076 46980
rect 20128 46968 20134 46980
rect 31018 46968 31024 46980
rect 20128 46940 20173 46968
rect 20364 46940 31024 46968
rect 20128 46928 20134 46940
rect 20364 46900 20392 46940
rect 31018 46928 31024 46940
rect 31076 46928 31082 46980
rect 48133 46971 48191 46977
rect 48133 46968 48145 46971
rect 47964 46940 48145 46968
rect 47964 46912 47992 46940
rect 48133 46937 48145 46940
rect 48179 46937 48191 46971
rect 48133 46931 48191 46937
rect 19904 46872 20392 46900
rect 1581 46863 1639 46869
rect 47946 46860 47952 46912
rect 48004 46860 48010 46912
rect 1104 46810 48852 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 48852 46810
rect 1104 46736 48852 46758
rect 44634 46696 44640 46708
rect 44595 46668 44640 46696
rect 44634 46656 44640 46668
rect 44692 46656 44698 46708
rect 47670 46696 47676 46708
rect 47631 46668 47676 46696
rect 47670 46656 47676 46668
rect 47728 46656 47734 46708
rect 2774 46628 2780 46640
rect 1964 46600 2780 46628
rect 1964 46569 1992 46600
rect 2774 46588 2780 46600
rect 2832 46588 2838 46640
rect 3786 46628 3792 46640
rect 3747 46600 3792 46628
rect 3786 46588 3792 46600
rect 3844 46588 3850 46640
rect 18230 46628 18236 46640
rect 18191 46600 18236 46628
rect 18230 46588 18236 46600
rect 18288 46588 18294 46640
rect 22922 46588 22928 46640
rect 22980 46628 22986 46640
rect 22980 46600 47624 46628
rect 22980 46588 22986 46600
rect 1949 46563 2007 46569
rect 1949 46529 1961 46563
rect 1995 46529 2007 46563
rect 1949 46523 2007 46529
rect 17957 46563 18015 46569
rect 17957 46529 17969 46563
rect 18003 46560 18015 46563
rect 19061 46563 19119 46569
rect 19061 46560 19073 46563
rect 18003 46532 19073 46560
rect 18003 46529 18015 46532
rect 17957 46523 18015 46529
rect 19061 46529 19073 46532
rect 19107 46560 19119 46563
rect 19242 46560 19248 46572
rect 19107 46532 19248 46560
rect 19107 46529 19119 46532
rect 19061 46523 19119 46529
rect 19242 46520 19248 46532
rect 19300 46520 19306 46572
rect 42794 46560 42800 46572
rect 42755 46532 42800 46560
rect 42794 46520 42800 46532
rect 42852 46520 42858 46572
rect 44082 46560 44088 46572
rect 44043 46532 44088 46560
rect 44082 46520 44088 46532
rect 44140 46520 44146 46572
rect 44542 46560 44548 46572
rect 44503 46532 44548 46560
rect 44542 46520 44548 46532
rect 44600 46520 44606 46572
rect 47026 46560 47032 46572
rect 46987 46532 47032 46560
rect 47026 46520 47032 46532
rect 47084 46520 47090 46572
rect 47596 46569 47624 46600
rect 47581 46563 47639 46569
rect 47581 46529 47593 46563
rect 47627 46529 47639 46563
rect 47581 46523 47639 46529
rect 2133 46495 2191 46501
rect 2133 46461 2145 46495
rect 2179 46492 2191 46495
rect 2498 46492 2504 46504
rect 2179 46464 2504 46492
rect 2179 46461 2191 46464
rect 2133 46455 2191 46461
rect 2498 46452 2504 46464
rect 2556 46452 2562 46504
rect 20070 46492 20076 46504
rect 20031 46464 20076 46492
rect 20070 46452 20076 46464
rect 20128 46452 20134 46504
rect 43441 46495 43499 46501
rect 43441 46461 43453 46495
rect 43487 46492 43499 46495
rect 45189 46495 45247 46501
rect 45189 46492 45201 46495
rect 43487 46464 45201 46492
rect 43487 46461 43499 46464
rect 43441 46455 43499 46461
rect 45189 46461 45201 46464
rect 45235 46461 45247 46495
rect 45189 46455 45247 46461
rect 45373 46495 45431 46501
rect 45373 46461 45385 46495
rect 45419 46492 45431 46495
rect 46382 46492 46388 46504
rect 45419 46464 46388 46492
rect 45419 46461 45431 46464
rect 45373 46455 45431 46461
rect 46382 46452 46388 46464
rect 46440 46452 46446 46504
rect 1104 46266 48852 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 48852 46266
rect 1104 46192 48852 46214
rect 2498 46152 2504 46164
rect 2459 46124 2504 46152
rect 2498 46112 2504 46124
rect 2556 46112 2562 46164
rect 18601 46155 18659 46161
rect 18601 46121 18613 46155
rect 18647 46152 18659 46155
rect 19242 46152 19248 46164
rect 18647 46124 19248 46152
rect 18647 46121 18659 46124
rect 18601 46115 18659 46121
rect 19242 46112 19248 46124
rect 19300 46112 19306 46164
rect 44453 46155 44511 46161
rect 44453 46121 44465 46155
rect 44499 46152 44511 46155
rect 45002 46152 45008 46164
rect 44499 46124 45008 46152
rect 44499 46121 44511 46124
rect 44453 46115 44511 46121
rect 45002 46112 45008 46124
rect 45060 46112 45066 46164
rect 45189 46155 45247 46161
rect 45189 46121 45201 46155
rect 45235 46152 45247 46155
rect 45370 46152 45376 46164
rect 45235 46124 45376 46152
rect 45235 46121 45247 46124
rect 45189 46115 45247 46121
rect 45370 46112 45376 46124
rect 45428 46112 45434 46164
rect 46293 46019 46351 46025
rect 46293 45985 46305 46019
rect 46339 46016 46351 46019
rect 47762 46016 47768 46028
rect 46339 45988 47768 46016
rect 46339 45985 46351 45988
rect 46293 45979 46351 45985
rect 47762 45976 47768 45988
rect 47820 45976 47826 46028
rect 48130 46016 48136 46028
rect 48091 45988 48136 46016
rect 48130 45976 48136 45988
rect 48188 45976 48194 46028
rect 1394 45948 1400 45960
rect 1355 45920 1400 45948
rect 1394 45908 1400 45920
rect 1452 45908 1458 45960
rect 2409 45951 2467 45957
rect 2409 45917 2421 45951
rect 2455 45948 2467 45951
rect 2498 45948 2504 45960
rect 2455 45920 2504 45948
rect 2455 45917 2467 45920
rect 2409 45911 2467 45917
rect 2498 45908 2504 45920
rect 2556 45908 2562 45960
rect 3234 45948 3240 45960
rect 3195 45920 3240 45948
rect 3234 45908 3240 45920
rect 3292 45908 3298 45960
rect 3970 45948 3976 45960
rect 3931 45920 3976 45948
rect 3970 45908 3976 45920
rect 4028 45908 4034 45960
rect 13262 45948 13268 45960
rect 13175 45920 13268 45948
rect 13262 45908 13268 45920
rect 13320 45948 13326 45960
rect 18230 45948 18236 45960
rect 13320 45920 18236 45948
rect 13320 45908 13326 45920
rect 18230 45908 18236 45920
rect 18288 45908 18294 45960
rect 18414 45948 18420 45960
rect 18327 45920 18420 45948
rect 18414 45908 18420 45920
rect 18472 45948 18478 45960
rect 19242 45948 19248 45960
rect 18472 45920 18828 45948
rect 19203 45920 19248 45948
rect 18472 45908 18478 45920
rect 18800 45880 18828 45920
rect 19242 45908 19248 45920
rect 19300 45908 19306 45960
rect 44174 45908 44180 45960
rect 44232 45948 44238 45960
rect 45097 45951 45155 45957
rect 45097 45948 45109 45951
rect 44232 45920 45109 45948
rect 44232 45908 44238 45920
rect 45097 45917 45109 45920
rect 45143 45948 45155 45951
rect 45922 45948 45928 45960
rect 45143 45920 45928 45948
rect 45143 45917 45155 45920
rect 45097 45911 45155 45917
rect 45922 45908 45928 45920
rect 45980 45908 45986 45960
rect 19150 45880 19156 45892
rect 6886 45852 18736 45880
rect 18800 45852 19156 45880
rect 1581 45815 1639 45821
rect 1581 45781 1593 45815
rect 1627 45812 1639 45815
rect 6886 45812 6914 45852
rect 1627 45784 6914 45812
rect 1627 45781 1639 45784
rect 1581 45775 1639 45781
rect 13078 45772 13084 45824
rect 13136 45812 13142 45824
rect 13357 45815 13415 45821
rect 13357 45812 13369 45815
rect 13136 45784 13369 45812
rect 13136 45772 13142 45784
rect 13357 45781 13369 45784
rect 13403 45781 13415 45815
rect 18708 45812 18736 45852
rect 19150 45840 19156 45852
rect 19208 45840 19214 45892
rect 19978 45840 19984 45892
rect 20036 45880 20042 45892
rect 20073 45883 20131 45889
rect 20073 45880 20085 45883
rect 20036 45852 20085 45880
rect 20036 45840 20042 45852
rect 20073 45849 20085 45852
rect 20119 45880 20131 45883
rect 34514 45880 34520 45892
rect 20119 45852 34520 45880
rect 20119 45849 20131 45852
rect 20073 45843 20131 45849
rect 34514 45840 34520 45852
rect 34572 45840 34578 45892
rect 46477 45883 46535 45889
rect 46477 45849 46489 45883
rect 46523 45880 46535 45883
rect 47670 45880 47676 45892
rect 46523 45852 47676 45880
rect 46523 45849 46535 45852
rect 46477 45843 46535 45849
rect 47670 45840 47676 45852
rect 47728 45840 47734 45892
rect 22830 45812 22836 45824
rect 18708 45784 22836 45812
rect 13357 45775 13415 45781
rect 22830 45772 22836 45784
rect 22888 45772 22894 45824
rect 1104 45722 48852 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 48852 45722
rect 1104 45648 48852 45670
rect 2498 45608 2504 45620
rect 2411 45580 2504 45608
rect 2498 45568 2504 45580
rect 2556 45608 2562 45620
rect 2556 45580 3372 45608
rect 2556 45568 2562 45580
rect 2041 45475 2099 45481
rect 2041 45441 2053 45475
rect 2087 45472 2099 45475
rect 2516 45472 2544 45568
rect 3234 45540 3240 45552
rect 2700 45512 3240 45540
rect 2700 45481 2728 45512
rect 3234 45500 3240 45512
rect 3292 45500 3298 45552
rect 3344 45540 3372 45580
rect 20070 45568 20076 45620
rect 20128 45608 20134 45620
rect 28074 45608 28080 45620
rect 20128 45580 28080 45608
rect 20128 45568 20134 45580
rect 28074 45568 28080 45580
rect 28132 45608 28138 45620
rect 28810 45608 28816 45620
rect 28132 45580 28816 45608
rect 28132 45568 28138 45580
rect 28810 45568 28816 45580
rect 28868 45568 28874 45620
rect 13078 45540 13084 45552
rect 3344 45512 6914 45540
rect 13039 45512 13084 45540
rect 2087 45444 2544 45472
rect 2685 45475 2743 45481
rect 2087 45441 2099 45444
rect 2041 45435 2099 45441
rect 2685 45441 2697 45475
rect 2731 45441 2743 45475
rect 2685 45435 2743 45441
rect 2869 45407 2927 45413
rect 2869 45373 2881 45407
rect 2915 45404 2927 45407
rect 3878 45404 3884 45416
rect 2915 45376 3884 45404
rect 2915 45373 2927 45376
rect 2869 45367 2927 45373
rect 3878 45364 3884 45376
rect 3936 45364 3942 45416
rect 4062 45404 4068 45416
rect 4023 45376 4068 45404
rect 4062 45364 4068 45376
rect 4120 45364 4126 45416
rect 6886 45336 6914 45512
rect 13078 45500 13084 45512
rect 13136 45500 13142 45552
rect 47670 45540 47676 45552
rect 40696 45512 46980 45540
rect 47631 45512 47676 45540
rect 18969 45475 19027 45481
rect 18969 45441 18981 45475
rect 19015 45472 19027 45475
rect 19242 45472 19248 45484
rect 19015 45444 19248 45472
rect 19015 45441 19027 45444
rect 18969 45435 19027 45441
rect 19242 45432 19248 45444
rect 19300 45432 19306 45484
rect 12897 45407 12955 45413
rect 12897 45373 12909 45407
rect 12943 45404 12955 45407
rect 13170 45404 13176 45416
rect 12943 45376 13176 45404
rect 12943 45373 12955 45376
rect 12897 45367 12955 45373
rect 13170 45364 13176 45376
rect 13228 45364 13234 45416
rect 13814 45404 13820 45416
rect 13775 45376 13820 45404
rect 13814 45364 13820 45376
rect 13872 45364 13878 45416
rect 19337 45407 19395 45413
rect 19337 45373 19349 45407
rect 19383 45404 19395 45407
rect 21542 45404 21548 45416
rect 19383 45376 21548 45404
rect 19383 45373 19395 45376
rect 19337 45367 19395 45373
rect 19352 45336 19380 45367
rect 21542 45364 21548 45376
rect 21600 45404 21606 45416
rect 21600 45376 26234 45404
rect 21600 45364 21606 45376
rect 6886 45308 19380 45336
rect 26206 45336 26234 45376
rect 28810 45364 28816 45416
rect 28868 45404 28874 45416
rect 40696 45404 40724 45512
rect 42334 45432 42340 45484
rect 42392 45472 42398 45484
rect 44821 45475 44879 45481
rect 44821 45472 44833 45475
rect 42392 45444 44833 45472
rect 42392 45432 42398 45444
rect 44821 45441 44833 45444
rect 44867 45441 44879 45475
rect 45462 45472 45468 45484
rect 45423 45444 45468 45472
rect 44821 45435 44879 45441
rect 45462 45432 45468 45444
rect 45520 45432 45526 45484
rect 46290 45432 46296 45484
rect 46348 45472 46354 45484
rect 46385 45475 46443 45481
rect 46385 45472 46397 45475
rect 46348 45444 46397 45472
rect 46348 45432 46354 45444
rect 46385 45441 46397 45444
rect 46431 45441 46443 45475
rect 46385 45435 46443 45441
rect 46845 45475 46903 45481
rect 46845 45441 46857 45475
rect 46891 45441 46903 45475
rect 46952 45472 46980 45512
rect 47670 45500 47676 45512
rect 47728 45500 47734 45552
rect 47118 45472 47124 45484
rect 46952 45444 47124 45472
rect 46845 45435 46903 45441
rect 46750 45404 46756 45416
rect 28868 45376 40724 45404
rect 41386 45376 46756 45404
rect 28868 45364 28874 45376
rect 41386 45336 41414 45376
rect 46750 45364 46756 45376
rect 46808 45404 46814 45416
rect 46860 45404 46888 45435
rect 47118 45432 47124 45444
rect 47176 45472 47182 45484
rect 47581 45475 47639 45481
rect 47581 45472 47593 45475
rect 47176 45444 47593 45472
rect 47176 45432 47182 45444
rect 47581 45441 47593 45444
rect 47627 45441 47639 45475
rect 47581 45435 47639 45441
rect 46808 45376 46888 45404
rect 46808 45364 46814 45376
rect 26206 45308 41414 45336
rect 1394 45228 1400 45280
rect 1452 45268 1458 45280
rect 1581 45271 1639 45277
rect 1581 45268 1593 45271
rect 1452 45240 1593 45268
rect 1452 45228 1458 45240
rect 1581 45237 1593 45240
rect 1627 45237 1639 45271
rect 1581 45231 1639 45237
rect 2038 45228 2044 45280
rect 2096 45268 2102 45280
rect 2133 45271 2191 45277
rect 2133 45268 2145 45271
rect 2096 45240 2145 45268
rect 2096 45228 2102 45240
rect 2133 45237 2145 45240
rect 2179 45237 2191 45271
rect 2133 45231 2191 45237
rect 46474 45228 46480 45280
rect 46532 45268 46538 45280
rect 46937 45271 46995 45277
rect 46937 45268 46949 45271
rect 46532 45240 46949 45268
rect 46532 45228 46538 45240
rect 46937 45237 46949 45240
rect 46983 45237 46995 45271
rect 46937 45231 46995 45237
rect 1104 45178 48852 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 48852 45178
rect 1104 45104 48852 45126
rect 3878 45064 3884 45076
rect 3839 45036 3884 45064
rect 3878 45024 3884 45036
rect 3936 45024 3942 45076
rect 13170 45064 13176 45076
rect 13131 45036 13176 45064
rect 13170 45024 13176 45036
rect 13228 45024 13234 45076
rect 1394 44928 1400 44940
rect 1355 44900 1400 44928
rect 1394 44888 1400 44900
rect 1452 44888 1458 44940
rect 2774 44928 2780 44940
rect 2735 44900 2780 44928
rect 2774 44888 2780 44900
rect 2832 44888 2838 44940
rect 46474 44928 46480 44940
rect 46435 44900 46480 44928
rect 46474 44888 46480 44900
rect 46532 44888 46538 44940
rect 48130 44928 48136 44940
rect 48091 44900 48136 44928
rect 48130 44888 48136 44900
rect 48188 44888 48194 44940
rect 3786 44860 3792 44872
rect 3747 44832 3792 44860
rect 3786 44820 3792 44832
rect 3844 44820 3850 44872
rect 45186 44860 45192 44872
rect 45147 44832 45192 44860
rect 45186 44820 45192 44832
rect 45244 44820 45250 44872
rect 45833 44863 45891 44869
rect 45833 44829 45845 44863
rect 45879 44860 45891 44863
rect 46293 44863 46351 44869
rect 46293 44860 46305 44863
rect 45879 44832 46305 44860
rect 45879 44829 45891 44832
rect 45833 44823 45891 44829
rect 46293 44829 46305 44832
rect 46339 44829 46351 44863
rect 46293 44823 46351 44829
rect 1581 44795 1639 44801
rect 1581 44761 1593 44795
rect 1627 44792 1639 44795
rect 2774 44792 2780 44804
rect 1627 44764 2780 44792
rect 1627 44761 1639 44764
rect 1581 44755 1639 44761
rect 2774 44752 2780 44764
rect 2832 44752 2838 44804
rect 1104 44634 48852 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 48852 44634
rect 1104 44560 48852 44582
rect 3970 44520 3976 44532
rect 1872 44492 3976 44520
rect 1872 44393 1900 44492
rect 3970 44480 3976 44492
rect 4028 44480 4034 44532
rect 2038 44452 2044 44464
rect 1999 44424 2044 44452
rect 2038 44412 2044 44424
rect 2096 44412 2102 44464
rect 45373 44455 45431 44461
rect 45373 44421 45385 44455
rect 45419 44452 45431 44455
rect 47302 44452 47308 44464
rect 45419 44424 47308 44452
rect 45419 44421 45431 44424
rect 45373 44415 45431 44421
rect 47302 44412 47308 44424
rect 47360 44412 47366 44464
rect 1857 44387 1915 44393
rect 1857 44353 1869 44387
rect 1903 44353 1915 44387
rect 45186 44384 45192 44396
rect 45147 44356 45192 44384
rect 1857 44347 1915 44353
rect 45186 44344 45192 44356
rect 45244 44344 45250 44396
rect 47762 44384 47768 44396
rect 47723 44356 47768 44384
rect 47762 44344 47768 44356
rect 47820 44344 47826 44396
rect 2866 44316 2872 44328
rect 2827 44288 2872 44316
rect 2866 44276 2872 44288
rect 2924 44276 2930 44328
rect 46842 44316 46848 44328
rect 46803 44288 46848 44316
rect 46842 44276 46848 44288
rect 46900 44276 46906 44328
rect 1104 44090 48852 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 48852 44090
rect 1104 44016 48852 44038
rect 2774 43976 2780 43988
rect 2735 43948 2780 43976
rect 2774 43936 2780 43948
rect 2832 43936 2838 43988
rect 1854 43772 1860 43784
rect 1815 43744 1860 43772
rect 1854 43732 1860 43744
rect 1912 43732 1918 43784
rect 2130 43732 2136 43784
rect 2188 43772 2194 43784
rect 2685 43775 2743 43781
rect 2685 43772 2697 43775
rect 2188 43744 2697 43772
rect 2188 43732 2194 43744
rect 2685 43741 2697 43744
rect 2731 43741 2743 43775
rect 2685 43735 2743 43741
rect 45833 43775 45891 43781
rect 45833 43741 45845 43775
rect 45879 43772 45891 43775
rect 46293 43775 46351 43781
rect 46293 43772 46305 43775
rect 45879 43744 46305 43772
rect 45879 43741 45891 43744
rect 45833 43735 45891 43741
rect 46293 43741 46305 43744
rect 46339 43741 46351 43775
rect 46293 43735 46351 43741
rect 46477 43707 46535 43713
rect 46477 43673 46489 43707
rect 46523 43704 46535 43707
rect 46934 43704 46940 43716
rect 46523 43676 46940 43704
rect 46523 43673 46535 43676
rect 46477 43667 46535 43673
rect 46934 43664 46940 43676
rect 46992 43664 46998 43716
rect 48130 43704 48136 43716
rect 48091 43676 48136 43704
rect 48130 43664 48136 43676
rect 48188 43664 48194 43716
rect 1946 43636 1952 43648
rect 1907 43608 1952 43636
rect 1946 43596 1952 43608
rect 2004 43596 2010 43648
rect 1104 43546 48852 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 48852 43546
rect 1104 43472 48852 43494
rect 46934 43432 46940 43444
rect 46895 43404 46940 43432
rect 46934 43392 46940 43404
rect 46992 43392 46998 43444
rect 1854 43364 1860 43376
rect 1815 43336 1860 43364
rect 1854 43324 1860 43336
rect 1912 43324 1918 43376
rect 7926 43256 7932 43308
rect 7984 43296 7990 43308
rect 46845 43299 46903 43305
rect 46845 43296 46857 43299
rect 7984 43268 46857 43296
rect 7984 43256 7990 43268
rect 46845 43265 46857 43268
rect 46891 43265 46903 43299
rect 47854 43296 47860 43308
rect 47815 43268 47860 43296
rect 46845 43259 46903 43265
rect 47854 43256 47860 43268
rect 47912 43256 47918 43308
rect 2133 43095 2191 43101
rect 2133 43061 2145 43095
rect 2179 43092 2191 43095
rect 2222 43092 2228 43104
rect 2179 43064 2228 43092
rect 2179 43061 2191 43064
rect 2133 43055 2191 43061
rect 2222 43052 2228 43064
rect 2280 43052 2286 43104
rect 48041 43095 48099 43101
rect 48041 43061 48053 43095
rect 48087 43092 48099 43095
rect 48222 43092 48228 43104
rect 48087 43064 48228 43092
rect 48087 43061 48099 43064
rect 48041 43055 48099 43061
rect 48222 43052 48228 43064
rect 48280 43052 48286 43104
rect 1104 43002 48852 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 48852 43002
rect 1104 42928 48852 42950
rect 47302 42752 47308 42764
rect 47263 42724 47308 42752
rect 47302 42712 47308 42724
rect 47360 42712 47366 42764
rect 47210 42684 47216 42696
rect 47171 42656 47216 42684
rect 47210 42644 47216 42656
rect 47268 42644 47274 42696
rect 47946 42616 47952 42628
rect 26206 42588 47440 42616
rect 47907 42588 47952 42616
rect 22646 42508 22652 42560
rect 22704 42548 22710 42560
rect 26206 42548 26234 42588
rect 22704 42520 26234 42548
rect 47412 42548 47440 42588
rect 47946 42576 47952 42588
rect 48004 42576 48010 42628
rect 48041 42551 48099 42557
rect 48041 42548 48053 42551
rect 47412 42520 48053 42548
rect 22704 42508 22710 42520
rect 48041 42517 48053 42520
rect 48087 42517 48099 42551
rect 48041 42511 48099 42517
rect 1104 42458 48852 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 48852 42458
rect 1104 42384 48852 42406
rect 46750 42208 46756 42220
rect 46711 42180 46756 42208
rect 46750 42168 46756 42180
rect 46808 42168 46814 42220
rect 20438 42032 20444 42084
rect 20496 42072 20502 42084
rect 20622 42072 20628 42084
rect 20496 42044 20628 42072
rect 20496 42032 20502 42044
rect 20622 42032 20628 42044
rect 20680 42032 20686 42084
rect 1394 41964 1400 42016
rect 1452 42004 1458 42016
rect 2041 42007 2099 42013
rect 2041 42004 2053 42007
rect 1452 41976 2053 42004
rect 1452 41964 1458 41976
rect 2041 41973 2053 41976
rect 2087 41973 2099 42007
rect 2041 41967 2099 41973
rect 46474 41964 46480 42016
rect 46532 42004 46538 42016
rect 46845 42007 46903 42013
rect 46845 42004 46857 42007
rect 46532 41976 46857 42004
rect 46532 41964 46538 41976
rect 46845 41973 46857 41976
rect 46891 41973 46903 42007
rect 47762 42004 47768 42016
rect 47723 41976 47768 42004
rect 46845 41967 46903 41973
rect 47762 41964 47768 41976
rect 47820 41964 47826 42016
rect 1104 41914 48852 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 48852 41914
rect 1104 41840 48852 41862
rect 47762 41732 47768 41744
rect 46308 41704 47768 41732
rect 1394 41664 1400 41676
rect 1355 41636 1400 41664
rect 1394 41624 1400 41636
rect 1452 41624 1458 41676
rect 1854 41664 1860 41676
rect 1815 41636 1860 41664
rect 1854 41624 1860 41636
rect 1912 41624 1918 41676
rect 46308 41673 46336 41704
rect 47762 41692 47768 41704
rect 47820 41692 47826 41744
rect 46293 41667 46351 41673
rect 46293 41633 46305 41667
rect 46339 41633 46351 41667
rect 46474 41664 46480 41676
rect 46435 41636 46480 41664
rect 46293 41627 46351 41633
rect 46474 41624 46480 41636
rect 46532 41624 46538 41676
rect 21082 41556 21088 41608
rect 21140 41596 21146 41608
rect 24118 41596 24124 41608
rect 21140 41568 24124 41596
rect 21140 41556 21146 41568
rect 24118 41556 24124 41568
rect 24176 41556 24182 41608
rect 1578 41528 1584 41540
rect 1539 41500 1584 41528
rect 1578 41488 1584 41500
rect 1636 41488 1642 41540
rect 48130 41528 48136 41540
rect 48091 41500 48136 41528
rect 48130 41488 48136 41500
rect 48188 41488 48194 41540
rect 1104 41370 48852 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 48852 41370
rect 1104 41296 48852 41318
rect 1578 41216 1584 41268
rect 1636 41256 1642 41268
rect 2593 41259 2651 41265
rect 2593 41256 2605 41259
rect 1636 41228 2605 41256
rect 1636 41216 1642 41228
rect 2593 41225 2605 41228
rect 2639 41225 2651 41259
rect 2593 41219 2651 41225
rect 1854 41120 1860 41132
rect 1815 41092 1860 41120
rect 1854 41080 1860 41092
rect 1912 41080 1918 41132
rect 2501 41123 2559 41129
rect 2501 41089 2513 41123
rect 2547 41089 2559 41123
rect 2501 41083 2559 41089
rect 1486 41012 1492 41064
rect 1544 41052 1550 41064
rect 2516 41052 2544 41083
rect 45738 41080 45744 41132
rect 45796 41120 45802 41132
rect 46477 41123 46535 41129
rect 46477 41120 46489 41123
rect 45796 41092 46489 41120
rect 45796 41080 45802 41092
rect 46477 41089 46489 41092
rect 46523 41089 46535 41123
rect 46477 41083 46535 41089
rect 46198 41052 46204 41064
rect 1544 41024 2544 41052
rect 46159 41024 46204 41052
rect 1544 41012 1550 41024
rect 46198 41012 46204 41024
rect 46256 41012 46262 41064
rect 2041 40987 2099 40993
rect 2041 40953 2053 40987
rect 2087 40984 2099 40987
rect 2314 40984 2320 40996
rect 2087 40956 2320 40984
rect 2087 40953 2099 40956
rect 2041 40947 2099 40953
rect 2314 40944 2320 40956
rect 2372 40944 2378 40996
rect 46290 40876 46296 40928
rect 46348 40916 46354 40928
rect 47765 40919 47823 40925
rect 47765 40916 47777 40919
rect 46348 40888 47777 40916
rect 46348 40876 46354 40888
rect 47765 40885 47777 40888
rect 47811 40885 47823 40919
rect 47765 40879 47823 40885
rect 1104 40826 48852 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 48852 40826
rect 1104 40752 48852 40774
rect 21818 40536 21824 40588
rect 21876 40576 21882 40588
rect 23382 40576 23388 40588
rect 21876 40548 23388 40576
rect 21876 40536 21882 40548
rect 1394 40508 1400 40520
rect 1355 40480 1400 40508
rect 1394 40468 1400 40480
rect 1452 40468 1458 40520
rect 22646 40508 22652 40520
rect 22607 40480 22652 40508
rect 22646 40468 22652 40480
rect 22704 40468 22710 40520
rect 22756 40517 22784 40548
rect 23382 40536 23388 40548
rect 23440 40536 23446 40588
rect 46290 40576 46296 40588
rect 46251 40548 46296 40576
rect 46290 40536 46296 40548
rect 46348 40536 46354 40588
rect 22741 40511 22799 40517
rect 22741 40477 22753 40511
rect 22787 40477 22799 40511
rect 22741 40471 22799 40477
rect 22833 40511 22891 40517
rect 22833 40477 22845 40511
rect 22879 40477 22891 40511
rect 22833 40471 22891 40477
rect 23017 40511 23075 40517
rect 23017 40477 23029 40511
rect 23063 40508 23075 40511
rect 23842 40508 23848 40520
rect 23063 40480 23848 40508
rect 23063 40477 23075 40480
rect 23017 40471 23075 40477
rect 22462 40400 22468 40452
rect 22520 40440 22526 40452
rect 22848 40440 22876 40471
rect 23842 40468 23848 40480
rect 23900 40468 23906 40520
rect 22520 40412 22876 40440
rect 46477 40443 46535 40449
rect 22520 40400 22526 40412
rect 46477 40409 46489 40443
rect 46523 40440 46535 40443
rect 47670 40440 47676 40452
rect 46523 40412 47676 40440
rect 46523 40409 46535 40412
rect 46477 40403 46535 40409
rect 47670 40400 47676 40412
rect 47728 40400 47734 40452
rect 48130 40440 48136 40452
rect 48091 40412 48136 40440
rect 48130 40400 48136 40412
rect 48188 40400 48194 40452
rect 1578 40372 1584 40384
rect 1539 40344 1584 40372
rect 1578 40332 1584 40344
rect 1636 40332 1642 40384
rect 22370 40372 22376 40384
rect 22331 40344 22376 40372
rect 22370 40332 22376 40344
rect 22428 40332 22434 40384
rect 1104 40282 48852 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 48852 40282
rect 1104 40208 48852 40230
rect 21177 40171 21235 40177
rect 21177 40137 21189 40171
rect 21223 40168 21235 40171
rect 22646 40168 22652 40180
rect 21223 40140 22652 40168
rect 21223 40137 21235 40140
rect 21177 40131 21235 40137
rect 22646 40128 22652 40140
rect 22704 40128 22710 40180
rect 23201 40171 23259 40177
rect 23201 40137 23213 40171
rect 23247 40168 23259 40171
rect 24026 40168 24032 40180
rect 23247 40140 24032 40168
rect 23247 40137 23259 40140
rect 23201 40131 23259 40137
rect 24026 40128 24032 40140
rect 24084 40128 24090 40180
rect 22088 40103 22146 40109
rect 22088 40069 22100 40103
rect 22134 40100 22146 40103
rect 22370 40100 22376 40112
rect 22134 40072 22376 40100
rect 22134 40069 22146 40072
rect 22088 40063 22146 40069
rect 22370 40060 22376 40072
rect 22428 40060 22434 40112
rect 20990 40032 20996 40044
rect 20951 40004 20996 40032
rect 20990 39992 20996 40004
rect 21048 39992 21054 40044
rect 21266 40032 21272 40044
rect 21227 40004 21272 40032
rect 21266 39992 21272 40004
rect 21324 39992 21330 40044
rect 23106 39992 23112 40044
rect 23164 40032 23170 40044
rect 23917 40035 23975 40041
rect 23917 40032 23929 40035
rect 23164 40004 23929 40032
rect 23164 39992 23170 40004
rect 23917 40001 23929 40004
rect 23963 40001 23975 40035
rect 23917 39995 23975 40001
rect 44542 39992 44548 40044
rect 44600 40032 44606 40044
rect 47302 40032 47308 40044
rect 44600 40004 47308 40032
rect 44600 39992 44606 40004
rect 47302 39992 47308 40004
rect 47360 40032 47366 40044
rect 47581 40035 47639 40041
rect 47581 40032 47593 40035
rect 47360 40004 47593 40032
rect 47360 39992 47366 40004
rect 47581 40001 47593 40004
rect 47627 40001 47639 40035
rect 47581 39995 47639 40001
rect 47670 39992 47676 40044
rect 47728 40032 47734 40044
rect 47728 40004 47773 40032
rect 47728 39992 47734 40004
rect 20438 39924 20444 39976
rect 20496 39964 20502 39976
rect 21821 39967 21879 39973
rect 21821 39964 21833 39967
rect 20496 39936 21833 39964
rect 20496 39924 20502 39936
rect 21821 39933 21833 39936
rect 21867 39933 21879 39967
rect 23658 39964 23664 39976
rect 23619 39936 23664 39964
rect 21821 39927 21879 39933
rect 23658 39924 23664 39936
rect 23716 39924 23722 39976
rect 18874 39856 18880 39908
rect 18932 39896 18938 39908
rect 18932 39868 21036 39896
rect 18932 39856 18938 39868
rect 20809 39831 20867 39837
rect 20809 39797 20821 39831
rect 20855 39828 20867 39831
rect 20898 39828 20904 39840
rect 20855 39800 20904 39828
rect 20855 39797 20867 39800
rect 20809 39791 20867 39797
rect 20898 39788 20904 39800
rect 20956 39788 20962 39840
rect 21008 39828 21036 39868
rect 23124 39868 23336 39896
rect 23124 39828 23152 39868
rect 21008 39800 23152 39828
rect 23308 39828 23336 39868
rect 24394 39828 24400 39840
rect 23308 39800 24400 39828
rect 24394 39788 24400 39800
rect 24452 39788 24458 39840
rect 25038 39828 25044 39840
rect 24999 39800 25044 39828
rect 25038 39788 25044 39800
rect 25096 39788 25102 39840
rect 1104 39738 48852 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 48852 39738
rect 1104 39664 48852 39686
rect 23106 39624 23112 39636
rect 23067 39596 23112 39624
rect 23106 39584 23112 39596
rect 23164 39584 23170 39636
rect 23934 39624 23940 39636
rect 23216 39596 23940 39624
rect 23216 39556 23244 39596
rect 23934 39584 23940 39596
rect 23992 39584 23998 39636
rect 23124 39528 23244 39556
rect 20438 39488 20444 39500
rect 20399 39460 20444 39488
rect 20438 39448 20444 39460
rect 20496 39448 20502 39500
rect 2038 39380 2044 39432
rect 2096 39420 2102 39432
rect 2225 39423 2283 39429
rect 2225 39420 2237 39423
rect 2096 39392 2237 39420
rect 2096 39380 2102 39392
rect 2225 39389 2237 39392
rect 2271 39389 2283 39423
rect 2225 39383 2283 39389
rect 17405 39423 17463 39429
rect 17405 39389 17417 39423
rect 17451 39420 17463 39423
rect 18230 39420 18236 39432
rect 17451 39392 18236 39420
rect 17451 39389 17463 39392
rect 17405 39383 17463 39389
rect 18230 39380 18236 39392
rect 18288 39380 18294 39432
rect 18322 39380 18328 39432
rect 18380 39420 18386 39432
rect 18380 39392 18425 39420
rect 18380 39380 18386 39392
rect 20714 39361 20720 39364
rect 20708 39315 20720 39361
rect 20772 39352 20778 39364
rect 23124 39352 23152 39528
rect 23382 39516 23388 39568
rect 23440 39556 23446 39568
rect 23750 39556 23756 39568
rect 23440 39528 23756 39556
rect 23440 39516 23446 39528
rect 23492 39429 23520 39528
rect 23750 39516 23756 39528
rect 23808 39516 23814 39568
rect 23658 39448 23664 39500
rect 23716 39488 23722 39500
rect 23716 39460 24440 39488
rect 23716 39448 23722 39460
rect 23385 39423 23443 39429
rect 23385 39389 23397 39423
rect 23431 39389 23443 39423
rect 23385 39383 23443 39389
rect 23474 39423 23532 39429
rect 23474 39389 23486 39423
rect 23520 39389 23532 39423
rect 23474 39383 23532 39389
rect 23400 39352 23428 39383
rect 23566 39380 23572 39432
rect 23624 39420 23630 39432
rect 23753 39423 23811 39429
rect 23624 39392 23669 39420
rect 23624 39380 23630 39392
rect 23753 39389 23765 39423
rect 23799 39420 23811 39423
rect 23842 39420 23848 39432
rect 23799 39392 23848 39420
rect 23799 39389 23811 39392
rect 23753 39383 23811 39389
rect 23842 39380 23848 39392
rect 23900 39380 23906 39432
rect 24412 39429 24440 39460
rect 24397 39423 24455 39429
rect 24397 39389 24409 39423
rect 24443 39420 24455 39423
rect 26694 39420 26700 39432
rect 24443 39392 26700 39420
rect 24443 39389 24455 39392
rect 24397 39383 24455 39389
rect 26694 39380 26700 39392
rect 26752 39420 26758 39432
rect 26881 39423 26939 39429
rect 26881 39420 26893 39423
rect 26752 39392 26893 39420
rect 26752 39380 26758 39392
rect 26881 39389 26893 39392
rect 26927 39389 26939 39423
rect 47670 39420 47676 39432
rect 47631 39392 47676 39420
rect 26881 39383 26939 39389
rect 47670 39380 47676 39392
rect 47728 39380 47734 39432
rect 20772 39324 20808 39352
rect 23124 39324 23428 39352
rect 20714 39312 20720 39315
rect 20772 39312 20778 39324
rect 23658 39312 23664 39364
rect 23716 39352 23722 39364
rect 24642 39355 24700 39361
rect 24642 39352 24654 39355
rect 23716 39324 24654 39352
rect 23716 39312 23722 39324
rect 24642 39321 24654 39324
rect 24688 39321 24700 39355
rect 24642 39315 24700 39321
rect 26970 39312 26976 39364
rect 27028 39352 27034 39364
rect 27126 39355 27184 39361
rect 27126 39352 27138 39355
rect 27028 39324 27138 39352
rect 27028 39312 27034 39324
rect 27126 39321 27138 39324
rect 27172 39321 27184 39355
rect 27126 39315 27184 39321
rect 17218 39244 17224 39296
rect 17276 39284 17282 39296
rect 17589 39287 17647 39293
rect 17589 39284 17601 39287
rect 17276 39256 17601 39284
rect 17276 39244 17282 39256
rect 17589 39253 17601 39256
rect 17635 39253 17647 39287
rect 17589 39247 17647 39253
rect 18417 39287 18475 39293
rect 18417 39253 18429 39287
rect 18463 39284 18475 39287
rect 19426 39284 19432 39296
rect 18463 39256 19432 39284
rect 18463 39253 18475 39256
rect 18417 39247 18475 39253
rect 19426 39244 19432 39256
rect 19484 39244 19490 39296
rect 21266 39244 21272 39296
rect 21324 39284 21330 39296
rect 21821 39287 21879 39293
rect 21821 39284 21833 39287
rect 21324 39256 21833 39284
rect 21324 39244 21330 39256
rect 21821 39253 21833 39256
rect 21867 39284 21879 39287
rect 22002 39284 22008 39296
rect 21867 39256 22008 39284
rect 21867 39253 21879 39256
rect 21821 39247 21879 39253
rect 22002 39244 22008 39256
rect 22060 39244 22066 39296
rect 23014 39244 23020 39296
rect 23072 39284 23078 39296
rect 25038 39284 25044 39296
rect 23072 39256 25044 39284
rect 23072 39244 23078 39256
rect 25038 39244 25044 39256
rect 25096 39244 25102 39296
rect 25774 39284 25780 39296
rect 25735 39256 25780 39284
rect 25774 39244 25780 39256
rect 25832 39244 25838 39296
rect 28261 39287 28319 39293
rect 28261 39253 28273 39287
rect 28307 39284 28319 39287
rect 29270 39284 29276 39296
rect 28307 39256 29276 39284
rect 28307 39253 28319 39256
rect 28261 39247 28319 39253
rect 29270 39244 29276 39256
rect 29328 39244 29334 39296
rect 1104 39194 48852 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 48852 39194
rect 1104 39120 48852 39142
rect 20441 39083 20499 39089
rect 20441 39049 20453 39083
rect 20487 39080 20499 39083
rect 20714 39080 20720 39092
rect 20487 39052 20720 39080
rect 20487 39049 20499 39052
rect 20441 39043 20499 39049
rect 20714 39040 20720 39052
rect 20772 39040 20778 39092
rect 22646 39080 22652 39092
rect 22607 39052 22652 39080
rect 22646 39040 22652 39052
rect 22704 39040 22710 39092
rect 23201 39083 23259 39089
rect 23201 39049 23213 39083
rect 23247 39080 23259 39083
rect 23290 39080 23296 39092
rect 23247 39052 23296 39080
rect 23247 39049 23259 39052
rect 23201 39043 23259 39049
rect 23290 39040 23296 39052
rect 23348 39040 23354 39092
rect 23474 39040 23480 39092
rect 23532 39040 23538 39092
rect 26970 39080 26976 39092
rect 26931 39052 26976 39080
rect 26970 39040 26976 39052
rect 27028 39040 27034 39092
rect 48041 39083 48099 39089
rect 48041 39080 48053 39083
rect 31726 39052 48053 39080
rect 2958 38972 2964 39024
rect 3016 39012 3022 39024
rect 21818 39012 21824 39024
rect 3016 38984 20760 39012
rect 3016 38972 3022 38984
rect 2038 38944 2044 38956
rect 1999 38916 2044 38944
rect 2038 38904 2044 38916
rect 2096 38904 2102 38956
rect 17218 38944 17224 38956
rect 17179 38916 17224 38944
rect 17218 38904 17224 38916
rect 17276 38904 17282 38956
rect 18598 38944 18604 38956
rect 18559 38916 18604 38944
rect 18598 38904 18604 38916
rect 18656 38904 18662 38956
rect 20732 38953 20760 38984
rect 20824 38984 21824 39012
rect 20824 38953 20852 38984
rect 21818 38972 21824 38984
rect 21876 38972 21882 39024
rect 20717 38947 20775 38953
rect 20717 38913 20729 38947
rect 20763 38913 20775 38947
rect 20717 38907 20775 38913
rect 20809 38947 20867 38953
rect 20809 38913 20821 38947
rect 20855 38913 20867 38947
rect 20809 38907 20867 38913
rect 20898 38904 20904 38956
rect 20956 38944 20962 38956
rect 20956 38916 21001 38944
rect 20956 38904 20962 38916
rect 21082 38904 21088 38956
rect 21140 38944 21146 38956
rect 22465 38947 22523 38953
rect 21140 38916 21185 38944
rect 21140 38904 21146 38916
rect 22465 38913 22477 38947
rect 22511 38944 22523 38947
rect 22554 38944 22560 38956
rect 22511 38916 22560 38944
rect 22511 38913 22523 38916
rect 22465 38907 22523 38913
rect 22554 38904 22560 38916
rect 22612 38904 22618 38956
rect 22741 38947 22799 38953
rect 22741 38913 22753 38947
rect 22787 38944 22799 38947
rect 23014 38944 23020 38956
rect 22787 38916 23020 38944
rect 22787 38913 22799 38916
rect 22741 38907 22799 38913
rect 23014 38904 23020 38916
rect 23072 38904 23078 38956
rect 23492 38953 23520 39040
rect 23934 39012 23940 39024
rect 23768 38984 23940 39012
rect 23457 38947 23520 38953
rect 23457 38913 23469 38947
rect 23503 38916 23520 38947
rect 23569 38947 23627 38953
rect 23503 38913 23515 38916
rect 23457 38907 23515 38913
rect 23569 38913 23581 38947
rect 23615 38913 23627 38947
rect 23569 38907 23627 38913
rect 23661 38947 23719 38953
rect 23768 38947 23796 38984
rect 23934 38972 23940 38984
rect 23992 38972 23998 39024
rect 26694 39012 26700 39024
rect 25056 38984 26700 39012
rect 25056 38953 25084 38984
rect 26694 38972 26700 38984
rect 26752 38972 26758 39024
rect 26786 38972 26792 39024
rect 26844 39012 26850 39024
rect 31726 39012 31754 39052
rect 48041 39049 48053 39052
rect 48087 39049 48099 39083
rect 48041 39043 48099 39049
rect 26844 38984 31754 39012
rect 26844 38972 26850 38984
rect 23661 38913 23673 38947
rect 23707 38919 23796 38947
rect 23845 38947 23903 38953
rect 23707 38913 23719 38919
rect 23661 38907 23719 38913
rect 23845 38913 23857 38947
rect 23891 38913 23903 38947
rect 23845 38907 23903 38913
rect 25041 38947 25099 38953
rect 25041 38913 25053 38947
rect 25087 38913 25099 38947
rect 25041 38907 25099 38913
rect 2225 38879 2283 38885
rect 2225 38845 2237 38879
rect 2271 38876 2283 38879
rect 2958 38876 2964 38888
rect 2271 38848 2964 38876
rect 2271 38845 2283 38848
rect 2225 38839 2283 38845
rect 2958 38836 2964 38848
rect 3016 38836 3022 38888
rect 3050 38836 3056 38888
rect 3108 38876 3114 38888
rect 18874 38876 18880 38888
rect 3108 38848 3153 38876
rect 18835 38848 18880 38876
rect 3108 38836 3114 38848
rect 18874 38836 18880 38848
rect 18932 38836 18938 38888
rect 22281 38879 22339 38885
rect 22281 38845 22293 38879
rect 22327 38876 22339 38879
rect 23198 38876 23204 38888
rect 22327 38848 23204 38876
rect 22327 38845 22339 38848
rect 22281 38839 22339 38845
rect 23198 38836 23204 38848
rect 23256 38836 23262 38888
rect 23584 38876 23612 38907
rect 23750 38876 23756 38888
rect 23584 38848 23756 38876
rect 23750 38836 23756 38848
rect 23808 38836 23814 38888
rect 23860 38820 23888 38907
rect 25130 38904 25136 38956
rect 25188 38944 25194 38956
rect 25297 38947 25355 38953
rect 25297 38944 25309 38947
rect 25188 38916 25309 38944
rect 25188 38904 25194 38916
rect 25297 38913 25309 38916
rect 25343 38913 25355 38947
rect 27249 38947 27307 38953
rect 27249 38944 27261 38947
rect 25297 38907 25355 38913
rect 26068 38916 27261 38944
rect 13722 38768 13728 38820
rect 13780 38808 13786 38820
rect 13780 38780 20116 38808
rect 13780 38768 13786 38780
rect 17497 38743 17555 38749
rect 17497 38709 17509 38743
rect 17543 38740 17555 38743
rect 18322 38740 18328 38752
rect 17543 38712 18328 38740
rect 17543 38709 17555 38712
rect 17497 38703 17555 38709
rect 18322 38700 18328 38712
rect 18380 38700 18386 38752
rect 19978 38740 19984 38752
rect 19939 38712 19984 38740
rect 19978 38700 19984 38712
rect 20036 38700 20042 38752
rect 20088 38740 20116 38780
rect 21082 38768 21088 38820
rect 21140 38808 21146 38820
rect 23842 38808 23848 38820
rect 21140 38780 23848 38808
rect 21140 38768 21146 38780
rect 23842 38768 23848 38780
rect 23900 38768 23906 38820
rect 26068 38740 26096 38916
rect 27249 38913 27261 38916
rect 27295 38913 27307 38947
rect 27249 38907 27307 38913
rect 27341 38947 27399 38953
rect 27341 38913 27353 38947
rect 27387 38913 27399 38947
rect 27341 38907 27399 38913
rect 27433 38947 27491 38953
rect 27433 38913 27445 38947
rect 27479 38944 27491 38947
rect 27522 38944 27528 38956
rect 27479 38916 27528 38944
rect 27479 38913 27491 38916
rect 27433 38907 27491 38913
rect 26234 38836 26240 38888
rect 26292 38876 26298 38888
rect 27356 38876 27384 38907
rect 27522 38904 27528 38916
rect 27580 38904 27586 38956
rect 27617 38947 27675 38953
rect 27617 38913 27629 38947
rect 27663 38913 27675 38947
rect 27617 38907 27675 38913
rect 26292 38848 27384 38876
rect 26292 38836 26298 38848
rect 26142 38768 26148 38820
rect 26200 38808 26206 38820
rect 27632 38808 27660 38907
rect 30190 38904 30196 38956
rect 30248 38944 30254 38956
rect 30377 38947 30435 38953
rect 30377 38944 30389 38947
rect 30248 38916 30389 38944
rect 30248 38904 30254 38916
rect 30377 38913 30389 38916
rect 30423 38913 30435 38947
rect 30377 38907 30435 38913
rect 30561 38947 30619 38953
rect 30561 38913 30573 38947
rect 30607 38944 30619 38947
rect 30926 38944 30932 38956
rect 30607 38916 30932 38944
rect 30607 38913 30619 38916
rect 30561 38907 30619 38913
rect 30926 38904 30932 38916
rect 30984 38904 30990 38956
rect 47946 38944 47952 38956
rect 47907 38916 47952 38944
rect 47946 38904 47952 38916
rect 48004 38904 48010 38956
rect 26200 38780 27660 38808
rect 26200 38768 26206 38780
rect 26418 38740 26424 38752
rect 20088 38712 26096 38740
rect 26379 38712 26424 38740
rect 26418 38700 26424 38712
rect 26476 38700 26482 38752
rect 30745 38743 30803 38749
rect 30745 38709 30757 38743
rect 30791 38740 30803 38743
rect 31110 38740 31116 38752
rect 30791 38712 31116 38740
rect 30791 38709 30803 38712
rect 30745 38703 30803 38709
rect 31110 38700 31116 38712
rect 31168 38700 31174 38752
rect 1104 38650 48852 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 48852 38650
rect 1104 38576 48852 38598
rect 2958 38536 2964 38548
rect 2919 38508 2964 38536
rect 2958 38496 2964 38508
rect 3016 38496 3022 38548
rect 21818 38536 21824 38548
rect 21779 38508 21824 38536
rect 21818 38496 21824 38508
rect 21876 38496 21882 38548
rect 22373 38539 22431 38545
rect 22373 38505 22385 38539
rect 22419 38536 22431 38539
rect 22462 38536 22468 38548
rect 22419 38508 22468 38536
rect 22419 38505 22431 38508
rect 22373 38499 22431 38505
rect 22462 38496 22468 38508
rect 22520 38496 22526 38548
rect 38746 38536 38752 38548
rect 22664 38508 38752 38536
rect 22664 38468 22692 38508
rect 38746 38496 38752 38508
rect 38804 38496 38810 38548
rect 18156 38440 22692 38468
rect 23293 38471 23351 38477
rect 18156 38409 18184 38440
rect 23293 38437 23305 38471
rect 23339 38468 23351 38471
rect 23934 38468 23940 38480
rect 23339 38440 23940 38468
rect 23339 38437 23351 38440
rect 23293 38431 23351 38437
rect 23934 38428 23940 38440
rect 23992 38428 23998 38480
rect 24765 38471 24823 38477
rect 24765 38437 24777 38471
rect 24811 38468 24823 38471
rect 25130 38468 25136 38480
rect 24811 38440 25136 38468
rect 24811 38437 24823 38440
rect 24765 38431 24823 38437
rect 25130 38428 25136 38440
rect 25188 38428 25194 38480
rect 35158 38428 35164 38480
rect 35216 38468 35222 38480
rect 39298 38468 39304 38480
rect 35216 38440 39304 38468
rect 35216 38428 35222 38440
rect 39298 38428 39304 38440
rect 39356 38428 39362 38480
rect 18141 38403 18199 38409
rect 18141 38369 18153 38403
rect 18187 38369 18199 38403
rect 19426 38400 19432 38412
rect 19387 38372 19432 38400
rect 18141 38363 18199 38369
rect 19426 38360 19432 38372
rect 19484 38360 19490 38412
rect 20990 38360 20996 38412
rect 21048 38400 21054 38412
rect 21634 38400 21640 38412
rect 21048 38372 21640 38400
rect 21048 38360 21054 38372
rect 21634 38360 21640 38372
rect 21692 38400 21698 38412
rect 21692 38372 22600 38400
rect 21692 38360 21698 38372
rect 2869 38335 2927 38341
rect 2869 38301 2881 38335
rect 2915 38332 2927 38335
rect 8938 38332 8944 38344
rect 2915 38304 8944 38332
rect 2915 38301 2927 38304
rect 2869 38295 2927 38301
rect 8938 38292 8944 38304
rect 8996 38292 9002 38344
rect 15657 38335 15715 38341
rect 15657 38301 15669 38335
rect 15703 38301 15715 38335
rect 15657 38295 15715 38301
rect 6914 38224 6920 38276
rect 6972 38264 6978 38276
rect 15562 38264 15568 38276
rect 6972 38236 15568 38264
rect 6972 38224 6978 38236
rect 15562 38224 15568 38236
rect 15620 38224 15626 38276
rect 15672 38196 15700 38295
rect 16114 38292 16120 38344
rect 16172 38332 16178 38344
rect 16301 38335 16359 38341
rect 16301 38332 16313 38335
rect 16172 38304 16313 38332
rect 16172 38292 16178 38304
rect 16301 38301 16313 38304
rect 16347 38301 16359 38335
rect 19242 38332 19248 38344
rect 19203 38304 19248 38332
rect 16301 38295 16359 38301
rect 19242 38292 19248 38304
rect 19300 38292 19306 38344
rect 22572 38341 22600 38372
rect 22646 38360 22652 38412
rect 22704 38400 22710 38412
rect 22922 38400 22928 38412
rect 22704 38372 22928 38400
rect 22704 38360 22710 38372
rect 22922 38360 22928 38372
rect 22980 38360 22986 38412
rect 24026 38400 24032 38412
rect 23400 38372 24032 38400
rect 21085 38335 21143 38341
rect 21085 38301 21097 38335
rect 21131 38332 21143 38335
rect 22557 38335 22615 38341
rect 21131 38304 22508 38332
rect 21131 38301 21143 38304
rect 21085 38295 21143 38301
rect 15749 38267 15807 38273
rect 15749 38233 15761 38267
rect 15795 38264 15807 38267
rect 16485 38267 16543 38273
rect 16485 38264 16497 38267
rect 15795 38236 16497 38264
rect 15795 38233 15807 38236
rect 15749 38227 15807 38233
rect 16485 38233 16497 38236
rect 16531 38233 16543 38267
rect 16485 38227 16543 38233
rect 17402 38224 17408 38276
rect 17460 38264 17466 38276
rect 21729 38267 21787 38273
rect 17460 38236 18460 38264
rect 17460 38224 17466 38236
rect 18322 38196 18328 38208
rect 15672 38168 18328 38196
rect 18322 38156 18328 38168
rect 18380 38156 18386 38208
rect 18432 38196 18460 38236
rect 21729 38233 21741 38267
rect 21775 38264 21787 38267
rect 22370 38264 22376 38276
rect 21775 38236 22376 38264
rect 21775 38233 21787 38236
rect 21729 38227 21787 38233
rect 22370 38224 22376 38236
rect 22428 38224 22434 38276
rect 22480 38264 22508 38304
rect 22557 38301 22569 38335
rect 22603 38301 22615 38335
rect 22738 38332 22744 38344
rect 22699 38304 22744 38332
rect 22557 38295 22615 38301
rect 22738 38292 22744 38304
rect 22796 38292 22802 38344
rect 22833 38335 22891 38341
rect 22833 38301 22845 38335
rect 22879 38332 22891 38335
rect 23400 38332 23428 38372
rect 24026 38360 24032 38372
rect 24084 38360 24090 38412
rect 25774 38400 25780 38412
rect 24136 38372 25780 38400
rect 22879 38304 23428 38332
rect 22879 38301 22891 38304
rect 22833 38295 22891 38301
rect 23474 38292 23480 38344
rect 23532 38332 23538 38344
rect 23753 38335 23811 38341
rect 23532 38304 23577 38332
rect 23532 38292 23538 38304
rect 23753 38301 23765 38335
rect 23799 38332 23811 38335
rect 24136 38332 24164 38372
rect 25774 38360 25780 38372
rect 25832 38360 25838 38412
rect 31294 38360 31300 38412
rect 31352 38400 31358 38412
rect 46293 38403 46351 38409
rect 31352 38372 31791 38400
rect 31352 38360 31358 38372
rect 23799 38304 24164 38332
rect 23799 38301 23811 38304
rect 23753 38295 23811 38301
rect 24210 38292 24216 38344
rect 24268 38332 24274 38344
rect 25041 38335 25099 38341
rect 25041 38332 25053 38335
rect 24268 38304 25053 38332
rect 24268 38292 24274 38304
rect 25041 38301 25053 38304
rect 25087 38301 25099 38335
rect 25041 38295 25099 38301
rect 25133 38335 25191 38341
rect 25133 38301 25145 38335
rect 25179 38301 25191 38335
rect 25133 38295 25191 38301
rect 25148 38264 25176 38295
rect 25222 38292 25228 38344
rect 25280 38332 25286 38344
rect 25409 38335 25467 38341
rect 25280 38304 25325 38332
rect 25280 38292 25286 38304
rect 25409 38301 25421 38335
rect 25455 38332 25467 38335
rect 26142 38332 26148 38344
rect 25455 38304 26148 38332
rect 25455 38301 25467 38304
rect 25409 38295 25467 38301
rect 26142 38292 26148 38304
rect 26200 38292 26206 38344
rect 26418 38292 26424 38344
rect 26476 38332 26482 38344
rect 29454 38332 29460 38344
rect 26476 38304 29460 38332
rect 26476 38292 26482 38304
rect 29454 38292 29460 38304
rect 29512 38292 29518 38344
rect 29549 38335 29607 38341
rect 29549 38301 29561 38335
rect 29595 38332 29607 38335
rect 31478 38332 31484 38344
rect 29595 38304 31484 38332
rect 29595 38301 29607 38304
rect 29549 38295 29607 38301
rect 31478 38292 31484 38304
rect 31536 38292 31542 38344
rect 31662 38332 31668 38344
rect 31623 38304 31668 38332
rect 31662 38292 31668 38304
rect 31720 38292 31726 38344
rect 31763 38341 31791 38372
rect 46293 38369 46305 38403
rect 46339 38400 46351 38403
rect 47670 38400 47676 38412
rect 46339 38372 47676 38400
rect 46339 38369 46351 38372
rect 46293 38363 46351 38369
rect 47670 38360 47676 38372
rect 47728 38360 47734 38412
rect 48130 38400 48136 38412
rect 48091 38372 48136 38400
rect 48130 38360 48136 38372
rect 48188 38360 48194 38412
rect 31754 38335 31812 38341
rect 31754 38301 31766 38335
rect 31800 38301 31812 38335
rect 31754 38295 31812 38301
rect 31849 38335 31907 38341
rect 31849 38301 31861 38335
rect 31895 38332 31907 38335
rect 31938 38332 31944 38344
rect 31895 38304 31944 38332
rect 31895 38301 31907 38304
rect 31849 38295 31907 38301
rect 31938 38292 31944 38304
rect 31996 38292 32002 38344
rect 32033 38335 32091 38341
rect 32033 38301 32045 38335
rect 32079 38332 32091 38335
rect 32122 38332 32128 38344
rect 32079 38304 32128 38332
rect 32079 38301 32091 38304
rect 32033 38295 32091 38301
rect 32122 38292 32128 38304
rect 32180 38292 32186 38344
rect 25866 38264 25872 38276
rect 22480 38236 23796 38264
rect 25148 38236 25872 38264
rect 22646 38196 22652 38208
rect 18432 38168 22652 38196
rect 22646 38156 22652 38168
rect 22704 38156 22710 38208
rect 22738 38156 22744 38208
rect 22796 38196 22802 38208
rect 23661 38199 23719 38205
rect 23661 38196 23673 38199
rect 22796 38168 23673 38196
rect 22796 38156 22802 38168
rect 23661 38165 23673 38168
rect 23707 38165 23719 38199
rect 23768 38196 23796 38236
rect 25866 38224 25872 38236
rect 25924 38224 25930 38276
rect 27890 38224 27896 38276
rect 27948 38264 27954 38276
rect 29794 38267 29852 38273
rect 29794 38264 29806 38267
rect 27948 38236 29806 38264
rect 27948 38224 27954 38236
rect 29794 38233 29806 38236
rect 29840 38233 29852 38267
rect 31386 38264 31392 38276
rect 31347 38236 31392 38264
rect 29794 38227 29852 38233
rect 31386 38224 31392 38236
rect 31444 38224 31450 38276
rect 38930 38224 38936 38276
rect 38988 38264 38994 38276
rect 46477 38267 46535 38273
rect 46477 38264 46489 38267
rect 38988 38236 46489 38264
rect 38988 38224 38994 38236
rect 46477 38233 46489 38236
rect 46523 38233 46535 38267
rect 46477 38227 46535 38233
rect 29914 38196 29920 38208
rect 23768 38168 29920 38196
rect 23661 38159 23719 38165
rect 29914 38156 29920 38168
rect 29972 38156 29978 38208
rect 30006 38156 30012 38208
rect 30064 38196 30070 38208
rect 30929 38199 30987 38205
rect 30929 38196 30941 38199
rect 30064 38168 30941 38196
rect 30064 38156 30070 38168
rect 30929 38165 30941 38168
rect 30975 38165 30987 38199
rect 30929 38159 30987 38165
rect 32030 38156 32036 38208
rect 32088 38196 32094 38208
rect 46658 38196 46664 38208
rect 32088 38168 46664 38196
rect 32088 38156 32094 38168
rect 46658 38156 46664 38168
rect 46716 38156 46722 38208
rect 1104 38106 48852 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 48852 38106
rect 1104 38032 48852 38054
rect 5258 37952 5264 38004
rect 5316 37992 5322 38004
rect 5316 37964 26280 37992
rect 5316 37952 5322 37964
rect 1486 37884 1492 37936
rect 1544 37924 1550 37936
rect 19702 37924 19708 37936
rect 1544 37896 19708 37924
rect 1544 37884 1550 37896
rect 19702 37884 19708 37896
rect 19760 37884 19766 37936
rect 21818 37884 21824 37936
rect 21876 37924 21882 37936
rect 21876 37896 22229 37924
rect 21876 37884 21882 37896
rect 1854 37856 1860 37868
rect 1815 37828 1860 37856
rect 1854 37816 1860 37828
rect 1912 37816 1918 37868
rect 8938 37856 8944 37868
rect 8899 37828 8944 37856
rect 8938 37816 8944 37828
rect 8996 37816 9002 37868
rect 15657 37859 15715 37865
rect 15657 37825 15669 37859
rect 15703 37856 15715 37859
rect 17218 37856 17224 37868
rect 15703 37828 17224 37856
rect 15703 37825 15715 37828
rect 15657 37819 15715 37825
rect 17218 37816 17224 37828
rect 17276 37816 17282 37868
rect 18598 37856 18604 37868
rect 17328 37828 18000 37856
rect 18559 37828 18604 37856
rect 1670 37748 1676 37800
rect 1728 37788 1734 37800
rect 1728 37760 12434 37788
rect 1728 37748 1734 37760
rect 2041 37723 2099 37729
rect 2041 37689 2053 37723
rect 2087 37720 2099 37723
rect 12406 37720 12434 37760
rect 15562 37748 15568 37800
rect 15620 37788 15626 37800
rect 15841 37791 15899 37797
rect 15841 37788 15853 37791
rect 15620 37760 15853 37788
rect 15620 37748 15626 37760
rect 15841 37757 15853 37760
rect 15887 37757 15899 37791
rect 17328 37788 17356 37828
rect 15841 37751 15899 37757
rect 15948 37760 17356 37788
rect 13998 37720 14004 37732
rect 2087 37692 9251 37720
rect 12406 37692 14004 37720
rect 2087 37689 2099 37692
rect 2041 37683 2099 37689
rect 9033 37655 9091 37661
rect 9033 37621 9045 37655
rect 9079 37652 9091 37655
rect 9122 37652 9128 37664
rect 9079 37624 9128 37652
rect 9079 37621 9091 37624
rect 9033 37615 9091 37621
rect 9122 37612 9128 37624
rect 9180 37612 9186 37664
rect 9223 37652 9251 37692
rect 13998 37680 14004 37692
rect 14056 37680 14062 37732
rect 14090 37680 14096 37732
rect 14148 37720 14154 37732
rect 15948 37720 15976 37760
rect 17402 37748 17408 37800
rect 17460 37788 17466 37800
rect 17972 37788 18000 37828
rect 18598 37816 18604 37828
rect 18656 37856 18662 37868
rect 22201 37865 22229 37896
rect 20441 37859 20499 37865
rect 22077 37859 22135 37865
rect 20441 37856 20453 37859
rect 18656 37828 20453 37856
rect 18656 37816 18662 37828
rect 20441 37825 20453 37828
rect 20487 37825 20499 37859
rect 21928 37856 22048 37859
rect 22077 37856 22089 37859
rect 20441 37819 20499 37825
rect 20548 37831 22089 37856
rect 20548 37828 21956 37831
rect 22020 37828 22089 37831
rect 20548 37788 20576 37828
rect 22077 37825 22089 37828
rect 22123 37825 22135 37859
rect 22077 37819 22135 37825
rect 22170 37859 22229 37865
rect 22170 37825 22182 37859
rect 22216 37828 22229 37859
rect 22216 37825 22228 37828
rect 22170 37819 22228 37825
rect 22278 37816 22284 37868
rect 22336 37856 22342 37868
rect 22336 37828 22381 37856
rect 22336 37816 22342 37828
rect 22462 37816 22468 37868
rect 22520 37856 22526 37868
rect 23014 37856 23020 37868
rect 22520 37828 22565 37856
rect 22975 37828 23020 37856
rect 22520 37816 22526 37828
rect 23014 37816 23020 37828
rect 23072 37816 23078 37868
rect 23198 37856 23204 37868
rect 23159 37828 23204 37856
rect 23198 37816 23204 37828
rect 23256 37856 23262 37868
rect 24854 37856 24860 37868
rect 23256 37828 24860 37856
rect 23256 37816 23262 37828
rect 24854 37816 24860 37828
rect 24912 37816 24918 37868
rect 25406 37856 25412 37868
rect 25367 37828 25412 37856
rect 25406 37816 25412 37828
rect 25464 37816 25470 37868
rect 25593 37859 25651 37865
rect 25593 37825 25605 37859
rect 25639 37825 25651 37859
rect 26252 37856 26280 37964
rect 26326 37952 26332 38004
rect 26384 37992 26390 38004
rect 26384 37964 41414 37992
rect 26384 37952 26390 37964
rect 27890 37924 27896 37936
rect 27851 37896 27896 37924
rect 27890 37884 27896 37896
rect 27948 37884 27954 37936
rect 30653 37927 30711 37933
rect 28000 37896 29500 37924
rect 28000 37856 28028 37896
rect 26252 37828 28028 37856
rect 28169 37859 28227 37865
rect 25593 37819 25651 37825
rect 28169 37825 28181 37859
rect 28215 37825 28227 37859
rect 28169 37819 28227 37825
rect 28258 37859 28316 37865
rect 28258 37825 28270 37859
rect 28304 37825 28316 37859
rect 28258 37819 28316 37825
rect 28353 37859 28411 37865
rect 28353 37825 28365 37859
rect 28399 37825 28411 37859
rect 28353 37819 28411 37825
rect 28537 37859 28595 37865
rect 28537 37825 28549 37859
rect 28583 37856 28595 37859
rect 28902 37856 28908 37868
rect 28583 37828 28908 37856
rect 28583 37825 28595 37828
rect 28537 37819 28595 37825
rect 20714 37788 20720 37800
rect 17460 37760 17505 37788
rect 17972 37760 20576 37788
rect 20675 37760 20720 37788
rect 17460 37748 17466 37760
rect 20714 37748 20720 37760
rect 20772 37748 20778 37800
rect 22554 37748 22560 37800
rect 22612 37788 22618 37800
rect 23382 37788 23388 37800
rect 22612 37760 23388 37788
rect 22612 37748 22618 37760
rect 23382 37748 23388 37760
rect 23440 37748 23446 37800
rect 24872 37788 24900 37816
rect 25608 37788 25636 37819
rect 26050 37788 26056 37800
rect 24872 37760 26056 37788
rect 26050 37748 26056 37760
rect 26108 37748 26114 37800
rect 28184 37720 28212 37819
rect 14148 37692 15976 37720
rect 17052 37692 22232 37720
rect 14148 37680 14154 37692
rect 17052 37652 17080 37692
rect 21818 37652 21824 37664
rect 9223 37624 17080 37652
rect 21779 37624 21824 37652
rect 21818 37612 21824 37624
rect 21876 37612 21882 37664
rect 22204 37652 22232 37692
rect 23216 37692 28212 37720
rect 28273 37720 28301 37819
rect 28368 37788 28396 37819
rect 28902 37816 28908 37828
rect 28960 37816 28966 37868
rect 29362 37856 29368 37868
rect 29323 37828 29368 37856
rect 29362 37816 29368 37828
rect 29420 37816 29426 37868
rect 29472 37856 29500 37896
rect 30653 37893 30665 37927
rect 30699 37924 30711 37927
rect 41386 37924 41414 37964
rect 47026 37924 47032 37936
rect 30699 37896 31432 37924
rect 41386 37896 47032 37924
rect 30699 37893 30711 37896
rect 30653 37887 30711 37893
rect 30929 37859 30987 37865
rect 30929 37856 30941 37859
rect 29472 37828 30941 37856
rect 30929 37825 30941 37828
rect 30975 37825 30987 37859
rect 30929 37819 30987 37825
rect 31021 37859 31079 37865
rect 31021 37825 31033 37859
rect 31067 37825 31079 37859
rect 31021 37819 31079 37825
rect 29178 37788 29184 37800
rect 28368 37760 29184 37788
rect 29178 37748 29184 37760
rect 29236 37748 29242 37800
rect 29454 37788 29460 37800
rect 29415 37760 29460 37788
rect 29454 37748 29460 37760
rect 29512 37748 29518 37800
rect 29641 37791 29699 37797
rect 29641 37757 29653 37791
rect 29687 37788 29699 37791
rect 30282 37788 30288 37800
rect 29687 37760 30288 37788
rect 29687 37757 29699 37760
rect 29641 37751 29699 37757
rect 30282 37748 30288 37760
rect 30340 37748 30346 37800
rect 31036 37788 31064 37819
rect 31110 37816 31116 37868
rect 31168 37856 31174 37868
rect 31297 37859 31355 37865
rect 31168 37828 31213 37856
rect 31168 37816 31174 37828
rect 31297 37825 31309 37859
rect 31343 37825 31355 37859
rect 31404 37856 31432 37896
rect 47026 37884 47032 37896
rect 47084 37924 47090 37936
rect 47210 37924 47216 37936
rect 47084 37896 47216 37924
rect 47084 37884 47090 37896
rect 47210 37884 47216 37896
rect 47268 37884 47274 37936
rect 32381 37859 32439 37865
rect 32381 37856 32393 37859
rect 31404 37828 32393 37856
rect 31297 37819 31355 37825
rect 32381 37825 32393 37828
rect 32427 37825 32439 37859
rect 47854 37856 47860 37868
rect 47815 37828 47860 37856
rect 32381 37819 32439 37825
rect 31202 37788 31208 37800
rect 31036 37760 31208 37788
rect 31202 37748 31208 37760
rect 31260 37748 31266 37800
rect 28350 37720 28356 37732
rect 28273 37692 28356 37720
rect 23216 37652 23244 37692
rect 28350 37680 28356 37692
rect 28408 37680 28414 37732
rect 28902 37680 28908 37732
rect 28960 37720 28966 37732
rect 31312 37720 31340 37819
rect 47854 37816 47860 37828
rect 47912 37816 47918 37868
rect 31478 37748 31484 37800
rect 31536 37788 31542 37800
rect 32125 37791 32183 37797
rect 32125 37788 32137 37791
rect 31536 37760 32137 37788
rect 31536 37748 31542 37760
rect 32125 37757 32137 37760
rect 32171 37757 32183 37791
rect 32125 37751 32183 37757
rect 31570 37720 31576 37732
rect 28960 37692 31576 37720
rect 28960 37680 28966 37692
rect 31570 37680 31576 37692
rect 31628 37720 31634 37732
rect 32030 37720 32036 37732
rect 31628 37692 32036 37720
rect 31628 37680 31634 37692
rect 32030 37680 32036 37692
rect 32088 37680 32094 37732
rect 23382 37652 23388 37664
rect 22204 37624 23244 37652
rect 23343 37624 23388 37652
rect 23382 37612 23388 37624
rect 23440 37612 23446 37664
rect 25777 37655 25835 37661
rect 25777 37621 25789 37655
rect 25823 37652 25835 37655
rect 26786 37652 26792 37664
rect 25823 37624 26792 37652
rect 25823 37621 25835 37624
rect 25777 37615 25835 37621
rect 26786 37612 26792 37624
rect 26844 37612 26850 37664
rect 28994 37652 29000 37664
rect 28955 37624 29000 37652
rect 28994 37612 29000 37624
rect 29052 37612 29058 37664
rect 29362 37612 29368 37664
rect 29420 37652 29426 37664
rect 30006 37652 30012 37664
rect 29420 37624 30012 37652
rect 29420 37612 29426 37624
rect 30006 37612 30012 37624
rect 30064 37612 30070 37664
rect 30558 37612 30564 37664
rect 30616 37652 30622 37664
rect 33505 37655 33563 37661
rect 33505 37652 33517 37655
rect 30616 37624 33517 37652
rect 30616 37612 30622 37624
rect 33505 37621 33517 37624
rect 33551 37652 33563 37655
rect 35618 37652 35624 37664
rect 33551 37624 35624 37652
rect 33551 37621 33563 37624
rect 33505 37615 33563 37621
rect 35618 37612 35624 37624
rect 35676 37612 35682 37664
rect 47486 37612 47492 37664
rect 47544 37652 47550 37664
rect 48041 37655 48099 37661
rect 48041 37652 48053 37655
rect 47544 37624 48053 37652
rect 47544 37612 47550 37624
rect 48041 37621 48053 37624
rect 48087 37621 48099 37655
rect 48041 37615 48099 37621
rect 1104 37562 48852 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 48852 37562
rect 1104 37488 48852 37510
rect 8938 37408 8944 37460
rect 8996 37448 9002 37460
rect 20714 37448 20720 37460
rect 8996 37420 20720 37448
rect 8996 37408 9002 37420
rect 20714 37408 20720 37420
rect 20772 37448 20778 37460
rect 21450 37448 21456 37460
rect 20772 37420 21456 37448
rect 20772 37408 20778 37420
rect 21450 37408 21456 37420
rect 21508 37408 21514 37460
rect 23014 37408 23020 37460
rect 23072 37448 23078 37460
rect 23109 37451 23167 37457
rect 23109 37448 23121 37451
rect 23072 37420 23121 37448
rect 23072 37408 23078 37420
rect 23109 37417 23121 37420
rect 23155 37417 23167 37451
rect 25041 37451 25099 37457
rect 23109 37411 23167 37417
rect 23216 37420 24992 37448
rect 4062 37340 4068 37392
rect 4120 37380 4126 37392
rect 4120 37352 9444 37380
rect 4120 37340 4126 37352
rect 1394 37312 1400 37324
rect 1355 37284 1400 37312
rect 1394 37272 1400 37284
rect 1452 37272 1458 37324
rect 9122 37312 9128 37324
rect 9083 37284 9128 37312
rect 9122 37272 9128 37284
rect 9180 37272 9186 37324
rect 9416 37321 9444 37352
rect 13998 37340 14004 37392
rect 14056 37380 14062 37392
rect 17402 37380 17408 37392
rect 14056 37352 17408 37380
rect 14056 37340 14062 37352
rect 17402 37340 17408 37352
rect 17460 37340 17466 37392
rect 22370 37340 22376 37392
rect 22428 37380 22434 37392
rect 23216 37380 23244 37420
rect 22428 37352 23244 37380
rect 24964 37380 24992 37420
rect 25041 37417 25053 37451
rect 25087 37448 25099 37451
rect 25222 37448 25228 37460
rect 25087 37420 25228 37448
rect 25087 37417 25099 37420
rect 25041 37411 25099 37417
rect 25222 37408 25228 37420
rect 25280 37408 25286 37460
rect 27430 37448 27436 37460
rect 26068 37420 27436 37448
rect 26068 37380 26096 37420
rect 27430 37408 27436 37420
rect 27488 37408 27494 37460
rect 28997 37451 29055 37457
rect 28997 37417 29009 37451
rect 29043 37448 29055 37451
rect 29178 37448 29184 37460
rect 29043 37420 29184 37448
rect 29043 37417 29055 37420
rect 28997 37411 29055 37417
rect 29178 37408 29184 37420
rect 29236 37408 29242 37460
rect 24964 37352 26096 37380
rect 22428 37340 22434 37352
rect 26142 37340 26148 37392
rect 26200 37340 26206 37392
rect 28350 37340 28356 37392
rect 28408 37380 28414 37392
rect 31294 37380 31300 37392
rect 28408 37352 31300 37380
rect 28408 37340 28414 37352
rect 31294 37340 31300 37352
rect 31352 37340 31358 37392
rect 32861 37383 32919 37389
rect 32861 37349 32873 37383
rect 32907 37349 32919 37383
rect 32861 37343 32919 37349
rect 9401 37315 9459 37321
rect 9401 37281 9413 37315
rect 9447 37281 9459 37315
rect 9401 37275 9459 37281
rect 15286 37272 15292 37324
rect 15344 37312 15350 37324
rect 15565 37315 15623 37321
rect 15565 37312 15577 37315
rect 15344 37284 15577 37312
rect 15344 37272 15350 37284
rect 15565 37281 15577 37284
rect 15611 37281 15623 37315
rect 23566 37312 23572 37324
rect 23527 37284 23572 37312
rect 15565 37275 15623 37281
rect 23566 37272 23572 37284
rect 23624 37272 23630 37324
rect 23753 37315 23811 37321
rect 23753 37281 23765 37315
rect 23799 37312 23811 37315
rect 25682 37312 25688 37324
rect 23799 37284 25688 37312
rect 23799 37281 23811 37284
rect 23753 37275 23811 37281
rect 25682 37272 25688 37284
rect 25740 37272 25746 37324
rect 25866 37272 25872 37324
rect 25924 37312 25930 37324
rect 26160 37312 26188 37340
rect 25924 37284 26096 37312
rect 26160 37284 26372 37312
rect 25924 37272 25930 37284
rect 1670 37244 1676 37256
rect 1631 37216 1676 37244
rect 1670 37204 1676 37216
rect 1728 37204 1734 37256
rect 8938 37244 8944 37256
rect 8899 37216 8944 37244
rect 8938 37204 8944 37216
rect 8996 37204 9002 37256
rect 15102 37244 15108 37256
rect 15063 37216 15108 37244
rect 15102 37204 15108 37216
rect 15160 37204 15166 37256
rect 17218 37204 17224 37256
rect 17276 37244 17282 37256
rect 17405 37247 17463 37253
rect 17405 37244 17417 37247
rect 17276 37216 17417 37244
rect 17276 37204 17282 37216
rect 17405 37213 17417 37216
rect 17451 37213 17463 37247
rect 17405 37207 17463 37213
rect 17788 37216 18552 37244
rect 15286 37176 15292 37188
rect 15247 37148 15292 37176
rect 15286 37136 15292 37148
rect 15344 37136 15350 37188
rect 3602 37068 3608 37120
rect 3660 37108 3666 37120
rect 17788 37108 17816 37216
rect 18138 37136 18144 37188
rect 18196 37176 18202 37188
rect 18233 37179 18291 37185
rect 18233 37176 18245 37179
rect 18196 37148 18245 37176
rect 18196 37136 18202 37148
rect 18233 37145 18245 37148
rect 18279 37145 18291 37179
rect 18524 37176 18552 37216
rect 18598 37204 18604 37256
rect 18656 37244 18662 37256
rect 19245 37247 19303 37253
rect 19245 37244 19257 37247
rect 18656 37216 19257 37244
rect 18656 37204 18662 37216
rect 19245 37213 19257 37216
rect 19291 37213 19303 37247
rect 19245 37207 19303 37213
rect 20438 37204 20444 37256
rect 20496 37244 20502 37256
rect 21085 37247 21143 37253
rect 21085 37244 21097 37247
rect 20496 37216 21097 37244
rect 20496 37204 20502 37216
rect 21085 37213 21097 37216
rect 21131 37213 21143 37247
rect 21085 37207 21143 37213
rect 21352 37247 21410 37253
rect 21352 37213 21364 37247
rect 21398 37244 21410 37247
rect 21818 37244 21824 37256
rect 21398 37216 21824 37244
rect 21398 37213 21410 37216
rect 21352 37207 21410 37213
rect 21818 37204 21824 37216
rect 21876 37204 21882 37256
rect 21910 37204 21916 37256
rect 21968 37244 21974 37256
rect 22462 37244 22468 37256
rect 21968 37216 22468 37244
rect 21968 37204 21974 37216
rect 22462 37204 22468 37216
rect 22520 37204 22526 37256
rect 24854 37244 24860 37256
rect 24815 37216 24860 37244
rect 24854 37204 24860 37216
rect 24912 37204 24918 37256
rect 25222 37204 25228 37256
rect 25280 37244 25286 37256
rect 26068 37253 26096 37284
rect 25961 37247 26019 37253
rect 25961 37244 25973 37247
rect 25280 37216 25973 37244
rect 25280 37204 25286 37216
rect 25961 37213 25973 37216
rect 26007 37213 26019 37247
rect 25961 37207 26019 37213
rect 26053 37247 26111 37253
rect 26053 37213 26065 37247
rect 26099 37213 26111 37247
rect 26053 37207 26111 37213
rect 26145 37247 26203 37253
rect 26145 37213 26157 37247
rect 26191 37244 26203 37247
rect 26234 37244 26240 37256
rect 26191 37216 26240 37244
rect 26191 37213 26203 37216
rect 26145 37207 26203 37213
rect 26234 37204 26240 37216
rect 26292 37204 26298 37256
rect 26344 37253 26372 37284
rect 30282 37272 30288 37324
rect 30340 37312 30346 37324
rect 30745 37315 30803 37321
rect 30745 37312 30757 37315
rect 30340 37284 30757 37312
rect 30340 37272 30346 37284
rect 30745 37281 30757 37284
rect 30791 37281 30803 37315
rect 30745 37275 30803 37281
rect 31386 37272 31392 37324
rect 31444 37312 31450 37324
rect 32876 37312 32904 37343
rect 31444 37284 31616 37312
rect 31444 37272 31450 37284
rect 26329 37247 26387 37253
rect 26329 37213 26341 37247
rect 26375 37213 26387 37247
rect 26329 37207 26387 37213
rect 26694 37204 26700 37256
rect 26752 37244 26758 37256
rect 26789 37247 26847 37253
rect 26789 37244 26801 37247
rect 26752 37216 26801 37244
rect 26752 37204 26758 37216
rect 26789 37213 26801 37216
rect 26835 37213 26847 37247
rect 26789 37207 26847 37213
rect 28629 37247 28687 37253
rect 28629 37213 28641 37247
rect 28675 37244 28687 37247
rect 28994 37244 29000 37256
rect 28675 37216 29000 37244
rect 28675 37213 28687 37216
rect 28629 37207 28687 37213
rect 28994 37204 29000 37216
rect 29052 37204 29058 37256
rect 29914 37204 29920 37256
rect 29972 37244 29978 37256
rect 30653 37247 30711 37253
rect 30653 37244 30665 37247
rect 29972 37216 30665 37244
rect 29972 37204 29978 37216
rect 30653 37213 30665 37216
rect 30699 37213 30711 37247
rect 31478 37244 31484 37256
rect 31439 37216 31484 37244
rect 30653 37207 30711 37213
rect 31478 37204 31484 37216
rect 31536 37204 31542 37256
rect 31588 37244 31616 37284
rect 32692 37284 32904 37312
rect 31737 37247 31795 37253
rect 31737 37244 31749 37247
rect 31588 37216 31749 37244
rect 31737 37213 31749 37216
rect 31783 37213 31795 37247
rect 31737 37207 31795 37213
rect 20346 37176 20352 37188
rect 18524 37148 20352 37176
rect 18233 37139 18291 37145
rect 3660 37080 17816 37108
rect 18248 37108 18276 37139
rect 20346 37136 20352 37148
rect 20404 37136 20410 37188
rect 22370 37176 22376 37188
rect 22066 37148 22376 37176
rect 22066 37108 22094 37148
rect 22370 37136 22376 37148
rect 22428 37136 22434 37188
rect 23566 37176 23572 37188
rect 22480 37148 23572 37176
rect 22480 37120 22508 37148
rect 23566 37136 23572 37148
rect 23624 37136 23630 37188
rect 24670 37176 24676 37188
rect 24631 37148 24676 37176
rect 24670 37136 24676 37148
rect 24728 37136 24734 37188
rect 25685 37179 25743 37185
rect 25685 37145 25697 37179
rect 25731 37176 25743 37179
rect 27034 37179 27092 37185
rect 27034 37176 27046 37179
rect 25731 37148 27046 37176
rect 25731 37145 25743 37148
rect 25685 37139 25743 37145
rect 27034 37145 27046 37148
rect 27080 37145 27092 37179
rect 28810 37176 28816 37188
rect 28723 37148 28816 37176
rect 27034 37139 27092 37145
rect 28810 37136 28816 37148
rect 28868 37176 28874 37188
rect 30558 37176 30564 37188
rect 28868 37148 30420 37176
rect 30519 37148 30564 37176
rect 28868 37136 28874 37148
rect 22462 37108 22468 37120
rect 18248 37080 22094 37108
rect 22375 37080 22468 37108
rect 3660 37068 3666 37080
rect 22462 37068 22468 37080
rect 22520 37068 22526 37120
rect 23477 37111 23535 37117
rect 23477 37077 23489 37111
rect 23523 37108 23535 37111
rect 24854 37108 24860 37120
rect 23523 37080 24860 37108
rect 23523 37077 23535 37080
rect 23477 37071 23535 37077
rect 24854 37068 24860 37080
rect 24912 37068 24918 37120
rect 25498 37068 25504 37120
rect 25556 37108 25562 37120
rect 28169 37111 28227 37117
rect 28169 37108 28181 37111
rect 25556 37080 28181 37108
rect 25556 37068 25562 37080
rect 28169 37077 28181 37080
rect 28215 37108 28227 37111
rect 30006 37108 30012 37120
rect 28215 37080 30012 37108
rect 28215 37077 28227 37080
rect 28169 37071 28227 37077
rect 30006 37068 30012 37080
rect 30064 37068 30070 37120
rect 30190 37108 30196 37120
rect 30151 37080 30196 37108
rect 30190 37068 30196 37080
rect 30248 37068 30254 37120
rect 30392 37108 30420 37148
rect 30558 37136 30564 37148
rect 30616 37136 30622 37188
rect 31202 37136 31208 37188
rect 31260 37176 31266 37188
rect 32692 37176 32720 37284
rect 46842 37204 46848 37256
rect 46900 37244 46906 37256
rect 47121 37247 47179 37253
rect 47121 37244 47133 37247
rect 46900 37216 47133 37244
rect 46900 37204 46906 37216
rect 47121 37213 47133 37216
rect 47167 37213 47179 37247
rect 47946 37244 47952 37256
rect 47907 37216 47952 37244
rect 47121 37207 47179 37213
rect 47946 37204 47952 37216
rect 48004 37204 48010 37256
rect 31260 37148 32720 37176
rect 31260 37136 31266 37148
rect 30926 37108 30932 37120
rect 30392 37080 30932 37108
rect 30926 37068 30932 37080
rect 30984 37068 30990 37120
rect 46474 37068 46480 37120
rect 46532 37108 46538 37120
rect 47213 37111 47271 37117
rect 47213 37108 47225 37111
rect 46532 37080 47225 37108
rect 46532 37068 46538 37080
rect 47213 37077 47225 37080
rect 47259 37077 47271 37111
rect 47213 37071 47271 37077
rect 1104 37018 48852 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 48852 37018
rect 1104 36944 48852 36966
rect 8938 36864 8944 36916
rect 8996 36904 9002 36916
rect 9585 36907 9643 36913
rect 9585 36904 9597 36907
rect 8996 36876 9597 36904
rect 8996 36864 9002 36876
rect 9585 36873 9597 36876
rect 9631 36873 9643 36907
rect 9585 36867 9643 36873
rect 11532 36876 15056 36904
rect 1670 36796 1676 36848
rect 1728 36836 1734 36848
rect 1728 36808 9251 36836
rect 1728 36796 1734 36808
rect 8205 36771 8263 36777
rect 8205 36737 8217 36771
rect 8251 36768 8263 36771
rect 8294 36768 8300 36780
rect 8251 36740 8300 36768
rect 8251 36737 8263 36740
rect 8205 36731 8263 36737
rect 8294 36728 8300 36740
rect 8352 36728 8358 36780
rect 8472 36771 8530 36777
rect 8472 36737 8484 36771
rect 8518 36768 8530 36771
rect 9030 36768 9036 36780
rect 8518 36740 9036 36768
rect 8518 36737 8530 36740
rect 8472 36731 8530 36737
rect 9030 36728 9036 36740
rect 9088 36728 9094 36780
rect 1670 36660 1676 36712
rect 1728 36700 1734 36712
rect 1946 36700 1952 36712
rect 1728 36672 1952 36700
rect 1728 36660 1734 36672
rect 1946 36660 1952 36672
rect 2004 36660 2010 36712
rect 9223 36632 9251 36808
rect 11532 36777 11560 36876
rect 13354 36836 13360 36848
rect 13315 36808 13360 36836
rect 13354 36796 13360 36808
rect 13412 36796 13418 36848
rect 15028 36836 15056 36876
rect 15102 36864 15108 36916
rect 15160 36904 15166 36916
rect 15565 36907 15623 36913
rect 15565 36904 15577 36907
rect 15160 36876 15577 36904
rect 15160 36864 15166 36876
rect 15565 36873 15577 36876
rect 15611 36873 15623 36907
rect 21726 36904 21732 36916
rect 15565 36867 15623 36873
rect 19352 36876 21732 36904
rect 16482 36836 16488 36848
rect 15028 36808 16488 36836
rect 16482 36796 16488 36808
rect 16540 36796 16546 36848
rect 18782 36796 18788 36848
rect 18840 36836 18846 36848
rect 19352 36845 19380 36876
rect 21726 36864 21732 36876
rect 21784 36864 21790 36916
rect 21821 36907 21879 36913
rect 21821 36873 21833 36907
rect 21867 36904 21879 36907
rect 22278 36904 22284 36916
rect 21867 36876 22284 36904
rect 21867 36873 21879 36876
rect 21821 36867 21879 36873
rect 22278 36864 22284 36876
rect 22336 36864 22342 36916
rect 22370 36864 22376 36916
rect 22428 36904 22434 36916
rect 24670 36904 24676 36916
rect 22428 36876 22876 36904
rect 24631 36876 24676 36904
rect 22428 36864 22434 36876
rect 19337 36839 19395 36845
rect 19337 36836 19349 36839
rect 18840 36808 19349 36836
rect 18840 36796 18846 36808
rect 19337 36805 19349 36808
rect 19383 36805 19395 36839
rect 19337 36799 19395 36805
rect 20438 36796 20444 36848
rect 20496 36836 20502 36848
rect 22848 36836 22876 36876
rect 24670 36864 24676 36876
rect 24728 36864 24734 36916
rect 26234 36904 26240 36916
rect 26195 36876 26240 36904
rect 26234 36864 26240 36876
rect 26292 36864 26298 36916
rect 29549 36907 29607 36913
rect 29549 36873 29561 36907
rect 29595 36904 29607 36907
rect 31113 36907 31171 36913
rect 29595 36876 30788 36904
rect 29595 36873 29607 36876
rect 29549 36867 29607 36873
rect 30760 36845 30788 36876
rect 31113 36873 31125 36907
rect 31159 36904 31171 36907
rect 31938 36904 31944 36916
rect 31159 36876 31944 36904
rect 31159 36873 31171 36876
rect 31113 36867 31171 36873
rect 31938 36864 31944 36876
rect 31996 36864 32002 36916
rect 30745 36839 30803 36845
rect 20496 36808 22784 36836
rect 22848 36808 30052 36836
rect 20496 36796 20502 36808
rect 14458 36777 14464 36780
rect 11517 36771 11575 36777
rect 11517 36737 11529 36771
rect 11563 36737 11575 36771
rect 11517 36731 11575 36737
rect 14452 36731 14464 36777
rect 14516 36768 14522 36780
rect 17218 36768 17224 36780
rect 14516 36740 14552 36768
rect 17179 36740 17224 36768
rect 14458 36728 14464 36731
rect 14516 36728 14522 36740
rect 17218 36728 17224 36740
rect 17276 36728 17282 36780
rect 18598 36768 18604 36780
rect 18559 36740 18604 36768
rect 18598 36728 18604 36740
rect 18656 36728 18662 36780
rect 20717 36771 20775 36777
rect 20717 36737 20729 36771
rect 20763 36768 20775 36771
rect 21082 36768 21088 36780
rect 20763 36740 21088 36768
rect 20763 36737 20775 36740
rect 20717 36731 20775 36737
rect 21082 36728 21088 36740
rect 21140 36768 21146 36780
rect 21910 36768 21916 36780
rect 21140 36740 21916 36768
rect 21140 36728 21146 36740
rect 21910 36728 21916 36740
rect 21968 36728 21974 36780
rect 22005 36771 22063 36777
rect 22005 36737 22017 36771
rect 22051 36737 22063 36771
rect 22005 36731 22063 36737
rect 22189 36771 22247 36777
rect 22189 36737 22201 36771
rect 22235 36737 22247 36771
rect 22189 36731 22247 36737
rect 22281 36771 22339 36777
rect 22281 36737 22293 36771
rect 22327 36768 22339 36771
rect 22462 36768 22468 36780
rect 22327 36740 22468 36768
rect 22327 36737 22339 36740
rect 22281 36731 22339 36737
rect 11698 36700 11704 36712
rect 11659 36672 11704 36700
rect 11698 36660 11704 36672
rect 11756 36660 11762 36712
rect 14185 36703 14243 36709
rect 14185 36669 14197 36703
rect 14231 36669 14243 36703
rect 14185 36663 14243 36669
rect 14090 36632 14096 36644
rect 9223 36604 14096 36632
rect 14090 36592 14096 36604
rect 14148 36592 14154 36644
rect 2317 36567 2375 36573
rect 2317 36533 2329 36567
rect 2363 36564 2375 36567
rect 2498 36564 2504 36576
rect 2363 36536 2504 36564
rect 2363 36533 2375 36536
rect 2317 36527 2375 36533
rect 2498 36524 2504 36536
rect 2556 36524 2562 36576
rect 12710 36524 12716 36576
rect 12768 36564 12774 36576
rect 13814 36564 13820 36576
rect 12768 36536 13820 36564
rect 12768 36524 12774 36536
rect 13814 36524 13820 36536
rect 13872 36524 13878 36576
rect 14200 36564 14228 36663
rect 16850 36660 16856 36712
rect 16908 36700 16914 36712
rect 17405 36703 17463 36709
rect 17405 36700 17417 36703
rect 16908 36672 17417 36700
rect 16908 36660 16914 36672
rect 17405 36669 17417 36672
rect 17451 36700 17463 36703
rect 17862 36700 17868 36712
rect 17451 36672 17868 36700
rect 17451 36669 17463 36672
rect 17405 36663 17463 36669
rect 17862 36660 17868 36672
rect 17920 36660 17926 36712
rect 20346 36660 20352 36712
rect 20404 36700 20410 36712
rect 20441 36703 20499 36709
rect 20441 36700 20453 36703
rect 20404 36672 20453 36700
rect 20404 36660 20410 36672
rect 20441 36669 20453 36672
rect 20487 36669 20499 36703
rect 22020 36700 22048 36731
rect 22204 36700 22232 36731
rect 22462 36728 22468 36740
rect 22520 36728 22526 36780
rect 22756 36777 22784 36808
rect 23014 36777 23020 36780
rect 22741 36771 22799 36777
rect 22741 36737 22753 36771
rect 22787 36737 22799 36771
rect 22741 36731 22799 36737
rect 23008 36731 23020 36777
rect 23072 36768 23078 36780
rect 25041 36771 25099 36777
rect 23072 36740 23108 36768
rect 23014 36728 23020 36731
rect 23072 36728 23078 36740
rect 25041 36737 25053 36771
rect 25087 36768 25099 36771
rect 25866 36768 25872 36780
rect 25087 36740 25268 36768
rect 25827 36740 25872 36768
rect 25087 36737 25099 36740
rect 25041 36731 25099 36737
rect 22646 36700 22652 36712
rect 22020 36672 22094 36700
rect 22204 36672 22652 36700
rect 20441 36663 20499 36669
rect 22066 36632 22094 36672
rect 22646 36660 22652 36672
rect 22704 36660 22710 36712
rect 24302 36660 24308 36712
rect 24360 36700 24366 36712
rect 25133 36703 25191 36709
rect 25133 36700 25145 36703
rect 24360 36672 25145 36700
rect 24360 36660 24366 36672
rect 25133 36669 25145 36672
rect 25179 36669 25191 36703
rect 25133 36663 25191 36669
rect 22370 36632 22376 36644
rect 22066 36604 22376 36632
rect 22370 36592 22376 36604
rect 22428 36592 22434 36644
rect 25240 36632 25268 36740
rect 25866 36728 25872 36740
rect 25924 36728 25930 36780
rect 26050 36768 26056 36780
rect 26011 36740 26056 36768
rect 26050 36728 26056 36740
rect 26108 36728 26114 36780
rect 26326 36728 26332 36780
rect 26384 36768 26390 36780
rect 27229 36771 27287 36777
rect 27229 36768 27241 36771
rect 26384 36740 27241 36768
rect 26384 36728 26390 36740
rect 27229 36737 27241 36740
rect 27275 36737 27287 36771
rect 27229 36731 27287 36737
rect 27798 36728 27804 36780
rect 27856 36768 27862 36780
rect 29917 36771 29975 36777
rect 29917 36768 29929 36771
rect 27856 36740 29929 36768
rect 27856 36728 27862 36740
rect 25317 36703 25375 36709
rect 25317 36669 25329 36703
rect 25363 36700 25375 36703
rect 25682 36700 25688 36712
rect 25363 36672 25688 36700
rect 25363 36669 25375 36672
rect 25317 36663 25375 36669
rect 25682 36660 25688 36672
rect 25740 36660 25746 36712
rect 26694 36660 26700 36712
rect 26752 36700 26758 36712
rect 26973 36703 27031 36709
rect 26973 36700 26985 36703
rect 26752 36672 26985 36700
rect 26752 36660 26758 36672
rect 26973 36669 26985 36672
rect 27019 36669 27031 36703
rect 26973 36663 27031 36669
rect 26418 36632 26424 36644
rect 25240 36604 26424 36632
rect 26418 36592 26424 36604
rect 26476 36592 26482 36644
rect 29840 36632 29868 36740
rect 29917 36737 29929 36740
rect 29963 36737 29975 36771
rect 30024 36768 30052 36808
rect 30745 36805 30757 36839
rect 30791 36805 30803 36839
rect 45830 36836 45836 36848
rect 30745 36799 30803 36805
rect 30852 36808 45836 36836
rect 30852 36768 30880 36808
rect 45830 36796 45836 36808
rect 45888 36836 45894 36848
rect 46750 36836 46756 36848
rect 45888 36808 46756 36836
rect 45888 36796 45894 36808
rect 46750 36796 46756 36808
rect 46808 36796 46814 36848
rect 30024 36740 30880 36768
rect 29917 36731 29975 36737
rect 30926 36728 30932 36780
rect 30984 36768 30990 36780
rect 30984 36740 31029 36768
rect 30984 36728 30990 36740
rect 30006 36700 30012 36712
rect 29967 36672 30012 36700
rect 30006 36660 30012 36672
rect 30064 36660 30070 36712
rect 30193 36703 30251 36709
rect 30193 36669 30205 36703
rect 30239 36700 30251 36703
rect 30282 36700 30288 36712
rect 30239 36672 30288 36700
rect 30239 36669 30251 36672
rect 30193 36663 30251 36669
rect 30282 36660 30288 36672
rect 30340 36660 30346 36712
rect 31202 36632 31208 36644
rect 29840 36604 31208 36632
rect 31202 36592 31208 36604
rect 31260 36592 31266 36644
rect 15194 36564 15200 36576
rect 14200 36536 15200 36564
rect 15194 36524 15200 36536
rect 15252 36524 15258 36576
rect 24121 36567 24179 36573
rect 24121 36533 24133 36567
rect 24167 36564 24179 36567
rect 24854 36564 24860 36576
rect 24167 36536 24860 36564
rect 24167 36533 24179 36536
rect 24121 36527 24179 36533
rect 24854 36524 24860 36536
rect 24912 36564 24918 36576
rect 25958 36564 25964 36576
rect 24912 36536 25964 36564
rect 24912 36524 24918 36536
rect 25958 36524 25964 36536
rect 26016 36524 26022 36576
rect 28353 36567 28411 36573
rect 28353 36533 28365 36567
rect 28399 36564 28411 36567
rect 28902 36564 28908 36576
rect 28399 36536 28908 36564
rect 28399 36533 28411 36536
rect 28353 36527 28411 36533
rect 28902 36524 28908 36536
rect 28960 36524 28966 36576
rect 46842 36524 46848 36576
rect 46900 36564 46906 36576
rect 47765 36567 47823 36573
rect 47765 36564 47777 36567
rect 46900 36536 47777 36564
rect 46900 36524 46906 36536
rect 47765 36533 47777 36536
rect 47811 36533 47823 36567
rect 47765 36527 47823 36533
rect 1104 36474 48852 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 48852 36474
rect 1104 36400 48852 36422
rect 11517 36363 11575 36369
rect 11517 36329 11529 36363
rect 11563 36360 11575 36363
rect 11698 36360 11704 36372
rect 11563 36332 11704 36360
rect 11563 36329 11575 36332
rect 11517 36323 11575 36329
rect 11698 36320 11704 36332
rect 11756 36320 11762 36372
rect 16482 36360 16488 36372
rect 12406 36332 16344 36360
rect 16443 36332 16488 36360
rect 2130 36184 2136 36236
rect 2188 36224 2194 36236
rect 2498 36224 2504 36236
rect 2188 36196 2504 36224
rect 2188 36184 2194 36196
rect 2498 36184 2504 36196
rect 2556 36184 2562 36236
rect 2961 36159 3019 36165
rect 2961 36125 2973 36159
rect 3007 36156 3019 36159
rect 3694 36156 3700 36168
rect 3007 36128 3700 36156
rect 3007 36125 3019 36128
rect 2961 36119 3019 36125
rect 3694 36116 3700 36128
rect 3752 36116 3758 36168
rect 3786 36116 3792 36168
rect 3844 36156 3850 36168
rect 11425 36159 11483 36165
rect 11425 36156 11437 36159
rect 3844 36128 11437 36156
rect 3844 36116 3850 36128
rect 11425 36125 11437 36128
rect 11471 36156 11483 36159
rect 12406 36156 12434 36332
rect 16316 36292 16344 36332
rect 16482 36320 16488 36332
rect 16540 36320 16546 36372
rect 18598 36360 18604 36372
rect 18559 36332 18604 36360
rect 18598 36320 18604 36332
rect 18656 36320 18662 36372
rect 25133 36363 25191 36369
rect 25133 36329 25145 36363
rect 25179 36360 25191 36363
rect 25866 36360 25872 36372
rect 25179 36332 25872 36360
rect 25179 36329 25191 36332
rect 25133 36323 25191 36329
rect 25866 36320 25872 36332
rect 25924 36320 25930 36372
rect 26326 36360 26332 36372
rect 26287 36332 26332 36360
rect 26326 36320 26332 36332
rect 26384 36320 26390 36372
rect 26620 36332 27016 36360
rect 18138 36292 18144 36304
rect 16316 36264 18144 36292
rect 18138 36252 18144 36264
rect 18196 36252 18202 36304
rect 24673 36295 24731 36301
rect 24673 36261 24685 36295
rect 24719 36292 24731 36295
rect 24854 36292 24860 36304
rect 24719 36264 24860 36292
rect 24719 36261 24731 36264
rect 24673 36255 24731 36261
rect 24854 36252 24860 36264
rect 24912 36292 24918 36304
rect 26142 36292 26148 36304
rect 24912 36264 26148 36292
rect 24912 36252 24918 36264
rect 26142 36252 26148 36264
rect 26200 36292 26206 36304
rect 26620 36292 26648 36332
rect 26200 36264 26648 36292
rect 26200 36252 26206 36264
rect 19978 36184 19984 36236
rect 20036 36224 20042 36236
rect 20073 36227 20131 36233
rect 20073 36224 20085 36227
rect 20036 36196 20085 36224
rect 20036 36184 20042 36196
rect 20073 36193 20085 36196
rect 20119 36193 20131 36227
rect 22646 36224 22652 36236
rect 22607 36196 22652 36224
rect 20073 36187 20131 36193
rect 22646 36184 22652 36196
rect 22704 36184 22710 36236
rect 25682 36224 25688 36236
rect 25643 36196 25688 36224
rect 25682 36184 25688 36196
rect 25740 36184 25746 36236
rect 11471 36128 12434 36156
rect 15105 36159 15163 36165
rect 11471 36125 11483 36128
rect 11425 36119 11483 36125
rect 15105 36125 15117 36159
rect 15151 36156 15163 36159
rect 15194 36156 15200 36168
rect 15151 36128 15200 36156
rect 15151 36125 15163 36128
rect 15105 36119 15163 36125
rect 15194 36116 15200 36128
rect 15252 36156 15258 36168
rect 17221 36159 17279 36165
rect 17221 36156 17233 36159
rect 15252 36128 16068 36156
rect 15252 36116 15258 36128
rect 16040 36100 16068 36128
rect 16132 36128 17233 36156
rect 15372 36091 15430 36097
rect 15372 36057 15384 36091
rect 15418 36088 15430 36091
rect 15838 36088 15844 36100
rect 15418 36060 15844 36088
rect 15418 36057 15430 36060
rect 15372 36051 15430 36057
rect 15838 36048 15844 36060
rect 15896 36048 15902 36100
rect 16022 36048 16028 36100
rect 16080 36048 16086 36100
rect 3050 36020 3056 36032
rect 3011 35992 3056 36020
rect 3050 35980 3056 35992
rect 3108 35980 3114 36032
rect 15010 35980 15016 36032
rect 15068 36020 15074 36032
rect 16132 36020 16160 36128
rect 17221 36125 17233 36128
rect 17267 36125 17279 36159
rect 17221 36119 17279 36125
rect 17313 36159 17371 36165
rect 17313 36125 17325 36159
rect 17359 36125 17371 36159
rect 17313 36119 17371 36125
rect 17034 36048 17040 36100
rect 17092 36088 17098 36100
rect 17328 36088 17356 36119
rect 17402 36116 17408 36168
rect 17460 36156 17466 36168
rect 17460 36128 17505 36156
rect 17460 36116 17466 36128
rect 17586 36116 17592 36168
rect 17644 36156 17650 36168
rect 17644 36128 17689 36156
rect 17644 36116 17650 36128
rect 18138 36116 18144 36168
rect 18196 36156 18202 36168
rect 19150 36156 19156 36168
rect 18196 36128 19156 36156
rect 18196 36116 18202 36128
rect 19150 36116 19156 36128
rect 19208 36156 19214 36168
rect 19245 36159 19303 36165
rect 19245 36156 19257 36159
rect 19208 36128 19257 36156
rect 19208 36116 19214 36128
rect 19245 36125 19257 36128
rect 19291 36125 19303 36159
rect 19245 36119 19303 36125
rect 22186 36116 22192 36168
rect 22244 36156 22250 36168
rect 22373 36159 22431 36165
rect 22373 36156 22385 36159
rect 22244 36128 22385 36156
rect 22244 36116 22250 36128
rect 22373 36125 22385 36128
rect 22419 36125 22431 36159
rect 22373 36119 22431 36125
rect 23290 36116 23296 36168
rect 23348 36156 23354 36168
rect 25498 36156 25504 36168
rect 23348 36128 25360 36156
rect 25459 36128 25504 36156
rect 23348 36116 23354 36128
rect 17092 36060 17356 36088
rect 17092 36048 17098 36060
rect 18230 36048 18236 36100
rect 18288 36088 18294 36100
rect 18325 36091 18383 36097
rect 18325 36088 18337 36091
rect 18288 36060 18337 36088
rect 18288 36048 18294 36060
rect 18325 36057 18337 36060
rect 18371 36088 18383 36091
rect 20257 36091 20315 36097
rect 18371 36060 19472 36088
rect 18371 36057 18383 36060
rect 18325 36051 18383 36057
rect 19168 36032 19196 36060
rect 16942 36020 16948 36032
rect 15068 35992 16160 36020
rect 16903 35992 16948 36020
rect 15068 35980 15074 35992
rect 16942 35980 16948 35992
rect 17000 35980 17006 36032
rect 19150 35980 19156 36032
rect 19208 35980 19214 36032
rect 19444 36029 19472 36060
rect 20257 36057 20269 36091
rect 20303 36088 20315 36091
rect 21726 36088 21732 36100
rect 20303 36060 21732 36088
rect 20303 36057 20315 36060
rect 20257 36051 20315 36057
rect 21726 36048 21732 36060
rect 21784 36048 21790 36100
rect 21910 36088 21916 36100
rect 21871 36060 21916 36088
rect 21910 36048 21916 36060
rect 21968 36048 21974 36100
rect 24489 36091 24547 36097
rect 24489 36057 24501 36091
rect 24535 36057 24547 36091
rect 25332 36088 25360 36128
rect 25498 36116 25504 36128
rect 25556 36116 25562 36168
rect 25593 36159 25651 36165
rect 25593 36125 25605 36159
rect 25639 36156 25651 36159
rect 25774 36156 25780 36168
rect 25639 36128 25780 36156
rect 25639 36125 25651 36128
rect 25593 36119 25651 36125
rect 25774 36116 25780 36128
rect 25832 36116 25838 36168
rect 26234 36116 26240 36168
rect 26292 36156 26298 36168
rect 26559 36159 26617 36165
rect 26559 36156 26571 36159
rect 26292 36128 26571 36156
rect 26292 36116 26298 36128
rect 26559 36125 26571 36128
rect 26605 36125 26617 36159
rect 26559 36119 26617 36125
rect 26697 36159 26755 36165
rect 26697 36125 26709 36159
rect 26743 36125 26755 36159
rect 26697 36119 26755 36125
rect 26050 36088 26056 36100
rect 25332 36060 26056 36088
rect 24489 36051 24547 36057
rect 19429 36023 19487 36029
rect 19429 35989 19441 36023
rect 19475 35989 19487 36023
rect 19429 35983 19487 35989
rect 21266 35980 21272 36032
rect 21324 36020 21330 36032
rect 24504 36020 24532 36051
rect 26050 36048 26056 36060
rect 26108 36088 26114 36100
rect 26712 36088 26740 36119
rect 26786 36116 26792 36168
rect 26844 36156 26850 36168
rect 26988 36165 27016 36332
rect 31294 36292 31300 36304
rect 31220 36264 31300 36292
rect 26973 36159 27031 36165
rect 26844 36128 26889 36156
rect 26844 36116 26850 36128
rect 26973 36125 26985 36159
rect 27019 36125 27031 36159
rect 27709 36159 27767 36165
rect 27709 36156 27721 36159
rect 26973 36119 27031 36125
rect 27080 36128 27721 36156
rect 27080 36088 27108 36128
rect 27709 36125 27721 36128
rect 27755 36125 27767 36159
rect 31110 36156 31116 36168
rect 31071 36128 31116 36156
rect 27709 36119 27767 36125
rect 31110 36116 31116 36128
rect 31168 36116 31174 36168
rect 31220 36165 31248 36264
rect 31294 36252 31300 36264
rect 31352 36252 31358 36304
rect 47946 36292 47952 36304
rect 46308 36264 47952 36292
rect 31846 36224 31852 36236
rect 31404 36196 31852 36224
rect 31205 36159 31263 36165
rect 31205 36125 31217 36159
rect 31251 36125 31263 36159
rect 31205 36119 31263 36125
rect 31318 36159 31376 36165
rect 31318 36125 31330 36159
rect 31364 36156 31376 36159
rect 31404 36156 31432 36196
rect 31846 36184 31852 36196
rect 31904 36184 31910 36236
rect 46308 36233 46336 36264
rect 47946 36252 47952 36264
rect 48004 36252 48010 36304
rect 46293 36227 46351 36233
rect 46293 36193 46305 36227
rect 46339 36193 46351 36227
rect 46474 36224 46480 36236
rect 46435 36196 46480 36224
rect 46293 36187 46351 36193
rect 46474 36184 46480 36196
rect 46532 36184 46538 36236
rect 48130 36224 48136 36236
rect 48091 36196 48136 36224
rect 48130 36184 48136 36196
rect 48188 36184 48194 36236
rect 31364 36128 31432 36156
rect 31481 36159 31539 36165
rect 31364 36125 31376 36128
rect 31318 36119 31376 36125
rect 31481 36125 31493 36159
rect 31527 36156 31539 36159
rect 31570 36156 31576 36168
rect 31527 36128 31576 36156
rect 31527 36125 31539 36128
rect 31481 36119 31539 36125
rect 26108 36060 27108 36088
rect 26108 36048 26114 36060
rect 27154 36048 27160 36100
rect 27212 36088 27218 36100
rect 27430 36088 27436 36100
rect 27212 36060 27436 36088
rect 27212 36048 27218 36060
rect 27430 36048 27436 36060
rect 27488 36088 27494 36100
rect 27525 36091 27583 36097
rect 27525 36088 27537 36091
rect 27488 36060 27537 36088
rect 27488 36048 27494 36060
rect 27525 36057 27537 36060
rect 27571 36057 27583 36091
rect 27525 36051 27583 36057
rect 29178 36048 29184 36100
rect 29236 36088 29242 36100
rect 29730 36088 29736 36100
rect 29236 36060 29736 36088
rect 29236 36048 29242 36060
rect 29730 36048 29736 36060
rect 29788 36048 29794 36100
rect 31220 36088 31248 36119
rect 31570 36116 31576 36128
rect 31628 36116 31634 36168
rect 31662 36088 31668 36100
rect 31220 36060 31668 36088
rect 31662 36048 31668 36060
rect 31720 36048 31726 36100
rect 27890 36020 27896 36032
rect 21324 35992 27896 36020
rect 21324 35980 21330 35992
rect 27890 35980 27896 35992
rect 27948 35980 27954 36032
rect 30837 36023 30895 36029
rect 30837 35989 30849 36023
rect 30883 36020 30895 36023
rect 32030 36020 32036 36032
rect 30883 35992 32036 36020
rect 30883 35989 30895 35992
rect 30837 35983 30895 35989
rect 32030 35980 32036 35992
rect 32088 35980 32094 36032
rect 1104 35930 48852 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 48852 35930
rect 1104 35856 48852 35878
rect 9030 35816 9036 35828
rect 8991 35788 9036 35816
rect 9030 35776 9036 35788
rect 9088 35776 9094 35828
rect 15197 35819 15255 35825
rect 15197 35785 15209 35819
rect 15243 35816 15255 35819
rect 15286 35816 15292 35828
rect 15243 35788 15292 35816
rect 15243 35785 15255 35788
rect 15197 35779 15255 35785
rect 15286 35776 15292 35788
rect 15344 35776 15350 35828
rect 15856 35788 17908 35816
rect 2225 35751 2283 35757
rect 2225 35717 2237 35751
rect 2271 35748 2283 35751
rect 3050 35748 3056 35760
rect 2271 35720 3056 35748
rect 2271 35717 2283 35720
rect 2225 35711 2283 35717
rect 3050 35708 3056 35720
rect 3108 35708 3114 35760
rect 3694 35708 3700 35760
rect 3752 35748 3758 35760
rect 12066 35748 12072 35760
rect 3752 35720 12072 35748
rect 3752 35708 3758 35720
rect 12066 35708 12072 35720
rect 12124 35748 12130 35760
rect 15856 35748 15884 35788
rect 12124 35720 15884 35748
rect 15933 35751 15991 35757
rect 12124 35708 12130 35720
rect 15933 35717 15945 35751
rect 15979 35748 15991 35751
rect 16482 35748 16488 35760
rect 15979 35720 16488 35748
rect 15979 35717 15991 35720
rect 15933 35711 15991 35717
rect 16482 35708 16488 35720
rect 16540 35708 16546 35760
rect 16942 35708 16948 35760
rect 17000 35748 17006 35760
rect 17098 35751 17156 35757
rect 17098 35748 17110 35751
rect 17000 35720 17110 35748
rect 17000 35708 17006 35720
rect 17098 35717 17110 35720
rect 17144 35717 17156 35751
rect 17880 35748 17908 35788
rect 17954 35776 17960 35828
rect 18012 35816 18018 35828
rect 18233 35819 18291 35825
rect 18233 35816 18245 35819
rect 18012 35788 18245 35816
rect 18012 35776 18018 35788
rect 18233 35785 18245 35788
rect 18279 35816 18291 35819
rect 19242 35816 19248 35828
rect 18279 35788 19248 35816
rect 18279 35785 18291 35788
rect 18233 35779 18291 35785
rect 19242 35776 19248 35788
rect 19300 35776 19306 35828
rect 21082 35816 21088 35828
rect 19904 35788 21088 35816
rect 19904 35748 19932 35788
rect 21082 35776 21088 35788
rect 21140 35816 21146 35828
rect 21140 35788 21588 35816
rect 21140 35776 21146 35788
rect 17880 35720 19932 35748
rect 19981 35751 20039 35757
rect 17098 35711 17156 35717
rect 19981 35717 19993 35751
rect 20027 35748 20039 35751
rect 20254 35748 20260 35760
rect 20027 35720 20260 35748
rect 20027 35717 20039 35720
rect 19981 35711 20039 35717
rect 20254 35708 20260 35720
rect 20312 35708 20318 35760
rect 21560 35748 21588 35788
rect 21726 35776 21732 35828
rect 21784 35816 21790 35828
rect 21913 35819 21971 35825
rect 21913 35816 21925 35819
rect 21784 35788 21925 35816
rect 21784 35776 21790 35788
rect 21913 35785 21925 35788
rect 21959 35785 21971 35819
rect 21913 35779 21971 35785
rect 22925 35819 22983 35825
rect 22925 35785 22937 35819
rect 22971 35816 22983 35819
rect 23014 35816 23020 35828
rect 22971 35788 23020 35816
rect 22971 35785 22983 35788
rect 22925 35779 22983 35785
rect 23014 35776 23020 35788
rect 23072 35776 23078 35828
rect 24854 35816 24860 35828
rect 23584 35788 24860 35816
rect 22278 35748 22284 35760
rect 21192 35720 21496 35748
rect 21560 35720 22284 35748
rect 2038 35680 2044 35692
rect 1999 35652 2044 35680
rect 2038 35640 2044 35652
rect 2096 35640 2102 35692
rect 9217 35683 9275 35689
rect 9217 35649 9229 35683
rect 9263 35680 9275 35683
rect 9398 35680 9404 35692
rect 9263 35652 9404 35680
rect 9263 35649 9275 35652
rect 9217 35643 9275 35649
rect 9398 35640 9404 35652
rect 9456 35640 9462 35692
rect 14826 35640 14832 35692
rect 14884 35680 14890 35692
rect 15105 35683 15163 35689
rect 15105 35680 15117 35683
rect 14884 35652 15117 35680
rect 14884 35640 14890 35652
rect 15105 35649 15117 35652
rect 15151 35649 15163 35683
rect 15105 35643 15163 35649
rect 15749 35683 15807 35689
rect 15749 35649 15761 35683
rect 15795 35680 15807 35683
rect 16758 35680 16764 35692
rect 15795 35652 16764 35680
rect 15795 35649 15807 35652
rect 15749 35643 15807 35649
rect 16758 35640 16764 35652
rect 16816 35640 16822 35692
rect 19242 35680 19248 35692
rect 19203 35652 19248 35680
rect 19242 35640 19248 35652
rect 19300 35640 19306 35692
rect 20622 35640 20628 35692
rect 20680 35680 20686 35692
rect 20855 35683 20913 35689
rect 20855 35680 20867 35683
rect 20680 35652 20867 35680
rect 20680 35640 20686 35652
rect 20855 35649 20867 35652
rect 20901 35649 20913 35683
rect 20990 35680 20996 35692
rect 20951 35652 20996 35680
rect 20855 35643 20913 35649
rect 20990 35640 20996 35652
rect 21048 35640 21054 35692
rect 21106 35683 21164 35689
rect 21106 35649 21118 35683
rect 21152 35680 21164 35683
rect 21192 35680 21220 35720
rect 21152 35652 21220 35680
rect 21269 35683 21327 35689
rect 21152 35649 21164 35652
rect 21106 35643 21164 35649
rect 21269 35649 21281 35683
rect 21315 35649 21327 35683
rect 21269 35643 21327 35649
rect 2774 35572 2780 35624
rect 2832 35612 2838 35624
rect 2832 35584 2877 35612
rect 2832 35572 2838 35584
rect 16022 35572 16028 35624
rect 16080 35612 16086 35624
rect 16853 35615 16911 35621
rect 16853 35612 16865 35615
rect 16080 35584 16865 35612
rect 16080 35572 16086 35584
rect 16853 35581 16865 35584
rect 16899 35581 16911 35615
rect 16853 35575 16911 35581
rect 20714 35572 20720 35624
rect 20772 35612 20778 35624
rect 21284 35612 21312 35643
rect 20772 35584 21312 35612
rect 21468 35612 21496 35720
rect 22278 35708 22284 35720
rect 22336 35708 22342 35760
rect 21542 35640 21548 35692
rect 21600 35680 21606 35692
rect 21821 35683 21879 35689
rect 21821 35680 21833 35683
rect 21600 35652 21833 35680
rect 21600 35640 21606 35652
rect 21821 35649 21833 35652
rect 21867 35649 21879 35683
rect 23155 35683 23213 35689
rect 23155 35680 23167 35683
rect 21821 35643 21879 35649
rect 22020 35652 23167 35680
rect 21726 35612 21732 35624
rect 21468 35584 21732 35612
rect 20772 35572 20778 35584
rect 21726 35572 21732 35584
rect 21784 35572 21790 35624
rect 22020 35544 22048 35652
rect 23155 35649 23167 35652
rect 23201 35649 23213 35683
rect 23290 35680 23296 35692
rect 23251 35652 23296 35680
rect 23155 35643 23213 35649
rect 23290 35640 23296 35652
rect 23348 35640 23354 35692
rect 23382 35640 23388 35692
rect 23440 35680 23446 35692
rect 23584 35689 23612 35788
rect 24854 35776 24860 35788
rect 24912 35776 24918 35828
rect 25041 35819 25099 35825
rect 25041 35785 25053 35819
rect 25087 35816 25099 35819
rect 25406 35816 25412 35828
rect 25087 35788 25412 35816
rect 25087 35785 25099 35788
rect 25041 35779 25099 35785
rect 25406 35776 25412 35788
rect 25464 35776 25470 35828
rect 28350 35816 28356 35828
rect 28311 35788 28356 35816
rect 28350 35776 28356 35788
rect 28408 35776 28414 35828
rect 28994 35776 29000 35828
rect 29052 35816 29058 35828
rect 29089 35819 29147 35825
rect 29089 35816 29101 35819
rect 29052 35788 29101 35816
rect 29052 35776 29058 35788
rect 29089 35785 29101 35788
rect 29135 35785 29147 35819
rect 30469 35819 30527 35825
rect 30469 35816 30481 35819
rect 29089 35779 29147 35785
rect 29656 35788 30481 35816
rect 28902 35748 28908 35760
rect 25424 35720 28908 35748
rect 23569 35683 23627 35689
rect 23440 35652 23485 35680
rect 23440 35640 23446 35652
rect 23569 35649 23581 35683
rect 23615 35649 23627 35683
rect 24026 35680 24032 35692
rect 23987 35652 24032 35680
rect 23569 35643 23627 35649
rect 24026 35640 24032 35652
rect 24084 35640 24090 35692
rect 24136 35678 24256 35680
rect 24302 35678 24308 35692
rect 24136 35652 24308 35678
rect 23750 35572 23756 35624
rect 23808 35612 23814 35624
rect 24136 35612 24164 35652
rect 24228 35650 24308 35652
rect 24302 35640 24308 35650
rect 24360 35680 24366 35692
rect 25424 35689 25452 35720
rect 28902 35708 28908 35720
rect 28960 35708 28966 35760
rect 29656 35757 29684 35788
rect 30469 35785 30481 35788
rect 30515 35785 30527 35819
rect 30469 35779 30527 35785
rect 30837 35819 30895 35825
rect 30837 35785 30849 35819
rect 30883 35816 30895 35819
rect 32858 35816 32864 35828
rect 30883 35788 32864 35816
rect 30883 35785 30895 35788
rect 30837 35779 30895 35785
rect 32858 35776 32864 35788
rect 32916 35776 32922 35828
rect 29641 35751 29699 35757
rect 29641 35717 29653 35751
rect 29687 35717 29699 35751
rect 29641 35711 29699 35717
rect 30009 35751 30067 35757
rect 30009 35717 30021 35751
rect 30055 35748 30067 35751
rect 31846 35748 31852 35760
rect 30055 35720 31852 35748
rect 30055 35717 30067 35720
rect 30009 35711 30067 35717
rect 31846 35708 31852 35720
rect 31904 35708 31910 35760
rect 32030 35708 32036 35760
rect 32088 35748 32094 35760
rect 32370 35751 32428 35757
rect 32370 35748 32382 35751
rect 32088 35720 32382 35748
rect 32088 35708 32094 35720
rect 32370 35717 32382 35720
rect 32416 35717 32428 35751
rect 32370 35711 32428 35717
rect 25409 35683 25467 35689
rect 24360 35652 24405 35680
rect 24360 35640 24366 35652
rect 25409 35649 25421 35683
rect 25455 35649 25467 35683
rect 25409 35643 25467 35649
rect 25590 35640 25596 35692
rect 25648 35680 25654 35692
rect 26237 35683 26295 35689
rect 26237 35680 26249 35683
rect 25648 35652 26249 35680
rect 25648 35640 25654 35652
rect 26237 35649 26249 35652
rect 26283 35649 26295 35683
rect 26237 35643 26295 35649
rect 23808 35584 24164 35612
rect 24213 35615 24271 35621
rect 23808 35572 23814 35584
rect 24213 35581 24225 35615
rect 24259 35612 24271 35615
rect 25038 35612 25044 35624
rect 24259 35584 25044 35612
rect 24259 35581 24271 35584
rect 24213 35575 24271 35581
rect 25038 35572 25044 35584
rect 25096 35612 25102 35624
rect 25501 35615 25559 35621
rect 25501 35612 25513 35615
rect 25096 35584 25513 35612
rect 25096 35572 25102 35584
rect 25501 35581 25513 35584
rect 25547 35581 25559 35615
rect 25682 35612 25688 35624
rect 25643 35584 25688 35612
rect 25501 35575 25559 35581
rect 25682 35572 25688 35584
rect 25740 35572 25746 35624
rect 26252 35612 26280 35643
rect 26326 35640 26332 35692
rect 26384 35680 26390 35692
rect 26384 35652 26429 35680
rect 26384 35640 26390 35652
rect 27706 35640 27712 35692
rect 27764 35680 27770 35692
rect 28261 35683 28319 35689
rect 28261 35680 28273 35683
rect 27764 35652 28273 35680
rect 27764 35640 27770 35652
rect 28261 35649 28273 35652
rect 28307 35649 28319 35683
rect 28261 35643 28319 35649
rect 28718 35640 28724 35692
rect 28776 35680 28782 35692
rect 28997 35683 29055 35689
rect 28997 35680 29009 35683
rect 28776 35652 29009 35680
rect 28776 35640 28782 35652
rect 28997 35649 29009 35652
rect 29043 35649 29055 35683
rect 28997 35643 29055 35649
rect 29825 35683 29883 35689
rect 29825 35649 29837 35683
rect 29871 35649 29883 35683
rect 34790 35680 34796 35692
rect 29825 35643 29883 35649
rect 29932 35652 34796 35680
rect 28350 35612 28356 35624
rect 26252 35584 28356 35612
rect 28350 35572 28356 35584
rect 28408 35572 28414 35624
rect 28810 35572 28816 35624
rect 28868 35612 28874 35624
rect 29840 35612 29868 35643
rect 28868 35584 29868 35612
rect 28868 35572 28874 35584
rect 2746 35516 16896 35544
rect 1946 35436 1952 35488
rect 2004 35476 2010 35488
rect 2746 35476 2774 35516
rect 2004 35448 2774 35476
rect 16117 35479 16175 35485
rect 2004 35436 2010 35448
rect 16117 35445 16129 35479
rect 16163 35476 16175 35479
rect 16298 35476 16304 35488
rect 16163 35448 16304 35476
rect 16163 35445 16175 35448
rect 16117 35439 16175 35445
rect 16298 35436 16304 35448
rect 16356 35436 16362 35488
rect 16868 35476 16896 35516
rect 17788 35516 22048 35544
rect 17788 35476 17816 35516
rect 22278 35504 22284 35556
rect 22336 35544 22342 35556
rect 29932 35544 29960 35652
rect 34790 35640 34796 35652
rect 34848 35640 34854 35692
rect 45922 35640 45928 35692
rect 45980 35680 45986 35692
rect 46658 35680 46664 35692
rect 45980 35652 46664 35680
rect 45980 35640 45986 35652
rect 46658 35640 46664 35652
rect 46716 35680 46722 35692
rect 46845 35683 46903 35689
rect 46845 35680 46857 35683
rect 46716 35652 46857 35680
rect 46716 35640 46722 35652
rect 46845 35649 46857 35652
rect 46891 35649 46903 35683
rect 47854 35680 47860 35692
rect 47815 35652 47860 35680
rect 46845 35643 46903 35649
rect 47854 35640 47860 35652
rect 47912 35640 47918 35692
rect 30929 35615 30987 35621
rect 30929 35612 30941 35615
rect 22336 35516 29960 35544
rect 30024 35584 30941 35612
rect 22336 35504 22342 35516
rect 20622 35476 20628 35488
rect 16868 35448 17816 35476
rect 20583 35448 20628 35476
rect 20622 35436 20628 35448
rect 20680 35436 20686 35488
rect 23566 35436 23572 35488
rect 23624 35476 23630 35488
rect 24029 35479 24087 35485
rect 24029 35476 24041 35479
rect 23624 35448 24041 35476
rect 23624 35436 23630 35448
rect 24029 35445 24041 35448
rect 24075 35445 24087 35479
rect 24486 35476 24492 35488
rect 24447 35448 24492 35476
rect 24029 35439 24087 35445
rect 24486 35436 24492 35448
rect 24544 35436 24550 35488
rect 24578 35436 24584 35488
rect 24636 35476 24642 35488
rect 29178 35476 29184 35488
rect 24636 35448 29184 35476
rect 24636 35436 24642 35448
rect 29178 35436 29184 35448
rect 29236 35436 29242 35488
rect 29270 35436 29276 35488
rect 29328 35476 29334 35488
rect 30024 35476 30052 35584
rect 30929 35581 30941 35584
rect 30975 35581 30987 35615
rect 30929 35575 30987 35581
rect 31021 35615 31079 35621
rect 31021 35581 31033 35615
rect 31067 35581 31079 35615
rect 31021 35575 31079 35581
rect 32125 35615 32183 35621
rect 32125 35581 32137 35615
rect 32171 35581 32183 35615
rect 32125 35575 32183 35581
rect 30282 35504 30288 35556
rect 30340 35544 30346 35556
rect 31036 35544 31064 35575
rect 30340 35516 31064 35544
rect 30340 35504 30346 35516
rect 29328 35448 30052 35476
rect 29328 35436 29334 35448
rect 31478 35436 31484 35488
rect 31536 35476 31542 35488
rect 32140 35476 32168 35575
rect 32490 35476 32496 35488
rect 31536 35448 32496 35476
rect 31536 35436 31542 35448
rect 32490 35436 32496 35448
rect 32548 35436 32554 35488
rect 32858 35436 32864 35488
rect 32916 35476 32922 35488
rect 33505 35479 33563 35485
rect 33505 35476 33517 35479
rect 32916 35448 33517 35476
rect 32916 35436 32922 35448
rect 33505 35445 33517 35448
rect 33551 35445 33563 35479
rect 46934 35476 46940 35488
rect 46895 35448 46940 35476
rect 33505 35439 33563 35445
rect 46934 35436 46940 35448
rect 46992 35436 46998 35488
rect 47578 35436 47584 35488
rect 47636 35476 47642 35488
rect 48041 35479 48099 35485
rect 48041 35476 48053 35479
rect 47636 35448 48053 35476
rect 47636 35436 47642 35448
rect 48041 35445 48053 35448
rect 48087 35445 48099 35479
rect 48041 35439 48099 35445
rect 1104 35386 48852 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 48852 35386
rect 1104 35312 48852 35334
rect 1946 35272 1952 35284
rect 1907 35244 1952 35272
rect 1946 35232 1952 35244
rect 2004 35232 2010 35284
rect 15838 35272 15844 35284
rect 15799 35244 15844 35272
rect 15838 35232 15844 35244
rect 15896 35232 15902 35284
rect 17402 35232 17408 35284
rect 17460 35272 17466 35284
rect 17497 35275 17555 35281
rect 17497 35272 17509 35275
rect 17460 35244 17509 35272
rect 17460 35232 17466 35244
rect 17497 35241 17509 35244
rect 17543 35241 17555 35275
rect 20438 35272 20444 35284
rect 17497 35235 17555 35241
rect 20088 35244 20444 35272
rect 11514 35096 11520 35148
rect 11572 35136 11578 35148
rect 18325 35139 18383 35145
rect 18325 35136 18337 35139
rect 11572 35108 12296 35136
rect 11572 35096 11578 35108
rect 12158 35068 12164 35080
rect 12119 35040 12164 35068
rect 12158 35028 12164 35040
rect 12216 35028 12222 35080
rect 12268 35068 12296 35108
rect 16040 35108 18337 35136
rect 16040 35068 16068 35108
rect 18325 35105 18337 35108
rect 18371 35105 18383 35139
rect 18325 35099 18383 35105
rect 12268 35040 16068 35068
rect 16117 35071 16175 35077
rect 16117 35037 16129 35071
rect 16163 35037 16175 35071
rect 16117 35031 16175 35037
rect 16209 35071 16267 35077
rect 16209 35037 16221 35071
rect 16255 35037 16267 35071
rect 16209 35031 16267 35037
rect 1854 35000 1860 35012
rect 1815 34972 1860 35000
rect 1854 34960 1860 34972
rect 1912 34960 1918 35012
rect 12250 34960 12256 35012
rect 12308 35000 12314 35012
rect 12406 35003 12464 35009
rect 12406 35000 12418 35003
rect 12308 34972 12418 35000
rect 12308 34960 12314 34972
rect 12406 34969 12418 34972
rect 12452 34969 12464 35003
rect 12406 34963 12464 34969
rect 15102 34960 15108 35012
rect 15160 35000 15166 35012
rect 16132 35000 16160 35031
rect 15160 34972 16160 35000
rect 15160 34960 15166 34972
rect 13541 34935 13599 34941
rect 13541 34901 13553 34935
rect 13587 34932 13599 34935
rect 14182 34932 14188 34944
rect 13587 34904 14188 34932
rect 13587 34901 13599 34904
rect 13541 34895 13599 34901
rect 14182 34892 14188 34904
rect 14240 34892 14246 34944
rect 16224 34932 16252 35031
rect 16298 35028 16304 35080
rect 16356 35068 16362 35080
rect 16485 35071 16543 35077
rect 16356 35040 16401 35068
rect 16356 35028 16362 35040
rect 16485 35037 16497 35071
rect 16531 35037 16543 35071
rect 16485 35031 16543 35037
rect 16500 35000 16528 35031
rect 16758 35028 16764 35080
rect 16816 35068 16822 35080
rect 17129 35071 17187 35077
rect 17129 35068 17141 35071
rect 16816 35040 17141 35068
rect 16816 35028 16822 35040
rect 17129 35037 17141 35040
rect 17175 35037 17187 35071
rect 17129 35031 17187 35037
rect 17313 35071 17371 35077
rect 17313 35037 17325 35071
rect 17359 35068 17371 35071
rect 17954 35068 17960 35080
rect 17359 35040 17960 35068
rect 17359 35037 17371 35040
rect 17313 35031 17371 35037
rect 17954 35028 17960 35040
rect 18012 35028 18018 35080
rect 18049 35071 18107 35077
rect 18049 35037 18061 35071
rect 18095 35068 18107 35071
rect 18095 35040 18276 35068
rect 18095 35037 18107 35040
rect 18049 35031 18107 35037
rect 17586 35000 17592 35012
rect 16500 34972 17592 35000
rect 17586 34960 17592 34972
rect 17644 34960 17650 35012
rect 17034 34932 17040 34944
rect 16224 34904 17040 34932
rect 17034 34892 17040 34904
rect 17092 34892 17098 34944
rect 18248 34932 18276 35040
rect 18340 35000 18368 35099
rect 19978 35096 19984 35148
rect 20036 35136 20042 35148
rect 20088 35145 20116 35244
rect 20438 35232 20444 35244
rect 20496 35232 20502 35284
rect 45922 35272 45928 35284
rect 22066 35244 45928 35272
rect 22066 35204 22094 35244
rect 45922 35232 45928 35244
rect 45980 35232 45986 35284
rect 27614 35204 27620 35216
rect 21100 35176 22094 35204
rect 27575 35176 27620 35204
rect 20073 35139 20131 35145
rect 20073 35136 20085 35139
rect 20036 35108 20085 35136
rect 20036 35096 20042 35108
rect 20073 35105 20085 35108
rect 20119 35105 20131 35139
rect 20073 35099 20131 35105
rect 18414 35028 18420 35080
rect 18472 35068 18478 35080
rect 19150 35068 19156 35080
rect 18472 35040 19156 35068
rect 18472 35028 18478 35040
rect 19150 35028 19156 35040
rect 19208 35068 19214 35080
rect 19245 35071 19303 35077
rect 19245 35068 19257 35071
rect 19208 35040 19257 35068
rect 19208 35028 19214 35040
rect 19245 35037 19257 35040
rect 19291 35037 19303 35071
rect 19245 35031 19303 35037
rect 20340 35071 20398 35077
rect 20340 35037 20352 35071
rect 20386 35068 20398 35071
rect 20622 35068 20628 35080
rect 20386 35040 20628 35068
rect 20386 35037 20398 35040
rect 20340 35031 20398 35037
rect 20622 35028 20628 35040
rect 20680 35028 20686 35080
rect 21100 35000 21128 35176
rect 27614 35164 27620 35176
rect 27672 35164 27678 35216
rect 28077 35207 28135 35213
rect 28077 35173 28089 35207
rect 28123 35204 28135 35207
rect 28810 35204 28816 35216
rect 28123 35176 28816 35204
rect 28123 35173 28135 35176
rect 28077 35167 28135 35173
rect 28810 35164 28816 35176
rect 28868 35164 28874 35216
rect 28997 35207 29055 35213
rect 28997 35173 29009 35207
rect 29043 35204 29055 35207
rect 30282 35204 30288 35216
rect 29043 35176 30288 35204
rect 29043 35173 29055 35176
rect 28997 35167 29055 35173
rect 30282 35164 30288 35176
rect 30340 35204 30346 35216
rect 30340 35176 30420 35204
rect 30340 35164 30346 35176
rect 22554 35136 22560 35148
rect 22467 35108 22560 35136
rect 22554 35096 22560 35108
rect 22612 35136 22618 35148
rect 24578 35136 24584 35148
rect 22612 35108 24584 35136
rect 22612 35096 22618 35108
rect 24578 35096 24584 35108
rect 24636 35096 24642 35148
rect 30392 35145 30420 35176
rect 31018 35164 31024 35216
rect 31076 35204 31082 35216
rect 31205 35207 31263 35213
rect 31205 35204 31217 35207
rect 31076 35176 31217 35204
rect 31076 35164 31082 35176
rect 31205 35173 31217 35176
rect 31251 35173 31263 35207
rect 31205 35167 31263 35173
rect 30377 35139 30435 35145
rect 26620 35108 30328 35136
rect 22005 35071 22063 35077
rect 22005 35068 22017 35071
rect 18340 34972 21128 35000
rect 21192 35040 22017 35068
rect 19242 34932 19248 34944
rect 18248 34904 19248 34932
rect 19242 34892 19248 34904
rect 19300 34932 19306 34944
rect 19429 34935 19487 34941
rect 19429 34932 19441 34935
rect 19300 34904 19441 34932
rect 19300 34892 19306 34904
rect 19429 34901 19441 34904
rect 19475 34932 19487 34935
rect 20806 34932 20812 34944
rect 19475 34904 20812 34932
rect 19475 34901 19487 34904
rect 19429 34895 19487 34901
rect 20806 34892 20812 34904
rect 20864 34932 20870 34944
rect 21192 34932 21220 35040
rect 22005 35037 22017 35040
rect 22051 35037 22063 35071
rect 22005 35031 22063 35037
rect 23290 35028 23296 35080
rect 23348 35068 23354 35080
rect 26620 35077 26648 35108
rect 23385 35071 23443 35077
rect 23385 35068 23397 35071
rect 23348 35040 23397 35068
rect 23348 35028 23354 35040
rect 23385 35037 23397 35040
rect 23431 35068 23443 35071
rect 26605 35071 26663 35077
rect 23431 35040 25728 35068
rect 23431 35037 23443 35040
rect 23385 35031 23443 35037
rect 23934 34960 23940 35012
rect 23992 35000 23998 35012
rect 24857 35003 24915 35009
rect 24857 35000 24869 35003
rect 23992 34972 24869 35000
rect 23992 34960 23998 34972
rect 24857 34969 24869 34972
rect 24903 34969 24915 35003
rect 24857 34963 24915 34969
rect 25041 35003 25099 35009
rect 25041 34969 25053 35003
rect 25087 35000 25099 35003
rect 25590 35000 25596 35012
rect 25087 34972 25596 35000
rect 25087 34969 25099 34972
rect 25041 34963 25099 34969
rect 25590 34960 25596 34972
rect 25648 34960 25654 35012
rect 25700 35000 25728 35040
rect 26605 35037 26617 35071
rect 26651 35037 26663 35071
rect 26605 35031 26663 35037
rect 26786 35028 26792 35080
rect 26844 35068 26850 35080
rect 28261 35071 28319 35077
rect 28261 35068 28273 35071
rect 26844 35040 28273 35068
rect 26844 35028 26850 35040
rect 28261 35037 28273 35040
rect 28307 35037 28319 35071
rect 28261 35031 28319 35037
rect 28350 35028 28356 35080
rect 28408 35068 28414 35080
rect 28813 35071 28871 35077
rect 28813 35068 28825 35071
rect 28408 35040 28825 35068
rect 28408 35028 28414 35040
rect 28813 35037 28825 35040
rect 28859 35068 28871 35071
rect 29730 35068 29736 35080
rect 28859 35040 29736 35068
rect 28859 35037 28871 35040
rect 28813 35031 28871 35037
rect 29730 35028 29736 35040
rect 29788 35028 29794 35080
rect 30300 35068 30328 35108
rect 30377 35105 30389 35139
rect 30423 35105 30435 35139
rect 30377 35099 30435 35105
rect 30742 35068 30748 35080
rect 30300 35040 30748 35068
rect 30742 35028 30748 35040
rect 30800 35028 30806 35080
rect 31220 35068 31248 35167
rect 31570 35164 31576 35216
rect 31628 35204 31634 35216
rect 31628 35176 32260 35204
rect 31628 35164 31634 35176
rect 31662 35096 31668 35148
rect 31720 35136 31726 35148
rect 31720 35108 31984 35136
rect 31720 35096 31726 35108
rect 31956 35077 31984 35108
rect 32232 35077 32260 35176
rect 31849 35071 31907 35077
rect 31849 35068 31861 35071
rect 31220 35040 31861 35068
rect 31844 35037 31861 35040
rect 31895 35037 31907 35071
rect 31849 35031 31907 35037
rect 31941 35071 31999 35077
rect 31941 35037 31953 35071
rect 31987 35037 31999 35071
rect 31941 35031 31999 35037
rect 32033 35071 32091 35077
rect 32033 35037 32045 35071
rect 32079 35037 32091 35071
rect 32033 35031 32091 35037
rect 32217 35071 32275 35077
rect 32217 35037 32229 35071
rect 32263 35037 32275 35071
rect 32217 35031 32275 35037
rect 26804 35000 26832 35028
rect 27246 35000 27252 35012
rect 25700 34972 26832 35000
rect 27207 34972 27252 35000
rect 27246 34960 27252 34972
rect 27304 34960 27310 35012
rect 27338 34960 27344 35012
rect 27396 35000 27402 35012
rect 27433 35003 27491 35009
rect 27433 35000 27445 35003
rect 27396 34972 27445 35000
rect 27396 34960 27402 34972
rect 27433 34969 27445 34972
rect 27479 34969 27491 35003
rect 27433 34963 27491 34969
rect 27890 34960 27896 35012
rect 27948 35000 27954 35012
rect 28718 35000 28724 35012
rect 27948 34972 28724 35000
rect 27948 34960 27954 34972
rect 28718 34960 28724 34972
rect 28776 34960 28782 35012
rect 28902 34960 28908 35012
rect 28960 35000 28966 35012
rect 30285 35003 30343 35009
rect 30285 35000 30297 35003
rect 28960 34972 30297 35000
rect 28960 34960 28966 34972
rect 30285 34969 30297 34972
rect 30331 34969 30343 35003
rect 31570 35000 31576 35012
rect 31531 34972 31576 35000
rect 30285 34963 30343 34969
rect 31570 34960 31576 34972
rect 31628 34960 31634 35012
rect 31662 34960 31668 35012
rect 31720 35000 31726 35012
rect 32048 35000 32076 35031
rect 32490 35028 32496 35080
rect 32548 35068 32554 35080
rect 32769 35071 32827 35077
rect 32769 35068 32781 35071
rect 32548 35040 32781 35068
rect 32548 35028 32554 35040
rect 32769 35037 32781 35040
rect 32815 35037 32827 35071
rect 32769 35031 32827 35037
rect 45833 35071 45891 35077
rect 45833 35037 45845 35071
rect 45879 35068 45891 35071
rect 46293 35071 46351 35077
rect 46293 35068 46305 35071
rect 45879 35040 46305 35068
rect 45879 35037 45891 35040
rect 45833 35031 45891 35037
rect 46293 35037 46305 35040
rect 46339 35037 46351 35071
rect 46293 35031 46351 35037
rect 33042 35009 33048 35012
rect 33036 35000 33048 35009
rect 31720 34972 32076 35000
rect 33003 34972 33048 35000
rect 31720 34960 31726 34972
rect 33036 34963 33048 34972
rect 33042 34960 33048 34963
rect 33100 34960 33106 35012
rect 46477 35003 46535 35009
rect 46477 34969 46489 35003
rect 46523 35000 46535 35003
rect 47670 35000 47676 35012
rect 46523 34972 47676 35000
rect 46523 34969 46535 34972
rect 46477 34963 46535 34969
rect 47670 34960 47676 34972
rect 47728 34960 47734 35012
rect 48130 35000 48136 35012
rect 48091 34972 48136 35000
rect 48130 34960 48136 34972
rect 48188 34960 48194 35012
rect 20864 34904 21220 34932
rect 21453 34935 21511 34941
rect 20864 34892 20870 34904
rect 21453 34901 21465 34935
rect 21499 34932 21511 34935
rect 22278 34932 22284 34944
rect 21499 34904 22284 34932
rect 21499 34901 21511 34904
rect 21453 34895 21511 34901
rect 22278 34892 22284 34904
rect 22336 34892 22342 34944
rect 22922 34892 22928 34944
rect 22980 34932 22986 34944
rect 23198 34932 23204 34944
rect 22980 34904 23204 34932
rect 22980 34892 22986 34904
rect 23198 34892 23204 34904
rect 23256 34892 23262 34944
rect 24394 34892 24400 34944
rect 24452 34932 24458 34944
rect 25682 34932 25688 34944
rect 24452 34904 25688 34932
rect 24452 34892 24458 34904
rect 25682 34892 25688 34904
rect 25740 34892 25746 34944
rect 26694 34932 26700 34944
rect 26655 34904 26700 34932
rect 26694 34892 26700 34904
rect 26752 34892 26758 34944
rect 29822 34932 29828 34944
rect 29783 34904 29828 34932
rect 29822 34892 29828 34904
rect 29880 34892 29886 34944
rect 30190 34932 30196 34944
rect 30151 34904 30196 34932
rect 30190 34892 30196 34904
rect 30248 34892 30254 34944
rect 34149 34935 34207 34941
rect 34149 34901 34161 34935
rect 34195 34932 34207 34935
rect 34238 34932 34244 34944
rect 34195 34904 34244 34932
rect 34195 34901 34207 34904
rect 34149 34895 34207 34901
rect 34238 34892 34244 34904
rect 34296 34892 34302 34944
rect 1104 34842 48852 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 48852 34842
rect 1104 34768 48852 34790
rect 12161 34731 12219 34737
rect 12161 34697 12173 34731
rect 12207 34728 12219 34731
rect 12250 34728 12256 34740
rect 12207 34700 12256 34728
rect 12207 34697 12219 34700
rect 12161 34691 12219 34697
rect 12250 34688 12256 34700
rect 12308 34688 12314 34740
rect 12526 34688 12532 34740
rect 12584 34688 12590 34740
rect 14737 34731 14795 34737
rect 14737 34697 14749 34731
rect 14783 34728 14795 34731
rect 14783 34700 19104 34728
rect 14783 34697 14795 34700
rect 14737 34691 14795 34697
rect 2038 34592 2044 34604
rect 1951 34564 2044 34592
rect 2038 34552 2044 34564
rect 2096 34592 2102 34604
rect 2498 34592 2504 34604
rect 2096 34564 2504 34592
rect 2096 34552 2102 34564
rect 2498 34552 2504 34564
rect 2556 34552 2562 34604
rect 12544 34601 12572 34688
rect 15841 34663 15899 34669
rect 15841 34629 15853 34663
rect 15887 34660 15899 34663
rect 18141 34663 18199 34669
rect 18141 34660 18153 34663
rect 15887 34632 18153 34660
rect 15887 34629 15899 34632
rect 15841 34623 15899 34629
rect 18141 34629 18153 34632
rect 18187 34660 18199 34663
rect 18966 34660 18972 34672
rect 18187 34632 18972 34660
rect 18187 34629 18199 34632
rect 18141 34623 18199 34629
rect 18966 34620 18972 34632
rect 19024 34620 19030 34672
rect 19076 34660 19104 34700
rect 21726 34688 21732 34740
rect 21784 34728 21790 34740
rect 21821 34731 21879 34737
rect 21821 34728 21833 34731
rect 21784 34700 21833 34728
rect 21784 34688 21790 34700
rect 21821 34697 21833 34700
rect 21867 34697 21879 34731
rect 21821 34691 21879 34697
rect 27246 34688 27252 34740
rect 27304 34728 27310 34740
rect 27433 34731 27491 34737
rect 27433 34728 27445 34731
rect 27304 34700 27445 34728
rect 27304 34688 27310 34700
rect 27433 34697 27445 34700
rect 27479 34697 27491 34731
rect 27433 34691 27491 34697
rect 27801 34731 27859 34737
rect 27801 34697 27813 34731
rect 27847 34728 27859 34731
rect 29270 34728 29276 34740
rect 27847 34700 29276 34728
rect 27847 34697 27859 34700
rect 27801 34691 27859 34697
rect 29270 34688 29276 34700
rect 29328 34688 29334 34740
rect 30006 34728 30012 34740
rect 29472 34700 30012 34728
rect 23842 34660 23848 34672
rect 19076 34632 23848 34660
rect 23842 34620 23848 34632
rect 23900 34620 23906 34672
rect 29472 34669 29500 34700
rect 30006 34688 30012 34700
rect 30064 34688 30070 34740
rect 41046 34688 41052 34740
rect 41104 34728 41110 34740
rect 47670 34728 47676 34740
rect 41104 34700 47532 34728
rect 47631 34700 47676 34728
rect 41104 34688 41110 34700
rect 27893 34663 27951 34669
rect 27893 34660 27905 34663
rect 24780 34632 25176 34660
rect 12437 34595 12495 34601
rect 12437 34561 12449 34595
rect 12483 34561 12495 34595
rect 12437 34555 12495 34561
rect 12529 34595 12587 34601
rect 12529 34561 12541 34595
rect 12575 34561 12587 34595
rect 12529 34555 12587 34561
rect 12621 34595 12679 34601
rect 12621 34561 12633 34595
rect 12667 34561 12679 34595
rect 12621 34555 12679 34561
rect 12805 34595 12863 34601
rect 12805 34561 12817 34595
rect 12851 34592 12863 34595
rect 12986 34592 12992 34604
rect 12851 34564 12992 34592
rect 12851 34561 12863 34564
rect 12805 34555 12863 34561
rect 1854 34484 1860 34536
rect 1912 34524 1918 34536
rect 2685 34527 2743 34533
rect 2685 34524 2697 34527
rect 1912 34496 2697 34524
rect 1912 34484 1918 34496
rect 2685 34493 2697 34496
rect 2731 34493 2743 34527
rect 2685 34487 2743 34493
rect 12443 34468 12471 34555
rect 12636 34524 12664 34555
rect 12986 34552 12992 34564
rect 13044 34552 13050 34604
rect 13630 34592 13636 34604
rect 13591 34564 13636 34592
rect 13630 34552 13636 34564
rect 13688 34552 13694 34604
rect 13814 34592 13820 34604
rect 13775 34564 13820 34592
rect 13814 34552 13820 34564
rect 13872 34552 13878 34604
rect 14458 34592 14464 34604
rect 14419 34564 14464 34592
rect 14458 34552 14464 34564
rect 14516 34552 14522 34604
rect 14642 34592 14648 34604
rect 14603 34564 14648 34592
rect 14642 34552 14648 34564
rect 14700 34552 14706 34604
rect 16899 34595 16957 34601
rect 16899 34592 16911 34595
rect 14752 34564 16911 34592
rect 12894 34524 12900 34536
rect 12636 34496 12900 34524
rect 12894 34484 12900 34496
rect 12952 34484 12958 34536
rect 13725 34527 13783 34533
rect 13725 34493 13737 34527
rect 13771 34524 13783 34527
rect 13906 34524 13912 34536
rect 13771 34496 13912 34524
rect 13771 34493 13783 34496
rect 13725 34487 13783 34493
rect 13906 34484 13912 34496
rect 13964 34484 13970 34536
rect 14182 34484 14188 34536
rect 14240 34524 14246 34536
rect 14752 34524 14780 34564
rect 16899 34561 16911 34564
rect 16945 34561 16957 34595
rect 17034 34592 17040 34604
rect 16995 34564 17040 34592
rect 16899 34555 16957 34561
rect 17034 34552 17040 34564
rect 17092 34552 17098 34604
rect 17129 34595 17187 34601
rect 17129 34561 17141 34595
rect 17175 34592 17187 34595
rect 17218 34592 17224 34604
rect 17175 34564 17224 34592
rect 17175 34561 17187 34564
rect 17129 34555 17187 34561
rect 17218 34552 17224 34564
rect 17276 34552 17282 34604
rect 17313 34595 17371 34601
rect 17313 34561 17325 34595
rect 17359 34561 17371 34595
rect 17954 34592 17960 34604
rect 17915 34564 17960 34592
rect 17313 34555 17371 34561
rect 16022 34524 16028 34536
rect 14240 34496 14780 34524
rect 15983 34496 16028 34524
rect 14240 34484 14246 34496
rect 16022 34484 16028 34496
rect 16080 34484 16086 34536
rect 17328 34524 17356 34555
rect 17954 34552 17960 34564
rect 18012 34552 18018 34604
rect 19429 34595 19487 34601
rect 19429 34561 19441 34595
rect 19475 34592 19487 34595
rect 20806 34592 20812 34604
rect 19475 34564 20812 34592
rect 19475 34561 19487 34564
rect 19429 34555 19487 34561
rect 20806 34552 20812 34564
rect 20864 34552 20870 34604
rect 21174 34592 21180 34604
rect 21135 34564 21180 34592
rect 21174 34552 21180 34564
rect 21232 34552 21238 34604
rect 21634 34552 21640 34604
rect 21692 34592 21698 34604
rect 22005 34595 22063 34601
rect 22005 34592 22017 34595
rect 21692 34564 22017 34592
rect 21692 34552 21698 34564
rect 22005 34561 22017 34564
rect 22051 34561 22063 34595
rect 22186 34592 22192 34604
rect 22147 34564 22192 34592
rect 22005 34555 22063 34561
rect 22186 34552 22192 34564
rect 22244 34552 22250 34604
rect 22278 34552 22284 34604
rect 22336 34592 22342 34604
rect 23385 34595 23443 34601
rect 22336 34564 23336 34592
rect 22336 34552 22342 34564
rect 17586 34524 17592 34536
rect 17328 34496 17592 34524
rect 17586 34484 17592 34496
rect 17644 34524 17650 34536
rect 19702 34524 19708 34536
rect 17644 34496 19708 34524
rect 17644 34484 17650 34496
rect 19702 34484 19708 34496
rect 19760 34484 19766 34536
rect 20073 34527 20131 34533
rect 20073 34493 20085 34527
rect 20119 34524 20131 34527
rect 21082 34524 21088 34536
rect 20119 34496 21088 34524
rect 20119 34493 20131 34496
rect 20073 34487 20131 34493
rect 21082 34484 21088 34496
rect 21140 34484 21146 34536
rect 12434 34416 12440 34468
rect 12492 34416 12498 34468
rect 1394 34348 1400 34400
rect 1452 34388 1458 34400
rect 1581 34391 1639 34397
rect 1581 34388 1593 34391
rect 1452 34360 1593 34388
rect 1452 34348 1458 34360
rect 1581 34357 1593 34360
rect 1627 34357 1639 34391
rect 2130 34388 2136 34400
rect 2091 34360 2136 34388
rect 1581 34351 1639 34357
rect 2130 34348 2136 34360
rect 2188 34348 2194 34400
rect 8478 34348 8484 34400
rect 8536 34388 8542 34400
rect 15654 34388 15660 34400
rect 8536 34360 15660 34388
rect 8536 34348 8542 34360
rect 15654 34348 15660 34360
rect 15712 34348 15718 34400
rect 16669 34391 16727 34397
rect 16669 34357 16681 34391
rect 16715 34388 16727 34391
rect 17310 34388 17316 34400
rect 16715 34360 17316 34388
rect 16715 34357 16727 34360
rect 16669 34351 16727 34357
rect 17310 34348 17316 34360
rect 17368 34348 17374 34400
rect 23014 34388 23020 34400
rect 22975 34360 23020 34388
rect 23014 34348 23020 34360
rect 23072 34348 23078 34400
rect 23308 34388 23336 34564
rect 23385 34561 23397 34595
rect 23431 34592 23443 34595
rect 23566 34592 23572 34604
rect 23431 34564 23572 34592
rect 23431 34561 23443 34564
rect 23385 34555 23443 34561
rect 23566 34552 23572 34564
rect 23624 34552 23630 34604
rect 24210 34592 24216 34604
rect 24171 34564 24216 34592
rect 24210 34552 24216 34564
rect 24268 34552 24274 34604
rect 24397 34595 24455 34601
rect 24397 34561 24409 34595
rect 24443 34592 24455 34595
rect 24578 34592 24584 34604
rect 24443 34564 24584 34592
rect 24443 34561 24455 34564
rect 24397 34555 24455 34561
rect 24578 34552 24584 34564
rect 24636 34552 24642 34604
rect 23474 34524 23480 34536
rect 23435 34496 23480 34524
rect 23474 34484 23480 34496
rect 23532 34484 23538 34536
rect 23661 34527 23719 34533
rect 23661 34493 23673 34527
rect 23707 34493 23719 34527
rect 24780 34524 24808 34632
rect 25038 34592 25044 34604
rect 24999 34564 25044 34592
rect 25038 34552 25044 34564
rect 25096 34552 25102 34604
rect 25148 34601 25176 34632
rect 25240 34632 27905 34660
rect 25133 34595 25191 34601
rect 25133 34561 25145 34595
rect 25179 34561 25191 34595
rect 25133 34555 25191 34561
rect 23661 34487 23719 34493
rect 24596 34496 24808 34524
rect 23676 34456 23704 34487
rect 24394 34456 24400 34468
rect 23676 34428 24400 34456
rect 24394 34416 24400 34428
rect 24452 34416 24458 34468
rect 24596 34465 24624 34496
rect 24854 34484 24860 34536
rect 24912 34524 24918 34536
rect 25240 34524 25268 34632
rect 27893 34629 27905 34632
rect 27939 34629 27951 34663
rect 27893 34623 27951 34629
rect 29457 34663 29515 34669
rect 29457 34629 29469 34663
rect 29503 34629 29515 34663
rect 29457 34623 29515 34629
rect 29822 34620 29828 34672
rect 29880 34660 29886 34672
rect 30377 34663 30435 34669
rect 30377 34660 30389 34663
rect 29880 34632 30389 34660
rect 29880 34620 29886 34632
rect 30377 34629 30389 34632
rect 30423 34629 30435 34663
rect 30377 34623 30435 34629
rect 30561 34663 30619 34669
rect 30561 34629 30573 34663
rect 30607 34660 30619 34663
rect 30926 34660 30932 34672
rect 30607 34632 30932 34660
rect 30607 34629 30619 34632
rect 30561 34623 30619 34629
rect 30926 34620 30932 34632
rect 30984 34620 30990 34672
rect 47394 34660 47400 34672
rect 45204 34632 47400 34660
rect 25958 34592 25964 34604
rect 25919 34564 25964 34592
rect 25958 34552 25964 34564
rect 26016 34552 26022 34604
rect 26237 34595 26295 34601
rect 26237 34561 26249 34595
rect 26283 34592 26295 34595
rect 26418 34592 26424 34604
rect 26283 34564 26424 34592
rect 26283 34561 26295 34564
rect 26237 34555 26295 34561
rect 26418 34552 26424 34564
rect 26476 34552 26482 34604
rect 28902 34592 28908 34604
rect 27908 34564 28908 34592
rect 24912 34496 25268 34524
rect 26145 34527 26203 34533
rect 24912 34484 24918 34496
rect 26145 34493 26157 34527
rect 26191 34524 26203 34527
rect 27908 34524 27936 34564
rect 28902 34552 28908 34564
rect 28960 34552 28966 34604
rect 29733 34595 29791 34601
rect 29733 34561 29745 34595
rect 29779 34592 29791 34595
rect 30098 34592 30104 34604
rect 29779 34564 30104 34592
rect 29779 34561 29791 34564
rect 29733 34555 29791 34561
rect 30098 34552 30104 34564
rect 30156 34552 30162 34604
rect 45204 34601 45232 34632
rect 47394 34620 47400 34632
rect 47452 34620 47458 34672
rect 45189 34595 45247 34601
rect 45189 34561 45201 34595
rect 45235 34561 45247 34595
rect 47504 34592 47532 34700
rect 47670 34688 47676 34700
rect 47728 34688 47734 34740
rect 47581 34595 47639 34601
rect 47581 34592 47593 34595
rect 47504 34564 47593 34592
rect 45189 34555 45247 34561
rect 47581 34561 47593 34564
rect 47627 34592 47639 34595
rect 47854 34592 47860 34604
rect 47627 34564 47860 34592
rect 47627 34561 47639 34564
rect 47581 34555 47639 34561
rect 47854 34552 47860 34564
rect 47912 34552 47918 34604
rect 26191 34496 27936 34524
rect 28077 34527 28135 34533
rect 26191 34493 26203 34496
rect 26145 34487 26203 34493
rect 28077 34493 28089 34527
rect 28123 34493 28135 34527
rect 28077 34487 28135 34493
rect 29641 34527 29699 34533
rect 29641 34493 29653 34527
rect 29687 34524 29699 34527
rect 29914 34524 29920 34536
rect 29687 34496 29920 34524
rect 29687 34493 29699 34496
rect 29641 34487 29699 34493
rect 24581 34459 24639 34465
rect 24581 34425 24593 34459
rect 24627 34425 24639 34459
rect 24581 34419 24639 34425
rect 25866 34416 25872 34468
rect 25924 34456 25930 34468
rect 28092 34456 28120 34487
rect 29914 34484 29920 34496
rect 29972 34484 29978 34536
rect 45373 34527 45431 34533
rect 45373 34493 45385 34527
rect 45419 34524 45431 34527
rect 46382 34524 46388 34536
rect 45419 34496 46388 34524
rect 45419 34493 45431 34496
rect 45373 34487 45431 34493
rect 46382 34484 46388 34496
rect 46440 34484 46446 34536
rect 46845 34527 46903 34533
rect 46845 34493 46857 34527
rect 46891 34493 46903 34527
rect 46845 34487 46903 34493
rect 28442 34456 28448 34468
rect 25924 34428 26556 34456
rect 28092 34428 28448 34456
rect 25924 34416 25930 34428
rect 24302 34388 24308 34400
rect 23308 34360 24308 34388
rect 24302 34348 24308 34360
rect 24360 34348 24366 34400
rect 24486 34348 24492 34400
rect 24544 34388 24550 34400
rect 25041 34391 25099 34397
rect 25041 34388 25053 34391
rect 24544 34360 25053 34388
rect 24544 34348 24550 34360
rect 25041 34357 25053 34360
rect 25087 34357 25099 34391
rect 25041 34351 25099 34357
rect 25409 34391 25467 34397
rect 25409 34357 25421 34391
rect 25455 34388 25467 34391
rect 25498 34388 25504 34400
rect 25455 34360 25504 34388
rect 25455 34357 25467 34360
rect 25409 34351 25467 34357
rect 25498 34348 25504 34360
rect 25556 34348 25562 34400
rect 26142 34388 26148 34400
rect 26103 34360 26148 34388
rect 26142 34348 26148 34360
rect 26200 34348 26206 34400
rect 26418 34388 26424 34400
rect 26379 34360 26424 34388
rect 26418 34348 26424 34360
rect 26476 34348 26482 34400
rect 26528 34388 26556 34428
rect 28442 34416 28448 34428
rect 28500 34416 28506 34468
rect 28552 34428 29960 34456
rect 28552 34388 28580 34428
rect 26528 34360 28580 34388
rect 29270 34348 29276 34400
rect 29328 34388 29334 34400
rect 29932 34397 29960 34428
rect 46860 34400 46888 34487
rect 29457 34391 29515 34397
rect 29457 34388 29469 34391
rect 29328 34360 29469 34388
rect 29328 34348 29334 34360
rect 29457 34357 29469 34360
rect 29503 34357 29515 34391
rect 29457 34351 29515 34357
rect 29917 34391 29975 34397
rect 29917 34357 29929 34391
rect 29963 34357 29975 34391
rect 29917 34351 29975 34357
rect 30745 34391 30803 34397
rect 30745 34357 30757 34391
rect 30791 34388 30803 34391
rect 30834 34388 30840 34400
rect 30791 34360 30840 34388
rect 30791 34357 30803 34360
rect 30745 34351 30803 34357
rect 30834 34348 30840 34360
rect 30892 34348 30898 34400
rect 46842 34348 46848 34400
rect 46900 34348 46906 34400
rect 1104 34298 48852 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 48852 34298
rect 1104 34224 48852 34246
rect 12158 34184 12164 34196
rect 10336 34156 12164 34184
rect 8294 34076 8300 34128
rect 8352 34116 8358 34128
rect 10336 34116 10364 34156
rect 12158 34144 12164 34156
rect 12216 34144 12222 34196
rect 14093 34187 14151 34193
rect 14093 34184 14105 34187
rect 12406 34156 14105 34184
rect 8352 34088 10364 34116
rect 8352 34076 8358 34088
rect 1394 34048 1400 34060
rect 1355 34020 1400 34048
rect 1394 34008 1400 34020
rect 1452 34008 1458 34060
rect 1581 34051 1639 34057
rect 1581 34017 1593 34051
rect 1627 34048 1639 34051
rect 2130 34048 2136 34060
rect 1627 34020 2136 34048
rect 1627 34017 1639 34020
rect 1581 34011 1639 34017
rect 2130 34008 2136 34020
rect 2188 34008 2194 34060
rect 2774 34008 2780 34060
rect 2832 34048 2838 34060
rect 9585 34051 9643 34057
rect 2832 34020 2877 34048
rect 2832 34008 2838 34020
rect 9585 34017 9597 34051
rect 9631 34048 9643 34051
rect 10226 34048 10232 34060
rect 9631 34020 10232 34048
rect 9631 34017 9643 34020
rect 9585 34011 9643 34017
rect 10226 34008 10232 34020
rect 10284 34008 10290 34060
rect 10336 34057 10364 34088
rect 10321 34051 10379 34057
rect 10321 34017 10333 34051
rect 10367 34017 10379 34051
rect 10321 34011 10379 34017
rect 9214 33940 9220 33992
rect 9272 33980 9278 33992
rect 9493 33983 9551 33989
rect 9493 33980 9505 33983
rect 9272 33952 9505 33980
rect 9272 33940 9278 33952
rect 9493 33949 9505 33952
rect 9539 33980 9551 33983
rect 9539 33952 10732 33980
rect 9539 33949 9551 33952
rect 9493 33943 9551 33949
rect 10318 33872 10324 33924
rect 10376 33912 10382 33924
rect 10566 33915 10624 33921
rect 10566 33912 10578 33915
rect 10376 33884 10578 33912
rect 10376 33872 10382 33884
rect 10566 33881 10578 33884
rect 10612 33881 10624 33915
rect 10704 33912 10732 33952
rect 10870 33940 10876 33992
rect 10928 33980 10934 33992
rect 12406 33980 12434 34156
rect 14093 34153 14105 34156
rect 14139 34153 14151 34187
rect 14093 34147 14151 34153
rect 14553 34187 14611 34193
rect 14553 34153 14565 34187
rect 14599 34184 14611 34187
rect 14642 34184 14648 34196
rect 14599 34156 14648 34184
rect 14599 34153 14611 34156
rect 14553 34147 14611 34153
rect 14642 34144 14648 34156
rect 14700 34144 14706 34196
rect 21266 34184 21272 34196
rect 17052 34156 21272 34184
rect 17052 34116 17080 34156
rect 21266 34144 21272 34156
rect 21324 34184 21330 34196
rect 21818 34184 21824 34196
rect 21324 34156 21824 34184
rect 21324 34144 21330 34156
rect 21818 34144 21824 34156
rect 21876 34144 21882 34196
rect 22002 34144 22008 34196
rect 22060 34184 22066 34196
rect 23474 34184 23480 34196
rect 22060 34156 23480 34184
rect 22060 34144 22066 34156
rect 23474 34144 23480 34156
rect 23532 34184 23538 34196
rect 24578 34184 24584 34196
rect 23532 34156 24584 34184
rect 23532 34144 23538 34156
rect 24578 34144 24584 34156
rect 24636 34144 24642 34196
rect 24765 34187 24823 34193
rect 24765 34153 24777 34187
rect 24811 34184 24823 34187
rect 24854 34184 24860 34196
rect 24811 34156 24860 34184
rect 24811 34153 24823 34156
rect 24765 34147 24823 34153
rect 24854 34144 24860 34156
rect 24912 34144 24918 34196
rect 25038 34184 25044 34196
rect 24999 34156 25044 34184
rect 25038 34144 25044 34156
rect 25096 34144 25102 34196
rect 26602 34184 26608 34196
rect 26563 34156 26608 34184
rect 26602 34144 26608 34156
rect 26660 34144 26666 34196
rect 26896 34156 28994 34184
rect 12728 34088 17080 34116
rect 12728 34057 12756 34088
rect 23842 34076 23848 34128
rect 23900 34116 23906 34128
rect 26896 34116 26924 34156
rect 27062 34116 27068 34128
rect 23900 34088 26924 34116
rect 27023 34088 27068 34116
rect 23900 34076 23906 34088
rect 27062 34076 27068 34088
rect 27120 34076 27126 34128
rect 28966 34116 28994 34156
rect 46750 34116 46756 34128
rect 28966 34088 31754 34116
rect 12713 34051 12771 34057
rect 12713 34017 12725 34051
rect 12759 34017 12771 34051
rect 12986 34048 12992 34060
rect 12947 34020 12992 34048
rect 12713 34011 12771 34017
rect 12986 34008 12992 34020
rect 13044 34008 13050 34060
rect 14182 34048 14188 34060
rect 14143 34020 14188 34048
rect 14182 34008 14188 34020
rect 14240 34008 14246 34060
rect 15102 34048 15108 34060
rect 14292 34020 15108 34048
rect 10928 33952 12434 33980
rect 10928 33940 10934 33952
rect 13814 33940 13820 33992
rect 13872 33980 13878 33992
rect 14093 33983 14151 33989
rect 14093 33980 14105 33983
rect 13872 33952 14105 33980
rect 13872 33940 13878 33952
rect 14093 33949 14105 33952
rect 14139 33980 14151 33983
rect 14292 33980 14320 34020
rect 15102 34008 15108 34020
rect 15160 34048 15166 34060
rect 15473 34051 15531 34057
rect 15473 34048 15485 34051
rect 15160 34020 15485 34048
rect 15160 34008 15166 34020
rect 15473 34017 15485 34020
rect 15519 34017 15531 34051
rect 15473 34011 15531 34017
rect 16022 34008 16028 34060
rect 16080 34048 16086 34060
rect 17037 34051 17095 34057
rect 17037 34048 17049 34051
rect 16080 34020 17049 34048
rect 16080 34008 16086 34020
rect 17037 34017 17049 34020
rect 17083 34017 17095 34051
rect 17310 34048 17316 34060
rect 17271 34020 17316 34048
rect 17037 34011 17095 34017
rect 17310 34008 17316 34020
rect 17368 34008 17374 34060
rect 19429 34051 19487 34057
rect 19429 34017 19441 34051
rect 19475 34048 19487 34051
rect 20346 34048 20352 34060
rect 19475 34020 20352 34048
rect 19475 34017 19487 34020
rect 19429 34011 19487 34017
rect 20346 34008 20352 34020
rect 20404 34008 20410 34060
rect 25961 34051 26019 34057
rect 25961 34017 25973 34051
rect 26007 34048 26019 34051
rect 26050 34048 26056 34060
rect 26007 34020 26056 34048
rect 26007 34017 26019 34020
rect 25961 34011 26019 34017
rect 26050 34008 26056 34020
rect 26108 34008 26114 34060
rect 26789 34051 26847 34057
rect 26789 34017 26801 34051
rect 26835 34048 26847 34051
rect 27430 34048 27436 34060
rect 26835 34020 27436 34048
rect 26835 34017 26847 34020
rect 26789 34011 26847 34017
rect 27430 34008 27436 34020
rect 27488 34008 27494 34060
rect 28442 34048 28448 34060
rect 28403 34020 28448 34048
rect 28442 34008 28448 34020
rect 28500 34048 28506 34060
rect 28994 34048 29000 34060
rect 28500 34020 29000 34048
rect 28500 34008 28506 34020
rect 28994 34008 29000 34020
rect 29052 34048 29058 34060
rect 30193 34051 30251 34057
rect 30193 34048 30205 34051
rect 29052 34020 30205 34048
rect 29052 34008 29058 34020
rect 30193 34017 30205 34020
rect 30239 34048 30251 34051
rect 30282 34048 30288 34060
rect 30239 34020 30288 34048
rect 30239 34017 30251 34020
rect 30193 34011 30251 34017
rect 30282 34008 30288 34020
rect 30340 34008 30346 34060
rect 31726 34048 31754 34088
rect 46308 34088 46756 34116
rect 35805 34051 35863 34057
rect 35805 34048 35817 34051
rect 31726 34020 35817 34048
rect 35805 34017 35817 34020
rect 35851 34017 35863 34051
rect 37642 34048 37648 34060
rect 37603 34020 37648 34048
rect 35805 34011 35863 34017
rect 37642 34008 37648 34020
rect 37700 34008 37706 34060
rect 46308 34057 46336 34088
rect 46750 34076 46756 34088
rect 46808 34076 46814 34128
rect 46293 34051 46351 34057
rect 46293 34017 46305 34051
rect 46339 34017 46351 34051
rect 46293 34011 46351 34017
rect 46477 34051 46535 34057
rect 46477 34017 46489 34051
rect 46523 34048 46535 34051
rect 46934 34048 46940 34060
rect 46523 34020 46940 34048
rect 46523 34017 46535 34020
rect 46477 34011 46535 34017
rect 46934 34008 46940 34020
rect 46992 34008 46998 34060
rect 48133 34051 48191 34057
rect 48133 34017 48145 34051
rect 48179 34048 48191 34051
rect 48222 34048 48228 34060
rect 48179 34020 48228 34048
rect 48179 34017 48191 34020
rect 48133 34011 48191 34017
rect 48222 34008 48228 34020
rect 48280 34008 48286 34060
rect 14139 33952 14320 33980
rect 14369 33983 14427 33989
rect 14139 33949 14151 33952
rect 14093 33943 14151 33949
rect 14369 33949 14381 33983
rect 14415 33949 14427 33983
rect 14369 33943 14427 33949
rect 15197 33983 15255 33989
rect 15197 33949 15209 33983
rect 15243 33980 15255 33983
rect 15378 33980 15384 33992
rect 15243 33952 15384 33980
rect 15243 33949 15255 33952
rect 15197 33943 15255 33949
rect 10704 33884 11744 33912
rect 10566 33875 10624 33881
rect 9861 33847 9919 33853
rect 9861 33813 9873 33847
rect 9907 33844 9919 33847
rect 10778 33844 10784 33856
rect 9907 33816 10784 33844
rect 9907 33813 9919 33816
rect 9861 33807 9919 33813
rect 10778 33804 10784 33816
rect 10836 33804 10842 33856
rect 11716 33853 11744 33884
rect 11701 33847 11759 33853
rect 11701 33813 11713 33847
rect 11747 33844 11759 33847
rect 14384 33844 14412 33943
rect 15378 33940 15384 33952
rect 15436 33940 15442 33992
rect 19702 33980 19708 33992
rect 19615 33952 19708 33980
rect 19702 33940 19708 33952
rect 19760 33980 19766 33992
rect 20622 33980 20628 33992
rect 19760 33952 20628 33980
rect 19760 33940 19766 33952
rect 20622 33940 20628 33952
rect 20680 33940 20686 33992
rect 22741 33983 22799 33989
rect 22741 33949 22753 33983
rect 22787 33980 22799 33983
rect 23014 33980 23020 33992
rect 22787 33952 23020 33980
rect 22787 33949 22799 33952
rect 22741 33943 22799 33949
rect 23014 33940 23020 33952
rect 23072 33940 23078 33992
rect 24762 33980 24768 33992
rect 24723 33952 24768 33980
rect 24762 33940 24768 33952
rect 24820 33940 24826 33992
rect 24857 33983 24915 33989
rect 24857 33949 24869 33983
rect 24903 33980 24915 33983
rect 25038 33980 25044 33992
rect 24903 33952 25044 33980
rect 24903 33949 24915 33952
rect 24857 33943 24915 33949
rect 25038 33940 25044 33952
rect 25096 33940 25102 33992
rect 25498 33980 25504 33992
rect 25459 33952 25504 33980
rect 25498 33940 25504 33952
rect 25556 33940 25562 33992
rect 25866 33980 25872 33992
rect 25827 33952 25872 33980
rect 25866 33940 25872 33952
rect 25924 33940 25930 33992
rect 26418 33940 26424 33992
rect 26476 33980 26482 33992
rect 26605 33983 26663 33989
rect 26605 33980 26617 33983
rect 26476 33952 26617 33980
rect 26476 33940 26482 33952
rect 26605 33949 26617 33952
rect 26651 33949 26663 33983
rect 26605 33943 26663 33949
rect 26878 33940 26884 33992
rect 26936 33980 26942 33992
rect 28261 33983 28319 33989
rect 26936 33952 26981 33980
rect 26936 33940 26942 33952
rect 28261 33949 28273 33983
rect 28307 33980 28319 33983
rect 29822 33980 29828 33992
rect 28307 33952 29828 33980
rect 28307 33949 28319 33952
rect 28261 33943 28319 33949
rect 29822 33940 29828 33952
rect 29880 33940 29886 33992
rect 30742 33980 30748 33992
rect 30703 33952 30748 33980
rect 30742 33940 30748 33952
rect 30800 33940 30806 33992
rect 22922 33912 22928 33924
rect 22883 33884 22928 33912
rect 22922 33872 22928 33884
rect 22980 33872 22986 33924
rect 24581 33915 24639 33921
rect 24581 33881 24593 33915
rect 24627 33912 24639 33915
rect 25774 33912 25780 33924
rect 24627 33884 25780 33912
rect 24627 33881 24639 33884
rect 24581 33875 24639 33881
rect 25774 33872 25780 33884
rect 25832 33872 25838 33924
rect 28350 33912 28356 33924
rect 28311 33884 28356 33912
rect 28350 33872 28356 33884
rect 28408 33872 28414 33924
rect 30006 33872 30012 33924
rect 30064 33912 30070 33924
rect 35986 33912 35992 33924
rect 30064 33884 30109 33912
rect 35947 33884 35992 33912
rect 30064 33872 30070 33884
rect 35986 33872 35992 33884
rect 36044 33872 36050 33924
rect 18598 33844 18604 33856
rect 11747 33816 14412 33844
rect 18559 33816 18604 33844
rect 11747 33813 11759 33816
rect 11701 33807 11759 33813
rect 18598 33804 18604 33816
rect 18656 33804 18662 33856
rect 22462 33804 22468 33856
rect 22520 33844 22526 33856
rect 23109 33847 23167 33853
rect 23109 33844 23121 33847
rect 22520 33816 23121 33844
rect 22520 33804 22526 33816
rect 23109 33813 23121 33816
rect 23155 33813 23167 33847
rect 25590 33844 25596 33856
rect 25551 33816 25596 33844
rect 23109 33807 23167 33813
rect 25590 33804 25596 33816
rect 25648 33804 25654 33856
rect 27522 33804 27528 33856
rect 27580 33844 27586 33856
rect 27893 33847 27951 33853
rect 27893 33844 27905 33847
rect 27580 33816 27905 33844
rect 27580 33804 27586 33816
rect 27893 33813 27905 33816
rect 27939 33813 27951 33847
rect 27893 33807 27951 33813
rect 30558 33804 30564 33856
rect 30616 33844 30622 33856
rect 30837 33847 30895 33853
rect 30837 33844 30849 33847
rect 30616 33816 30849 33844
rect 30616 33804 30622 33816
rect 30837 33813 30849 33816
rect 30883 33813 30895 33847
rect 30837 33807 30895 33813
rect 1104 33754 48852 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 48852 33754
rect 1104 33680 48852 33702
rect 10318 33640 10324 33652
rect 10279 33612 10324 33640
rect 10318 33600 10324 33612
rect 10376 33600 10382 33652
rect 11977 33643 12035 33649
rect 11977 33640 11989 33643
rect 10612 33612 11989 33640
rect 10226 33532 10232 33584
rect 10284 33572 10290 33584
rect 10612 33572 10640 33612
rect 11977 33609 11989 33612
rect 12023 33609 12035 33643
rect 12802 33640 12808 33652
rect 11977 33603 12035 33609
rect 12084 33612 12808 33640
rect 10284 33544 10640 33572
rect 10284 33532 10290 33544
rect 11238 33532 11244 33584
rect 11296 33572 11302 33584
rect 11885 33575 11943 33581
rect 11885 33572 11897 33575
rect 11296 33544 11897 33572
rect 11296 33532 11302 33544
rect 11885 33541 11897 33544
rect 11931 33541 11943 33575
rect 11885 33535 11943 33541
rect 1854 33504 1860 33516
rect 1815 33476 1860 33504
rect 1854 33464 1860 33476
rect 1912 33464 1918 33516
rect 8294 33464 8300 33516
rect 8352 33504 8358 33516
rect 8389 33507 8447 33513
rect 8389 33504 8401 33507
rect 8352 33476 8401 33504
rect 8352 33464 8358 33476
rect 8389 33473 8401 33476
rect 8435 33473 8447 33507
rect 8389 33467 8447 33473
rect 8656 33507 8714 33513
rect 8656 33473 8668 33507
rect 8702 33504 8714 33507
rect 8702 33476 9674 33504
rect 8702 33473 8714 33476
rect 8656 33467 8714 33473
rect 2041 33439 2099 33445
rect 2041 33405 2053 33439
rect 2087 33405 2099 33439
rect 2041 33399 2099 33405
rect 2056 33300 2084 33399
rect 2774 33396 2780 33448
rect 2832 33436 2838 33448
rect 2832 33408 2877 33436
rect 2832 33396 2838 33408
rect 9646 33368 9674 33476
rect 10502 33464 10508 33516
rect 10560 33513 10566 33516
rect 10560 33507 10609 33513
rect 10560 33473 10563 33507
rect 10597 33473 10609 33507
rect 10686 33504 10692 33516
rect 10647 33476 10692 33504
rect 10560 33467 10609 33473
rect 10560 33464 10566 33467
rect 10686 33464 10692 33476
rect 10744 33464 10750 33516
rect 10778 33464 10784 33516
rect 10836 33513 10842 33516
rect 10836 33504 10844 33513
rect 10962 33504 10968 33516
rect 10836 33476 10881 33504
rect 10923 33476 10968 33504
rect 10836 33467 10844 33476
rect 10836 33464 10842 33467
rect 10962 33464 10968 33476
rect 11020 33464 11026 33516
rect 11793 33507 11851 33513
rect 11793 33473 11805 33507
rect 11839 33504 11851 33507
rect 11974 33504 11980 33516
rect 11839 33476 11980 33504
rect 11839 33473 11851 33476
rect 11793 33467 11851 33473
rect 11974 33464 11980 33476
rect 12032 33464 12038 33516
rect 12084 33436 12112 33612
rect 12802 33600 12808 33612
rect 12860 33600 12866 33652
rect 12894 33600 12900 33652
rect 12952 33640 12958 33652
rect 12989 33643 13047 33649
rect 12989 33640 13001 33643
rect 12952 33612 13001 33640
rect 12952 33600 12958 33612
rect 12989 33609 13001 33612
rect 13035 33609 13047 33643
rect 12989 33603 13047 33609
rect 17218 33600 17224 33652
rect 17276 33640 17282 33652
rect 17497 33643 17555 33649
rect 17497 33640 17509 33643
rect 17276 33612 17509 33640
rect 17276 33600 17282 33612
rect 17497 33609 17509 33612
rect 17543 33609 17555 33643
rect 17497 33603 17555 33609
rect 26602 33600 26608 33652
rect 26660 33640 26666 33652
rect 27246 33640 27252 33652
rect 26660 33612 27252 33640
rect 26660 33600 26666 33612
rect 27246 33600 27252 33612
rect 27304 33640 27310 33652
rect 27798 33640 27804 33652
rect 27304 33612 27804 33640
rect 27304 33600 27310 33612
rect 27798 33600 27804 33612
rect 27856 33600 27862 33652
rect 29733 33643 29791 33649
rect 29733 33609 29745 33643
rect 29779 33640 29791 33643
rect 29822 33640 29828 33652
rect 29779 33612 29828 33640
rect 29779 33609 29791 33612
rect 29733 33603 29791 33609
rect 29822 33600 29828 33612
rect 29880 33600 29886 33652
rect 30098 33600 30104 33652
rect 30156 33640 30162 33652
rect 32950 33640 32956 33652
rect 30156 33612 32956 33640
rect 30156 33600 30162 33612
rect 32950 33600 32956 33612
rect 33008 33640 33014 33652
rect 33873 33643 33931 33649
rect 33873 33640 33885 33643
rect 33008 33612 33885 33640
rect 33008 33600 33014 33612
rect 33873 33609 33885 33612
rect 33919 33609 33931 33643
rect 33873 33603 33931 33609
rect 35897 33643 35955 33649
rect 35897 33609 35909 33643
rect 35943 33640 35955 33643
rect 35986 33640 35992 33652
rect 35943 33612 35992 33640
rect 35943 33609 35955 33612
rect 35897 33603 35955 33609
rect 35986 33600 35992 33612
rect 36044 33600 36050 33652
rect 46382 33600 46388 33652
rect 46440 33640 46446 33652
rect 46937 33643 46995 33649
rect 46937 33640 46949 33643
rect 46440 33612 46949 33640
rect 46440 33600 46446 33612
rect 46937 33609 46949 33612
rect 46983 33609 46995 33643
rect 46937 33603 46995 33609
rect 12158 33532 12164 33584
rect 12216 33572 12222 33584
rect 16022 33572 16028 33584
rect 12216 33544 16028 33572
rect 12216 33532 12222 33544
rect 12342 33464 12348 33516
rect 12400 33504 12406 33516
rect 12713 33507 12771 33513
rect 12713 33504 12725 33507
rect 12400 33476 12725 33504
rect 12400 33464 12406 33476
rect 12713 33473 12725 33476
rect 12759 33473 12771 33507
rect 12713 33467 12771 33473
rect 13078 33464 13084 33516
rect 13136 33504 13142 33516
rect 14292 33513 14320 33544
rect 16022 33532 16028 33544
rect 16080 33532 16086 33584
rect 18966 33572 18972 33584
rect 18927 33544 18972 33572
rect 18966 33532 18972 33544
rect 19024 33532 19030 33584
rect 22186 33572 22192 33584
rect 22099 33544 22192 33572
rect 22186 33532 22192 33544
rect 22244 33572 22250 33584
rect 26237 33575 26295 33581
rect 22244 33544 23980 33572
rect 22244 33532 22250 33544
rect 14550 33513 14556 33516
rect 13633 33507 13691 33513
rect 13633 33504 13645 33507
rect 13136 33476 13645 33504
rect 13136 33464 13142 33476
rect 13633 33473 13645 33476
rect 13679 33473 13691 33507
rect 13633 33467 13691 33473
rect 14277 33507 14335 33513
rect 14277 33473 14289 33507
rect 14323 33473 14335 33507
rect 14277 33467 14335 33473
rect 14544 33467 14556 33513
rect 14608 33504 14614 33516
rect 14608 33476 14644 33504
rect 14550 33464 14556 33467
rect 14608 33464 14614 33476
rect 16758 33464 16764 33516
rect 16816 33504 16822 33516
rect 17129 33507 17187 33513
rect 17129 33504 17141 33507
rect 16816 33476 17141 33504
rect 16816 33464 16822 33476
rect 17129 33473 17141 33476
rect 17175 33473 17187 33507
rect 17129 33467 17187 33473
rect 17313 33507 17371 33513
rect 17313 33473 17325 33507
rect 17359 33504 17371 33507
rect 18598 33504 18604 33516
rect 17359 33476 18604 33504
rect 17359 33473 17371 33476
rect 17313 33467 17371 33473
rect 18598 33464 18604 33476
rect 18656 33464 18662 33516
rect 19153 33507 19211 33513
rect 19153 33473 19165 33507
rect 19199 33504 19211 33507
rect 19889 33507 19947 33513
rect 19889 33504 19901 33507
rect 19199 33476 19901 33504
rect 19199 33473 19211 33476
rect 19153 33467 19211 33473
rect 19889 33473 19901 33476
rect 19935 33504 19947 33507
rect 19978 33504 19984 33516
rect 19935 33476 19984 33504
rect 19935 33473 19947 33476
rect 19889 33467 19947 33473
rect 19978 33464 19984 33476
rect 20036 33464 20042 33516
rect 20156 33507 20214 33513
rect 20156 33473 20168 33507
rect 20202 33504 20214 33507
rect 20438 33504 20444 33516
rect 20202 33476 20444 33504
rect 20202 33473 20214 33476
rect 20156 33467 20214 33473
rect 20438 33464 20444 33476
rect 20496 33464 20502 33516
rect 21634 33464 21640 33516
rect 21692 33504 21698 33516
rect 22005 33507 22063 33513
rect 22005 33504 22017 33507
rect 21692 33476 22017 33504
rect 21692 33464 21698 33476
rect 22005 33473 22017 33476
rect 22051 33473 22063 33507
rect 22005 33467 22063 33473
rect 22281 33507 22339 33513
rect 22281 33473 22293 33507
rect 22327 33473 22339 33507
rect 22281 33467 22339 33473
rect 12161 33439 12219 33445
rect 12161 33436 12173 33439
rect 12084 33408 12173 33436
rect 12161 33405 12173 33408
rect 12207 33405 12219 33439
rect 12161 33399 12219 33405
rect 12250 33396 12256 33448
rect 12308 33436 12314 33448
rect 12986 33436 12992 33448
rect 12308 33408 12353 33436
rect 12947 33408 12992 33436
rect 12308 33396 12314 33408
rect 12986 33396 12992 33408
rect 13044 33396 13050 33448
rect 13449 33439 13507 33445
rect 13449 33405 13461 33439
rect 13495 33436 13507 33439
rect 13814 33436 13820 33448
rect 13495 33408 13820 33436
rect 13495 33405 13507 33408
rect 13449 33399 13507 33405
rect 13814 33396 13820 33408
rect 13872 33396 13878 33448
rect 22296 33436 22324 33467
rect 22646 33464 22652 33516
rect 22704 33504 22710 33516
rect 23661 33507 23719 33513
rect 23661 33504 23673 33507
rect 22704 33476 23673 33504
rect 22704 33464 22710 33476
rect 23661 33473 23673 33476
rect 23707 33473 23719 33507
rect 23952 33504 23980 33544
rect 26237 33541 26249 33575
rect 26283 33572 26295 33575
rect 26326 33572 26332 33584
rect 26283 33544 26332 33572
rect 26283 33541 26295 33544
rect 26237 33535 26295 33541
rect 26326 33532 26332 33544
rect 26384 33572 26390 33584
rect 26878 33572 26884 33584
rect 26384 33544 26884 33572
rect 26384 33532 26390 33544
rect 26878 33532 26884 33544
rect 26936 33532 26942 33584
rect 27522 33572 27528 33584
rect 27483 33544 27528 33572
rect 27522 33532 27528 33544
rect 27580 33532 27586 33584
rect 30558 33572 30564 33584
rect 28368 33544 30564 33572
rect 28368 33513 28396 33544
rect 30558 33532 30564 33544
rect 30616 33572 30622 33584
rect 30616 33544 32536 33572
rect 30616 33532 30622 33544
rect 27709 33507 27767 33513
rect 23952 33476 26464 33504
rect 23661 33467 23719 33473
rect 24210 33436 24216 33448
rect 21284 33408 24216 33436
rect 21284 33377 21312 33408
rect 24210 33396 24216 33408
rect 24268 33396 24274 33448
rect 11517 33371 11575 33377
rect 11517 33368 11529 33371
rect 9646 33340 11529 33368
rect 11517 33337 11529 33340
rect 11563 33337 11575 33371
rect 11517 33331 11575 33337
rect 21269 33371 21327 33377
rect 21269 33337 21281 33371
rect 21315 33337 21327 33371
rect 23842 33368 23848 33380
rect 23755 33340 23848 33368
rect 21269 33331 21327 33337
rect 23842 33328 23848 33340
rect 23900 33368 23906 33380
rect 26050 33368 26056 33380
rect 23900 33340 26056 33368
rect 23900 33328 23906 33340
rect 26050 33328 26056 33340
rect 26108 33328 26114 33380
rect 26436 33377 26464 33476
rect 27709 33473 27721 33507
rect 27755 33473 27767 33507
rect 27709 33467 27767 33473
rect 28353 33507 28411 33513
rect 28353 33473 28365 33507
rect 28399 33473 28411 33507
rect 28353 33467 28411 33473
rect 27338 33396 27344 33448
rect 27396 33436 27402 33448
rect 27522 33436 27528 33448
rect 27396 33408 27528 33436
rect 27396 33396 27402 33408
rect 27522 33396 27528 33408
rect 27580 33436 27586 33448
rect 27724 33436 27752 33467
rect 28442 33464 28448 33516
rect 28500 33504 28506 33516
rect 28609 33507 28667 33513
rect 28609 33504 28621 33507
rect 28500 33476 28621 33504
rect 28500 33464 28506 33476
rect 28609 33473 28621 33476
rect 28655 33473 28667 33507
rect 30650 33504 30656 33516
rect 30611 33476 30656 33504
rect 28609 33467 28667 33473
rect 30650 33464 30656 33476
rect 30708 33464 30714 33516
rect 30745 33507 30803 33513
rect 30745 33473 30757 33507
rect 30791 33473 30803 33507
rect 30745 33467 30803 33473
rect 27580 33408 27752 33436
rect 30760 33436 30788 33467
rect 30834 33464 30840 33516
rect 30892 33504 30898 33516
rect 30892 33476 30937 33504
rect 30892 33464 30898 33476
rect 31018 33464 31024 33516
rect 31076 33504 31082 33516
rect 31076 33476 31121 33504
rect 31076 33464 31082 33476
rect 32508 33448 32536 33544
rect 32760 33507 32818 33513
rect 32760 33473 32772 33507
rect 32806 33504 32818 33507
rect 33042 33504 33048 33516
rect 32806 33476 33048 33504
rect 32806 33473 32818 33476
rect 32760 33467 32818 33473
rect 33042 33464 33048 33476
rect 33100 33464 33106 33516
rect 35805 33507 35863 33513
rect 35805 33473 35817 33507
rect 35851 33504 35863 33507
rect 35894 33504 35900 33516
rect 35851 33476 35900 33504
rect 35851 33473 35863 33476
rect 35805 33467 35863 33473
rect 35894 33464 35900 33476
rect 35952 33464 35958 33516
rect 46658 33464 46664 33516
rect 46716 33504 46722 33516
rect 46845 33507 46903 33513
rect 46845 33504 46857 33507
rect 46716 33476 46857 33504
rect 46716 33464 46722 33476
rect 46845 33473 46857 33476
rect 46891 33473 46903 33507
rect 47946 33504 47952 33516
rect 47907 33476 47952 33504
rect 46845 33467 46903 33473
rect 47946 33464 47952 33476
rect 48004 33464 48010 33516
rect 32306 33436 32312 33448
rect 30760 33408 32312 33436
rect 27580 33396 27586 33408
rect 26421 33371 26479 33377
rect 26421 33337 26433 33371
rect 26467 33368 26479 33371
rect 26602 33368 26608 33380
rect 26467 33340 26608 33368
rect 26467 33337 26479 33340
rect 26421 33331 26479 33337
rect 26602 33328 26608 33340
rect 26660 33328 26666 33380
rect 27893 33371 27951 33377
rect 27893 33337 27905 33371
rect 27939 33368 27951 33371
rect 28258 33368 28264 33380
rect 27939 33340 28264 33368
rect 27939 33337 27951 33340
rect 27893 33331 27951 33337
rect 28258 33328 28264 33340
rect 28316 33328 28322 33380
rect 30760 33368 30788 33408
rect 32306 33396 32312 33408
rect 32364 33396 32370 33448
rect 32490 33436 32496 33448
rect 32451 33408 32496 33436
rect 32490 33396 32496 33408
rect 32548 33396 32554 33448
rect 29288 33340 30788 33368
rect 2774 33300 2780 33312
rect 2056 33272 2780 33300
rect 2774 33260 2780 33272
rect 2832 33260 2838 33312
rect 9766 33300 9772 33312
rect 9679 33272 9772 33300
rect 9766 33260 9772 33272
rect 9824 33300 9830 33312
rect 10870 33300 10876 33312
rect 9824 33272 10876 33300
rect 9824 33260 9830 33272
rect 10870 33260 10876 33272
rect 10928 33260 10934 33312
rect 12802 33300 12808 33312
rect 12715 33272 12808 33300
rect 12802 33260 12808 33272
rect 12860 33300 12866 33312
rect 13630 33300 13636 33312
rect 12860 33272 13636 33300
rect 12860 33260 12866 33272
rect 13630 33260 13636 33272
rect 13688 33260 13694 33312
rect 13817 33303 13875 33309
rect 13817 33269 13829 33303
rect 13863 33300 13875 33303
rect 14274 33300 14280 33312
rect 13863 33272 14280 33300
rect 13863 33269 13875 33272
rect 13817 33263 13875 33269
rect 14274 33260 14280 33272
rect 14332 33260 14338 33312
rect 15378 33260 15384 33312
rect 15436 33300 15442 33312
rect 15657 33303 15715 33309
rect 15657 33300 15669 33303
rect 15436 33272 15669 33300
rect 15436 33260 15442 33272
rect 15657 33269 15669 33272
rect 15703 33269 15715 33303
rect 15657 33263 15715 33269
rect 18874 33260 18880 33312
rect 18932 33300 18938 33312
rect 19058 33300 19064 33312
rect 18932 33272 19064 33300
rect 18932 33260 18938 33272
rect 19058 33260 19064 33272
rect 19116 33260 19122 33312
rect 20990 33260 20996 33312
rect 21048 33300 21054 33312
rect 21821 33303 21879 33309
rect 21821 33300 21833 33303
rect 21048 33272 21833 33300
rect 21048 33260 21054 33272
rect 21821 33269 21833 33272
rect 21867 33269 21879 33303
rect 21821 33263 21879 33269
rect 26234 33260 26240 33312
rect 26292 33300 26298 33312
rect 26510 33300 26516 33312
rect 26292 33272 26516 33300
rect 26292 33260 26298 33272
rect 26510 33260 26516 33272
rect 26568 33260 26574 33312
rect 28166 33260 28172 33312
rect 28224 33300 28230 33312
rect 29288 33300 29316 33340
rect 30374 33300 30380 33312
rect 28224 33272 29316 33300
rect 30335 33272 30380 33300
rect 28224 33260 28230 33272
rect 30374 33260 30380 33272
rect 30432 33260 30438 33312
rect 46934 33260 46940 33312
rect 46992 33300 46998 33312
rect 48041 33303 48099 33309
rect 48041 33300 48053 33303
rect 46992 33272 48053 33300
rect 46992 33260 46998 33272
rect 48041 33269 48053 33272
rect 48087 33269 48099 33303
rect 48041 33263 48099 33269
rect 1104 33210 48852 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 48852 33210
rect 1104 33136 48852 33158
rect 2774 33056 2780 33108
rect 2832 33096 2838 33108
rect 2832 33068 2877 33096
rect 2832 33056 2838 33068
rect 10226 33056 10232 33108
rect 10284 33096 10290 33108
rect 10321 33099 10379 33105
rect 10321 33096 10333 33099
rect 10284 33068 10333 33096
rect 10284 33056 10290 33068
rect 10321 33065 10333 33068
rect 10367 33065 10379 33099
rect 11238 33096 11244 33108
rect 11199 33068 11244 33096
rect 10321 33059 10379 33065
rect 11238 33056 11244 33068
rect 11296 33056 11302 33108
rect 12158 33056 12164 33108
rect 12216 33096 12222 33108
rect 12526 33096 12532 33108
rect 12216 33068 12532 33096
rect 12216 33056 12222 33068
rect 12526 33056 12532 33068
rect 12584 33096 12590 33108
rect 13449 33099 13507 33105
rect 13449 33096 13461 33099
rect 12584 33068 13461 33096
rect 12584 33056 12590 33068
rect 13449 33065 13461 33068
rect 13495 33065 13507 33099
rect 20438 33096 20444 33108
rect 20399 33068 20444 33096
rect 13449 33059 13507 33065
rect 20438 33056 20444 33068
rect 20496 33056 20502 33108
rect 27801 33099 27859 33105
rect 20548 33068 22140 33096
rect 12342 32988 12348 33040
rect 12400 33028 12406 33040
rect 13722 33028 13728 33040
rect 12400 33000 13728 33028
rect 12400 32988 12406 33000
rect 13722 32988 13728 33000
rect 13780 32988 13786 33040
rect 19978 32988 19984 33040
rect 20036 33028 20042 33040
rect 20548 33028 20576 33068
rect 20036 33000 20576 33028
rect 20036 32988 20042 33000
rect 20622 32988 20628 33040
rect 20680 33028 20686 33040
rect 20680 33000 21128 33028
rect 20680 32988 20686 33000
rect 11054 32960 11060 32972
rect 10244 32932 11060 32960
rect 2038 32852 2044 32904
rect 2096 32892 2102 32904
rect 2225 32895 2283 32901
rect 2225 32892 2237 32895
rect 2096 32864 2237 32892
rect 2096 32852 2102 32864
rect 2225 32861 2237 32864
rect 2271 32861 2283 32895
rect 2682 32892 2688 32904
rect 2643 32864 2688 32892
rect 2225 32855 2283 32861
rect 2682 32852 2688 32864
rect 2740 32852 2746 32904
rect 10244 32901 10272 32932
rect 11054 32920 11060 32932
rect 11112 32920 11118 32972
rect 12253 32963 12311 32969
rect 12253 32929 12265 32963
rect 12299 32960 12311 32963
rect 12434 32960 12440 32972
rect 12299 32932 12440 32960
rect 12299 32929 12311 32932
rect 12253 32923 12311 32929
rect 12434 32920 12440 32932
rect 12492 32920 12498 32972
rect 20990 32960 20996 32972
rect 20916 32932 20996 32960
rect 10229 32895 10287 32901
rect 10229 32861 10241 32895
rect 10275 32861 10287 32895
rect 10229 32855 10287 32861
rect 10413 32895 10471 32901
rect 10413 32861 10425 32895
rect 10459 32892 10471 32895
rect 10873 32895 10931 32901
rect 10459 32864 10824 32892
rect 10459 32861 10471 32864
rect 10413 32855 10471 32861
rect 10796 32836 10824 32864
rect 10873 32861 10885 32895
rect 10919 32892 10931 32895
rect 11072 32892 11100 32920
rect 10919 32864 11100 32892
rect 11977 32895 12035 32901
rect 10919 32861 10931 32864
rect 10873 32855 10931 32861
rect 11977 32861 11989 32895
rect 12023 32892 12035 32895
rect 13170 32892 13176 32904
rect 12023 32864 13176 32892
rect 12023 32861 12035 32864
rect 11977 32855 12035 32861
rect 12268 32836 12296 32864
rect 13170 32852 13176 32864
rect 13228 32852 13234 32904
rect 13538 32852 13544 32904
rect 13596 32892 13602 32904
rect 14182 32892 14188 32904
rect 13596 32864 14188 32892
rect 13596 32852 13602 32864
rect 14182 32852 14188 32864
rect 14240 32892 14246 32904
rect 14461 32895 14519 32901
rect 14461 32892 14473 32895
rect 14240 32864 14473 32892
rect 14240 32852 14246 32864
rect 14461 32861 14473 32864
rect 14507 32892 14519 32895
rect 14734 32892 14740 32904
rect 14507 32864 14740 32892
rect 14507 32861 14519 32864
rect 14461 32855 14519 32861
rect 14734 32852 14740 32864
rect 14792 32852 14798 32904
rect 14921 32895 14979 32901
rect 14921 32861 14933 32895
rect 14967 32892 14979 32895
rect 15378 32892 15384 32904
rect 14967 32864 15384 32892
rect 14967 32861 14979 32864
rect 14921 32855 14979 32861
rect 15378 32852 15384 32864
rect 15436 32852 15442 32904
rect 20803 32901 20809 32904
rect 18509 32895 18567 32901
rect 18509 32861 18521 32895
rect 18555 32892 18567 32895
rect 19245 32895 19303 32901
rect 19245 32892 19257 32895
rect 18555 32864 19257 32892
rect 18555 32861 18567 32864
rect 18509 32855 18567 32861
rect 19245 32861 19257 32864
rect 19291 32861 19303 32895
rect 19245 32855 19303 32861
rect 20697 32895 20755 32901
rect 20697 32861 20709 32895
rect 20743 32892 20755 32895
rect 20790 32895 20809 32901
rect 20743 32861 20760 32892
rect 20697 32855 20760 32861
rect 20790 32861 20802 32895
rect 20790 32855 20809 32861
rect 10778 32784 10784 32836
rect 10836 32824 10842 32836
rect 11057 32827 11115 32833
rect 11057 32824 11069 32827
rect 10836 32796 11069 32824
rect 10836 32784 10842 32796
rect 11057 32793 11069 32796
rect 11103 32793 11115 32827
rect 11057 32787 11115 32793
rect 12250 32784 12256 32836
rect 12308 32784 12314 32836
rect 13078 32784 13084 32836
rect 13136 32824 13142 32836
rect 13357 32827 13415 32833
rect 13357 32824 13369 32827
rect 13136 32796 13369 32824
rect 13136 32784 13142 32796
rect 13357 32793 13369 32796
rect 13403 32793 13415 32827
rect 18322 32824 18328 32836
rect 13357 32787 13415 32793
rect 13648 32796 18328 32824
rect 7650 32716 7656 32768
rect 7708 32756 7714 32768
rect 13648 32756 13676 32796
rect 18322 32784 18328 32796
rect 18380 32824 18386 32836
rect 18524 32824 18552 32855
rect 18380 32796 18552 32824
rect 18380 32784 18386 32796
rect 7708 32728 13676 32756
rect 7708 32716 7714 32728
rect 13722 32716 13728 32768
rect 13780 32756 13786 32768
rect 15289 32759 15347 32765
rect 15289 32756 15301 32759
rect 13780 32728 15301 32756
rect 13780 32716 13786 32728
rect 15289 32725 15301 32728
rect 15335 32725 15347 32759
rect 15289 32719 15347 32725
rect 18601 32759 18659 32765
rect 18601 32725 18613 32759
rect 18647 32756 18659 32759
rect 18874 32756 18880 32768
rect 18647 32728 18880 32756
rect 18647 32725 18659 32728
rect 18601 32719 18659 32725
rect 18874 32716 18880 32728
rect 18932 32716 18938 32768
rect 19337 32759 19395 32765
rect 19337 32725 19349 32759
rect 19383 32756 19395 32759
rect 19426 32756 19432 32768
rect 19383 32728 19432 32756
rect 19383 32725 19395 32728
rect 19337 32719 19395 32725
rect 19426 32716 19432 32728
rect 19484 32716 19490 32768
rect 20732 32756 20760 32855
rect 20803 32852 20809 32855
rect 20861 32852 20867 32904
rect 20916 32898 20944 32932
rect 20990 32920 20996 32932
rect 21048 32920 21054 32972
rect 21100 32901 21128 33000
rect 20901 32892 20959 32898
rect 20901 32858 20913 32892
rect 20947 32858 20959 32892
rect 20901 32852 20959 32858
rect 21085 32895 21143 32901
rect 21085 32861 21097 32895
rect 21131 32861 21143 32895
rect 21085 32855 21143 32861
rect 22002 32852 22008 32904
rect 22060 32892 22066 32904
rect 22112 32892 22140 33068
rect 27801 33065 27813 33099
rect 27847 33096 27859 33099
rect 28442 33096 28448 33108
rect 27847 33068 28448 33096
rect 27847 33065 27859 33068
rect 27801 33059 27859 33065
rect 28442 33056 28448 33068
rect 28500 33056 28506 33108
rect 30650 33056 30656 33108
rect 30708 33096 30714 33108
rect 30926 33096 30932 33108
rect 30708 33068 30932 33096
rect 30708 33056 30714 33068
rect 30926 33056 30932 33068
rect 30984 33056 30990 33108
rect 31018 33056 31024 33108
rect 31076 33096 31082 33108
rect 32398 33096 32404 33108
rect 31076 33068 32404 33096
rect 31076 33056 31082 33068
rect 32398 33056 32404 33068
rect 32456 33056 32462 33108
rect 33042 33096 33048 33108
rect 33003 33068 33048 33096
rect 33042 33056 33048 33068
rect 33100 33056 33106 33108
rect 47394 33056 47400 33108
rect 47452 33096 47458 33108
rect 47673 33099 47731 33105
rect 47673 33096 47685 33099
rect 47452 33068 47685 33096
rect 47452 33056 47458 33068
rect 47673 33065 47685 33068
rect 47719 33065 47731 33099
rect 47673 33059 47731 33065
rect 26237 33031 26295 33037
rect 26237 32997 26249 33031
rect 26283 33028 26295 33031
rect 27522 33028 27528 33040
rect 26283 33000 27528 33028
rect 26283 32997 26295 33000
rect 26237 32991 26295 32997
rect 27522 32988 27528 33000
rect 27580 32988 27586 33040
rect 28626 33028 28632 33040
rect 28460 33000 28632 33028
rect 27157 32963 27215 32969
rect 27157 32929 27169 32963
rect 27203 32960 27215 32963
rect 27203 32932 28212 32960
rect 27203 32929 27215 32932
rect 27157 32923 27215 32929
rect 28184 32904 28212 32932
rect 22189 32895 22247 32901
rect 22189 32892 22201 32895
rect 22060 32864 22201 32892
rect 22060 32852 22066 32864
rect 22189 32861 22201 32864
rect 22235 32861 22247 32895
rect 22189 32855 22247 32861
rect 26421 32895 26479 32901
rect 26421 32861 26433 32895
rect 26467 32892 26479 32895
rect 26786 32892 26792 32904
rect 26467 32864 26792 32892
rect 26467 32861 26479 32864
rect 26421 32855 26479 32861
rect 26786 32852 26792 32864
rect 26844 32852 26850 32904
rect 28031 32895 28089 32901
rect 28031 32892 28043 32895
rect 26896 32864 28043 32892
rect 22278 32784 22284 32836
rect 22336 32824 22342 32836
rect 22434 32827 22492 32833
rect 22434 32824 22446 32827
rect 22336 32796 22446 32824
rect 22336 32784 22342 32796
rect 22434 32793 22446 32796
rect 22480 32793 22492 32827
rect 26896 32824 26924 32864
rect 28031 32861 28043 32864
rect 28077 32861 28089 32895
rect 28166 32892 28172 32904
rect 28127 32864 28172 32892
rect 28031 32855 28089 32861
rect 28166 32852 28172 32864
rect 28224 32852 28230 32904
rect 28258 32852 28264 32904
rect 28316 32901 28322 32904
rect 28460 32901 28488 33000
rect 28626 32988 28632 33000
rect 28684 33028 28690 33040
rect 31036 33028 31064 33056
rect 28684 33000 31064 33028
rect 32416 33028 32444 33056
rect 32416 33000 33732 33028
rect 28684 32988 28690 33000
rect 30282 32960 30288 32972
rect 30243 32932 30288 32960
rect 30282 32920 30288 32932
rect 30340 32920 30346 32972
rect 30558 32920 30564 32972
rect 30616 32960 30622 32972
rect 31205 32963 31263 32969
rect 31205 32960 31217 32963
rect 30616 32932 31217 32960
rect 30616 32920 30622 32932
rect 31205 32929 31217 32932
rect 31251 32929 31263 32963
rect 31205 32923 31263 32929
rect 28316 32892 28324 32901
rect 28445 32895 28503 32901
rect 28316 32864 28361 32892
rect 28316 32855 28324 32864
rect 28445 32861 28457 32895
rect 28491 32861 28503 32895
rect 30098 32892 30104 32904
rect 30059 32864 30104 32892
rect 28445 32855 28503 32861
rect 28316 32852 28322 32855
rect 30098 32852 30104 32864
rect 30156 32852 30162 32904
rect 30190 32852 30196 32904
rect 30248 32852 30254 32904
rect 30374 32852 30380 32904
rect 30432 32892 30438 32904
rect 31461 32895 31519 32901
rect 31461 32892 31473 32895
rect 30432 32864 31473 32892
rect 30432 32852 30438 32864
rect 31461 32861 31473 32864
rect 31507 32861 31519 32895
rect 33318 32892 33324 32904
rect 33279 32864 33324 32892
rect 31461 32855 31519 32861
rect 33318 32852 33324 32864
rect 33376 32852 33382 32904
rect 33413 32895 33471 32901
rect 33413 32861 33425 32895
rect 33459 32861 33471 32895
rect 33413 32855 33471 32861
rect 22434 32787 22492 32793
rect 23446 32796 26924 32824
rect 26973 32827 27031 32833
rect 21726 32756 21732 32768
rect 20732 32728 21732 32756
rect 21726 32716 21732 32728
rect 21784 32716 21790 32768
rect 22094 32716 22100 32768
rect 22152 32756 22158 32768
rect 23446 32756 23474 32796
rect 26973 32793 26985 32827
rect 27019 32824 27031 32827
rect 27154 32824 27160 32836
rect 27019 32796 27160 32824
rect 27019 32793 27031 32796
rect 26973 32787 27031 32793
rect 27154 32784 27160 32796
rect 27212 32784 27218 32836
rect 30208 32824 30236 32852
rect 28966 32796 29868 32824
rect 30208 32796 30696 32824
rect 22152 32728 23474 32756
rect 22152 32716 22158 32728
rect 23566 32716 23572 32768
rect 23624 32756 23630 32768
rect 25038 32756 25044 32768
rect 23624 32728 25044 32756
rect 23624 32716 23630 32728
rect 25038 32716 25044 32728
rect 25096 32756 25102 32768
rect 28966 32756 28994 32796
rect 29730 32756 29736 32768
rect 25096 32728 28994 32756
rect 29691 32728 29736 32756
rect 25096 32716 25102 32728
rect 29730 32716 29736 32728
rect 29788 32716 29794 32768
rect 29840 32756 29868 32796
rect 30193 32759 30251 32765
rect 30193 32756 30205 32759
rect 29840 32728 30205 32756
rect 30193 32725 30205 32728
rect 30239 32725 30251 32759
rect 30668 32756 30696 32796
rect 32306 32784 32312 32836
rect 32364 32824 32370 32836
rect 33428 32824 33456 32855
rect 33502 32852 33508 32904
rect 33560 32892 33566 32904
rect 33704 32901 33732 33000
rect 33689 32895 33747 32901
rect 33560 32864 33605 32892
rect 33560 32852 33566 32864
rect 33689 32861 33701 32895
rect 33735 32861 33747 32895
rect 33689 32855 33747 32861
rect 32364 32796 33456 32824
rect 32364 32784 32370 32796
rect 32582 32756 32588 32768
rect 30668 32728 32588 32756
rect 30193 32719 30251 32725
rect 32582 32716 32588 32728
rect 32640 32716 32646 32768
rect 1104 32666 48852 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 48852 32666
rect 1104 32592 48852 32614
rect 12986 32512 12992 32564
rect 13044 32552 13050 32564
rect 13173 32555 13231 32561
rect 13173 32552 13185 32555
rect 13044 32524 13185 32552
rect 13044 32512 13050 32524
rect 13173 32521 13185 32524
rect 13219 32521 13231 32555
rect 13173 32515 13231 32521
rect 14461 32555 14519 32561
rect 14461 32521 14473 32555
rect 14507 32552 14519 32555
rect 14550 32552 14556 32564
rect 14507 32524 14556 32552
rect 14507 32521 14519 32524
rect 14461 32515 14519 32521
rect 14550 32512 14556 32524
rect 14608 32512 14614 32564
rect 17954 32512 17960 32564
rect 18012 32552 18018 32564
rect 18969 32555 19027 32561
rect 18969 32552 18981 32555
rect 18012 32524 18981 32552
rect 18012 32512 18018 32524
rect 18969 32521 18981 32524
rect 19015 32521 19027 32555
rect 18969 32515 19027 32521
rect 23385 32555 23443 32561
rect 23385 32521 23397 32555
rect 23431 32552 23443 32555
rect 23431 32524 24256 32552
rect 23431 32521 23443 32524
rect 23385 32515 23443 32521
rect 10686 32484 10692 32496
rect 10520 32456 10692 32484
rect 2038 32416 2044 32428
rect 1999 32388 2044 32416
rect 2038 32376 2044 32388
rect 2096 32376 2102 32428
rect 10318 32376 10324 32428
rect 10376 32425 10382 32428
rect 10520 32425 10548 32456
rect 10686 32444 10692 32456
rect 10744 32484 10750 32496
rect 12158 32484 12164 32496
rect 10744 32456 12164 32484
rect 10744 32444 10750 32456
rect 12158 32444 12164 32456
rect 12216 32444 12222 32496
rect 13538 32444 13544 32496
rect 13596 32444 13602 32496
rect 18877 32487 18935 32493
rect 13740 32456 18828 32484
rect 10376 32419 10425 32425
rect 10376 32385 10379 32419
rect 10413 32385 10425 32419
rect 10376 32379 10425 32385
rect 10505 32419 10563 32425
rect 10505 32385 10517 32419
rect 10551 32385 10563 32419
rect 10505 32379 10563 32385
rect 10376 32376 10382 32379
rect 10594 32376 10600 32428
rect 10652 32425 10658 32428
rect 10652 32416 10660 32425
rect 10781 32419 10839 32425
rect 10652 32388 10697 32416
rect 10652 32379 10660 32388
rect 10781 32385 10793 32419
rect 10827 32416 10839 32419
rect 10962 32416 10968 32428
rect 10827 32388 10968 32416
rect 10827 32385 10839 32388
rect 10781 32379 10839 32385
rect 10652 32376 10658 32379
rect 10962 32376 10968 32388
rect 11020 32376 11026 32428
rect 11790 32376 11796 32428
rect 11848 32416 11854 32428
rect 12069 32419 12127 32425
rect 12069 32416 12081 32419
rect 11848 32388 12081 32416
rect 11848 32376 11854 32388
rect 12069 32385 12081 32388
rect 12115 32385 12127 32419
rect 12250 32416 12256 32428
rect 12211 32388 12256 32416
rect 12069 32379 12127 32385
rect 2225 32351 2283 32357
rect 2225 32317 2237 32351
rect 2271 32348 2283 32351
rect 2774 32348 2780 32360
rect 2271 32320 2780 32348
rect 2271 32317 2283 32320
rect 2225 32311 2283 32317
rect 2774 32308 2780 32320
rect 2832 32308 2838 32360
rect 2866 32308 2872 32360
rect 2924 32348 2930 32360
rect 12084 32348 12112 32379
rect 12250 32376 12256 32388
rect 12308 32376 12314 32428
rect 13078 32416 13084 32428
rect 13039 32388 13084 32416
rect 13078 32376 13084 32388
rect 13136 32376 13142 32428
rect 13265 32419 13323 32425
rect 13265 32385 13277 32419
rect 13311 32416 13323 32419
rect 13556 32416 13584 32444
rect 13740 32425 13768 32456
rect 13311 32388 13584 32416
rect 13725 32419 13783 32425
rect 13311 32385 13323 32388
rect 13265 32379 13323 32385
rect 13725 32385 13737 32419
rect 13771 32385 13783 32419
rect 13725 32379 13783 32385
rect 13814 32376 13820 32428
rect 13872 32416 13878 32428
rect 13913 32419 13971 32425
rect 13913 32416 13925 32419
rect 13872 32388 13925 32416
rect 13872 32376 13878 32388
rect 13913 32385 13925 32388
rect 13959 32385 13971 32419
rect 13913 32379 13971 32385
rect 14001 32419 14059 32425
rect 14001 32385 14013 32419
rect 14047 32416 14059 32419
rect 14277 32419 14335 32425
rect 14047 32388 14228 32416
rect 14047 32385 14059 32388
rect 14001 32379 14059 32385
rect 13538 32348 13544 32360
rect 2924 32320 2969 32348
rect 12084 32320 13544 32348
rect 2924 32308 2930 32320
rect 13538 32308 13544 32320
rect 13596 32308 13602 32360
rect 13630 32308 13636 32360
rect 13688 32348 13694 32360
rect 14093 32351 14151 32357
rect 14093 32348 14105 32351
rect 13688 32320 14105 32348
rect 13688 32308 13694 32320
rect 14093 32317 14105 32320
rect 14139 32317 14151 32351
rect 14200 32348 14228 32388
rect 14277 32385 14289 32419
rect 14323 32416 14335 32419
rect 14323 32388 14412 32416
rect 14323 32385 14335 32388
rect 14277 32379 14335 32385
rect 14200 32320 14320 32348
rect 14093 32311 14151 32317
rect 14292 32292 14320 32320
rect 11606 32240 11612 32292
rect 11664 32280 11670 32292
rect 12986 32280 12992 32292
rect 11664 32252 12992 32280
rect 11664 32240 11670 32252
rect 12986 32240 12992 32252
rect 13044 32240 13050 32292
rect 14274 32240 14280 32292
rect 14332 32240 14338 32292
rect 8294 32172 8300 32224
rect 8352 32212 8358 32224
rect 10137 32215 10195 32221
rect 10137 32212 10149 32215
rect 8352 32184 10149 32212
rect 8352 32172 8358 32184
rect 10137 32181 10149 32184
rect 10183 32181 10195 32215
rect 10137 32175 10195 32181
rect 10226 32172 10232 32224
rect 10284 32212 10290 32224
rect 11054 32212 11060 32224
rect 10284 32184 11060 32212
rect 10284 32172 10290 32184
rect 11054 32172 11060 32184
rect 11112 32172 11118 32224
rect 12161 32215 12219 32221
rect 12161 32181 12173 32215
rect 12207 32212 12219 32215
rect 12802 32212 12808 32224
rect 12207 32184 12808 32212
rect 12207 32181 12219 32184
rect 12161 32175 12219 32181
rect 12802 32172 12808 32184
rect 12860 32172 12866 32224
rect 13170 32172 13176 32224
rect 13228 32212 13234 32224
rect 14384 32212 14412 32388
rect 14734 32376 14740 32428
rect 14792 32416 14798 32428
rect 14921 32419 14979 32425
rect 14921 32416 14933 32419
rect 14792 32388 14933 32416
rect 14792 32376 14798 32388
rect 14921 32385 14933 32388
rect 14967 32385 14979 32419
rect 15102 32416 15108 32428
rect 15063 32388 15108 32416
rect 14921 32379 14979 32385
rect 15102 32376 15108 32388
rect 15160 32376 15166 32428
rect 16022 32376 16028 32428
rect 16080 32416 16086 32428
rect 17218 32425 17224 32428
rect 16945 32419 17003 32425
rect 16945 32416 16957 32419
rect 16080 32388 16957 32416
rect 16080 32376 16086 32388
rect 16945 32385 16957 32388
rect 16991 32385 17003 32419
rect 16945 32379 17003 32385
rect 17212 32379 17224 32425
rect 17276 32416 17282 32428
rect 17276 32388 17312 32416
rect 17218 32376 17224 32379
rect 17276 32376 17282 32388
rect 13228 32184 14412 32212
rect 13228 32172 13234 32184
rect 15102 32172 15108 32224
rect 15160 32212 15166 32224
rect 15289 32215 15347 32221
rect 15289 32212 15301 32215
rect 15160 32184 15301 32212
rect 15160 32172 15166 32184
rect 15289 32181 15301 32184
rect 15335 32181 15347 32215
rect 15289 32175 15347 32181
rect 18325 32215 18383 32221
rect 18325 32181 18337 32215
rect 18371 32212 18383 32215
rect 18690 32212 18696 32224
rect 18371 32184 18696 32212
rect 18371 32181 18383 32184
rect 18325 32175 18383 32181
rect 18690 32172 18696 32184
rect 18748 32172 18754 32224
rect 18800 32212 18828 32456
rect 18877 32453 18889 32487
rect 18923 32484 18935 32487
rect 23842 32484 23848 32496
rect 18923 32456 23848 32484
rect 18923 32453 18935 32456
rect 18877 32447 18935 32453
rect 23842 32444 23848 32456
rect 23900 32444 23906 32496
rect 19889 32419 19947 32425
rect 19889 32385 19901 32419
rect 19935 32416 19947 32419
rect 20162 32416 20168 32428
rect 19935 32388 20168 32416
rect 19935 32385 19947 32388
rect 19889 32379 19947 32385
rect 20162 32376 20168 32388
rect 20220 32416 20226 32428
rect 20346 32416 20352 32428
rect 20220 32388 20352 32416
rect 20220 32376 20226 32388
rect 20346 32376 20352 32388
rect 20404 32376 20410 32428
rect 22002 32416 22008 32428
rect 21963 32388 22008 32416
rect 22002 32376 22008 32388
rect 22060 32376 22066 32428
rect 22272 32419 22330 32425
rect 22272 32385 22284 32419
rect 22318 32416 22330 32419
rect 23106 32416 23112 32428
rect 22318 32388 23112 32416
rect 22318 32385 22330 32388
rect 22272 32379 22330 32385
rect 23106 32376 23112 32388
rect 23164 32376 23170 32428
rect 24228 32425 24256 32524
rect 24854 32512 24860 32564
rect 24912 32552 24918 32564
rect 25406 32552 25412 32564
rect 24912 32524 25412 32552
rect 24912 32512 24918 32524
rect 25406 32512 25412 32524
rect 25464 32512 25470 32564
rect 27985 32555 28043 32561
rect 27985 32521 27997 32555
rect 28031 32521 28043 32555
rect 27985 32515 28043 32521
rect 31297 32555 31355 32561
rect 31297 32521 31309 32555
rect 31343 32552 31355 32555
rect 33502 32552 33508 32564
rect 31343 32524 33508 32552
rect 31343 32521 31355 32524
rect 31297 32515 31355 32521
rect 24302 32444 24308 32496
rect 24360 32484 24366 32496
rect 25501 32487 25559 32493
rect 25501 32484 25513 32487
rect 24360 32456 25513 32484
rect 24360 32444 24366 32456
rect 25501 32453 25513 32456
rect 25547 32453 25559 32487
rect 25501 32447 25559 32453
rect 27157 32487 27215 32493
rect 27157 32453 27169 32487
rect 27203 32484 27215 32487
rect 28000 32484 28028 32515
rect 33502 32512 33508 32524
rect 33560 32512 33566 32564
rect 29178 32484 29184 32496
rect 27203 32456 28028 32484
rect 28276 32456 29184 32484
rect 27203 32453 27215 32456
rect 27157 32447 27215 32453
rect 24213 32419 24271 32425
rect 24213 32385 24225 32419
rect 24259 32416 24271 32419
rect 25958 32416 25964 32428
rect 24259 32388 25964 32416
rect 24259 32385 24271 32388
rect 24213 32379 24271 32385
rect 25958 32376 25964 32388
rect 26016 32376 26022 32428
rect 27341 32419 27399 32425
rect 27341 32385 27353 32419
rect 27387 32416 27399 32419
rect 27522 32416 27528 32428
rect 27387 32388 27528 32416
rect 27387 32385 27399 32388
rect 27341 32379 27399 32385
rect 27522 32376 27528 32388
rect 27580 32416 27586 32428
rect 28276 32416 28304 32456
rect 29178 32444 29184 32456
rect 29236 32444 29242 32496
rect 29730 32444 29736 32496
rect 29788 32484 29794 32496
rect 30929 32487 30987 32493
rect 30929 32484 30941 32487
rect 29788 32456 30941 32484
rect 29788 32444 29794 32456
rect 30929 32453 30941 32456
rect 30975 32453 30987 32487
rect 30929 32447 30987 32453
rect 27580 32388 28304 32416
rect 28353 32419 28411 32425
rect 27580 32376 27586 32388
rect 28353 32385 28365 32419
rect 28399 32416 28411 32419
rect 29914 32416 29920 32428
rect 28399 32388 29920 32416
rect 28399 32385 28411 32388
rect 28353 32379 28411 32385
rect 29914 32376 29920 32388
rect 29972 32376 29978 32428
rect 30006 32376 30012 32428
rect 30064 32416 30070 32428
rect 30101 32419 30159 32425
rect 30101 32416 30113 32419
rect 30064 32388 30113 32416
rect 30064 32376 30070 32388
rect 30101 32385 30113 32388
rect 30147 32416 30159 32419
rect 30147 32388 30604 32416
rect 30147 32385 30159 32388
rect 30101 32379 30159 32385
rect 24026 32308 24032 32360
rect 24084 32348 24090 32360
rect 24305 32351 24363 32357
rect 24305 32348 24317 32351
rect 24084 32320 24317 32348
rect 24084 32308 24090 32320
rect 24305 32317 24317 32320
rect 24351 32317 24363 32351
rect 24305 32311 24363 32317
rect 24489 32351 24547 32357
rect 24489 32317 24501 32351
rect 24535 32317 24547 32351
rect 24489 32311 24547 32317
rect 25593 32351 25651 32357
rect 25593 32317 25605 32351
rect 25639 32317 25651 32351
rect 25593 32311 25651 32317
rect 24504 32280 24532 32311
rect 24762 32280 24768 32292
rect 24504 32252 24768 32280
rect 24762 32240 24768 32252
rect 24820 32280 24826 32292
rect 25608 32280 25636 32311
rect 24820 32252 25636 32280
rect 25976 32280 26004 32376
rect 26142 32308 26148 32360
rect 26200 32348 26206 32360
rect 28445 32351 28503 32357
rect 28445 32348 28457 32351
rect 26200 32320 28457 32348
rect 26200 32308 26206 32320
rect 28445 32317 28457 32320
rect 28491 32317 28503 32351
rect 28445 32311 28503 32317
rect 28629 32351 28687 32357
rect 28629 32317 28641 32351
rect 28675 32348 28687 32351
rect 28994 32348 29000 32360
rect 28675 32320 29000 32348
rect 28675 32317 28687 32320
rect 28629 32311 28687 32317
rect 28994 32308 29000 32320
rect 29052 32308 29058 32360
rect 30193 32351 30251 32357
rect 30193 32348 30205 32351
rect 29104 32320 30205 32348
rect 29104 32280 29132 32320
rect 30193 32317 30205 32320
rect 30239 32317 30251 32351
rect 30193 32311 30251 32317
rect 30282 32308 30288 32360
rect 30340 32348 30346 32360
rect 30576 32348 30604 32388
rect 30650 32376 30656 32428
rect 30708 32416 30714 32428
rect 31113 32419 31171 32425
rect 31113 32416 31125 32419
rect 30708 32388 31125 32416
rect 30708 32376 30714 32388
rect 31113 32385 31125 32388
rect 31159 32385 31171 32419
rect 31113 32379 31171 32385
rect 32490 32376 32496 32428
rect 32548 32416 32554 32428
rect 32677 32419 32735 32425
rect 32677 32416 32689 32419
rect 32548 32388 32689 32416
rect 32548 32376 32554 32388
rect 32677 32385 32689 32388
rect 32723 32385 32735 32419
rect 32677 32379 32735 32385
rect 32766 32376 32772 32428
rect 32824 32416 32830 32428
rect 32933 32419 32991 32425
rect 32933 32416 32945 32419
rect 32824 32388 32945 32416
rect 32824 32376 32830 32388
rect 32933 32385 32945 32388
rect 32979 32385 32991 32419
rect 32933 32379 32991 32385
rect 33318 32376 33324 32428
rect 33376 32416 33382 32428
rect 33870 32416 33876 32428
rect 33376 32388 33876 32416
rect 33376 32376 33382 32388
rect 33870 32376 33876 32388
rect 33928 32376 33934 32428
rect 47670 32416 47676 32428
rect 47631 32388 47676 32416
rect 47670 32376 47676 32388
rect 47728 32376 47734 32428
rect 30340 32320 30385 32348
rect 30576 32320 30788 32348
rect 30340 32308 30346 32320
rect 25976 32252 29132 32280
rect 24820 32240 24826 32252
rect 29178 32240 29184 32292
rect 29236 32280 29242 32292
rect 30650 32280 30656 32292
rect 29236 32252 30656 32280
rect 29236 32240 29242 32252
rect 30650 32240 30656 32252
rect 30708 32240 30714 32292
rect 20073 32215 20131 32221
rect 20073 32212 20085 32215
rect 18800 32184 20085 32212
rect 20073 32181 20085 32184
rect 20119 32212 20131 32215
rect 20346 32212 20352 32224
rect 20119 32184 20352 32212
rect 20119 32181 20131 32184
rect 20073 32175 20131 32181
rect 20346 32172 20352 32184
rect 20404 32172 20410 32224
rect 21358 32172 21364 32224
rect 21416 32212 21422 32224
rect 23382 32212 23388 32224
rect 21416 32184 23388 32212
rect 21416 32172 21422 32184
rect 23382 32172 23388 32184
rect 23440 32172 23446 32224
rect 23474 32172 23480 32224
rect 23532 32212 23538 32224
rect 23845 32215 23903 32221
rect 23845 32212 23857 32215
rect 23532 32184 23857 32212
rect 23532 32172 23538 32184
rect 23845 32181 23857 32184
rect 23891 32181 23903 32215
rect 23845 32175 23903 32181
rect 24486 32172 24492 32224
rect 24544 32212 24550 32224
rect 25041 32215 25099 32221
rect 25041 32212 25053 32215
rect 24544 32184 25053 32212
rect 24544 32172 24550 32184
rect 25041 32181 25053 32184
rect 25087 32181 25099 32215
rect 25041 32175 25099 32181
rect 27525 32215 27583 32221
rect 27525 32181 27537 32215
rect 27571 32212 27583 32215
rect 28534 32212 28540 32224
rect 27571 32184 28540 32212
rect 27571 32181 27583 32184
rect 27525 32175 27583 32181
rect 28534 32172 28540 32184
rect 28592 32172 28598 32224
rect 29733 32215 29791 32221
rect 29733 32181 29745 32215
rect 29779 32212 29791 32215
rect 30466 32212 30472 32224
rect 29779 32184 30472 32212
rect 29779 32181 29791 32184
rect 29733 32175 29791 32181
rect 30466 32172 30472 32184
rect 30524 32172 30530 32224
rect 30760 32212 30788 32320
rect 46842 32308 46848 32360
rect 46900 32348 46906 32360
rect 47857 32351 47915 32357
rect 47857 32348 47869 32351
rect 46900 32320 47869 32348
rect 46900 32308 46906 32320
rect 47857 32317 47869 32320
rect 47903 32317 47915 32351
rect 47857 32311 47915 32317
rect 34054 32212 34060 32224
rect 30760 32184 34060 32212
rect 34054 32172 34060 32184
rect 34112 32172 34118 32224
rect 1104 32122 48852 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 48852 32122
rect 1104 32048 48852 32070
rect 2774 31968 2780 32020
rect 2832 32008 2838 32020
rect 2961 32011 3019 32017
rect 2961 32008 2973 32011
rect 2832 31980 2973 32008
rect 2832 31968 2838 31980
rect 2961 31977 2973 31980
rect 3007 31977 3019 32011
rect 2961 31971 3019 31977
rect 9677 32011 9735 32017
rect 9677 31977 9689 32011
rect 9723 32008 9735 32011
rect 10594 32008 10600 32020
rect 9723 31980 10600 32008
rect 9723 31977 9735 31980
rect 9677 31971 9735 31977
rect 10594 31968 10600 31980
rect 10652 31968 10658 32020
rect 12526 32008 12532 32020
rect 10701 31980 12532 32008
rect 10502 31900 10508 31952
rect 10560 31940 10566 31952
rect 10701 31940 10729 31980
rect 12526 31968 12532 31980
rect 12584 31968 12590 32020
rect 15841 32011 15899 32017
rect 15841 31977 15853 32011
rect 15887 32008 15899 32011
rect 17218 32008 17224 32020
rect 15887 31980 17224 32008
rect 15887 31977 15899 31980
rect 15841 31971 15899 31977
rect 17218 31968 17224 31980
rect 17276 31968 17282 32020
rect 17310 31968 17316 32020
rect 17368 32008 17374 32020
rect 22005 32011 22063 32017
rect 17368 31980 19564 32008
rect 17368 31968 17374 31980
rect 11514 31940 11520 31952
rect 10560 31912 10729 31940
rect 11475 31912 11520 31940
rect 10560 31900 10566 31912
rect 1854 31804 1860 31816
rect 1815 31776 1860 31804
rect 1854 31764 1860 31776
rect 1912 31764 1918 31816
rect 2038 31804 2044 31816
rect 1999 31776 2044 31804
rect 2038 31764 2044 31776
rect 2096 31764 2102 31816
rect 2869 31807 2927 31813
rect 2869 31773 2881 31807
rect 2915 31804 2927 31807
rect 7650 31804 7656 31816
rect 2915 31776 7656 31804
rect 2915 31773 2927 31776
rect 2869 31767 2927 31773
rect 7650 31764 7656 31776
rect 7708 31764 7714 31816
rect 9674 31804 9680 31816
rect 9635 31776 9680 31804
rect 9674 31764 9680 31776
rect 9732 31764 9738 31816
rect 9861 31807 9919 31813
rect 9861 31773 9873 31807
rect 9907 31804 9919 31807
rect 10226 31804 10232 31816
rect 9907 31776 10232 31804
rect 9907 31773 9919 31776
rect 9861 31767 9919 31773
rect 10226 31764 10232 31776
rect 10284 31764 10290 31816
rect 10612 31813 10640 31912
rect 11514 31900 11520 31912
rect 11572 31900 11578 31952
rect 11698 31900 11704 31952
rect 11756 31940 11762 31952
rect 12894 31940 12900 31952
rect 11756 31912 12900 31940
rect 11756 31900 11762 31912
rect 12894 31900 12900 31912
rect 12952 31900 12958 31952
rect 12986 31900 12992 31952
rect 13044 31940 13050 31952
rect 13044 31912 14320 31940
rect 13044 31900 13050 31912
rect 12253 31875 12311 31881
rect 12253 31841 12265 31875
rect 12299 31872 12311 31875
rect 12434 31872 12440 31884
rect 12299 31844 12440 31872
rect 12299 31841 12311 31844
rect 12253 31835 12311 31841
rect 12434 31832 12440 31844
rect 12492 31832 12498 31884
rect 13449 31875 13507 31881
rect 13449 31872 13461 31875
rect 12728 31844 13461 31872
rect 10597 31807 10655 31813
rect 10781 31807 10839 31813
rect 10597 31773 10609 31807
rect 10643 31773 10655 31807
rect 10597 31767 10655 31773
rect 10686 31801 10744 31807
rect 10686 31767 10698 31801
rect 10732 31767 10744 31801
rect 10781 31773 10793 31807
rect 10827 31804 10839 31807
rect 10870 31804 10876 31816
rect 10827 31776 10876 31804
rect 10827 31773 10839 31776
rect 10781 31767 10839 31773
rect 10686 31761 10744 31767
rect 10870 31764 10876 31776
rect 10928 31764 10934 31816
rect 10962 31764 10968 31816
rect 11020 31804 11026 31816
rect 11698 31804 11704 31816
rect 11020 31776 11704 31804
rect 11020 31764 11026 31776
rect 11698 31764 11704 31776
rect 11756 31764 11762 31816
rect 11790 31764 11796 31816
rect 11848 31804 11854 31816
rect 12526 31804 12532 31816
rect 11848 31776 11893 31804
rect 12487 31776 12532 31804
rect 11848 31764 11854 31776
rect 12526 31764 12532 31776
rect 12584 31764 12590 31816
rect 12728 31813 12756 31844
rect 13449 31841 13461 31844
rect 13495 31841 13507 31875
rect 13449 31835 13507 31841
rect 14292 31816 14320 31912
rect 15286 31900 15292 31952
rect 15344 31940 15350 31952
rect 18322 31940 18328 31952
rect 15344 31912 16988 31940
rect 18235 31912 18328 31940
rect 15344 31900 15350 31912
rect 16960 31881 16988 31912
rect 18322 31900 18328 31912
rect 18380 31940 18386 31952
rect 18380 31912 19288 31940
rect 18380 31900 18386 31912
rect 19260 31881 19288 31912
rect 16945 31875 17003 31881
rect 16945 31841 16957 31875
rect 16991 31841 17003 31875
rect 16945 31835 17003 31841
rect 19245 31875 19303 31881
rect 19245 31841 19257 31875
rect 19291 31841 19303 31875
rect 19426 31872 19432 31884
rect 19387 31844 19432 31872
rect 19245 31835 19303 31841
rect 19426 31832 19432 31844
rect 19484 31832 19490 31884
rect 19536 31872 19564 31980
rect 22005 31977 22017 32011
rect 22051 32008 22063 32011
rect 22278 32008 22284 32020
rect 22051 31980 22284 32008
rect 22051 31977 22063 31980
rect 22005 31971 22063 31977
rect 22278 31968 22284 31980
rect 22336 31968 22342 32020
rect 23106 32008 23112 32020
rect 23067 31980 23112 32008
rect 23106 31968 23112 31980
rect 23164 31968 23170 32020
rect 25406 31968 25412 32020
rect 25464 32008 25470 32020
rect 26789 32011 26847 32017
rect 26789 32008 26801 32011
rect 25464 31980 26801 32008
rect 25464 31968 25470 31980
rect 26789 31977 26801 31980
rect 26835 31977 26847 32011
rect 26789 31971 26847 31977
rect 29914 31968 29920 32020
rect 29972 32008 29978 32020
rect 30009 32011 30067 32017
rect 30009 32008 30021 32011
rect 29972 31980 30021 32008
rect 29972 31968 29978 31980
rect 30009 31977 30021 31980
rect 30055 31977 30067 32011
rect 30009 31971 30067 31977
rect 31297 32011 31355 32017
rect 31297 31977 31309 32011
rect 31343 32008 31355 32011
rect 31662 32008 31668 32020
rect 31343 31980 31668 32008
rect 31343 31977 31355 31980
rect 31297 31971 31355 31977
rect 31662 31968 31668 31980
rect 31720 31968 31726 32020
rect 31757 32011 31815 32017
rect 31757 31977 31769 32011
rect 31803 32008 31815 32011
rect 32766 32008 32772 32020
rect 31803 31980 32772 32008
rect 31803 31977 31815 31980
rect 31757 31971 31815 31977
rect 32766 31968 32772 31980
rect 32824 31968 32830 32020
rect 27430 31900 27436 31952
rect 27488 31940 27494 31952
rect 27488 31912 28994 31940
rect 27488 31900 27494 31912
rect 22922 31872 22928 31884
rect 19536 31844 22324 31872
rect 12621 31807 12679 31813
rect 12621 31773 12633 31807
rect 12667 31773 12679 31807
rect 12621 31767 12679 31773
rect 12713 31807 12771 31813
rect 12713 31773 12725 31807
rect 12759 31773 12771 31807
rect 12894 31804 12900 31816
rect 12855 31776 12900 31804
rect 12713 31767 12771 31773
rect 10704 31680 10732 31761
rect 11517 31739 11575 31745
rect 11517 31705 11529 31739
rect 11563 31736 11575 31739
rect 11606 31736 11612 31748
rect 11563 31708 11612 31736
rect 11563 31705 11575 31708
rect 11517 31699 11575 31705
rect 11606 31696 11612 31708
rect 11664 31696 11670 31748
rect 12158 31696 12164 31748
rect 12216 31736 12222 31748
rect 12636 31736 12664 31767
rect 12894 31764 12900 31776
rect 12952 31764 12958 31816
rect 13357 31807 13415 31813
rect 13357 31773 13369 31807
rect 13403 31804 13415 31807
rect 13403 31776 13492 31804
rect 13403 31773 13415 31776
rect 13357 31767 13415 31773
rect 12216 31708 12664 31736
rect 13464 31736 13492 31776
rect 13538 31764 13544 31816
rect 13596 31804 13602 31816
rect 13596 31776 13641 31804
rect 13596 31764 13602 31776
rect 14274 31764 14280 31816
rect 14332 31804 14338 31816
rect 16117 31807 16175 31813
rect 16117 31804 16129 31807
rect 14332 31776 16129 31804
rect 14332 31764 14338 31776
rect 16117 31773 16129 31776
rect 16163 31773 16175 31807
rect 16117 31767 16175 31773
rect 16209 31807 16267 31813
rect 16209 31773 16221 31807
rect 16255 31773 16267 31807
rect 16209 31767 16267 31773
rect 16301 31807 16359 31813
rect 16301 31773 16313 31807
rect 16347 31804 16359 31807
rect 16485 31807 16543 31813
rect 16347 31776 16436 31804
rect 16347 31773 16359 31776
rect 16301 31767 16359 31773
rect 14918 31736 14924 31748
rect 13464 31708 14924 31736
rect 12216 31696 12222 31708
rect 14918 31696 14924 31708
rect 14976 31696 14982 31748
rect 10318 31668 10324 31680
rect 10279 31640 10324 31668
rect 10318 31628 10324 31640
rect 10376 31628 10382 31680
rect 10686 31628 10692 31680
rect 10744 31628 10750 31680
rect 11701 31671 11759 31677
rect 11701 31637 11713 31671
rect 11747 31668 11759 31671
rect 12250 31668 12256 31680
rect 11747 31640 12256 31668
rect 11747 31637 11759 31640
rect 11701 31631 11759 31637
rect 12250 31628 12256 31640
rect 12308 31628 12314 31680
rect 14826 31628 14832 31680
rect 14884 31668 14890 31680
rect 15010 31668 15016 31680
rect 14884 31640 15016 31668
rect 14884 31628 14890 31640
rect 15010 31628 15016 31640
rect 15068 31628 15074 31680
rect 16224 31668 16252 31767
rect 16408 31736 16436 31776
rect 16485 31773 16497 31807
rect 16531 31804 16543 31807
rect 21082 31804 21088 31816
rect 16531 31776 17356 31804
rect 21043 31776 21088 31804
rect 16531 31773 16543 31776
rect 16485 31767 16543 31773
rect 17328 31748 17356 31776
rect 21082 31764 21088 31776
rect 21140 31764 21146 31816
rect 22296 31813 22324 31844
rect 22388 31844 22928 31872
rect 22388 31813 22416 31844
rect 22922 31832 22928 31844
rect 22980 31872 22986 31884
rect 22980 31844 23520 31872
rect 22980 31832 22986 31844
rect 22281 31807 22339 31813
rect 22281 31773 22293 31807
rect 22327 31773 22339 31807
rect 22281 31767 22339 31773
rect 22373 31807 22431 31813
rect 22373 31773 22385 31807
rect 22419 31773 22431 31807
rect 22373 31767 22431 31773
rect 22462 31764 22468 31816
rect 22520 31804 22526 31816
rect 22649 31807 22707 31813
rect 22520 31776 22565 31804
rect 22520 31764 22526 31776
rect 22649 31773 22661 31807
rect 22695 31804 22707 31807
rect 23382 31804 23388 31816
rect 22695 31776 22729 31804
rect 23343 31776 23388 31804
rect 22695 31773 22707 31776
rect 22649 31767 22707 31773
rect 16574 31736 16580 31748
rect 16408 31708 16580 31736
rect 16574 31696 16580 31708
rect 16632 31696 16638 31748
rect 16666 31696 16672 31748
rect 16724 31736 16730 31748
rect 17190 31739 17248 31745
rect 17190 31736 17202 31739
rect 16724 31708 17202 31736
rect 16724 31696 16730 31708
rect 17190 31705 17202 31708
rect 17236 31705 17248 31739
rect 17190 31699 17248 31705
rect 17310 31696 17316 31748
rect 17368 31696 17374 31748
rect 22094 31696 22100 31748
rect 22152 31736 22158 31748
rect 22664 31736 22692 31767
rect 23382 31764 23388 31776
rect 23440 31764 23446 31816
rect 23492 31813 23520 31844
rect 28166 31832 28172 31884
rect 28224 31872 28230 31884
rect 28534 31872 28540 31884
rect 28224 31844 28396 31872
rect 28224 31832 28230 31844
rect 23477 31807 23535 31813
rect 23477 31773 23489 31807
rect 23523 31773 23535 31807
rect 23477 31767 23535 31773
rect 23566 31764 23572 31816
rect 23624 31804 23630 31816
rect 23753 31807 23811 31813
rect 23624 31776 23669 31804
rect 23624 31764 23630 31776
rect 23753 31773 23765 31807
rect 23799 31773 23811 31807
rect 24486 31804 24492 31816
rect 24447 31776 24492 31804
rect 23753 31767 23811 31773
rect 23768 31736 23796 31767
rect 24486 31764 24492 31776
rect 24544 31764 24550 31816
rect 25409 31807 25467 31813
rect 25409 31773 25421 31807
rect 25455 31804 25467 31807
rect 26694 31804 26700 31816
rect 25455 31776 26700 31804
rect 25455 31773 25467 31776
rect 25409 31767 25467 31773
rect 26694 31764 26700 31776
rect 26752 31764 26758 31816
rect 28368 31813 28396 31844
rect 28460 31844 28540 31872
rect 28460 31813 28488 31844
rect 28534 31832 28540 31844
rect 28592 31832 28598 31884
rect 28966 31872 28994 31912
rect 29362 31900 29368 31952
rect 29420 31940 29426 31952
rect 29546 31940 29552 31952
rect 29420 31912 29552 31940
rect 29420 31900 29426 31912
rect 29546 31900 29552 31912
rect 29604 31940 29610 31952
rect 30469 31943 30527 31949
rect 29604 31912 30328 31940
rect 29604 31900 29610 31912
rect 30190 31872 30196 31884
rect 28966 31844 29868 31872
rect 30151 31844 30196 31872
rect 28261 31807 28319 31813
rect 28261 31773 28273 31807
rect 28307 31773 28319 31807
rect 28261 31767 28319 31773
rect 28353 31807 28411 31813
rect 28353 31773 28365 31807
rect 28399 31773 28411 31807
rect 28353 31767 28411 31773
rect 28445 31807 28503 31813
rect 28445 31773 28457 31807
rect 28491 31773 28503 31807
rect 28445 31767 28503 31773
rect 24026 31736 24032 31748
rect 22152 31708 24032 31736
rect 22152 31696 22158 31708
rect 24026 31696 24032 31708
rect 24084 31696 24090 31748
rect 24578 31696 24584 31748
rect 24636 31736 24642 31748
rect 24673 31739 24731 31745
rect 24673 31736 24685 31739
rect 24636 31708 24685 31736
rect 24636 31696 24642 31708
rect 24673 31705 24685 31708
rect 24719 31705 24731 31739
rect 24673 31699 24731 31705
rect 25314 31696 25320 31748
rect 25372 31736 25378 31748
rect 25654 31739 25712 31745
rect 25654 31736 25666 31739
rect 25372 31708 25666 31736
rect 25372 31696 25378 31708
rect 25654 31705 25666 31708
rect 25700 31705 25712 31739
rect 25654 31699 25712 31705
rect 28276 31680 28304 31767
rect 28626 31764 28632 31816
rect 28684 31804 28690 31816
rect 28684 31776 28729 31804
rect 28684 31764 28690 31776
rect 29840 31736 29868 31844
rect 30190 31832 30196 31844
rect 30248 31832 30254 31884
rect 30006 31804 30012 31816
rect 29967 31776 30012 31804
rect 30006 31764 30012 31776
rect 30064 31764 30070 31816
rect 30300 31813 30328 31912
rect 30469 31909 30481 31943
rect 30515 31909 30527 31943
rect 32953 31943 33011 31949
rect 32953 31940 32965 31943
rect 30469 31903 30527 31909
rect 30944 31912 32965 31940
rect 30484 31872 30512 31903
rect 30392 31844 30512 31872
rect 30285 31807 30343 31813
rect 30285 31773 30297 31807
rect 30331 31773 30343 31807
rect 30285 31767 30343 31773
rect 30392 31736 30420 31844
rect 30944 31813 30972 31912
rect 32953 31909 32965 31912
rect 32999 31909 33011 31943
rect 32953 31903 33011 31909
rect 32306 31872 32312 31884
rect 32140 31844 32312 31872
rect 30929 31807 30987 31813
rect 30929 31773 30941 31807
rect 30975 31773 30987 31807
rect 30929 31767 30987 31773
rect 31113 31807 31171 31813
rect 31113 31773 31125 31807
rect 31159 31804 31171 31807
rect 31202 31804 31208 31816
rect 31159 31776 31208 31804
rect 31159 31773 31171 31776
rect 31113 31767 31171 31773
rect 31202 31764 31208 31776
rect 31260 31764 31266 31816
rect 31846 31764 31852 31816
rect 31904 31804 31910 31816
rect 32140 31813 32168 31844
rect 32306 31832 32312 31844
rect 32364 31832 32370 31884
rect 33502 31872 33508 31884
rect 33463 31844 33508 31872
rect 33502 31832 33508 31844
rect 33560 31832 33566 31884
rect 37829 31875 37887 31881
rect 37829 31841 37841 31875
rect 37875 31872 37887 31875
rect 46106 31872 46112 31884
rect 37875 31844 46112 31872
rect 37875 31841 37887 31844
rect 37829 31835 37887 31841
rect 46106 31832 46112 31844
rect 46164 31832 46170 31884
rect 31987 31807 32045 31813
rect 31987 31804 31999 31807
rect 31904 31776 31999 31804
rect 31904 31764 31910 31776
rect 31987 31773 31999 31776
rect 32033 31773 32045 31807
rect 31987 31767 32045 31773
rect 32125 31807 32183 31813
rect 32125 31773 32137 31807
rect 32171 31773 32183 31807
rect 32125 31767 32183 31773
rect 32214 31764 32220 31816
rect 32272 31813 32278 31816
rect 32272 31804 32280 31813
rect 32272 31776 32317 31804
rect 32272 31767 32280 31776
rect 32272 31764 32278 31767
rect 32398 31764 32404 31816
rect 32456 31804 32462 31816
rect 33413 31807 33471 31813
rect 32456 31776 32501 31804
rect 32456 31764 32462 31776
rect 33413 31773 33425 31807
rect 33459 31804 33471 31807
rect 34054 31804 34060 31816
rect 33459 31776 34060 31804
rect 33459 31773 33471 31776
rect 33413 31767 33471 31773
rect 34054 31764 34060 31776
rect 34112 31764 34118 31816
rect 35986 31804 35992 31816
rect 35947 31776 35992 31804
rect 35986 31764 35992 31776
rect 36044 31764 36050 31816
rect 47946 31804 47952 31816
rect 47907 31776 47952 31804
rect 47946 31764 47952 31776
rect 48004 31764 48010 31816
rect 36170 31736 36176 31748
rect 29840 31708 30420 31736
rect 36131 31708 36176 31736
rect 36170 31696 36176 31708
rect 36228 31696 36234 31748
rect 17034 31668 17040 31680
rect 16224 31640 17040 31668
rect 17034 31628 17040 31640
rect 17092 31628 17098 31680
rect 24857 31671 24915 31677
rect 24857 31637 24869 31671
rect 24903 31668 24915 31671
rect 25774 31668 25780 31680
rect 24903 31640 25780 31668
rect 24903 31637 24915 31640
rect 24857 31631 24915 31637
rect 25774 31628 25780 31640
rect 25832 31628 25838 31680
rect 27982 31668 27988 31680
rect 27943 31640 27988 31668
rect 27982 31628 27988 31640
rect 28040 31628 28046 31680
rect 28258 31628 28264 31680
rect 28316 31628 28322 31680
rect 33321 31671 33379 31677
rect 33321 31637 33333 31671
rect 33367 31668 33379 31671
rect 34238 31668 34244 31680
rect 33367 31640 34244 31668
rect 33367 31637 33379 31640
rect 33321 31631 33379 31637
rect 34238 31628 34244 31640
rect 34296 31628 34302 31680
rect 48038 31668 48044 31680
rect 47999 31640 48044 31668
rect 48038 31628 48044 31640
rect 48096 31628 48102 31680
rect 1104 31578 48852 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 48852 31578
rect 1104 31504 48852 31526
rect 1578 31424 1584 31476
rect 1636 31464 1642 31476
rect 1636 31436 12434 31464
rect 1636 31424 1642 31436
rect 9208 31399 9266 31405
rect 7116 31368 8248 31396
rect 7116 31337 7144 31368
rect 7101 31331 7159 31337
rect 7101 31297 7113 31331
rect 7147 31297 7159 31331
rect 7101 31291 7159 31297
rect 7368 31331 7426 31337
rect 7368 31297 7380 31331
rect 7414 31328 7426 31331
rect 7414 31300 8156 31328
rect 7414 31297 7426 31300
rect 7368 31291 7426 31297
rect 1946 31260 1952 31272
rect 1907 31232 1952 31260
rect 1946 31220 1952 31232
rect 2004 31220 2010 31272
rect 2133 31263 2191 31269
rect 2133 31229 2145 31263
rect 2179 31260 2191 31263
rect 2866 31260 2872 31272
rect 2179 31232 2872 31260
rect 2179 31229 2191 31232
rect 2133 31223 2191 31229
rect 2866 31220 2872 31232
rect 2924 31220 2930 31272
rect 3050 31260 3056 31272
rect 3011 31232 3056 31260
rect 3050 31220 3056 31232
rect 3108 31220 3114 31272
rect 8128 31192 8156 31300
rect 8220 31272 8248 31368
rect 9208 31365 9220 31399
rect 9254 31396 9266 31399
rect 10318 31396 10324 31408
rect 9254 31368 10324 31396
rect 9254 31365 9266 31368
rect 9208 31359 9266 31365
rect 10318 31356 10324 31368
rect 10376 31356 10382 31408
rect 10870 31396 10876 31408
rect 10831 31368 10876 31396
rect 10870 31356 10876 31368
rect 10928 31356 10934 31408
rect 12406 31396 12434 31436
rect 12986 31424 12992 31476
rect 13044 31464 13050 31476
rect 13262 31464 13268 31476
rect 13044 31436 13268 31464
rect 13044 31424 13050 31436
rect 13262 31424 13268 31436
rect 13320 31424 13326 31476
rect 13449 31467 13507 31473
rect 13449 31433 13461 31467
rect 13495 31464 13507 31467
rect 13630 31464 13636 31476
rect 13495 31436 13636 31464
rect 13495 31433 13507 31436
rect 13449 31427 13507 31433
rect 13630 31424 13636 31436
rect 13688 31424 13694 31476
rect 14458 31464 14464 31476
rect 14419 31436 14464 31464
rect 14458 31424 14464 31436
rect 14516 31424 14522 31476
rect 23477 31467 23535 31473
rect 14568 31436 22094 31464
rect 14568 31396 14596 31436
rect 16666 31396 16672 31408
rect 12406 31368 14596 31396
rect 14660 31368 15415 31396
rect 16627 31368 16672 31396
rect 10781 31331 10839 31337
rect 10781 31297 10793 31331
rect 10827 31297 10839 31331
rect 10962 31328 10968 31340
rect 10923 31300 10968 31328
rect 10781 31291 10839 31297
rect 8202 31220 8208 31272
rect 8260 31260 8266 31272
rect 8941 31263 8999 31269
rect 8941 31260 8953 31263
rect 8260 31232 8953 31260
rect 8260 31220 8266 31232
rect 8941 31229 8953 31232
rect 8987 31229 8999 31263
rect 10796 31260 10824 31291
rect 10962 31288 10968 31300
rect 11020 31288 11026 31340
rect 11790 31288 11796 31340
rect 11848 31328 11854 31340
rect 11974 31328 11980 31340
rect 11848 31300 11980 31328
rect 11848 31288 11854 31300
rect 11974 31288 11980 31300
rect 12032 31288 12038 31340
rect 12161 31331 12219 31337
rect 12161 31297 12173 31331
rect 12207 31297 12219 31331
rect 12161 31291 12219 31297
rect 11514 31260 11520 31272
rect 10796 31232 11520 31260
rect 8941 31223 8999 31229
rect 11514 31220 11520 31232
rect 11572 31220 11578 31272
rect 12176 31260 12204 31291
rect 13078 31288 13084 31340
rect 13136 31328 13142 31340
rect 13354 31328 13360 31340
rect 13136 31300 13360 31328
rect 13136 31288 13142 31300
rect 13354 31288 13360 31300
rect 13412 31288 13418 31340
rect 14001 31331 14059 31337
rect 14001 31297 14013 31331
rect 14047 31328 14059 31331
rect 14277 31331 14335 31337
rect 14047 31300 14228 31328
rect 14047 31297 14059 31300
rect 14001 31291 14059 31297
rect 13262 31260 13268 31272
rect 12176 31232 13268 31260
rect 8294 31192 8300 31204
rect 8128 31164 8300 31192
rect 8294 31152 8300 31164
rect 8352 31152 8358 31204
rect 10410 31152 10416 31204
rect 10468 31192 10474 31204
rect 12176 31192 12204 31232
rect 13262 31220 13268 31232
rect 13320 31260 13326 31272
rect 14093 31263 14151 31269
rect 14093 31260 14105 31263
rect 13320 31232 14105 31260
rect 13320 31220 13326 31232
rect 14093 31229 14105 31232
rect 14139 31229 14151 31263
rect 14200 31260 14228 31300
rect 14277 31297 14289 31331
rect 14323 31328 14335 31331
rect 14458 31328 14464 31340
rect 14323 31300 14464 31328
rect 14323 31297 14335 31300
rect 14277 31291 14335 31297
rect 14458 31288 14464 31300
rect 14516 31328 14522 31340
rect 14660 31328 14688 31368
rect 14516 31300 14688 31328
rect 14516 31288 14522 31300
rect 14826 31288 14832 31340
rect 14884 31328 14890 31340
rect 14921 31331 14979 31337
rect 14921 31328 14933 31331
rect 14884 31300 14933 31328
rect 14884 31288 14890 31300
rect 14921 31297 14933 31300
rect 14967 31297 14979 31331
rect 14921 31291 14979 31297
rect 15010 31288 15016 31340
rect 15068 31328 15074 31340
rect 15105 31331 15163 31337
rect 15105 31328 15117 31331
rect 15068 31300 15117 31328
rect 15068 31288 15074 31300
rect 15105 31297 15117 31300
rect 15151 31297 15163 31331
rect 15105 31291 15163 31297
rect 15194 31288 15200 31340
rect 15252 31328 15258 31340
rect 15252 31300 15297 31328
rect 15252 31288 15258 31300
rect 14844 31260 14872 31288
rect 14200 31232 14872 31260
rect 14093 31223 14151 31229
rect 14458 31192 14464 31204
rect 10468 31164 12204 31192
rect 12268 31164 14464 31192
rect 10468 31152 10474 31164
rect 8481 31127 8539 31133
rect 8481 31093 8493 31127
rect 8527 31124 8539 31127
rect 10134 31124 10140 31136
rect 8527 31096 10140 31124
rect 8527 31093 8539 31096
rect 8481 31087 8539 31093
rect 10134 31084 10140 31096
rect 10192 31084 10198 31136
rect 10321 31127 10379 31133
rect 10321 31093 10333 31127
rect 10367 31124 10379 31127
rect 10778 31124 10784 31136
rect 10367 31096 10784 31124
rect 10367 31093 10379 31096
rect 10321 31087 10379 31093
rect 10778 31084 10784 31096
rect 10836 31084 10842 31136
rect 11698 31084 11704 31136
rect 11756 31124 11762 31136
rect 12268 31124 12296 31164
rect 14458 31152 14464 31164
rect 14516 31152 14522 31204
rect 14918 31192 14924 31204
rect 14879 31164 14924 31192
rect 14918 31152 14924 31164
rect 14976 31152 14982 31204
rect 15387 31192 15415 31368
rect 16666 31356 16672 31368
rect 16724 31356 16730 31408
rect 16758 31356 16764 31408
rect 16816 31396 16822 31408
rect 17773 31399 17831 31405
rect 17773 31396 17785 31399
rect 16816 31368 17785 31396
rect 16816 31356 16822 31368
rect 17773 31365 17785 31368
rect 17819 31365 17831 31399
rect 17773 31359 17831 31365
rect 17957 31399 18015 31405
rect 17957 31365 17969 31399
rect 18003 31396 18015 31399
rect 18322 31396 18328 31408
rect 18003 31368 18328 31396
rect 18003 31365 18015 31368
rect 17957 31359 18015 31365
rect 18322 31356 18328 31368
rect 18380 31356 18386 31408
rect 18874 31396 18880 31408
rect 18835 31368 18880 31396
rect 18874 31356 18880 31368
rect 18932 31356 18938 31408
rect 20162 31356 20168 31408
rect 20220 31396 20226 31408
rect 20220 31368 21864 31396
rect 20220 31356 20226 31368
rect 16022 31288 16028 31340
rect 16080 31328 16086 31340
rect 16899 31331 16957 31337
rect 16899 31328 16911 31331
rect 16080 31300 16911 31328
rect 16080 31288 16086 31300
rect 16899 31297 16911 31300
rect 16945 31297 16957 31331
rect 17034 31328 17040 31340
rect 16995 31300 17040 31328
rect 16899 31291 16957 31297
rect 17034 31288 17040 31300
rect 17092 31288 17098 31340
rect 17129 31331 17187 31337
rect 17129 31297 17141 31331
rect 17175 31297 17187 31331
rect 17129 31291 17187 31297
rect 17144 31260 17172 31291
rect 17218 31288 17224 31340
rect 17276 31328 17282 31340
rect 21836 31337 21864 31368
rect 17313 31331 17371 31337
rect 17313 31328 17325 31331
rect 17276 31300 17325 31328
rect 17276 31288 17282 31300
rect 17313 31297 17325 31300
rect 17359 31297 17371 31331
rect 17313 31291 17371 31297
rect 21085 31331 21143 31337
rect 21085 31297 21097 31331
rect 21131 31297 21143 31331
rect 21085 31291 21143 31297
rect 21821 31331 21879 31337
rect 21821 31297 21833 31331
rect 21867 31297 21879 31331
rect 22066 31328 22094 31436
rect 23477 31433 23489 31467
rect 23523 31464 23535 31467
rect 23566 31464 23572 31476
rect 23523 31436 23572 31464
rect 23523 31433 23535 31436
rect 23477 31427 23535 31433
rect 23566 31424 23572 31436
rect 23624 31424 23630 31476
rect 24394 31424 24400 31476
rect 24452 31464 24458 31476
rect 25314 31464 25320 31476
rect 24452 31436 24532 31464
rect 25275 31436 25320 31464
rect 24452 31424 24458 31436
rect 23109 31399 23167 31405
rect 23109 31365 23121 31399
rect 23155 31396 23167 31399
rect 24504 31396 24532 31436
rect 25314 31424 25320 31436
rect 25372 31424 25378 31476
rect 28077 31467 28135 31473
rect 28077 31433 28089 31467
rect 28123 31464 28135 31467
rect 28626 31464 28632 31476
rect 28123 31436 28632 31464
rect 28123 31433 28135 31436
rect 28077 31427 28135 31433
rect 28626 31424 28632 31436
rect 28684 31424 28690 31476
rect 30837 31467 30895 31473
rect 30837 31433 30849 31467
rect 30883 31464 30895 31467
rect 32214 31464 32220 31476
rect 30883 31436 32220 31464
rect 30883 31433 30895 31436
rect 30837 31427 30895 31433
rect 32214 31424 32220 31436
rect 32272 31424 32278 31476
rect 36081 31467 36139 31473
rect 36081 31433 36093 31467
rect 36127 31464 36139 31467
rect 36170 31464 36176 31476
rect 36127 31436 36176 31464
rect 36127 31433 36139 31436
rect 36081 31427 36139 31433
rect 36170 31424 36176 31436
rect 36228 31424 36234 31476
rect 24581 31399 24639 31405
rect 24581 31396 24593 31399
rect 23155 31368 23520 31396
rect 24504 31368 24593 31396
rect 23155 31365 23167 31368
rect 23109 31359 23167 31365
rect 23492 31340 23520 31368
rect 24581 31365 24593 31368
rect 24627 31365 24639 31399
rect 24581 31359 24639 31365
rect 25038 31356 25044 31408
rect 25096 31396 25102 31408
rect 25096 31368 25697 31396
rect 25096 31356 25102 31368
rect 23293 31331 23351 31337
rect 22066 31300 23244 31328
rect 21821 31291 21879 31297
rect 18141 31263 18199 31269
rect 18141 31260 18153 31263
rect 17144 31232 18153 31260
rect 18141 31229 18153 31232
rect 18187 31229 18199 31263
rect 18690 31260 18696 31272
rect 18651 31232 18696 31260
rect 18141 31223 18199 31229
rect 18690 31220 18696 31232
rect 18748 31220 18754 31272
rect 20530 31260 20536 31272
rect 20491 31232 20536 31260
rect 20530 31220 20536 31232
rect 20588 31220 20594 31272
rect 17678 31192 17684 31204
rect 15387 31164 17684 31192
rect 17678 31152 17684 31164
rect 17736 31152 17742 31204
rect 21100 31192 21128 31291
rect 22094 31220 22100 31272
rect 22152 31260 22158 31272
rect 23216 31260 23244 31300
rect 23293 31297 23305 31331
rect 23339 31328 23351 31331
rect 23382 31328 23388 31340
rect 23339 31300 23388 31328
rect 23339 31297 23351 31300
rect 23293 31291 23351 31297
rect 23382 31288 23388 31300
rect 23440 31288 23446 31340
rect 23474 31288 23480 31340
rect 23532 31288 23538 31340
rect 24489 31331 24547 31337
rect 24489 31297 24501 31331
rect 24535 31328 24547 31331
rect 24670 31328 24676 31340
rect 24535 31300 24676 31328
rect 24535 31297 24547 31300
rect 24489 31291 24547 31297
rect 24670 31288 24676 31300
rect 24728 31288 24734 31340
rect 25669 31337 25697 31368
rect 26050 31356 26056 31408
rect 26108 31396 26114 31408
rect 28721 31399 28779 31405
rect 28721 31396 28733 31399
rect 26108 31368 28733 31396
rect 26108 31356 26114 31368
rect 28721 31365 28733 31368
rect 28767 31365 28779 31399
rect 28721 31359 28779 31365
rect 29641 31399 29699 31405
rect 29641 31365 29653 31399
rect 29687 31396 29699 31399
rect 30742 31396 30748 31408
rect 29687 31368 30748 31396
rect 29687 31365 29699 31368
rect 29641 31359 29699 31365
rect 30742 31356 30748 31368
rect 30800 31356 30806 31408
rect 48038 31396 48044 31408
rect 31036 31368 48044 31396
rect 25573 31331 25631 31337
rect 25666 31331 25724 31337
rect 25516 31303 25585 31331
rect 24762 31260 24768 31272
rect 22152 31232 22197 31260
rect 23216 31232 24624 31260
rect 24723 31232 24768 31260
rect 22152 31220 22158 31232
rect 22738 31192 22744 31204
rect 21100 31164 22744 31192
rect 22738 31152 22744 31164
rect 22796 31192 22802 31204
rect 23290 31192 23296 31204
rect 22796 31164 23296 31192
rect 22796 31152 22802 31164
rect 23290 31152 23296 31164
rect 23348 31152 23354 31204
rect 24596 31192 24624 31232
rect 24762 31220 24768 31232
rect 24820 31220 24826 31272
rect 25516 31260 25544 31303
rect 25573 31297 25585 31303
rect 25619 31300 25636 31331
rect 25619 31297 25631 31300
rect 25573 31291 25631 31297
rect 25666 31297 25678 31331
rect 25712 31297 25724 31331
rect 25666 31291 25724 31297
rect 25774 31288 25780 31340
rect 25832 31337 25838 31340
rect 25832 31328 25840 31337
rect 25832 31300 25877 31328
rect 25832 31291 25840 31300
rect 25832 31288 25838 31291
rect 25958 31288 25964 31340
rect 26016 31328 26022 31340
rect 26016 31300 26061 31328
rect 26016 31288 26022 31300
rect 27890 31288 27896 31340
rect 27948 31328 27954 31340
rect 27985 31331 28043 31337
rect 27985 31328 27997 31331
rect 27948 31300 27997 31328
rect 27948 31288 27954 31300
rect 27985 31297 27997 31300
rect 28031 31297 28043 31331
rect 27985 31291 28043 31297
rect 28810 31288 28816 31340
rect 28868 31328 28874 31340
rect 29457 31331 29515 31337
rect 29457 31328 29469 31331
rect 28868 31300 29469 31328
rect 28868 31288 28874 31300
rect 29457 31297 29469 31300
rect 29503 31297 29515 31331
rect 30466 31328 30472 31340
rect 30427 31300 30472 31328
rect 29457 31291 29515 31297
rect 30466 31288 30472 31300
rect 30524 31288 30530 31340
rect 30650 31328 30656 31340
rect 30611 31300 30656 31328
rect 30650 31288 30656 31300
rect 30708 31288 30714 31340
rect 31036 31260 31064 31368
rect 48038 31356 48044 31368
rect 48096 31356 48102 31408
rect 32122 31328 32128 31340
rect 32083 31300 32128 31328
rect 32122 31288 32128 31300
rect 32180 31288 32186 31340
rect 32309 31331 32367 31337
rect 32309 31297 32321 31331
rect 32355 31297 32367 31331
rect 32309 31291 32367 31297
rect 25516 31232 31064 31260
rect 31202 31220 31208 31272
rect 31260 31260 31266 31272
rect 32324 31260 32352 31291
rect 35894 31288 35900 31340
rect 35952 31328 35958 31340
rect 35989 31331 36047 31337
rect 35989 31328 36001 31331
rect 35952 31300 36001 31328
rect 35952 31288 35958 31300
rect 35989 31297 36001 31300
rect 36035 31297 36047 31331
rect 35989 31291 36047 31297
rect 31260 31232 32352 31260
rect 31260 31220 31266 31232
rect 30466 31192 30472 31204
rect 23400 31164 24532 31192
rect 24596 31164 30472 31192
rect 23400 31136 23428 31164
rect 11756 31096 12296 31124
rect 12345 31127 12403 31133
rect 11756 31084 11762 31096
rect 12345 31093 12357 31127
rect 12391 31124 12403 31127
rect 12710 31124 12716 31136
rect 12391 31096 12716 31124
rect 12391 31093 12403 31096
rect 12345 31087 12403 31093
rect 12710 31084 12716 31096
rect 12768 31084 12774 31136
rect 14274 31124 14280 31136
rect 14235 31096 14280 31124
rect 14274 31084 14280 31096
rect 14332 31084 14338 31136
rect 21177 31127 21235 31133
rect 21177 31093 21189 31127
rect 21223 31124 21235 31127
rect 21634 31124 21640 31136
rect 21223 31096 21640 31124
rect 21223 31093 21235 31096
rect 21177 31087 21235 31093
rect 21634 31084 21640 31096
rect 21692 31084 21698 31136
rect 23382 31084 23388 31136
rect 23440 31084 23446 31136
rect 24121 31127 24179 31133
rect 24121 31093 24133 31127
rect 24167 31124 24179 31127
rect 24394 31124 24400 31136
rect 24167 31096 24400 31124
rect 24167 31093 24179 31096
rect 24121 31087 24179 31093
rect 24394 31084 24400 31096
rect 24452 31084 24458 31136
rect 24504 31124 24532 31164
rect 30466 31152 30472 31164
rect 30524 31152 30530 31204
rect 27154 31124 27160 31136
rect 24504 31096 27160 31124
rect 27154 31084 27160 31096
rect 27212 31084 27218 31136
rect 28810 31124 28816 31136
rect 28771 31096 28816 31124
rect 28810 31084 28816 31096
rect 28868 31084 28874 31136
rect 31294 31084 31300 31136
rect 31352 31124 31358 31136
rect 32493 31127 32551 31133
rect 32493 31124 32505 31127
rect 31352 31096 32505 31124
rect 31352 31084 31358 31096
rect 32493 31093 32505 31096
rect 32539 31093 32551 31127
rect 32493 31087 32551 31093
rect 1104 31034 48852 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 48852 31034
rect 1104 30960 48852 30982
rect 1946 30880 1952 30932
rect 2004 30920 2010 30932
rect 2225 30923 2283 30929
rect 2225 30920 2237 30923
rect 2004 30892 2237 30920
rect 2004 30880 2010 30892
rect 2225 30889 2237 30892
rect 2271 30889 2283 30923
rect 2866 30920 2872 30932
rect 2827 30892 2872 30920
rect 2225 30883 2283 30889
rect 2866 30880 2872 30892
rect 2924 30880 2930 30932
rect 10410 30920 10416 30932
rect 10371 30892 10416 30920
rect 10410 30880 10416 30892
rect 10468 30880 10474 30932
rect 10502 30880 10508 30932
rect 10560 30920 10566 30932
rect 10597 30923 10655 30929
rect 10597 30920 10609 30923
rect 10560 30892 10609 30920
rect 10560 30880 10566 30892
rect 10597 30889 10609 30892
rect 10643 30920 10655 30923
rect 10962 30920 10968 30932
rect 10643 30892 10968 30920
rect 10643 30889 10655 30892
rect 10597 30883 10655 30889
rect 10962 30880 10968 30892
rect 11020 30880 11026 30932
rect 12989 30923 13047 30929
rect 12989 30889 13001 30923
rect 13035 30920 13047 30923
rect 13630 30920 13636 30932
rect 13035 30892 13636 30920
rect 13035 30889 13047 30892
rect 12989 30883 13047 30889
rect 13630 30880 13636 30892
rect 13688 30880 13694 30932
rect 14277 30923 14335 30929
rect 14277 30889 14289 30923
rect 14323 30920 14335 30923
rect 15194 30920 15200 30932
rect 14323 30892 15200 30920
rect 14323 30889 14335 30892
rect 14277 30883 14335 30889
rect 15194 30880 15200 30892
rect 15252 30880 15258 30932
rect 16485 30923 16543 30929
rect 16485 30889 16497 30923
rect 16531 30920 16543 30923
rect 16758 30920 16764 30932
rect 16531 30892 16764 30920
rect 16531 30889 16543 30892
rect 16485 30883 16543 30889
rect 16758 30880 16764 30892
rect 16816 30880 16822 30932
rect 24670 30880 24676 30932
rect 24728 30920 24734 30932
rect 26789 30923 26847 30929
rect 26789 30920 26801 30923
rect 24728 30892 26801 30920
rect 24728 30880 24734 30892
rect 26789 30889 26801 30892
rect 26835 30889 26847 30923
rect 30466 30920 30472 30932
rect 30427 30892 30472 30920
rect 26789 30883 26847 30889
rect 30466 30880 30472 30892
rect 30524 30880 30530 30932
rect 35986 30880 35992 30932
rect 36044 30920 36050 30932
rect 36081 30923 36139 30929
rect 36081 30920 36093 30923
rect 36044 30892 36093 30920
rect 36044 30880 36050 30892
rect 36081 30889 36093 30892
rect 36127 30889 36139 30923
rect 36081 30883 36139 30889
rect 11054 30812 11060 30864
rect 11112 30852 11118 30864
rect 12066 30852 12072 30864
rect 11112 30824 12072 30852
rect 11112 30812 11118 30824
rect 12066 30812 12072 30824
rect 12124 30812 12130 30864
rect 14366 30812 14372 30864
rect 14424 30852 14430 30864
rect 14918 30852 14924 30864
rect 14424 30824 14924 30852
rect 14424 30812 14430 30824
rect 14918 30812 14924 30824
rect 14976 30812 14982 30864
rect 15286 30852 15292 30864
rect 15247 30824 15292 30852
rect 15286 30812 15292 30824
rect 15344 30812 15350 30864
rect 16574 30812 16580 30864
rect 16632 30852 16638 30864
rect 17497 30855 17555 30861
rect 17497 30852 17509 30855
rect 16632 30824 17509 30852
rect 16632 30812 16638 30824
rect 17497 30821 17509 30824
rect 17543 30821 17555 30855
rect 17497 30815 17555 30821
rect 31294 30812 31300 30864
rect 31352 30812 31358 30864
rect 18233 30787 18291 30793
rect 18233 30784 18245 30787
rect 15120 30756 18245 30784
rect 2777 30719 2835 30725
rect 2777 30685 2789 30719
rect 2823 30716 2835 30719
rect 7650 30716 7656 30728
rect 2823 30688 7656 30716
rect 2823 30685 2835 30688
rect 2777 30679 2835 30685
rect 7650 30676 7656 30688
rect 7708 30676 7714 30728
rect 10778 30676 10784 30728
rect 10836 30716 10842 30728
rect 11057 30719 11115 30725
rect 11057 30716 11069 30719
rect 10836 30688 11069 30716
rect 10836 30676 10842 30688
rect 11057 30685 11069 30688
rect 11103 30685 11115 30719
rect 11057 30679 11115 30685
rect 11333 30719 11391 30725
rect 11333 30685 11345 30719
rect 11379 30685 11391 30719
rect 11333 30679 11391 30685
rect 10229 30651 10287 30657
rect 10229 30617 10241 30651
rect 10275 30648 10287 30651
rect 11348 30648 11376 30679
rect 12158 30676 12164 30728
rect 12216 30716 12222 30728
rect 12621 30719 12679 30725
rect 12621 30716 12633 30719
rect 12216 30688 12633 30716
rect 12216 30676 12222 30688
rect 11606 30648 11612 30660
rect 10275 30620 11612 30648
rect 10275 30617 10287 30620
rect 10229 30611 10287 30617
rect 11606 30608 11612 30620
rect 11664 30648 11670 30660
rect 11790 30648 11796 30660
rect 11664 30620 11796 30648
rect 11664 30608 11670 30620
rect 11790 30608 11796 30620
rect 11848 30608 11854 30660
rect 10439 30583 10497 30589
rect 10439 30549 10451 30583
rect 10485 30580 10497 30583
rect 11974 30580 11980 30592
rect 10485 30552 11980 30580
rect 10485 30549 10497 30552
rect 10439 30543 10497 30549
rect 11974 30540 11980 30552
rect 12032 30540 12038 30592
rect 12342 30580 12348 30592
rect 12303 30552 12348 30580
rect 12342 30540 12348 30552
rect 12400 30540 12406 30592
rect 12544 30580 12572 30688
rect 12621 30685 12633 30688
rect 12667 30685 12679 30719
rect 12802 30716 12808 30728
rect 12763 30688 12808 30716
rect 12621 30679 12679 30685
rect 12802 30676 12808 30688
rect 12860 30676 12866 30728
rect 13078 30716 13084 30728
rect 13039 30688 13084 30716
rect 13078 30676 13084 30688
rect 13136 30676 13142 30728
rect 13354 30676 13360 30728
rect 13412 30716 13418 30728
rect 14185 30719 14243 30725
rect 14185 30716 14197 30719
rect 13412 30688 14197 30716
rect 13412 30676 13418 30688
rect 14185 30685 14197 30688
rect 14231 30716 14243 30719
rect 14366 30716 14372 30728
rect 14231 30688 14372 30716
rect 14231 30685 14243 30688
rect 14185 30679 14243 30685
rect 14366 30676 14372 30688
rect 14424 30676 14430 30728
rect 15120 30725 15148 30756
rect 18233 30753 18245 30756
rect 18279 30784 18291 30787
rect 18414 30784 18420 30796
rect 18279 30756 18420 30784
rect 18279 30753 18291 30756
rect 18233 30747 18291 30753
rect 18414 30744 18420 30756
rect 18472 30744 18478 30796
rect 21177 30787 21235 30793
rect 21177 30784 21189 30787
rect 20180 30756 21189 30784
rect 20180 30728 20208 30756
rect 21177 30753 21189 30756
rect 21223 30753 21235 30787
rect 22922 30784 22928 30796
rect 22883 30756 22928 30784
rect 21177 30747 21235 30753
rect 22922 30744 22928 30756
rect 22980 30744 22986 30796
rect 24026 30744 24032 30796
rect 24084 30784 24090 30796
rect 27706 30784 27712 30796
rect 24084 30756 25544 30784
rect 24084 30744 24090 30756
rect 25516 30728 25544 30756
rect 27540 30756 27712 30784
rect 15105 30719 15163 30725
rect 15105 30685 15117 30719
rect 15151 30685 15163 30719
rect 16666 30716 16672 30728
rect 16627 30688 16672 30716
rect 15105 30679 15163 30685
rect 16666 30676 16672 30688
rect 16724 30676 16730 30728
rect 16758 30676 16764 30728
rect 16816 30716 16822 30728
rect 17129 30719 17187 30725
rect 17129 30716 17141 30719
rect 16816 30688 17141 30716
rect 16816 30676 16822 30688
rect 17129 30685 17141 30688
rect 17175 30685 17187 30719
rect 17129 30679 17187 30685
rect 17954 30676 17960 30728
rect 18012 30716 18018 30728
rect 18049 30719 18107 30725
rect 18049 30716 18061 30719
rect 18012 30688 18061 30716
rect 18012 30676 18018 30688
rect 18049 30685 18061 30688
rect 18095 30685 18107 30719
rect 18049 30679 18107 30685
rect 19705 30719 19763 30725
rect 19705 30685 19717 30719
rect 19751 30716 19763 30719
rect 20162 30716 20168 30728
rect 19751 30688 20168 30716
rect 19751 30685 19763 30688
rect 19705 30679 19763 30685
rect 20162 30676 20168 30688
rect 20220 30676 20226 30728
rect 20901 30719 20959 30725
rect 20901 30685 20913 30719
rect 20947 30716 20959 30719
rect 21910 30716 21916 30728
rect 20947 30688 21916 30716
rect 20947 30685 20959 30688
rect 20901 30679 20959 30685
rect 21910 30676 21916 30688
rect 21968 30676 21974 30728
rect 22462 30676 22468 30728
rect 22520 30716 22526 30728
rect 22649 30719 22707 30725
rect 22649 30716 22661 30719
rect 22520 30688 22661 30716
rect 22520 30676 22526 30688
rect 22649 30685 22661 30688
rect 22695 30716 22707 30719
rect 23382 30716 23388 30728
rect 22695 30688 23388 30716
rect 22695 30685 22707 30688
rect 22649 30679 22707 30685
rect 23382 30676 23388 30688
rect 23440 30676 23446 30728
rect 24394 30716 24400 30728
rect 24355 30688 24400 30716
rect 24394 30676 24400 30688
rect 24452 30676 24458 30728
rect 25406 30716 25412 30728
rect 25367 30688 25412 30716
rect 25406 30676 25412 30688
rect 25464 30676 25470 30728
rect 25498 30676 25504 30728
rect 25556 30716 25562 30728
rect 25958 30716 25964 30728
rect 25556 30688 25964 30716
rect 25556 30676 25562 30688
rect 25958 30676 25964 30688
rect 26016 30676 26022 30728
rect 27540 30725 27568 30756
rect 27706 30744 27712 30756
rect 27764 30744 27770 30796
rect 31018 30784 31024 30796
rect 28920 30756 31024 30784
rect 27525 30719 27583 30725
rect 27525 30685 27537 30719
rect 27571 30685 27583 30719
rect 27525 30679 27583 30685
rect 27890 30676 27896 30728
rect 27948 30716 27954 30728
rect 28261 30719 28319 30725
rect 28261 30716 28273 30719
rect 27948 30688 28273 30716
rect 27948 30676 27954 30688
rect 28261 30685 28273 30688
rect 28307 30685 28319 30719
rect 28261 30679 28319 30685
rect 12710 30648 12716 30660
rect 12671 30620 12716 30648
rect 12710 30608 12716 30620
rect 12768 30608 12774 30660
rect 17313 30651 17371 30657
rect 17313 30617 17325 30651
rect 17359 30648 17371 30651
rect 18690 30648 18696 30660
rect 17359 30620 18696 30648
rect 17359 30617 17371 30620
rect 17313 30611 17371 30617
rect 18690 30608 18696 30620
rect 18748 30608 18754 30660
rect 23474 30608 23480 30660
rect 23532 30648 23538 30660
rect 24578 30648 24584 30660
rect 23532 30620 24584 30648
rect 23532 30608 23538 30620
rect 24578 30608 24584 30620
rect 24636 30608 24642 30660
rect 24854 30608 24860 30660
rect 24912 30648 24918 30660
rect 25654 30651 25712 30657
rect 25654 30648 25666 30651
rect 24912 30620 25666 30648
rect 24912 30608 24918 30620
rect 25654 30617 25666 30620
rect 25700 30617 25712 30651
rect 28920 30648 28948 30756
rect 31018 30744 31024 30756
rect 31076 30784 31082 30796
rect 31076 30756 31248 30784
rect 31076 30744 31082 30756
rect 30466 30676 30472 30728
rect 30524 30716 30530 30728
rect 31220 30725 31248 30756
rect 31312 30725 31340 30812
rect 31404 30756 31754 30784
rect 31113 30719 31171 30725
rect 31113 30716 31125 30719
rect 30524 30688 31125 30716
rect 30524 30676 30530 30688
rect 31113 30685 31125 30688
rect 31159 30685 31171 30719
rect 31113 30679 31171 30685
rect 31205 30719 31263 30725
rect 31205 30685 31217 30719
rect 31251 30685 31263 30719
rect 31205 30679 31263 30685
rect 31297 30719 31355 30725
rect 31297 30685 31309 30719
rect 31343 30685 31355 30719
rect 31297 30679 31355 30685
rect 25654 30611 25712 30617
rect 27632 30620 28948 30648
rect 30837 30651 30895 30657
rect 13170 30580 13176 30592
rect 12544 30552 13176 30580
rect 13170 30540 13176 30552
rect 13228 30540 13234 30592
rect 17218 30540 17224 30592
rect 17276 30580 17282 30592
rect 19797 30583 19855 30589
rect 19797 30580 19809 30583
rect 17276 30552 19809 30580
rect 17276 30540 17282 30552
rect 19797 30549 19809 30552
rect 19843 30549 19855 30583
rect 19797 30543 19855 30549
rect 24765 30583 24823 30589
rect 24765 30549 24777 30583
rect 24811 30580 24823 30583
rect 25314 30580 25320 30592
rect 24811 30552 25320 30580
rect 24811 30549 24823 30552
rect 24765 30543 24823 30549
rect 25314 30540 25320 30552
rect 25372 30540 25378 30592
rect 26694 30540 26700 30592
rect 26752 30580 26758 30592
rect 27522 30580 27528 30592
rect 26752 30552 27528 30580
rect 26752 30540 26758 30552
rect 27522 30540 27528 30552
rect 27580 30580 27586 30592
rect 27632 30589 27660 30620
rect 30837 30617 30849 30651
rect 30883 30648 30895 30651
rect 31404 30648 31432 30756
rect 31481 30719 31539 30725
rect 31481 30685 31493 30719
rect 31527 30685 31539 30719
rect 31481 30679 31539 30685
rect 30883 30620 31432 30648
rect 30883 30617 30895 30620
rect 30837 30611 30895 30617
rect 27617 30583 27675 30589
rect 27617 30580 27629 30583
rect 27580 30552 27629 30580
rect 27580 30540 27586 30552
rect 27617 30549 27629 30552
rect 27663 30549 27675 30583
rect 27617 30543 27675 30549
rect 28166 30540 28172 30592
rect 28224 30580 28230 30592
rect 28353 30583 28411 30589
rect 28353 30580 28365 30583
rect 28224 30552 28365 30580
rect 28224 30540 28230 30552
rect 28353 30549 28365 30552
rect 28399 30580 28411 30583
rect 31496 30580 31524 30679
rect 31726 30648 31754 30756
rect 31938 30716 31944 30728
rect 31899 30688 31944 30716
rect 31938 30676 31944 30688
rect 31996 30676 32002 30728
rect 34701 30719 34759 30725
rect 34701 30685 34713 30719
rect 34747 30716 34759 30719
rect 35342 30716 35348 30728
rect 34747 30688 35348 30716
rect 34747 30685 34759 30688
rect 34701 30679 34759 30685
rect 35342 30676 35348 30688
rect 35400 30676 35406 30728
rect 32186 30651 32244 30657
rect 32186 30648 32198 30651
rect 31726 30620 32198 30648
rect 32186 30617 32198 30620
rect 32232 30617 32244 30651
rect 32186 30611 32244 30617
rect 34514 30608 34520 30660
rect 34572 30648 34578 30660
rect 34946 30651 35004 30657
rect 34946 30648 34958 30651
rect 34572 30620 34958 30648
rect 34572 30608 34578 30620
rect 34946 30617 34958 30620
rect 34992 30617 35004 30651
rect 34946 30611 35004 30617
rect 32306 30580 32312 30592
rect 28399 30552 32312 30580
rect 28399 30549 28411 30552
rect 28353 30543 28411 30549
rect 32306 30540 32312 30552
rect 32364 30540 32370 30592
rect 33318 30580 33324 30592
rect 33279 30552 33324 30580
rect 33318 30540 33324 30552
rect 33376 30540 33382 30592
rect 1104 30490 48852 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 48852 30490
rect 1104 30416 48852 30438
rect 11790 30376 11796 30388
rect 11751 30348 11796 30376
rect 11790 30336 11796 30348
rect 11848 30336 11854 30388
rect 12250 30336 12256 30388
rect 12308 30376 12314 30388
rect 13357 30379 13415 30385
rect 13357 30376 13369 30379
rect 12308 30348 13369 30376
rect 12308 30336 12314 30348
rect 13357 30345 13369 30348
rect 13403 30345 13415 30379
rect 14366 30376 14372 30388
rect 14327 30348 14372 30376
rect 13357 30339 13415 30345
rect 9674 30268 9680 30320
rect 9732 30308 9738 30320
rect 10597 30311 10655 30317
rect 10597 30308 10609 30311
rect 9732 30280 10609 30308
rect 9732 30268 9738 30280
rect 10597 30277 10609 30280
rect 10643 30277 10655 30311
rect 11609 30311 11667 30317
rect 11609 30308 11621 30311
rect 10597 30271 10655 30277
rect 10704 30280 11621 30308
rect 10502 30240 10508 30252
rect 10463 30212 10508 30240
rect 10502 30200 10508 30212
rect 10560 30200 10566 30252
rect 10704 30249 10732 30280
rect 11609 30277 11621 30280
rect 11655 30308 11667 30311
rect 11698 30308 11704 30320
rect 11655 30280 11704 30308
rect 11655 30277 11667 30280
rect 11609 30271 11667 30277
rect 11698 30268 11704 30280
rect 11756 30268 11762 30320
rect 12066 30268 12072 30320
rect 12124 30308 12130 30320
rect 12161 30311 12219 30317
rect 12161 30308 12173 30311
rect 12124 30280 12173 30308
rect 12124 30268 12130 30280
rect 12161 30277 12173 30280
rect 12207 30277 12219 30311
rect 13262 30308 13268 30320
rect 13223 30280 13268 30308
rect 12161 30271 12219 30277
rect 13262 30268 13268 30280
rect 13320 30268 13326 30320
rect 13372 30308 13400 30339
rect 14366 30336 14372 30348
rect 14424 30336 14430 30388
rect 19334 30336 19340 30388
rect 19392 30376 19398 30388
rect 20438 30376 20444 30388
rect 19392 30348 20444 30376
rect 19392 30336 19398 30348
rect 20438 30336 20444 30348
rect 20496 30336 20502 30388
rect 20898 30336 20904 30388
rect 20956 30376 20962 30388
rect 21177 30379 21235 30385
rect 21177 30376 21189 30379
rect 20956 30348 21189 30376
rect 20956 30336 20962 30348
rect 21177 30345 21189 30348
rect 21223 30345 21235 30379
rect 21177 30339 21235 30345
rect 22922 30336 22928 30388
rect 22980 30336 22986 30388
rect 24026 30336 24032 30388
rect 24084 30376 24090 30388
rect 24302 30376 24308 30388
rect 24084 30348 24308 30376
rect 24084 30336 24090 30348
rect 24302 30336 24308 30348
rect 24360 30336 24366 30388
rect 24854 30376 24860 30388
rect 24815 30348 24860 30376
rect 24854 30336 24860 30348
rect 24912 30336 24918 30388
rect 27982 30336 27988 30388
rect 28040 30336 28046 30388
rect 32122 30376 32128 30388
rect 32083 30348 32128 30376
rect 32122 30336 32128 30348
rect 32180 30336 32186 30388
rect 13372 30280 15240 30308
rect 10689 30243 10747 30249
rect 10689 30209 10701 30243
rect 10735 30209 10747 30243
rect 10689 30203 10747 30209
rect 11885 30243 11943 30249
rect 11885 30209 11897 30243
rect 11931 30209 11943 30243
rect 11885 30203 11943 30209
rect 11977 30243 12035 30249
rect 11977 30209 11989 30243
rect 12023 30240 12035 30243
rect 12526 30240 12532 30252
rect 12023 30238 12388 30240
rect 12421 30238 12532 30240
rect 12023 30212 12532 30238
rect 12023 30209 12035 30212
rect 12360 30210 12449 30212
rect 11977 30203 12035 30209
rect 1946 30172 1952 30184
rect 1907 30144 1952 30172
rect 1946 30132 1952 30144
rect 2004 30132 2010 30184
rect 2133 30175 2191 30181
rect 2133 30141 2145 30175
rect 2179 30172 2191 30175
rect 2774 30172 2780 30184
rect 2179 30144 2780 30172
rect 2179 30141 2191 30144
rect 2133 30135 2191 30141
rect 2774 30132 2780 30144
rect 2832 30132 2838 30184
rect 2866 30132 2872 30184
rect 2924 30172 2930 30184
rect 2924 30144 2969 30172
rect 2924 30132 2930 30144
rect 10226 30132 10232 30184
rect 10284 30172 10290 30184
rect 10704 30172 10732 30203
rect 10284 30144 10732 30172
rect 11900 30172 11928 30203
rect 12526 30200 12532 30212
rect 12584 30200 12590 30252
rect 14366 30240 14372 30252
rect 14327 30212 14372 30240
rect 14366 30200 14372 30212
rect 14424 30200 14430 30252
rect 15212 30249 15240 30280
rect 19518 30268 19524 30320
rect 19576 30308 19582 30320
rect 22940 30308 22968 30336
rect 25038 30308 25044 30320
rect 19576 30280 20300 30308
rect 22940 30280 25044 30308
rect 19576 30268 19582 30280
rect 15197 30243 15255 30249
rect 15197 30209 15209 30243
rect 15243 30240 15255 30243
rect 16022 30240 16028 30252
rect 15243 30212 16028 30240
rect 15243 30209 15255 30212
rect 15197 30203 15255 30209
rect 16022 30200 16028 30212
rect 16080 30200 16086 30252
rect 17034 30200 17040 30252
rect 17092 30240 17098 30252
rect 17405 30243 17463 30249
rect 17405 30240 17417 30243
rect 17092 30212 17417 30240
rect 17092 30200 17098 30212
rect 17405 30209 17417 30212
rect 17451 30209 17463 30243
rect 19702 30240 19708 30252
rect 19663 30212 19708 30240
rect 17405 30203 17463 30209
rect 19702 30200 19708 30212
rect 19760 30200 19766 30252
rect 19889 30243 19947 30249
rect 19889 30209 19901 30243
rect 19935 30240 19947 30243
rect 20162 30240 20168 30252
rect 19935 30212 20168 30240
rect 19935 30209 19947 30212
rect 19889 30203 19947 30209
rect 20162 30200 20168 30212
rect 20220 30200 20226 30252
rect 20272 30249 20300 30280
rect 20257 30243 20315 30249
rect 20257 30209 20269 30243
rect 20303 30209 20315 30243
rect 20257 30203 20315 30209
rect 20993 30243 21051 30249
rect 20993 30209 21005 30243
rect 21039 30209 21051 30243
rect 20993 30203 21051 30209
rect 21821 30243 21879 30249
rect 21821 30209 21833 30243
rect 21867 30240 21879 30243
rect 21910 30240 21916 30252
rect 21867 30212 21916 30240
rect 21867 30209 21879 30212
rect 21821 30203 21879 30209
rect 12250 30172 12256 30184
rect 11900 30144 12256 30172
rect 10284 30132 10290 30144
rect 12250 30132 12256 30144
rect 12308 30132 12314 30184
rect 14182 30172 14188 30184
rect 14143 30144 14188 30172
rect 14182 30132 14188 30144
rect 14240 30132 14246 30184
rect 14737 30175 14795 30181
rect 14737 30141 14749 30175
rect 14783 30172 14795 30175
rect 16666 30172 16672 30184
rect 14783 30144 16672 30172
rect 14783 30141 14795 30144
rect 14737 30135 14795 30141
rect 11716 30076 13952 30104
rect 8938 29996 8944 30048
rect 8996 30036 9002 30048
rect 11716 30036 11744 30076
rect 8996 30008 11744 30036
rect 13924 30036 13952 30076
rect 14752 30036 14780 30135
rect 16666 30132 16672 30144
rect 16724 30132 16730 30184
rect 17129 30175 17187 30181
rect 17129 30141 17141 30175
rect 17175 30172 17187 30175
rect 17494 30172 17500 30184
rect 17175 30144 17500 30172
rect 17175 30141 17187 30144
rect 17129 30135 17187 30141
rect 17494 30132 17500 30144
rect 17552 30132 17558 30184
rect 19978 30172 19984 30184
rect 19939 30144 19984 30172
rect 19978 30132 19984 30144
rect 20036 30132 20042 30184
rect 20073 30175 20131 30181
rect 20073 30141 20085 30175
rect 20119 30172 20131 30175
rect 20898 30172 20904 30184
rect 20119 30144 20904 30172
rect 20119 30141 20131 30144
rect 20073 30135 20131 30141
rect 20898 30132 20904 30144
rect 20956 30132 20962 30184
rect 21008 30172 21036 30203
rect 21910 30200 21916 30212
rect 21968 30200 21974 30252
rect 22925 30243 22983 30249
rect 22925 30209 22937 30243
rect 22971 30240 22983 30243
rect 23198 30240 23204 30252
rect 22971 30212 23204 30240
rect 22971 30209 22983 30212
rect 22925 30203 22983 30209
rect 23198 30200 23204 30212
rect 23256 30240 23262 30252
rect 23474 30240 23480 30252
rect 23256 30212 23480 30240
rect 23256 30200 23262 30212
rect 23474 30200 23480 30212
rect 23532 30200 23538 30252
rect 24044 30249 24072 30280
rect 25038 30268 25044 30280
rect 25096 30308 25102 30320
rect 26050 30308 26056 30320
rect 25096 30280 25268 30308
rect 26011 30280 26056 30308
rect 25096 30268 25102 30280
rect 23937 30243 23995 30249
rect 23937 30209 23949 30243
rect 23983 30209 23995 30243
rect 23937 30203 23995 30209
rect 24029 30243 24087 30249
rect 24029 30209 24041 30243
rect 24075 30209 24087 30243
rect 24029 30203 24087 30209
rect 22462 30172 22468 30184
rect 21008 30144 22468 30172
rect 22462 30132 22468 30144
rect 22520 30132 22526 30184
rect 23952 30172 23980 30203
rect 24118 30200 24124 30252
rect 24176 30240 24182 30252
rect 24176 30212 24221 30240
rect 24176 30200 24182 30212
rect 24302 30200 24308 30252
rect 24360 30240 24366 30252
rect 25240 30249 25268 30280
rect 26050 30268 26056 30280
rect 26108 30268 26114 30320
rect 28000 30308 28028 30336
rect 28782 30311 28840 30317
rect 28782 30308 28794 30311
rect 28000 30280 28794 30308
rect 28782 30277 28794 30280
rect 28828 30277 28840 30311
rect 28782 30271 28840 30277
rect 29822 30268 29828 30320
rect 29880 30308 29886 30320
rect 30469 30311 30527 30317
rect 30469 30308 30481 30311
rect 29880 30280 30481 30308
rect 29880 30268 29886 30280
rect 30469 30277 30481 30280
rect 30515 30277 30527 30311
rect 32582 30308 32588 30320
rect 32543 30280 32588 30308
rect 30469 30271 30527 30277
rect 32582 30268 32588 30280
rect 32640 30268 32646 30320
rect 33042 30268 33048 30320
rect 33100 30308 33106 30320
rect 34885 30311 34943 30317
rect 33100 30280 33916 30308
rect 33100 30268 33106 30280
rect 25133 30243 25191 30249
rect 24360 30212 24405 30240
rect 24360 30200 24366 30212
rect 25133 30209 25145 30243
rect 25179 30209 25191 30243
rect 25133 30203 25191 30209
rect 25225 30243 25283 30249
rect 25225 30209 25237 30243
rect 25271 30209 25283 30243
rect 25225 30203 25283 30209
rect 25038 30172 25044 30184
rect 23952 30144 25044 30172
rect 25038 30132 25044 30144
rect 25096 30132 25102 30184
rect 25148 30172 25176 30203
rect 25314 30200 25320 30252
rect 25372 30240 25378 30252
rect 25372 30212 25417 30240
rect 25372 30200 25378 30212
rect 25498 30200 25504 30252
rect 25556 30240 25562 30252
rect 25556 30212 25601 30240
rect 25556 30200 25562 30212
rect 27614 30200 27620 30252
rect 27672 30243 27678 30252
rect 27914 30249 27972 30255
rect 27709 30243 27767 30249
rect 27672 30215 27721 30243
rect 27672 30200 27678 30215
rect 27709 30209 27721 30215
rect 27755 30209 27767 30243
rect 27709 30203 27767 30209
rect 27814 30243 27872 30249
rect 27814 30209 27826 30243
rect 27860 30209 27872 30243
rect 27914 30215 27926 30249
rect 27960 30246 27972 30249
rect 27960 30218 28028 30246
rect 27960 30215 27972 30218
rect 27914 30209 27972 30215
rect 27814 30203 27872 30209
rect 25774 30172 25780 30184
rect 25148 30144 25780 30172
rect 25774 30132 25780 30144
rect 25832 30132 25838 30184
rect 26237 30175 26295 30181
rect 26237 30141 26249 30175
rect 26283 30172 26295 30175
rect 26326 30172 26332 30184
rect 26283 30144 26332 30172
rect 26283 30141 26295 30144
rect 26237 30135 26295 30141
rect 26326 30132 26332 30144
rect 26384 30132 26390 30184
rect 27522 30132 27528 30184
rect 27580 30172 27586 30184
rect 27829 30172 27857 30203
rect 27580 30144 27857 30172
rect 27580 30132 27586 30144
rect 21818 30064 21824 30116
rect 21876 30104 21882 30116
rect 22005 30107 22063 30113
rect 22005 30104 22017 30107
rect 21876 30076 22017 30104
rect 21876 30064 21882 30076
rect 22005 30073 22017 30076
rect 22051 30073 22063 30107
rect 22005 30067 22063 30073
rect 27798 30064 27804 30116
rect 27856 30104 27862 30116
rect 28000 30104 28028 30218
rect 28077 30243 28135 30249
rect 28077 30209 28089 30243
rect 28123 30240 28135 30243
rect 28166 30240 28172 30252
rect 28123 30212 28172 30240
rect 28123 30209 28135 30212
rect 28077 30203 28135 30209
rect 28166 30200 28172 30212
rect 28224 30200 28230 30252
rect 32493 30243 32551 30249
rect 32493 30209 32505 30243
rect 32539 30240 32551 30243
rect 33318 30240 33324 30252
rect 32539 30212 33324 30240
rect 32539 30209 32551 30212
rect 32493 30203 32551 30209
rect 33318 30200 33324 30212
rect 33376 30240 33382 30252
rect 33888 30249 33916 30280
rect 34885 30277 34897 30311
rect 34931 30308 34943 30311
rect 35986 30308 35992 30320
rect 34931 30280 35992 30308
rect 34931 30277 34943 30280
rect 34885 30271 34943 30277
rect 35986 30268 35992 30280
rect 36044 30268 36050 30320
rect 33873 30243 33931 30249
rect 33376 30212 33824 30240
rect 33376 30200 33382 30212
rect 28534 30172 28540 30184
rect 28495 30144 28540 30172
rect 28534 30132 28540 30144
rect 28592 30132 28598 30184
rect 32769 30175 32827 30181
rect 32769 30141 32781 30175
rect 32815 30172 32827 30175
rect 33502 30172 33508 30184
rect 32815 30144 33508 30172
rect 32815 30141 32827 30144
rect 32769 30135 32827 30141
rect 33502 30132 33508 30144
rect 33560 30132 33566 30184
rect 33796 30172 33824 30212
rect 33873 30209 33885 30243
rect 33919 30209 33931 30243
rect 33873 30203 33931 30209
rect 33965 30243 34023 30249
rect 33965 30209 33977 30243
rect 34011 30209 34023 30243
rect 33965 30203 34023 30209
rect 34057 30243 34115 30249
rect 34057 30209 34069 30243
rect 34103 30209 34115 30243
rect 34057 30203 34115 30209
rect 34241 30243 34299 30249
rect 34241 30209 34253 30243
rect 34287 30209 34299 30243
rect 34241 30203 34299 30209
rect 33980 30172 34008 30203
rect 33796 30144 34008 30172
rect 29914 30104 29920 30116
rect 27856 30076 28028 30104
rect 29875 30076 29920 30104
rect 27856 30064 27862 30076
rect 29914 30064 29920 30076
rect 29972 30064 29978 30116
rect 30098 30064 30104 30116
rect 30156 30104 30162 30116
rect 34072 30104 34100 30203
rect 34256 30172 34284 30203
rect 34606 30200 34612 30252
rect 34664 30240 34670 30252
rect 35069 30243 35127 30249
rect 35069 30240 35081 30243
rect 34664 30212 35081 30240
rect 34664 30200 34670 30212
rect 35069 30209 35081 30212
rect 35115 30209 35127 30243
rect 35069 30203 35127 30209
rect 35253 30175 35311 30181
rect 35253 30172 35265 30175
rect 34256 30144 35265 30172
rect 35253 30141 35265 30144
rect 35299 30141 35311 30175
rect 35253 30135 35311 30141
rect 30156 30076 34100 30104
rect 30156 30064 30162 30076
rect 35802 30064 35808 30116
rect 35860 30104 35866 30116
rect 46014 30104 46020 30116
rect 35860 30076 46020 30104
rect 35860 30064 35866 30076
rect 46014 30064 46020 30076
rect 46072 30064 46078 30116
rect 13924 30008 14780 30036
rect 8996 29996 9002 30008
rect 15194 29996 15200 30048
rect 15252 30036 15258 30048
rect 15289 30039 15347 30045
rect 15289 30036 15301 30039
rect 15252 30008 15301 30036
rect 15252 29996 15258 30008
rect 15289 30005 15301 30008
rect 15335 30005 15347 30039
rect 15289 29999 15347 30005
rect 16758 29996 16764 30048
rect 16816 30036 16822 30048
rect 17126 30036 17132 30048
rect 16816 30008 17132 30036
rect 16816 29996 16822 30008
rect 17126 29996 17132 30008
rect 17184 29996 17190 30048
rect 20438 30036 20444 30048
rect 20399 30008 20444 30036
rect 20438 29996 20444 30008
rect 20496 29996 20502 30048
rect 20530 29996 20536 30048
rect 20588 30036 20594 30048
rect 22370 30036 22376 30048
rect 20588 30008 22376 30036
rect 20588 29996 20594 30008
rect 22370 29996 22376 30008
rect 22428 30036 22434 30048
rect 23106 30036 23112 30048
rect 22428 30008 23112 30036
rect 22428 29996 22434 30008
rect 23106 29996 23112 30008
rect 23164 29996 23170 30048
rect 23658 30036 23664 30048
rect 23619 30008 23664 30036
rect 23658 29996 23664 30008
rect 23716 29996 23722 30048
rect 23750 29996 23756 30048
rect 23808 30036 23814 30048
rect 25682 30036 25688 30048
rect 23808 30008 25688 30036
rect 23808 29996 23814 30008
rect 25682 29996 25688 30008
rect 25740 29996 25746 30048
rect 27430 30036 27436 30048
rect 27391 30008 27436 30036
rect 27430 29996 27436 30008
rect 27488 29996 27494 30048
rect 30190 29996 30196 30048
rect 30248 30036 30254 30048
rect 30561 30039 30619 30045
rect 30561 30036 30573 30039
rect 30248 30008 30573 30036
rect 30248 29996 30254 30008
rect 30561 30005 30573 30008
rect 30607 30036 30619 30039
rect 33318 30036 33324 30048
rect 30607 30008 33324 30036
rect 30607 30005 30619 30008
rect 30561 29999 30619 30005
rect 33318 29996 33324 30008
rect 33376 29996 33382 30048
rect 33597 30039 33655 30045
rect 33597 30005 33609 30039
rect 33643 30036 33655 30039
rect 34514 30036 34520 30048
rect 33643 30008 34520 30036
rect 33643 30005 33655 30008
rect 33597 29999 33655 30005
rect 34514 29996 34520 30008
rect 34572 29996 34578 30048
rect 1104 29946 48852 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 48852 29946
rect 1104 29872 48852 29894
rect 1946 29792 1952 29844
rect 2004 29832 2010 29844
rect 2225 29835 2283 29841
rect 2225 29832 2237 29835
rect 2004 29804 2237 29832
rect 2004 29792 2010 29804
rect 2225 29801 2237 29804
rect 2271 29801 2283 29835
rect 2225 29795 2283 29801
rect 2774 29792 2780 29844
rect 2832 29832 2838 29844
rect 2869 29835 2927 29841
rect 2869 29832 2881 29835
rect 2832 29804 2881 29832
rect 2832 29792 2838 29804
rect 2869 29801 2881 29804
rect 2915 29801 2927 29835
rect 2869 29795 2927 29801
rect 14182 29792 14188 29844
rect 14240 29832 14246 29844
rect 15102 29832 15108 29844
rect 14240 29804 15108 29832
rect 14240 29792 14246 29804
rect 15102 29792 15108 29804
rect 15160 29832 15166 29844
rect 15289 29835 15347 29841
rect 15289 29832 15301 29835
rect 15160 29804 15301 29832
rect 15160 29792 15166 29804
rect 15289 29801 15301 29804
rect 15335 29801 15347 29835
rect 15289 29795 15347 29801
rect 15841 29835 15899 29841
rect 15841 29801 15853 29835
rect 15887 29832 15899 29835
rect 15930 29832 15936 29844
rect 15887 29804 15936 29832
rect 15887 29801 15899 29804
rect 15841 29795 15899 29801
rect 15930 29792 15936 29804
rect 15988 29792 15994 29844
rect 16574 29792 16580 29844
rect 16632 29832 16638 29844
rect 17218 29832 17224 29844
rect 16632 29804 17224 29832
rect 16632 29792 16638 29804
rect 17218 29792 17224 29804
rect 17276 29832 17282 29844
rect 19337 29835 19395 29841
rect 17276 29804 18552 29832
rect 17276 29792 17282 29804
rect 8938 29764 8944 29776
rect 8036 29736 8944 29764
rect 2777 29631 2835 29637
rect 2777 29597 2789 29631
rect 2823 29628 2835 29631
rect 2866 29628 2872 29640
rect 2823 29600 2872 29628
rect 2823 29597 2835 29600
rect 2777 29591 2835 29597
rect 2866 29588 2872 29600
rect 2924 29588 2930 29640
rect 8036 29637 8064 29736
rect 8938 29724 8944 29736
rect 8996 29724 9002 29776
rect 12526 29724 12532 29776
rect 12584 29764 12590 29776
rect 12584 29736 13400 29764
rect 12584 29724 12590 29736
rect 8202 29656 8208 29708
rect 8260 29656 8266 29708
rect 8389 29699 8447 29705
rect 8389 29665 8401 29699
rect 8435 29696 8447 29699
rect 9306 29696 9312 29708
rect 8435 29668 9312 29696
rect 8435 29665 8447 29668
rect 8389 29659 8447 29665
rect 9306 29656 9312 29668
rect 9364 29656 9370 29708
rect 12989 29699 13047 29705
rect 12989 29665 13001 29699
rect 13035 29696 13047 29699
rect 13262 29696 13268 29708
rect 13035 29668 13268 29696
rect 13035 29665 13047 29668
rect 12989 29659 13047 29665
rect 13262 29656 13268 29668
rect 13320 29656 13326 29708
rect 13372 29696 13400 29736
rect 17770 29724 17776 29776
rect 17828 29764 17834 29776
rect 17828 29736 18276 29764
rect 17828 29724 17834 29736
rect 14645 29699 14703 29705
rect 14645 29696 14657 29699
rect 13372 29668 14657 29696
rect 14645 29665 14657 29668
rect 14691 29665 14703 29699
rect 14645 29659 14703 29665
rect 15102 29656 15108 29708
rect 15160 29696 15166 29708
rect 15160 29668 16160 29696
rect 15160 29656 15166 29668
rect 8021 29631 8079 29637
rect 8021 29597 8033 29631
rect 8067 29597 8079 29631
rect 8220 29628 8248 29656
rect 10873 29631 10931 29637
rect 10873 29628 10885 29631
rect 8220 29600 10885 29628
rect 8021 29591 8079 29597
rect 10873 29597 10885 29600
rect 10919 29628 10931 29631
rect 12158 29628 12164 29640
rect 10919 29600 12164 29628
rect 10919 29597 10931 29600
rect 10873 29591 10931 29597
rect 12158 29588 12164 29600
rect 12216 29588 12222 29640
rect 12713 29631 12771 29637
rect 12713 29597 12725 29631
rect 12759 29597 12771 29631
rect 12713 29591 12771 29597
rect 8205 29563 8263 29569
rect 8205 29529 8217 29563
rect 8251 29560 8263 29563
rect 8294 29560 8300 29572
rect 8251 29532 8300 29560
rect 8251 29529 8263 29532
rect 8205 29523 8263 29529
rect 8294 29520 8300 29532
rect 8352 29520 8358 29572
rect 8938 29560 8944 29572
rect 8899 29532 8944 29560
rect 8938 29520 8944 29532
rect 8996 29520 9002 29572
rect 9125 29563 9183 29569
rect 9125 29529 9137 29563
rect 9171 29529 9183 29563
rect 9125 29523 9183 29529
rect 11140 29563 11198 29569
rect 11140 29529 11152 29563
rect 11186 29560 11198 29563
rect 12342 29560 12348 29572
rect 11186 29532 12348 29560
rect 11186 29529 11198 29532
rect 11140 29523 11198 29529
rect 8478 29452 8484 29504
rect 8536 29492 8542 29504
rect 9140 29492 9168 29523
rect 12342 29520 12348 29532
rect 12400 29520 12406 29572
rect 8536 29464 9168 29492
rect 9309 29495 9367 29501
rect 8536 29452 8542 29464
rect 9309 29461 9321 29495
rect 9355 29492 9367 29495
rect 9490 29492 9496 29504
rect 9355 29464 9496 29492
rect 9355 29461 9367 29464
rect 9309 29455 9367 29461
rect 9490 29452 9496 29464
rect 9548 29452 9554 29504
rect 12250 29492 12256 29504
rect 12211 29464 12256 29492
rect 12250 29452 12256 29464
rect 12308 29492 12314 29504
rect 12728 29492 12756 29591
rect 14274 29588 14280 29640
rect 14332 29628 14338 29640
rect 14826 29628 14832 29640
rect 14332 29600 14832 29628
rect 14332 29588 14338 29600
rect 14826 29588 14832 29600
rect 14884 29628 14890 29640
rect 14921 29631 14979 29637
rect 14921 29628 14933 29631
rect 14884 29600 14933 29628
rect 14884 29588 14890 29600
rect 14921 29597 14933 29600
rect 14967 29597 14979 29631
rect 14921 29591 14979 29597
rect 15010 29588 15016 29640
rect 15068 29628 15074 29640
rect 15381 29631 15439 29637
rect 15068 29600 15113 29628
rect 15068 29588 15074 29600
rect 15381 29597 15393 29631
rect 15427 29628 15439 29631
rect 15562 29628 15568 29640
rect 15427 29600 15568 29628
rect 15427 29597 15439 29600
rect 15381 29591 15439 29597
rect 15562 29588 15568 29600
rect 15620 29588 15626 29640
rect 16022 29628 16028 29640
rect 15983 29600 16028 29628
rect 16022 29588 16028 29600
rect 16080 29588 16086 29640
rect 16132 29637 16160 29668
rect 16482 29656 16488 29708
rect 16540 29696 16546 29708
rect 17405 29699 17463 29705
rect 17405 29696 17417 29699
rect 16540 29668 17417 29696
rect 16540 29656 16546 29668
rect 17405 29665 17417 29668
rect 17451 29665 17463 29699
rect 17405 29659 17463 29665
rect 16117 29631 16175 29637
rect 16117 29597 16129 29631
rect 16163 29597 16175 29631
rect 17126 29628 17132 29640
rect 17087 29600 17132 29628
rect 16117 29591 16175 29597
rect 17126 29588 17132 29600
rect 17184 29588 17190 29640
rect 17221 29631 17279 29637
rect 17221 29597 17233 29631
rect 17267 29628 17279 29631
rect 17586 29628 17592 29640
rect 17267 29600 17592 29628
rect 17267 29597 17279 29600
rect 17221 29591 17279 29597
rect 17586 29588 17592 29600
rect 17644 29588 17650 29640
rect 17678 29588 17684 29640
rect 17736 29628 17742 29640
rect 18248 29637 18276 29736
rect 18141 29631 18199 29637
rect 18141 29628 18153 29631
rect 17736 29600 18153 29628
rect 17736 29588 17742 29600
rect 18141 29597 18153 29600
rect 18187 29597 18199 29631
rect 18141 29591 18199 29597
rect 18233 29631 18291 29637
rect 18233 29597 18245 29631
rect 18279 29597 18291 29631
rect 18233 29591 18291 29597
rect 18322 29588 18328 29640
rect 18380 29628 18386 29640
rect 18524 29637 18552 29804
rect 19337 29801 19349 29835
rect 19383 29832 19395 29835
rect 19518 29832 19524 29844
rect 19383 29804 19524 29832
rect 19383 29801 19395 29804
rect 19337 29795 19395 29801
rect 19518 29792 19524 29804
rect 19576 29792 19582 29844
rect 19978 29792 19984 29844
rect 20036 29832 20042 29844
rect 21542 29832 21548 29844
rect 20036 29804 21548 29832
rect 20036 29792 20042 29804
rect 21542 29792 21548 29804
rect 21600 29792 21606 29844
rect 22649 29835 22707 29841
rect 22649 29801 22661 29835
rect 22695 29832 22707 29835
rect 22738 29832 22744 29844
rect 22695 29804 22744 29832
rect 22695 29801 22707 29804
rect 22649 29795 22707 29801
rect 22738 29792 22744 29804
rect 22796 29792 22802 29844
rect 23385 29835 23443 29841
rect 23385 29801 23397 29835
rect 23431 29832 23443 29835
rect 24118 29832 24124 29844
rect 23431 29804 24124 29832
rect 23431 29801 23443 29804
rect 23385 29795 23443 29801
rect 24118 29792 24124 29804
rect 24176 29792 24182 29844
rect 25682 29792 25688 29844
rect 25740 29832 25746 29844
rect 25777 29835 25835 29841
rect 25777 29832 25789 29835
rect 25740 29804 25789 29832
rect 25740 29792 25746 29804
rect 25777 29801 25789 29804
rect 25823 29801 25835 29835
rect 25777 29795 25835 29801
rect 26881 29835 26939 29841
rect 26881 29801 26893 29835
rect 26927 29832 26939 29835
rect 27706 29832 27712 29844
rect 26927 29804 27712 29832
rect 26927 29801 26939 29804
rect 26881 29795 26939 29801
rect 27706 29792 27712 29804
rect 27764 29792 27770 29844
rect 27798 29792 27804 29844
rect 27856 29832 27862 29844
rect 27856 29804 27901 29832
rect 27856 29792 27862 29804
rect 27982 29792 27988 29844
rect 28040 29832 28046 29844
rect 46934 29832 46940 29844
rect 28040 29804 46940 29832
rect 28040 29792 28046 29804
rect 46934 29792 46940 29804
rect 46992 29792 46998 29844
rect 24026 29764 24032 29776
rect 22066 29736 24032 29764
rect 20438 29696 20444 29708
rect 19168 29668 20300 29696
rect 20399 29668 20444 29696
rect 18509 29631 18567 29637
rect 18380 29600 18425 29628
rect 18380 29588 18386 29600
rect 18509 29597 18521 29631
rect 18555 29597 18567 29631
rect 18509 29591 18567 29597
rect 12986 29520 12992 29572
rect 13044 29560 13050 29572
rect 15841 29563 15899 29569
rect 13044 29532 15608 29560
rect 13044 29520 13050 29532
rect 12308 29464 12756 29492
rect 15105 29495 15163 29501
rect 12308 29452 12314 29464
rect 15105 29461 15117 29495
rect 15151 29492 15163 29495
rect 15470 29492 15476 29504
rect 15151 29464 15476 29492
rect 15151 29461 15163 29464
rect 15105 29455 15163 29461
rect 15470 29452 15476 29464
rect 15528 29452 15534 29504
rect 15580 29492 15608 29532
rect 15841 29529 15853 29563
rect 15887 29560 15899 29563
rect 19168 29560 19196 29668
rect 19245 29631 19303 29637
rect 19245 29597 19257 29631
rect 19291 29597 19303 29631
rect 19245 29591 19303 29597
rect 15887 29532 19196 29560
rect 15887 29529 15899 29532
rect 15841 29523 15899 29529
rect 17218 29492 17224 29504
rect 15580 29464 17224 29492
rect 17218 29452 17224 29464
rect 17276 29452 17282 29504
rect 17402 29492 17408 29504
rect 17363 29464 17408 29492
rect 17402 29452 17408 29464
rect 17460 29452 17466 29504
rect 17862 29492 17868 29504
rect 17823 29464 17868 29492
rect 17862 29452 17868 29464
rect 17920 29452 17926 29504
rect 17954 29452 17960 29504
rect 18012 29492 18018 29504
rect 19260 29492 19288 29591
rect 19334 29588 19340 29640
rect 19392 29628 19398 29640
rect 20165 29631 20223 29637
rect 20165 29628 20177 29631
rect 19392 29600 20177 29628
rect 19392 29588 19398 29600
rect 20165 29597 20177 29600
rect 20211 29597 20223 29631
rect 20272 29628 20300 29668
rect 20438 29656 20444 29668
rect 20496 29656 20502 29708
rect 21634 29656 21640 29708
rect 21692 29696 21698 29708
rect 22066 29696 22094 29736
rect 24026 29724 24032 29736
rect 24084 29724 24090 29776
rect 25866 29724 25872 29776
rect 25924 29764 25930 29776
rect 35802 29764 35808 29776
rect 25924 29736 35808 29764
rect 25924 29724 25930 29736
rect 35802 29724 35808 29736
rect 35860 29724 35866 29776
rect 21692 29668 22094 29696
rect 21692 29656 21698 29668
rect 25498 29656 25504 29708
rect 25556 29696 25562 29708
rect 26602 29696 26608 29708
rect 25556 29668 26608 29696
rect 25556 29656 25562 29668
rect 26602 29656 26608 29668
rect 26660 29696 26666 29708
rect 26786 29696 26792 29708
rect 26660 29668 26792 29696
rect 26660 29656 26666 29668
rect 26786 29656 26792 29668
rect 26844 29656 26850 29708
rect 28534 29696 28540 29708
rect 26988 29668 28540 29696
rect 26988 29640 27016 29668
rect 28534 29656 28540 29668
rect 28592 29656 28598 29708
rect 29546 29656 29552 29708
rect 29604 29696 29610 29708
rect 30009 29699 30067 29705
rect 30009 29696 30021 29699
rect 29604 29668 30021 29696
rect 29604 29656 29610 29668
rect 30009 29665 30021 29668
rect 30055 29665 30067 29699
rect 30190 29696 30196 29708
rect 30151 29668 30196 29696
rect 30009 29659 30067 29665
rect 30190 29656 30196 29668
rect 30248 29656 30254 29708
rect 34790 29696 34796 29708
rect 31864 29668 34796 29696
rect 20530 29628 20536 29640
rect 20272 29600 20536 29628
rect 20165 29591 20223 29597
rect 20530 29588 20536 29600
rect 20588 29588 20594 29640
rect 22370 29628 22376 29640
rect 22331 29600 22376 29628
rect 22370 29588 22376 29600
rect 22428 29588 22434 29640
rect 22465 29631 22523 29637
rect 22465 29597 22477 29631
rect 22511 29597 22523 29631
rect 22465 29591 22523 29597
rect 21818 29520 21824 29572
rect 21876 29560 21882 29572
rect 22480 29560 22508 29591
rect 23106 29588 23112 29640
rect 23164 29628 23170 29640
rect 23569 29631 23627 29637
rect 23569 29628 23581 29631
rect 23164 29600 23581 29628
rect 23164 29588 23170 29600
rect 23569 29597 23581 29600
rect 23615 29597 23627 29631
rect 23569 29591 23627 29597
rect 23750 29588 23756 29640
rect 23808 29628 23814 29640
rect 23845 29631 23903 29637
rect 23845 29628 23857 29631
rect 23808 29600 23857 29628
rect 23808 29588 23814 29600
rect 23845 29597 23857 29600
rect 23891 29597 23903 29631
rect 23845 29591 23903 29597
rect 24397 29631 24455 29637
rect 24397 29597 24409 29631
rect 24443 29628 24455 29631
rect 25406 29628 25412 29640
rect 24443 29600 25412 29628
rect 24443 29597 24455 29600
rect 24397 29591 24455 29597
rect 25406 29588 25412 29600
rect 25464 29628 25470 29640
rect 26970 29628 26976 29640
rect 25464 29600 26976 29628
rect 25464 29588 25470 29600
rect 26970 29588 26976 29600
rect 27028 29588 27034 29640
rect 27617 29631 27675 29637
rect 27617 29628 27629 29631
rect 27080 29600 27629 29628
rect 21876 29532 22508 29560
rect 21876 29520 21882 29532
rect 23658 29520 23664 29572
rect 23716 29560 23722 29572
rect 24642 29563 24700 29569
rect 24642 29560 24654 29563
rect 23716 29532 24654 29560
rect 23716 29520 23722 29532
rect 24642 29529 24654 29532
rect 24688 29529 24700 29563
rect 26786 29560 26792 29572
rect 24642 29523 24700 29529
rect 24780 29532 26556 29560
rect 26747 29532 26792 29560
rect 18012 29464 19288 29492
rect 18012 29452 18018 29464
rect 21542 29452 21548 29504
rect 21600 29492 21606 29504
rect 23382 29492 23388 29504
rect 21600 29464 23388 29492
rect 21600 29452 21606 29464
rect 23382 29452 23388 29464
rect 23440 29452 23446 29504
rect 23750 29492 23756 29504
rect 23711 29464 23756 29492
rect 23750 29452 23756 29464
rect 23808 29452 23814 29504
rect 24026 29452 24032 29504
rect 24084 29492 24090 29504
rect 24780 29492 24808 29532
rect 24084 29464 24808 29492
rect 24084 29452 24090 29464
rect 24854 29452 24860 29504
rect 24912 29492 24918 29504
rect 26418 29492 26424 29504
rect 24912 29464 26424 29492
rect 24912 29452 24918 29464
rect 26418 29452 26424 29464
rect 26476 29452 26482 29504
rect 26528 29492 26556 29532
rect 26786 29520 26792 29532
rect 26844 29520 26850 29572
rect 27080 29492 27108 29600
rect 27617 29597 27629 29600
rect 27663 29597 27675 29631
rect 28810 29628 28816 29640
rect 28771 29600 28816 29628
rect 27617 29591 27675 29597
rect 28810 29588 28816 29600
rect 28868 29588 28874 29640
rect 31864 29637 31892 29668
rect 34790 29656 34796 29668
rect 34848 29656 34854 29708
rect 35176 29668 35388 29696
rect 31849 29631 31907 29637
rect 31849 29597 31861 29631
rect 31895 29597 31907 29631
rect 31849 29591 31907 29597
rect 31941 29631 31999 29637
rect 31941 29597 31953 29631
rect 31987 29597 31999 29631
rect 31941 29591 31999 29597
rect 27433 29563 27491 29569
rect 27433 29529 27445 29563
rect 27479 29529 27491 29563
rect 27433 29523 27491 29529
rect 26528 29464 27108 29492
rect 27448 29492 27476 29523
rect 27522 29520 27528 29572
rect 27580 29560 27586 29572
rect 28997 29563 29055 29569
rect 28997 29560 29009 29563
rect 27580 29532 29009 29560
rect 27580 29520 27586 29532
rect 28997 29529 29009 29532
rect 29043 29560 29055 29563
rect 30374 29560 30380 29572
rect 29043 29532 30380 29560
rect 29043 29529 29055 29532
rect 28997 29523 29055 29529
rect 30374 29520 30380 29532
rect 30432 29520 30438 29572
rect 31018 29520 31024 29572
rect 31076 29560 31082 29572
rect 31956 29560 31984 29591
rect 32030 29588 32036 29640
rect 32088 29628 32094 29640
rect 32217 29631 32275 29637
rect 32088 29600 32133 29628
rect 32088 29588 32094 29600
rect 32217 29597 32229 29631
rect 32263 29628 32275 29631
rect 32306 29628 32312 29640
rect 32263 29600 32312 29628
rect 32263 29597 32275 29600
rect 32217 29591 32275 29597
rect 32306 29588 32312 29600
rect 32364 29628 32370 29640
rect 32766 29628 32772 29640
rect 32364 29600 32772 29628
rect 32364 29588 32370 29600
rect 32766 29588 32772 29600
rect 32824 29588 32830 29640
rect 35066 29637 35072 29640
rect 35049 29631 35072 29637
rect 35049 29597 35061 29631
rect 35049 29591 35072 29597
rect 35066 29588 35072 29591
rect 35124 29588 35130 29640
rect 35176 29637 35204 29668
rect 35161 29631 35219 29637
rect 35161 29597 35173 29631
rect 35207 29597 35219 29631
rect 35161 29591 35219 29597
rect 35253 29631 35311 29637
rect 35253 29597 35265 29631
rect 35299 29597 35311 29631
rect 35253 29591 35311 29597
rect 32398 29560 32404 29572
rect 31076 29532 32404 29560
rect 31076 29520 31082 29532
rect 32398 29520 32404 29532
rect 32456 29520 32462 29572
rect 29549 29495 29607 29501
rect 29549 29492 29561 29495
rect 27448 29464 29561 29492
rect 29549 29461 29561 29464
rect 29595 29461 29607 29495
rect 29914 29492 29920 29504
rect 29875 29464 29920 29492
rect 29549 29455 29607 29461
rect 29914 29452 29920 29464
rect 29972 29452 29978 29504
rect 31570 29492 31576 29504
rect 31531 29464 31576 29492
rect 31570 29452 31576 29464
rect 31628 29452 31634 29504
rect 31754 29452 31760 29504
rect 31812 29492 31818 29504
rect 32122 29492 32128 29504
rect 31812 29464 32128 29492
rect 31812 29452 31818 29464
rect 32122 29452 32128 29464
rect 32180 29452 32186 29504
rect 34790 29492 34796 29504
rect 34751 29464 34796 29492
rect 34790 29452 34796 29464
rect 34848 29452 34854 29504
rect 35257 29492 35285 29591
rect 35360 29560 35388 29668
rect 35526 29656 35532 29708
rect 35584 29696 35590 29708
rect 47581 29699 47639 29705
rect 47581 29696 47593 29699
rect 35584 29668 47593 29696
rect 35584 29656 35590 29668
rect 47581 29665 47593 29668
rect 47627 29665 47639 29699
rect 47581 29659 47639 29665
rect 35431 29631 35489 29637
rect 35431 29597 35443 29631
rect 35477 29628 35489 29631
rect 35710 29628 35716 29640
rect 35477 29600 35716 29628
rect 35477 29597 35489 29600
rect 35431 29591 35489 29597
rect 35710 29588 35716 29600
rect 35768 29588 35774 29640
rect 47302 29628 47308 29640
rect 47263 29600 47308 29628
rect 47302 29588 47308 29600
rect 47360 29588 47366 29640
rect 35618 29560 35624 29572
rect 35360 29532 35624 29560
rect 35618 29520 35624 29532
rect 35676 29520 35682 29572
rect 35434 29492 35440 29504
rect 35257 29464 35440 29492
rect 35434 29452 35440 29464
rect 35492 29452 35498 29504
rect 1104 29402 48852 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 48852 29402
rect 1104 29328 48852 29350
rect 16574 29288 16580 29300
rect 9692 29260 16580 29288
rect 8202 29220 8208 29232
rect 7208 29192 8208 29220
rect 7006 29112 7012 29164
rect 7064 29152 7070 29164
rect 7208 29161 7236 29192
rect 8202 29180 8208 29192
rect 8260 29180 8266 29232
rect 9692 29164 9720 29260
rect 16574 29248 16580 29260
rect 16632 29248 16638 29300
rect 16666 29248 16672 29300
rect 16724 29288 16730 29300
rect 17218 29288 17224 29300
rect 16724 29260 17224 29288
rect 16724 29248 16730 29260
rect 17218 29248 17224 29260
rect 17276 29248 17282 29300
rect 17310 29248 17316 29300
rect 17368 29288 17374 29300
rect 17368 29260 18828 29288
rect 17368 29248 17374 29260
rect 12158 29180 12164 29232
rect 12216 29220 12222 29232
rect 15286 29220 15292 29232
rect 12216 29192 15292 29220
rect 12216 29180 12222 29192
rect 7193 29155 7251 29161
rect 7193 29152 7205 29155
rect 7064 29124 7205 29152
rect 7064 29112 7070 29124
rect 7193 29121 7205 29124
rect 7239 29121 7251 29155
rect 7193 29115 7251 29121
rect 7460 29155 7518 29161
rect 7460 29121 7472 29155
rect 7506 29152 7518 29155
rect 9263 29155 9321 29161
rect 9263 29152 9275 29155
rect 7506 29124 9076 29152
rect 7506 29121 7518 29124
rect 7460 29115 7518 29121
rect 9048 29093 9076 29124
rect 9140 29124 9275 29152
rect 9033 29087 9091 29093
rect 9033 29053 9045 29087
rect 9079 29053 9091 29087
rect 9140 29084 9168 29124
rect 9263 29121 9275 29124
rect 9309 29121 9321 29155
rect 9398 29152 9404 29164
rect 9359 29124 9404 29152
rect 9263 29115 9321 29121
rect 9398 29112 9404 29124
rect 9456 29112 9462 29164
rect 9490 29112 9496 29164
rect 9548 29152 9554 29164
rect 9548 29124 9593 29152
rect 9548 29112 9554 29124
rect 9674 29112 9680 29164
rect 9732 29152 9738 29164
rect 12526 29152 12532 29164
rect 9732 29124 9825 29152
rect 12487 29124 12532 29152
rect 9732 29112 9738 29124
rect 12526 29112 12532 29124
rect 12584 29112 12590 29164
rect 12989 29155 13047 29161
rect 12989 29121 13001 29155
rect 13035 29121 13047 29155
rect 12989 29115 13047 29121
rect 13173 29155 13231 29161
rect 13173 29121 13185 29155
rect 13219 29152 13231 29155
rect 13262 29152 13268 29164
rect 13219 29124 13268 29152
rect 13219 29121 13231 29124
rect 13173 29115 13231 29121
rect 9766 29084 9772 29096
rect 9140 29056 9772 29084
rect 9033 29047 9091 29053
rect 9766 29044 9772 29056
rect 9824 29084 9830 29096
rect 10318 29084 10324 29096
rect 9824 29056 10324 29084
rect 9824 29044 9830 29056
rect 10318 29044 10324 29056
rect 10376 29044 10382 29096
rect 13004 29084 13032 29115
rect 13262 29112 13268 29124
rect 13320 29112 13326 29164
rect 13832 29161 13860 29192
rect 15286 29180 15292 29192
rect 15344 29180 15350 29232
rect 15470 29180 15476 29232
rect 15528 29220 15534 29232
rect 15841 29223 15899 29229
rect 15841 29220 15853 29223
rect 15528 29192 15853 29220
rect 15528 29180 15534 29192
rect 15841 29189 15853 29192
rect 15887 29220 15899 29223
rect 17494 29220 17500 29232
rect 15887 29192 17500 29220
rect 15887 29189 15899 29192
rect 15841 29183 15899 29189
rect 17494 29180 17500 29192
rect 17552 29180 17558 29232
rect 17862 29180 17868 29232
rect 17920 29220 17926 29232
rect 18662 29223 18720 29229
rect 18662 29220 18674 29223
rect 17920 29192 18674 29220
rect 17920 29180 17926 29192
rect 18662 29189 18674 29192
rect 18708 29189 18720 29223
rect 18800 29220 18828 29260
rect 20162 29248 20168 29300
rect 20220 29288 20226 29300
rect 20441 29291 20499 29297
rect 20441 29288 20453 29291
rect 20220 29260 20453 29288
rect 20220 29248 20226 29260
rect 20441 29257 20453 29260
rect 20487 29257 20499 29291
rect 23198 29288 23204 29300
rect 23159 29260 23204 29288
rect 20441 29251 20499 29257
rect 23198 29248 23204 29260
rect 23256 29248 23262 29300
rect 25777 29291 25835 29297
rect 25777 29257 25789 29291
rect 25823 29288 25835 29291
rect 27062 29288 27068 29300
rect 25823 29260 27068 29288
rect 25823 29257 25835 29260
rect 25777 29251 25835 29257
rect 27062 29248 27068 29260
rect 27120 29288 27126 29300
rect 29549 29291 29607 29297
rect 27120 29260 29408 29288
rect 27120 29248 27126 29260
rect 20622 29220 20628 29232
rect 18800 29192 20484 29220
rect 20535 29192 20628 29220
rect 18662 29183 18720 29189
rect 14090 29161 14096 29164
rect 13817 29155 13875 29161
rect 13817 29121 13829 29155
rect 13863 29121 13875 29155
rect 13817 29115 13875 29121
rect 14084 29115 14096 29161
rect 14148 29152 14154 29164
rect 15657 29155 15715 29161
rect 14148 29124 14184 29152
rect 14090 29112 14096 29115
rect 14148 29112 14154 29124
rect 15657 29121 15669 29155
rect 15703 29152 15715 29155
rect 15746 29152 15752 29164
rect 15703 29124 15752 29152
rect 15703 29121 15715 29124
rect 15657 29115 15715 29121
rect 15746 29112 15752 29124
rect 15804 29112 15810 29164
rect 15930 29152 15936 29164
rect 15891 29124 15936 29152
rect 15930 29112 15936 29124
rect 15988 29112 15994 29164
rect 17126 29112 17132 29164
rect 17184 29152 17190 29164
rect 17678 29152 17684 29164
rect 17184 29124 17684 29152
rect 17184 29112 17190 29124
rect 17678 29112 17684 29124
rect 17736 29112 17742 29164
rect 17770 29112 17776 29164
rect 17828 29152 17834 29164
rect 19886 29152 19892 29164
rect 17828 29124 19892 29152
rect 17828 29112 17834 29124
rect 19886 29112 19892 29124
rect 19944 29152 19950 29164
rect 20349 29155 20407 29161
rect 20349 29152 20361 29155
rect 19944 29124 20361 29152
rect 19944 29112 19950 29124
rect 20349 29121 20361 29124
rect 20395 29121 20407 29155
rect 20349 29115 20407 29121
rect 13004 29056 13860 29084
rect 8478 28976 8484 29028
rect 8536 29016 8542 29028
rect 8573 29019 8631 29025
rect 8573 29016 8585 29019
rect 8536 28988 8585 29016
rect 8536 28976 8542 28988
rect 8573 28985 8585 28988
rect 8619 28985 8631 29019
rect 8573 28979 8631 28985
rect 11974 28976 11980 29028
rect 12032 29016 12038 29028
rect 12345 29019 12403 29025
rect 12345 29016 12357 29019
rect 12032 28988 12357 29016
rect 12032 28976 12038 28988
rect 12345 28985 12357 28988
rect 12391 28985 12403 29019
rect 12345 28979 12403 28985
rect 2038 28948 2044 28960
rect 1999 28920 2044 28948
rect 2038 28908 2044 28920
rect 2096 28908 2102 28960
rect 12986 28908 12992 28960
rect 13044 28948 13050 28960
rect 13081 28951 13139 28957
rect 13081 28948 13093 28951
rect 13044 28920 13093 28948
rect 13044 28908 13050 28920
rect 13081 28917 13093 28920
rect 13127 28917 13139 28951
rect 13832 28948 13860 29056
rect 15562 29044 15568 29096
rect 15620 29084 15626 29096
rect 16482 29084 16488 29096
rect 15620 29056 16488 29084
rect 15620 29044 15626 29056
rect 16482 29044 16488 29056
rect 16540 29084 16546 29096
rect 17405 29087 17463 29093
rect 17405 29084 17417 29087
rect 16540 29056 17417 29084
rect 16540 29044 16546 29056
rect 17405 29053 17417 29056
rect 17451 29053 17463 29087
rect 17405 29047 17463 29053
rect 17494 29044 17500 29096
rect 17552 29084 17558 29096
rect 17954 29084 17960 29096
rect 17552 29056 17960 29084
rect 17552 29044 17558 29056
rect 17954 29044 17960 29056
rect 18012 29044 18018 29096
rect 18417 29087 18475 29093
rect 18417 29053 18429 29087
rect 18463 29053 18475 29087
rect 20456 29084 20484 29192
rect 20548 29161 20576 29192
rect 20622 29180 20628 29192
rect 20680 29220 20686 29232
rect 22370 29220 22376 29232
rect 20680 29192 22376 29220
rect 20680 29180 20686 29192
rect 20533 29155 20591 29161
rect 20533 29121 20545 29155
rect 20579 29121 20591 29155
rect 20533 29115 20591 29121
rect 20898 29112 20904 29164
rect 20956 29152 20962 29164
rect 21818 29152 21824 29164
rect 20956 29124 21824 29152
rect 20956 29112 20962 29124
rect 21818 29112 21824 29124
rect 21876 29112 21882 29164
rect 22112 29161 22140 29192
rect 22370 29180 22376 29192
rect 22428 29180 22434 29232
rect 23937 29223 23995 29229
rect 23937 29189 23949 29223
rect 23983 29220 23995 29223
rect 25498 29220 25504 29232
rect 23983 29192 25504 29220
rect 23983 29189 23995 29192
rect 23937 29183 23995 29189
rect 25498 29180 25504 29192
rect 25556 29180 25562 29232
rect 27522 29220 27528 29232
rect 27483 29192 27528 29220
rect 27522 29180 27528 29192
rect 27580 29180 27586 29232
rect 22097 29155 22155 29161
rect 22097 29121 22109 29155
rect 22143 29152 22155 29155
rect 22143 29124 22177 29152
rect 22143 29121 22155 29124
rect 22097 29115 22155 29121
rect 22738 29112 22744 29164
rect 22796 29152 22802 29164
rect 23385 29155 23443 29161
rect 23385 29152 23397 29155
rect 22796 29124 23397 29152
rect 22796 29112 22802 29124
rect 23385 29121 23397 29124
rect 23431 29121 23443 29155
rect 23385 29115 23443 29121
rect 23750 29112 23756 29164
rect 23808 29152 23814 29164
rect 24121 29155 24179 29161
rect 24121 29152 24133 29155
rect 23808 29124 24133 29152
rect 23808 29112 23814 29124
rect 24121 29121 24133 29124
rect 24167 29152 24179 29155
rect 24762 29152 24768 29164
rect 24167 29124 24768 29152
rect 24167 29121 24179 29124
rect 24121 29115 24179 29121
rect 24762 29112 24768 29124
rect 24820 29112 24826 29164
rect 24854 29112 24860 29164
rect 24912 29152 24918 29164
rect 25593 29155 25651 29161
rect 25593 29152 25605 29155
rect 24912 29124 25605 29152
rect 24912 29112 24918 29124
rect 25593 29121 25605 29124
rect 25639 29121 25651 29155
rect 25593 29115 25651 29121
rect 27430 29112 27436 29164
rect 27488 29152 27494 29164
rect 28425 29155 28483 29161
rect 28425 29152 28437 29155
rect 27488 29124 28437 29152
rect 27488 29112 27494 29124
rect 28425 29121 28437 29124
rect 28471 29121 28483 29155
rect 29380 29152 29408 29260
rect 29549 29257 29561 29291
rect 29595 29288 29607 29291
rect 29914 29288 29920 29300
rect 29595 29260 29920 29288
rect 29595 29257 29607 29260
rect 29549 29251 29607 29257
rect 29914 29248 29920 29260
rect 29972 29248 29978 29300
rect 30006 29248 30012 29300
rect 30064 29288 30070 29300
rect 31297 29291 31355 29297
rect 31297 29288 31309 29291
rect 30064 29260 31309 29288
rect 30064 29248 30070 29260
rect 31297 29257 31309 29260
rect 31343 29257 31355 29291
rect 31297 29251 31355 29257
rect 31570 29248 31576 29300
rect 31628 29288 31634 29300
rect 31754 29288 31760 29300
rect 31628 29260 31760 29288
rect 31628 29248 31634 29260
rect 31754 29248 31760 29260
rect 31812 29248 31818 29300
rect 32950 29248 32956 29300
rect 33008 29288 33014 29300
rect 33137 29291 33195 29297
rect 33137 29288 33149 29291
rect 33008 29260 33149 29288
rect 33008 29248 33014 29260
rect 33137 29257 33149 29260
rect 33183 29257 33195 29291
rect 34698 29288 34704 29300
rect 34659 29260 34704 29288
rect 33137 29251 33195 29257
rect 34698 29248 34704 29260
rect 34756 29248 34762 29300
rect 36541 29291 36599 29297
rect 36541 29288 36553 29291
rect 34808 29260 36553 29288
rect 31205 29223 31263 29229
rect 31205 29189 31217 29223
rect 31251 29220 31263 29223
rect 33226 29220 33232 29232
rect 31251 29192 33232 29220
rect 31251 29189 31263 29192
rect 31205 29183 31263 29189
rect 33226 29180 33232 29192
rect 33284 29180 33290 29232
rect 33318 29180 33324 29232
rect 33376 29220 33382 29232
rect 34333 29223 34391 29229
rect 33376 29192 34100 29220
rect 33376 29180 33382 29192
rect 33045 29155 33103 29161
rect 29380 29124 31432 29152
rect 28425 29115 28483 29121
rect 22189 29087 22247 29093
rect 20456 29056 22094 29084
rect 18417 29047 18475 29053
rect 15102 28976 15108 29028
rect 15160 29016 15166 29028
rect 15657 29019 15715 29025
rect 15657 29016 15669 29019
rect 15160 28988 15669 29016
rect 15160 28976 15166 28988
rect 15657 28985 15669 28988
rect 15703 28985 15715 29019
rect 17586 29016 17592 29028
rect 17547 28988 17592 29016
rect 15657 28979 15715 28985
rect 17586 28976 17592 28988
rect 17644 28976 17650 29028
rect 14458 28948 14464 28960
rect 13832 28920 14464 28948
rect 13081 28911 13139 28917
rect 14458 28908 14464 28920
rect 14516 28908 14522 28960
rect 15010 28908 15016 28960
rect 15068 28948 15074 28960
rect 15197 28951 15255 28957
rect 15197 28948 15209 28951
rect 15068 28920 15209 28948
rect 15068 28908 15074 28920
rect 15197 28917 15209 28920
rect 15243 28917 15255 28951
rect 15197 28911 15255 28917
rect 16482 28908 16488 28960
rect 16540 28948 16546 28960
rect 18432 28948 18460 29047
rect 19797 29019 19855 29025
rect 19797 28985 19809 29019
rect 19843 28985 19855 29019
rect 22066 29016 22094 29056
rect 22189 29053 22201 29087
rect 22235 29084 22247 29087
rect 22462 29084 22468 29096
rect 22235 29056 22468 29084
rect 22235 29053 22247 29056
rect 22189 29047 22247 29053
rect 22462 29044 22468 29056
rect 22520 29044 22526 29096
rect 27614 29084 27620 29096
rect 23032 29056 27620 29084
rect 23032 29016 23060 29056
rect 27614 29044 27620 29056
rect 27672 29044 27678 29096
rect 31404 29093 31432 29124
rect 33045 29121 33057 29155
rect 33091 29152 33103 29155
rect 33962 29152 33968 29164
rect 33091 29124 33968 29152
rect 33091 29121 33103 29124
rect 33045 29115 33103 29121
rect 33962 29112 33968 29124
rect 34020 29112 34026 29164
rect 34072 29152 34100 29192
rect 34333 29189 34345 29223
rect 34379 29220 34391 29223
rect 34808 29220 34836 29260
rect 36541 29257 36553 29260
rect 36587 29288 36599 29291
rect 36630 29288 36636 29300
rect 36587 29260 36636 29288
rect 36587 29257 36599 29260
rect 36541 29251 36599 29257
rect 36630 29248 36636 29260
rect 36688 29248 36694 29300
rect 35406 29223 35464 29229
rect 35406 29220 35418 29223
rect 34379 29192 34836 29220
rect 35084 29192 35418 29220
rect 34379 29189 34391 29192
rect 34333 29183 34391 29189
rect 34517 29155 34575 29161
rect 34517 29152 34529 29155
rect 34072 29124 34529 29152
rect 34517 29121 34529 29124
rect 34563 29152 34575 29155
rect 34698 29152 34704 29164
rect 34563 29124 34704 29152
rect 34563 29121 34575 29124
rect 34517 29115 34575 29121
rect 34698 29112 34704 29124
rect 34756 29112 34762 29164
rect 34790 29112 34796 29164
rect 34848 29152 34854 29164
rect 35084 29152 35112 29192
rect 35406 29189 35418 29192
rect 35452 29189 35464 29223
rect 35406 29183 35464 29189
rect 46014 29180 46020 29232
rect 46072 29220 46078 29232
rect 46072 29192 47624 29220
rect 46072 29180 46078 29192
rect 34848 29124 35112 29152
rect 35161 29155 35219 29161
rect 34848 29112 34854 29124
rect 35161 29121 35173 29155
rect 35207 29152 35219 29155
rect 35250 29152 35256 29164
rect 35207 29124 35256 29152
rect 35207 29121 35219 29124
rect 35161 29115 35219 29121
rect 35250 29112 35256 29124
rect 35308 29112 35314 29164
rect 46293 29155 46351 29161
rect 46293 29121 46305 29155
rect 46339 29152 46351 29155
rect 46750 29152 46756 29164
rect 46339 29124 46756 29152
rect 46339 29121 46351 29124
rect 46293 29115 46351 29121
rect 46750 29112 46756 29124
rect 46808 29112 46814 29164
rect 47596 29161 47624 29192
rect 47581 29155 47639 29161
rect 47581 29121 47593 29155
rect 47627 29121 47639 29155
rect 47581 29115 47639 29121
rect 28169 29087 28227 29093
rect 28169 29053 28181 29087
rect 28215 29053 28227 29087
rect 28169 29047 28227 29053
rect 31389 29087 31447 29093
rect 31389 29053 31401 29087
rect 31435 29084 31447 29087
rect 33321 29087 33379 29093
rect 33321 29084 33333 29087
rect 31435 29056 33333 29084
rect 31435 29053 31447 29056
rect 31389 29047 31447 29053
rect 33321 29053 33333 29056
rect 33367 29084 33379 29087
rect 33502 29084 33508 29096
rect 33367 29056 33508 29084
rect 33367 29053 33379 29056
rect 33321 29047 33379 29053
rect 22066 28988 23060 29016
rect 23124 28988 23336 29016
rect 19797 28979 19855 28985
rect 19334 28948 19340 28960
rect 16540 28920 19340 28948
rect 16540 28908 16546 28920
rect 19334 28908 19340 28920
rect 19392 28908 19398 28960
rect 19610 28908 19616 28960
rect 19668 28948 19674 28960
rect 19812 28948 19840 28979
rect 23124 28948 23152 28988
rect 19668 28920 23152 28948
rect 23308 28948 23336 28988
rect 23952 28988 24164 29016
rect 23952 28948 23980 28988
rect 23308 28920 23980 28948
rect 24136 28948 24164 28988
rect 25700 28988 25912 29016
rect 25700 28948 25728 28988
rect 24136 28920 25728 28948
rect 25884 28948 25912 28988
rect 26970 28976 26976 29028
rect 27028 29016 27034 29028
rect 27709 29019 27767 29025
rect 27709 29016 27721 29019
rect 27028 28988 27721 29016
rect 27028 28976 27034 28988
rect 27709 28985 27721 28988
rect 27755 29016 27767 29019
rect 28184 29016 28212 29047
rect 33502 29044 33508 29056
rect 33560 29044 33566 29096
rect 32677 29019 32735 29025
rect 27755 28988 28212 29016
rect 30760 28988 31156 29016
rect 27755 28985 27767 28988
rect 27709 28979 27767 28985
rect 30760 28948 30788 28988
rect 25884 28920 30788 28948
rect 30837 28951 30895 28957
rect 19668 28908 19674 28920
rect 30837 28917 30849 28951
rect 30883 28948 30895 28951
rect 31018 28948 31024 28960
rect 30883 28920 31024 28948
rect 30883 28917 30895 28920
rect 30837 28911 30895 28917
rect 31018 28908 31024 28920
rect 31076 28908 31082 28960
rect 31128 28948 31156 28988
rect 32677 28985 32689 29019
rect 32723 29016 32735 29019
rect 33686 29016 33692 29028
rect 32723 28988 33692 29016
rect 32723 28985 32735 28988
rect 32677 28979 32735 28985
rect 33686 28976 33692 28988
rect 33744 28976 33750 29028
rect 34624 28988 34836 29016
rect 34624 28948 34652 28988
rect 31128 28920 34652 28948
rect 34808 28948 34836 28988
rect 36464 28988 36676 29016
rect 36464 28948 36492 28988
rect 34808 28920 36492 28948
rect 36648 28948 36676 28988
rect 46658 28976 46664 29028
rect 46716 29016 46722 29028
rect 47673 29019 47731 29025
rect 47673 29016 47685 29019
rect 46716 28988 47685 29016
rect 46716 28976 46722 28988
rect 47673 28985 47685 28988
rect 47719 28985 47731 29019
rect 47673 28979 47731 28985
rect 46290 28948 46296 28960
rect 36648 28920 46296 28948
rect 46290 28908 46296 28920
rect 46348 28908 46354 28960
rect 46385 28951 46443 28957
rect 46385 28917 46397 28951
rect 46431 28948 46443 28951
rect 46474 28948 46480 28960
rect 46431 28920 46480 28948
rect 46431 28917 46443 28920
rect 46385 28911 46443 28917
rect 46474 28908 46480 28920
rect 46532 28908 46538 28960
rect 1104 28858 48852 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 48852 28858
rect 1104 28784 48852 28806
rect 9398 28744 9404 28756
rect 9321 28716 9404 28744
rect 1397 28611 1455 28617
rect 1397 28577 1409 28611
rect 1443 28608 1455 28611
rect 2038 28608 2044 28620
rect 1443 28580 2044 28608
rect 1443 28577 1455 28580
rect 1397 28571 1455 28577
rect 2038 28568 2044 28580
rect 2096 28568 2102 28620
rect 2774 28568 2780 28620
rect 2832 28608 2838 28620
rect 7006 28608 7012 28620
rect 2832 28580 2877 28608
rect 6967 28580 7012 28608
rect 2832 28568 2838 28580
rect 7006 28568 7012 28580
rect 7064 28568 7070 28620
rect 9214 28540 9220 28552
rect 9175 28512 9220 28540
rect 9214 28500 9220 28512
rect 9272 28500 9278 28552
rect 9321 28549 9349 28716
rect 9398 28704 9404 28716
rect 9456 28704 9462 28756
rect 14090 28704 14096 28756
rect 14148 28744 14154 28756
rect 14185 28747 14243 28753
rect 14185 28744 14197 28747
rect 14148 28716 14197 28744
rect 14148 28704 14154 28716
rect 14185 28713 14197 28716
rect 14231 28713 14243 28747
rect 14185 28707 14243 28713
rect 15654 28704 15660 28756
rect 15712 28744 15718 28756
rect 23474 28744 23480 28756
rect 15712 28716 23480 28744
rect 15712 28704 15718 28716
rect 23474 28704 23480 28716
rect 23532 28704 23538 28756
rect 26326 28704 26332 28756
rect 26384 28744 26390 28756
rect 31202 28744 31208 28756
rect 26384 28716 31208 28744
rect 26384 28704 26390 28716
rect 31202 28704 31208 28716
rect 31260 28704 31266 28756
rect 31389 28747 31447 28753
rect 31389 28713 31401 28747
rect 31435 28744 31447 28747
rect 32030 28744 32036 28756
rect 31435 28716 32036 28744
rect 31435 28713 31447 28716
rect 31389 28707 31447 28713
rect 32030 28704 32036 28716
rect 32088 28704 32094 28756
rect 33226 28744 33232 28756
rect 33187 28716 33232 28744
rect 33226 28704 33232 28716
rect 33284 28704 33290 28756
rect 18322 28636 18328 28688
rect 18380 28676 18386 28688
rect 18693 28679 18751 28685
rect 18693 28676 18705 28679
rect 18380 28648 18705 28676
rect 18380 28636 18386 28648
rect 18693 28645 18705 28648
rect 18739 28645 18751 28679
rect 20162 28676 20168 28688
rect 20123 28648 20168 28676
rect 18693 28639 18751 28645
rect 20162 28636 20168 28648
rect 20220 28636 20226 28688
rect 22830 28636 22836 28688
rect 22888 28676 22894 28688
rect 24302 28676 24308 28688
rect 22888 28648 24308 28676
rect 22888 28636 22894 28648
rect 24302 28636 24308 28648
rect 24360 28636 24366 28688
rect 29546 28676 29552 28688
rect 27908 28648 29552 28676
rect 14458 28568 14464 28620
rect 14516 28608 14522 28620
rect 27062 28608 27068 28620
rect 14516 28580 16068 28608
rect 14516 28568 14522 28580
rect 16040 28552 16068 28580
rect 23032 28580 26648 28608
rect 27023 28580 27068 28608
rect 9306 28543 9364 28549
rect 9306 28509 9318 28543
rect 9352 28509 9364 28543
rect 9306 28503 9364 28509
rect 9398 28500 9404 28552
rect 9456 28540 9462 28552
rect 9585 28543 9643 28549
rect 9456 28512 9501 28540
rect 9456 28500 9462 28512
rect 9585 28509 9597 28543
rect 9631 28540 9643 28543
rect 9674 28540 9680 28552
rect 9631 28512 9680 28540
rect 9631 28509 9643 28512
rect 9585 28503 9643 28509
rect 9674 28500 9680 28512
rect 9732 28500 9738 28552
rect 10134 28540 10140 28552
rect 10095 28512 10140 28540
rect 10134 28500 10140 28512
rect 10192 28500 10198 28552
rect 14369 28543 14427 28549
rect 14369 28509 14381 28543
rect 14415 28509 14427 28543
rect 14369 28503 14427 28509
rect 14645 28543 14703 28549
rect 14645 28509 14657 28543
rect 14691 28540 14703 28543
rect 15010 28540 15016 28552
rect 14691 28512 15016 28540
rect 14691 28509 14703 28512
rect 14645 28503 14703 28509
rect 1581 28475 1639 28481
rect 1581 28441 1593 28475
rect 1627 28472 1639 28475
rect 2130 28472 2136 28484
rect 1627 28444 2136 28472
rect 1627 28441 1639 28444
rect 1581 28435 1639 28441
rect 2130 28432 2136 28444
rect 2188 28432 2194 28484
rect 7276 28475 7334 28481
rect 7276 28441 7288 28475
rect 7322 28472 7334 28475
rect 8941 28475 8999 28481
rect 8941 28472 8953 28475
rect 7322 28444 8953 28472
rect 7322 28441 7334 28444
rect 7276 28435 7334 28441
rect 8941 28441 8953 28444
rect 8987 28441 8999 28475
rect 8941 28435 8999 28441
rect 8386 28404 8392 28416
rect 8347 28376 8392 28404
rect 8386 28364 8392 28376
rect 8444 28364 8450 28416
rect 10226 28404 10232 28416
rect 10187 28376 10232 28404
rect 10226 28364 10232 28376
rect 10284 28364 10290 28416
rect 14384 28404 14412 28503
rect 15010 28500 15016 28512
rect 15068 28500 15074 28552
rect 15749 28543 15807 28549
rect 15749 28540 15761 28543
rect 15304 28512 15761 28540
rect 14553 28475 14611 28481
rect 14553 28441 14565 28475
rect 14599 28472 14611 28475
rect 15194 28472 15200 28484
rect 14599 28444 15200 28472
rect 14599 28441 14611 28444
rect 14553 28435 14611 28441
rect 15194 28432 15200 28444
rect 15252 28432 15258 28484
rect 15304 28404 15332 28512
rect 15749 28509 15761 28512
rect 15795 28540 15807 28543
rect 15838 28540 15844 28552
rect 15795 28512 15844 28540
rect 15795 28509 15807 28512
rect 15749 28503 15807 28509
rect 15838 28500 15844 28512
rect 15896 28500 15902 28552
rect 16022 28540 16028 28552
rect 15983 28512 16028 28540
rect 16022 28500 16028 28512
rect 16080 28500 16086 28552
rect 16482 28540 16488 28552
rect 16443 28512 16488 28540
rect 16482 28500 16488 28512
rect 16540 28500 16546 28552
rect 19886 28500 19892 28552
rect 19944 28540 19950 28552
rect 20349 28543 20407 28549
rect 20349 28540 20361 28543
rect 19944 28512 20361 28540
rect 19944 28500 19950 28512
rect 20349 28509 20361 28512
rect 20395 28509 20407 28543
rect 20349 28503 20407 28509
rect 20441 28543 20499 28549
rect 20441 28509 20453 28543
rect 20487 28540 20499 28543
rect 20714 28540 20720 28552
rect 20487 28512 20720 28540
rect 20487 28509 20499 28512
rect 20441 28503 20499 28509
rect 20714 28500 20720 28512
rect 20772 28500 20778 28552
rect 21174 28500 21180 28552
rect 21232 28540 21238 28552
rect 23032 28549 23060 28580
rect 23017 28543 23075 28549
rect 23017 28540 23029 28543
rect 21232 28512 23029 28540
rect 21232 28500 21238 28512
rect 23017 28509 23029 28512
rect 23063 28509 23075 28543
rect 23017 28503 23075 28509
rect 25685 28543 25743 28549
rect 25685 28509 25697 28543
rect 25731 28540 25743 28543
rect 25731 28512 26556 28540
rect 25731 28509 25743 28512
rect 25685 28503 25743 28509
rect 15565 28475 15623 28481
rect 15565 28441 15577 28475
rect 15611 28472 15623 28475
rect 16730 28475 16788 28481
rect 16730 28472 16742 28475
rect 15611 28444 16742 28472
rect 15611 28441 15623 28444
rect 15565 28435 15623 28441
rect 16730 28441 16742 28444
rect 16776 28441 16788 28475
rect 16730 28435 16788 28441
rect 17218 28432 17224 28484
rect 17276 28472 17282 28484
rect 18325 28475 18383 28481
rect 18325 28472 18337 28475
rect 17276 28444 18337 28472
rect 17276 28432 17282 28444
rect 18325 28441 18337 28444
rect 18371 28441 18383 28475
rect 18325 28435 18383 28441
rect 18509 28475 18567 28481
rect 18509 28441 18521 28475
rect 18555 28472 18567 28475
rect 19610 28472 19616 28484
rect 18555 28444 19616 28472
rect 18555 28441 18567 28444
rect 18509 28435 18567 28441
rect 19610 28432 19616 28444
rect 19668 28432 19674 28484
rect 20165 28475 20223 28481
rect 20165 28441 20177 28475
rect 20211 28472 20223 28475
rect 20530 28472 20536 28484
rect 20211 28444 20536 28472
rect 20211 28441 20223 28444
rect 20165 28435 20223 28441
rect 20530 28432 20536 28444
rect 20588 28432 20594 28484
rect 25869 28475 25927 28481
rect 25869 28441 25881 28475
rect 25915 28472 25927 28475
rect 26326 28472 26332 28484
rect 25915 28444 26332 28472
rect 25915 28441 25927 28444
rect 25869 28435 25927 28441
rect 26326 28432 26332 28444
rect 26384 28432 26390 28484
rect 14384 28376 15332 28404
rect 15933 28407 15991 28413
rect 15933 28373 15945 28407
rect 15979 28404 15991 28407
rect 17586 28404 17592 28416
rect 15979 28376 17592 28404
rect 15979 28373 15991 28376
rect 15933 28367 15991 28373
rect 17586 28364 17592 28376
rect 17644 28404 17650 28416
rect 17865 28407 17923 28413
rect 17865 28404 17877 28407
rect 17644 28376 17877 28404
rect 17644 28364 17650 28376
rect 17865 28373 17877 28376
rect 17911 28373 17923 28407
rect 17865 28367 17923 28373
rect 23109 28407 23167 28413
rect 23109 28373 23121 28407
rect 23155 28404 23167 28407
rect 23198 28404 23204 28416
rect 23155 28376 23204 28404
rect 23155 28373 23167 28376
rect 23109 28367 23167 28373
rect 23198 28364 23204 28376
rect 23256 28364 23262 28416
rect 26053 28407 26111 28413
rect 26053 28373 26065 28407
rect 26099 28404 26111 28407
rect 26234 28404 26240 28416
rect 26099 28376 26240 28404
rect 26099 28373 26111 28376
rect 26053 28367 26111 28373
rect 26234 28364 26240 28376
rect 26292 28364 26298 28416
rect 26528 28413 26556 28512
rect 26513 28407 26571 28413
rect 26513 28373 26525 28407
rect 26559 28373 26571 28407
rect 26620 28404 26648 28580
rect 27062 28568 27068 28580
rect 27120 28568 27126 28620
rect 27338 28568 27344 28620
rect 27396 28608 27402 28620
rect 27908 28608 27936 28648
rect 27396 28580 27936 28608
rect 27396 28568 27402 28580
rect 26973 28543 27031 28549
rect 26973 28509 26985 28543
rect 27019 28540 27031 28543
rect 27246 28540 27252 28552
rect 27019 28512 27252 28540
rect 27019 28509 27031 28512
rect 26973 28503 27031 28509
rect 27246 28500 27252 28512
rect 27304 28500 27310 28552
rect 27706 28500 27712 28552
rect 27764 28540 27770 28552
rect 28184 28549 28212 28648
rect 29546 28636 29552 28648
rect 29604 28676 29610 28688
rect 30098 28676 30104 28688
rect 29604 28648 30104 28676
rect 29604 28636 29610 28648
rect 30098 28636 30104 28648
rect 30156 28636 30162 28688
rect 34698 28608 34704 28620
rect 34659 28580 34704 28608
rect 34698 28568 34704 28580
rect 34756 28568 34762 28620
rect 36630 28608 36636 28620
rect 36591 28580 36636 28608
rect 36630 28568 36636 28580
rect 36688 28568 36694 28620
rect 46290 28608 46296 28620
rect 46251 28580 46296 28608
rect 46290 28568 46296 28580
rect 46348 28568 46354 28620
rect 46474 28608 46480 28620
rect 46435 28580 46480 28608
rect 46474 28568 46480 28580
rect 46532 28568 46538 28620
rect 47486 28568 47492 28620
rect 47544 28608 47550 28620
rect 47670 28608 47676 28620
rect 47544 28580 47676 28608
rect 47544 28568 47550 28580
rect 47670 28568 47676 28580
rect 47728 28568 47734 28620
rect 48130 28608 48136 28620
rect 48091 28580 48136 28608
rect 48130 28568 48136 28580
rect 48188 28568 48194 28620
rect 27985 28543 28043 28549
rect 27985 28540 27997 28543
rect 27764 28512 27997 28540
rect 27764 28500 27770 28512
rect 27985 28509 27997 28512
rect 28031 28509 28043 28543
rect 27985 28503 28043 28509
rect 28077 28543 28135 28549
rect 28077 28509 28089 28543
rect 28123 28509 28135 28543
rect 28077 28503 28135 28509
rect 28169 28543 28227 28549
rect 28169 28509 28181 28543
rect 28215 28509 28227 28543
rect 28350 28540 28356 28552
rect 28311 28512 28356 28540
rect 28169 28503 28227 28509
rect 26881 28475 26939 28481
rect 26881 28441 26893 28475
rect 26927 28472 26939 28475
rect 27338 28472 27344 28484
rect 26927 28444 27344 28472
rect 26927 28441 26939 28444
rect 26881 28435 26939 28441
rect 27338 28432 27344 28444
rect 27396 28472 27402 28484
rect 28092 28472 28120 28503
rect 28350 28500 28356 28512
rect 28408 28500 28414 28552
rect 30374 28540 30380 28552
rect 30335 28512 30380 28540
rect 30374 28500 30380 28512
rect 30432 28500 30438 28552
rect 30561 28543 30619 28549
rect 30561 28509 30573 28543
rect 30607 28540 30619 28543
rect 31849 28543 31907 28549
rect 31849 28540 31861 28543
rect 30607 28512 31861 28540
rect 30607 28509 30619 28512
rect 30561 28503 30619 28509
rect 31849 28509 31861 28512
rect 31895 28540 31907 28543
rect 31938 28540 31944 28552
rect 31895 28512 31944 28540
rect 31895 28509 31907 28512
rect 31849 28503 31907 28509
rect 31938 28500 31944 28512
rect 31996 28540 32002 28552
rect 32582 28540 32588 28552
rect 31996 28512 32588 28540
rect 31996 28500 32002 28512
rect 32582 28500 32588 28512
rect 32640 28500 32646 28552
rect 33686 28540 33692 28552
rect 33647 28512 33692 28540
rect 33686 28500 33692 28512
rect 33744 28500 33750 28552
rect 34514 28500 34520 28552
rect 34572 28540 34578 28552
rect 34977 28543 35035 28549
rect 34977 28540 34989 28543
rect 34572 28512 34989 28540
rect 34572 28500 34578 28512
rect 34977 28509 34989 28512
rect 35023 28509 35035 28543
rect 34977 28503 35035 28509
rect 35894 28500 35900 28552
rect 35952 28540 35958 28552
rect 35989 28543 36047 28549
rect 35989 28540 36001 28543
rect 35952 28512 36001 28540
rect 35952 28500 35958 28512
rect 35989 28509 36001 28512
rect 36035 28509 36047 28543
rect 35989 28503 36047 28509
rect 31018 28472 31024 28484
rect 27396 28444 28120 28472
rect 30979 28444 31024 28472
rect 27396 28432 27402 28444
rect 31018 28432 31024 28444
rect 31076 28432 31082 28484
rect 31202 28472 31208 28484
rect 31163 28444 31208 28472
rect 31202 28432 31208 28444
rect 31260 28432 31266 28484
rect 31754 28432 31760 28484
rect 31812 28472 31818 28484
rect 32094 28475 32152 28481
rect 32094 28472 32106 28475
rect 31812 28444 32106 28472
rect 31812 28432 31818 28444
rect 32094 28441 32106 28444
rect 32140 28441 32152 28475
rect 33873 28475 33931 28481
rect 33873 28472 33885 28475
rect 32094 28435 32152 28441
rect 32784 28444 33885 28472
rect 27430 28404 27436 28416
rect 26620 28376 27436 28404
rect 26513 28367 26571 28373
rect 27430 28364 27436 28376
rect 27488 28364 27494 28416
rect 27706 28404 27712 28416
rect 27667 28376 27712 28404
rect 27706 28364 27712 28376
rect 27764 28364 27770 28416
rect 31220 28404 31248 28432
rect 32784 28404 32812 28444
rect 33873 28441 33885 28444
rect 33919 28441 33931 28475
rect 33873 28435 33931 28441
rect 36081 28475 36139 28481
rect 36081 28441 36093 28475
rect 36127 28472 36139 28475
rect 36817 28475 36875 28481
rect 36817 28472 36829 28475
rect 36127 28444 36829 28472
rect 36127 28441 36139 28444
rect 36081 28435 36139 28441
rect 36817 28441 36829 28444
rect 36863 28441 36875 28475
rect 38470 28472 38476 28484
rect 38431 28444 38476 28472
rect 36817 28435 36875 28441
rect 38470 28432 38476 28444
rect 38528 28432 38534 28484
rect 34054 28404 34060 28416
rect 31220 28376 32812 28404
rect 34015 28376 34060 28404
rect 34054 28364 34060 28376
rect 34112 28364 34118 28416
rect 47578 28364 47584 28416
rect 47636 28404 47642 28416
rect 47854 28404 47860 28416
rect 47636 28376 47860 28404
rect 47636 28364 47642 28376
rect 47854 28364 47860 28376
rect 47912 28364 47918 28416
rect 1104 28314 48852 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 48852 28314
rect 1104 28240 48852 28262
rect 2130 28200 2136 28212
rect 2091 28172 2136 28200
rect 2130 28160 2136 28172
rect 2188 28160 2194 28212
rect 6362 28160 6368 28212
rect 6420 28200 6426 28212
rect 12529 28203 12587 28209
rect 6420 28172 12434 28200
rect 6420 28160 6426 28172
rect 9401 28135 9459 28141
rect 9401 28101 9413 28135
rect 9447 28132 9459 28135
rect 12406 28132 12434 28172
rect 12529 28169 12541 28203
rect 12575 28200 12587 28203
rect 13078 28200 13084 28212
rect 12575 28172 13084 28200
rect 12575 28169 12587 28172
rect 12529 28163 12587 28169
rect 13078 28160 13084 28172
rect 13136 28160 13142 28212
rect 16022 28160 16028 28212
rect 16080 28200 16086 28212
rect 16761 28203 16819 28209
rect 16761 28200 16773 28203
rect 16080 28172 16773 28200
rect 16080 28160 16086 28172
rect 16761 28169 16773 28172
rect 16807 28169 16819 28203
rect 17494 28200 17500 28212
rect 17455 28172 17500 28200
rect 16761 28163 16819 28169
rect 17494 28160 17500 28172
rect 17552 28160 17558 28212
rect 48041 28203 48099 28209
rect 48041 28200 48053 28203
rect 17604 28172 48053 28200
rect 17604 28132 17632 28172
rect 48041 28169 48053 28172
rect 48087 28169 48099 28203
rect 48041 28163 48099 28169
rect 18414 28132 18420 28144
rect 9447 28104 11836 28132
rect 12406 28104 17632 28132
rect 18375 28104 18420 28132
rect 9447 28101 9459 28104
rect 9401 28095 9459 28101
rect 2038 28064 2044 28076
rect 1999 28036 2044 28064
rect 2038 28024 2044 28036
rect 2096 28024 2102 28076
rect 9669 28067 9727 28073
rect 9577 28057 9635 28063
rect 9577 28054 9589 28057
rect 9508 28026 9589 28054
rect 9508 27860 9536 28026
rect 9577 28023 9589 28026
rect 9623 28023 9635 28057
rect 9669 28033 9681 28067
rect 9715 28033 9727 28067
rect 9669 28027 9727 28033
rect 9577 28017 9635 28023
rect 9692 27996 9720 28027
rect 9766 28024 9772 28076
rect 9824 28070 9830 28076
rect 9861 28070 9919 28073
rect 9824 28067 9919 28070
rect 9824 28042 9873 28067
rect 9824 28024 9830 28042
rect 9861 28033 9873 28042
rect 9907 28033 9919 28067
rect 9861 28027 9919 28033
rect 9950 28024 9956 28076
rect 10008 28064 10014 28076
rect 10008 28036 10053 28064
rect 10008 28024 10014 28036
rect 10318 28024 10324 28076
rect 10376 28064 10382 28076
rect 11701 28067 11759 28073
rect 11701 28064 11713 28067
rect 10376 28036 11713 28064
rect 10376 28024 10382 28036
rect 11701 28033 11713 28036
rect 11747 28033 11759 28067
rect 11808 28064 11836 28104
rect 18414 28092 18420 28104
rect 18472 28092 18478 28144
rect 20162 28141 20168 28144
rect 20156 28132 20168 28141
rect 20123 28104 20168 28132
rect 20156 28095 20168 28104
rect 20162 28092 20168 28095
rect 20220 28092 20226 28144
rect 23198 28132 23204 28144
rect 23159 28104 23204 28132
rect 23198 28092 23204 28104
rect 23256 28092 23262 28144
rect 27240 28135 27298 28141
rect 27240 28101 27252 28135
rect 27286 28132 27298 28135
rect 27706 28132 27712 28144
rect 27286 28104 27712 28132
rect 27286 28101 27298 28104
rect 27240 28095 27298 28101
rect 27706 28092 27712 28104
rect 27764 28092 27770 28144
rect 27798 28092 27804 28144
rect 27856 28132 27862 28144
rect 33042 28132 33048 28144
rect 27856 28104 33048 28132
rect 27856 28092 27862 28104
rect 12713 28067 12771 28073
rect 12713 28064 12725 28067
rect 11808 28036 12725 28064
rect 11701 28027 11759 28033
rect 12713 28033 12725 28036
rect 12759 28033 12771 28067
rect 12986 28064 12992 28076
rect 12947 28036 12992 28064
rect 12713 28027 12771 28033
rect 12986 28024 12992 28036
rect 13044 28024 13050 28076
rect 15562 28064 15568 28076
rect 15523 28036 15568 28064
rect 15562 28024 15568 28036
rect 15620 28064 15626 28076
rect 16669 28067 16727 28073
rect 16669 28064 16681 28067
rect 15620 28036 16681 28064
rect 15620 28024 15626 28036
rect 16669 28033 16681 28036
rect 16715 28064 16727 28067
rect 17313 28067 17371 28073
rect 17313 28064 17325 28067
rect 16715 28036 17325 28064
rect 16715 28033 16727 28036
rect 16669 28027 16727 28033
rect 17313 28033 17325 28036
rect 17359 28033 17371 28067
rect 17313 28027 17371 28033
rect 18601 28067 18659 28073
rect 18601 28033 18613 28067
rect 18647 28064 18659 28067
rect 19334 28064 19340 28076
rect 18647 28036 19340 28064
rect 18647 28033 18659 28036
rect 18601 28027 18659 28033
rect 19334 28024 19340 28036
rect 19392 28064 19398 28076
rect 19889 28067 19947 28073
rect 19889 28064 19901 28067
rect 19392 28036 19901 28064
rect 19392 28024 19398 28036
rect 19889 28033 19901 28036
rect 19935 28064 19947 28067
rect 19978 28064 19984 28076
rect 19935 28036 19984 28064
rect 19935 28033 19947 28036
rect 19889 28027 19947 28033
rect 19978 28024 19984 28036
rect 20036 28024 20042 28076
rect 26050 28064 26056 28076
rect 26011 28036 26056 28064
rect 26050 28024 26056 28036
rect 26108 28024 26114 28076
rect 26142 28067 26200 28073
rect 26142 28033 26154 28067
rect 26188 28033 26200 28067
rect 26142 28027 26200 28033
rect 9692 27968 9904 27996
rect 9766 27860 9772 27872
rect 9508 27832 9772 27860
rect 9766 27820 9772 27832
rect 9824 27820 9830 27872
rect 9876 27860 9904 27968
rect 11146 27956 11152 28008
rect 11204 27996 11210 28008
rect 11609 27999 11667 28005
rect 11609 27996 11621 27999
rect 11204 27968 11621 27996
rect 11204 27956 11210 27968
rect 11609 27965 11621 27968
rect 11655 27965 11667 27999
rect 11609 27959 11667 27965
rect 15194 27956 15200 28008
rect 15252 27996 15258 28008
rect 15289 27999 15347 28005
rect 15289 27996 15301 27999
rect 15252 27968 15301 27996
rect 15252 27956 15258 27968
rect 15289 27965 15301 27968
rect 15335 27965 15347 27999
rect 17678 27996 17684 28008
rect 17639 27968 17684 27996
rect 15289 27959 15347 27965
rect 17678 27956 17684 27968
rect 17736 27956 17742 28008
rect 23017 27999 23075 28005
rect 23017 27965 23029 27999
rect 23063 27965 23075 27999
rect 23474 27996 23480 28008
rect 23435 27968 23480 27996
rect 23017 27959 23075 27965
rect 12069 27931 12127 27937
rect 12069 27897 12081 27931
rect 12115 27928 12127 27931
rect 12805 27931 12863 27937
rect 12805 27928 12817 27931
rect 12115 27900 12817 27928
rect 12115 27897 12127 27900
rect 12069 27891 12127 27897
rect 12805 27897 12817 27900
rect 12851 27897 12863 27931
rect 12805 27891 12863 27897
rect 12894 27888 12900 27940
rect 12952 27928 12958 27940
rect 23032 27928 23060 27959
rect 23474 27956 23480 27968
rect 23532 27956 23538 28008
rect 26157 27996 26185 28027
rect 26234 28024 26240 28076
rect 26292 28073 26298 28076
rect 26292 28064 26300 28073
rect 26421 28067 26479 28073
rect 26292 28036 26337 28064
rect 26292 28027 26300 28036
rect 26421 28033 26433 28067
rect 26467 28064 26479 28067
rect 28166 28064 28172 28076
rect 26467 28036 28172 28064
rect 26467 28033 26479 28036
rect 26421 28027 26479 28033
rect 26292 28024 26298 28027
rect 28166 28024 28172 28036
rect 28224 28024 28230 28076
rect 29380 28073 29408 28104
rect 33042 28092 33048 28104
rect 33100 28092 33106 28144
rect 29365 28067 29423 28073
rect 29365 28033 29377 28067
rect 29411 28033 29423 28067
rect 29365 28027 29423 28033
rect 29454 28067 29512 28073
rect 29454 28033 29466 28067
rect 29500 28033 29512 28067
rect 29454 28027 29512 28033
rect 26694 27996 26700 28008
rect 26157 27968 26700 27996
rect 26694 27956 26700 27968
rect 26752 27956 26758 28008
rect 26970 27996 26976 28008
rect 26931 27968 26976 27996
rect 26970 27956 26976 27968
rect 27028 27956 27034 28008
rect 29472 27996 29500 28027
rect 29546 28024 29552 28076
rect 29604 28064 29610 28076
rect 29730 28064 29736 28076
rect 29604 28036 29649 28064
rect 29691 28036 29736 28064
rect 29604 28024 29610 28036
rect 29730 28024 29736 28036
rect 29788 28024 29794 28076
rect 32030 28024 32036 28076
rect 32088 28064 32094 28076
rect 32841 28067 32899 28073
rect 32841 28064 32853 28067
rect 32088 28036 32853 28064
rect 32088 28024 32094 28036
rect 32841 28033 32853 28036
rect 32887 28033 32899 28067
rect 32841 28027 32899 28033
rect 34790 28024 34796 28076
rect 34848 28064 34854 28076
rect 35253 28067 35311 28073
rect 35253 28064 35265 28067
rect 34848 28036 35265 28064
rect 34848 28024 34854 28036
rect 35253 28033 35265 28036
rect 35299 28033 35311 28067
rect 35253 28027 35311 28033
rect 35345 28067 35403 28073
rect 35345 28033 35357 28067
rect 35391 28033 35403 28067
rect 35345 28027 35403 28033
rect 29914 27996 29920 28008
rect 29472 27968 29920 27996
rect 29914 27956 29920 27968
rect 29972 27956 29978 28008
rect 32582 27996 32588 28008
rect 32543 27968 32588 27996
rect 32582 27956 32588 27968
rect 32640 27956 32646 28008
rect 35360 27996 35388 28027
rect 35434 28024 35440 28076
rect 35492 28064 35498 28076
rect 35618 28064 35624 28076
rect 35492 28036 35537 28064
rect 35579 28036 35624 28064
rect 35492 28024 35498 28036
rect 35618 28024 35624 28036
rect 35676 28024 35682 28076
rect 47118 28024 47124 28076
rect 47176 28024 47182 28076
rect 47854 28064 47860 28076
rect 47815 28036 47860 28064
rect 47854 28024 47860 28036
rect 47912 28024 47918 28076
rect 33980 27968 35388 27996
rect 33980 27940 34008 27968
rect 12952 27900 12997 27928
rect 23032 27900 27016 27928
rect 12952 27888 12958 27900
rect 9950 27860 9956 27872
rect 9876 27832 9956 27860
rect 9950 27820 9956 27832
rect 10008 27820 10014 27872
rect 17586 27820 17592 27872
rect 17644 27860 17650 27872
rect 17681 27863 17739 27869
rect 17681 27860 17693 27863
rect 17644 27832 17693 27860
rect 17644 27820 17650 27832
rect 17681 27829 17693 27832
rect 17727 27829 17739 27863
rect 17681 27823 17739 27829
rect 20622 27820 20628 27872
rect 20680 27860 20686 27872
rect 21269 27863 21327 27869
rect 21269 27860 21281 27863
rect 20680 27832 21281 27860
rect 20680 27820 20686 27832
rect 21269 27829 21281 27832
rect 21315 27829 21327 27863
rect 21269 27823 21327 27829
rect 25777 27863 25835 27869
rect 25777 27829 25789 27863
rect 25823 27860 25835 27863
rect 26234 27860 26240 27872
rect 25823 27832 26240 27860
rect 25823 27829 25835 27832
rect 25777 27823 25835 27829
rect 26234 27820 26240 27832
rect 26292 27820 26298 27872
rect 26988 27860 27016 27900
rect 28074 27888 28080 27940
rect 28132 27928 28138 27940
rect 33962 27928 33968 27940
rect 28132 27900 31754 27928
rect 33923 27900 33968 27928
rect 28132 27888 28138 27900
rect 27706 27860 27712 27872
rect 26988 27832 27712 27860
rect 27706 27820 27712 27832
rect 27764 27860 27770 27872
rect 28353 27863 28411 27869
rect 28353 27860 28365 27863
rect 27764 27832 28365 27860
rect 27764 27820 27770 27832
rect 28353 27829 28365 27832
rect 28399 27829 28411 27863
rect 28353 27823 28411 27829
rect 29089 27863 29147 27869
rect 29089 27829 29101 27863
rect 29135 27860 29147 27863
rect 29638 27860 29644 27872
rect 29135 27832 29644 27860
rect 29135 27829 29147 27832
rect 29089 27823 29147 27829
rect 29638 27820 29644 27832
rect 29696 27820 29702 27872
rect 31726 27860 31754 27900
rect 33962 27888 33968 27900
rect 34020 27888 34026 27940
rect 35894 27928 35900 27940
rect 34900 27900 35900 27928
rect 34900 27860 34928 27900
rect 35894 27888 35900 27900
rect 35952 27888 35958 27940
rect 47136 27872 47164 28024
rect 31726 27832 34928 27860
rect 34977 27863 35035 27869
rect 34977 27829 34989 27863
rect 35023 27860 35035 27863
rect 35986 27860 35992 27872
rect 35023 27832 35992 27860
rect 35023 27829 35035 27832
rect 34977 27823 35035 27829
rect 35986 27820 35992 27832
rect 36044 27820 36050 27872
rect 47026 27860 47032 27872
rect 46987 27832 47032 27860
rect 47026 27820 47032 27832
rect 47084 27820 47090 27872
rect 47118 27820 47124 27872
rect 47176 27820 47182 27872
rect 1104 27770 48852 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 48852 27770
rect 1104 27696 48852 27718
rect 2038 27616 2044 27668
rect 2096 27656 2102 27668
rect 2590 27656 2596 27668
rect 2096 27628 2596 27656
rect 2096 27616 2102 27628
rect 2590 27616 2596 27628
rect 2648 27656 2654 27668
rect 17034 27656 17040 27668
rect 2648 27628 17040 27656
rect 2648 27616 2654 27628
rect 17034 27616 17040 27628
rect 17092 27616 17098 27668
rect 20533 27659 20591 27665
rect 20533 27625 20545 27659
rect 20579 27656 20591 27659
rect 20898 27656 20904 27668
rect 20579 27628 20904 27656
rect 20579 27625 20591 27628
rect 20533 27619 20591 27625
rect 20898 27616 20904 27628
rect 20956 27616 20962 27668
rect 27338 27656 27344 27668
rect 27299 27628 27344 27656
rect 27338 27616 27344 27628
rect 27396 27616 27402 27668
rect 27430 27616 27436 27668
rect 27488 27656 27494 27668
rect 28074 27656 28080 27668
rect 27488 27628 28080 27656
rect 27488 27616 27494 27628
rect 28074 27616 28080 27628
rect 28132 27616 28138 27668
rect 28169 27659 28227 27665
rect 28169 27625 28181 27659
rect 28215 27656 28227 27659
rect 28350 27656 28356 27668
rect 28215 27628 28356 27656
rect 28215 27625 28227 27628
rect 28169 27619 28227 27625
rect 28350 27616 28356 27628
rect 28408 27616 28414 27668
rect 28997 27659 29055 27665
rect 28997 27625 29009 27659
rect 29043 27656 29055 27659
rect 29730 27656 29736 27668
rect 29043 27628 29736 27656
rect 29043 27625 29055 27628
rect 28997 27619 29055 27625
rect 29730 27616 29736 27628
rect 29788 27616 29794 27668
rect 32030 27656 32036 27668
rect 31991 27628 32036 27656
rect 32030 27616 32036 27628
rect 32088 27616 32094 27668
rect 32324 27628 32536 27656
rect 9674 27548 9680 27600
rect 9732 27588 9738 27600
rect 10137 27591 10195 27597
rect 10137 27588 10149 27591
rect 9732 27560 10149 27588
rect 9732 27548 9738 27560
rect 10137 27557 10149 27560
rect 10183 27557 10195 27591
rect 11146 27588 11152 27600
rect 11107 27560 11152 27588
rect 10137 27551 10195 27557
rect 11146 27548 11152 27560
rect 11204 27548 11210 27600
rect 17589 27591 17647 27597
rect 17589 27557 17601 27591
rect 17635 27588 17647 27591
rect 17770 27588 17776 27600
rect 17635 27560 17776 27588
rect 17635 27557 17647 27560
rect 17589 27551 17647 27557
rect 17770 27548 17776 27560
rect 17828 27548 17834 27600
rect 20714 27588 20720 27600
rect 20675 27560 20720 27588
rect 20714 27548 20720 27560
rect 20772 27548 20778 27600
rect 24489 27591 24547 27597
rect 24489 27557 24501 27591
rect 24535 27588 24547 27591
rect 24854 27588 24860 27600
rect 24535 27560 24860 27588
rect 24535 27557 24547 27560
rect 24489 27551 24547 27557
rect 24854 27548 24860 27560
rect 24912 27588 24918 27600
rect 25590 27588 25596 27600
rect 24912 27560 25596 27588
rect 24912 27548 24918 27560
rect 25590 27548 25596 27560
rect 25648 27548 25654 27600
rect 30558 27548 30564 27600
rect 30616 27588 30622 27600
rect 32324 27588 32352 27628
rect 30616 27560 32352 27588
rect 32508 27588 32536 27628
rect 33134 27616 33140 27668
rect 33192 27656 33198 27668
rect 33505 27659 33563 27665
rect 33505 27656 33517 27659
rect 33192 27628 33517 27656
rect 33192 27616 33198 27628
rect 33505 27625 33517 27628
rect 33551 27625 33563 27659
rect 33505 27619 33563 27625
rect 35437 27659 35495 27665
rect 35437 27625 35449 27659
rect 35483 27656 35495 27659
rect 35618 27656 35624 27668
rect 35483 27628 35624 27656
rect 35483 27625 35495 27628
rect 35437 27619 35495 27625
rect 35618 27616 35624 27628
rect 35676 27616 35682 27668
rect 34790 27588 34796 27600
rect 32508 27560 34796 27588
rect 30616 27548 30622 27560
rect 34790 27548 34796 27560
rect 34848 27588 34854 27600
rect 35066 27588 35072 27600
rect 34848 27560 35072 27588
rect 34848 27548 34854 27560
rect 35066 27548 35072 27560
rect 35124 27548 35130 27600
rect 37277 27591 37335 27597
rect 37277 27588 37289 27591
rect 36924 27560 37289 27588
rect 1854 27520 1860 27532
rect 1815 27492 1860 27520
rect 1854 27480 1860 27492
rect 1912 27480 1918 27532
rect 9306 27480 9312 27532
rect 9364 27520 9370 27532
rect 9953 27523 10011 27529
rect 9953 27520 9965 27523
rect 9364 27492 9965 27520
rect 9364 27480 9370 27492
rect 9953 27489 9965 27492
rect 9999 27489 10011 27523
rect 9953 27483 10011 27489
rect 10689 27523 10747 27529
rect 10689 27489 10701 27523
rect 10735 27489 10747 27523
rect 12158 27520 12164 27532
rect 12119 27492 12164 27520
rect 10689 27483 10747 27489
rect 1394 27452 1400 27464
rect 1355 27424 1400 27452
rect 1394 27412 1400 27424
rect 1452 27412 1458 27464
rect 9030 27412 9036 27464
rect 9088 27452 9094 27464
rect 9861 27455 9919 27461
rect 9861 27452 9873 27455
rect 9088 27424 9873 27452
rect 9088 27412 9094 27424
rect 9861 27421 9873 27424
rect 9907 27452 9919 27455
rect 10318 27452 10324 27464
rect 9907 27424 10324 27452
rect 9907 27421 9919 27424
rect 9861 27415 9919 27421
rect 10318 27412 10324 27424
rect 10376 27452 10382 27464
rect 10704 27452 10732 27483
rect 12158 27480 12164 27492
rect 12216 27480 12222 27532
rect 24578 27480 24584 27532
rect 24636 27520 24642 27532
rect 24673 27523 24731 27529
rect 24673 27520 24685 27523
rect 24636 27492 24685 27520
rect 24636 27480 24642 27492
rect 24673 27489 24685 27492
rect 24719 27489 24731 27523
rect 34054 27520 34060 27532
rect 24673 27483 24731 27489
rect 26988 27492 29592 27520
rect 26988 27464 27016 27492
rect 12434 27461 12440 27464
rect 10376 27424 10732 27452
rect 10781 27455 10839 27461
rect 10376 27412 10382 27424
rect 10781 27421 10793 27455
rect 10827 27421 10839 27455
rect 10781 27415 10839 27421
rect 12428 27415 12440 27461
rect 12492 27452 12498 27464
rect 14829 27455 14887 27461
rect 12492 27424 12528 27452
rect 1581 27387 1639 27393
rect 1581 27353 1593 27387
rect 1627 27384 1639 27387
rect 2130 27384 2136 27396
rect 1627 27356 2136 27384
rect 1627 27353 1639 27356
rect 1581 27347 1639 27353
rect 2130 27344 2136 27356
rect 2188 27344 2194 27396
rect 9493 27387 9551 27393
rect 9493 27353 9505 27387
rect 9539 27384 9551 27387
rect 10226 27384 10232 27396
rect 9539 27356 10232 27384
rect 9539 27353 9551 27356
rect 9493 27347 9551 27353
rect 10226 27344 10232 27356
rect 10284 27344 10290 27396
rect 10502 27344 10508 27396
rect 10560 27384 10566 27396
rect 10796 27384 10824 27415
rect 12434 27412 12440 27415
rect 12492 27412 12498 27424
rect 14829 27421 14841 27455
rect 14875 27452 14887 27455
rect 16482 27452 16488 27464
rect 14875 27424 16488 27452
rect 14875 27421 14887 27424
rect 14829 27415 14887 27421
rect 16482 27412 16488 27424
rect 16540 27412 16546 27464
rect 17402 27452 17408 27464
rect 17363 27424 17408 27452
rect 17402 27412 17408 27424
rect 17460 27412 17466 27464
rect 20257 27455 20315 27461
rect 20257 27421 20269 27455
rect 20303 27452 20315 27455
rect 20622 27452 20628 27464
rect 20303 27424 20628 27452
rect 20303 27421 20315 27424
rect 20257 27415 20315 27421
rect 20622 27412 20628 27424
rect 20680 27412 20686 27464
rect 22465 27455 22523 27461
rect 22465 27421 22477 27455
rect 22511 27452 22523 27455
rect 24397 27455 24455 27461
rect 22511 27424 24348 27452
rect 22511 27421 22523 27424
rect 22465 27415 22523 27421
rect 15102 27393 15108 27396
rect 15096 27384 15108 27393
rect 10560 27356 10824 27384
rect 15063 27356 15108 27384
rect 10560 27344 10566 27356
rect 15096 27347 15108 27356
rect 15102 27344 15108 27347
rect 15160 27344 15166 27396
rect 22732 27387 22790 27393
rect 22732 27353 22744 27387
rect 22778 27384 22790 27387
rect 22922 27384 22928 27396
rect 22778 27356 22928 27384
rect 22778 27353 22790 27356
rect 22732 27347 22790 27353
rect 22922 27344 22928 27356
rect 22980 27344 22986 27396
rect 24320 27384 24348 27424
rect 24397 27421 24409 27455
rect 24443 27452 24455 27455
rect 24762 27452 24768 27464
rect 24443 27424 24768 27452
rect 24443 27421 24455 27424
rect 24397 27415 24455 27421
rect 24762 27412 24768 27424
rect 24820 27412 24826 27464
rect 25961 27455 26019 27461
rect 25961 27421 25973 27455
rect 26007 27452 26019 27455
rect 26786 27452 26792 27464
rect 26007 27424 26792 27452
rect 26007 27421 26019 27424
rect 25961 27415 26019 27421
rect 25976 27384 26004 27415
rect 26786 27412 26792 27424
rect 26844 27452 26850 27464
rect 26970 27452 26976 27464
rect 26844 27424 26976 27452
rect 26844 27412 26850 27424
rect 26970 27412 26976 27424
rect 27028 27412 27034 27464
rect 27062 27412 27068 27464
rect 27120 27452 27126 27464
rect 28626 27452 28632 27464
rect 27120 27424 28632 27452
rect 27120 27412 27126 27424
rect 28626 27412 28632 27424
rect 28684 27412 28690 27464
rect 29564 27461 29592 27492
rect 32600 27492 34060 27520
rect 29549 27455 29607 27461
rect 29549 27421 29561 27455
rect 29595 27421 29607 27455
rect 29549 27415 29607 27421
rect 29638 27412 29644 27464
rect 29696 27452 29702 27464
rect 29805 27455 29863 27461
rect 29805 27452 29817 27455
rect 29696 27424 29817 27452
rect 29696 27412 29702 27424
rect 29805 27421 29817 27424
rect 29851 27421 29863 27455
rect 29805 27415 29863 27421
rect 32289 27455 32347 27461
rect 32514 27455 32572 27461
rect 32289 27421 32301 27455
rect 32335 27452 32347 27455
rect 32335 27421 32352 27452
rect 32289 27415 32352 27421
rect 26234 27393 26240 27396
rect 26228 27384 26240 27393
rect 24320 27356 26004 27384
rect 26195 27356 26240 27384
rect 26228 27347 26240 27356
rect 26234 27344 26240 27347
rect 26292 27344 26298 27396
rect 27706 27344 27712 27396
rect 27764 27384 27770 27396
rect 27801 27387 27859 27393
rect 27801 27384 27813 27387
rect 27764 27356 27813 27384
rect 27764 27344 27770 27356
rect 27801 27353 27813 27356
rect 27847 27353 27859 27387
rect 27801 27347 27859 27353
rect 27985 27387 28043 27393
rect 27985 27353 27997 27387
rect 28031 27384 28043 27387
rect 28813 27387 28871 27393
rect 28813 27384 28825 27387
rect 28031 27356 28825 27384
rect 28031 27353 28043 27356
rect 27985 27347 28043 27353
rect 28813 27353 28825 27356
rect 28859 27384 28871 27387
rect 31202 27384 31208 27396
rect 28859 27356 31208 27384
rect 28859 27353 28871 27356
rect 28813 27347 28871 27353
rect 31202 27344 31208 27356
rect 31260 27344 31266 27396
rect 9214 27276 9220 27328
rect 9272 27316 9278 27328
rect 10870 27316 10876 27328
rect 9272 27288 10876 27316
rect 9272 27276 9278 27288
rect 10870 27276 10876 27288
rect 10928 27276 10934 27328
rect 13541 27319 13599 27325
rect 13541 27285 13553 27319
rect 13587 27316 13599 27319
rect 14182 27316 14188 27328
rect 13587 27288 14188 27316
rect 13587 27285 13599 27288
rect 13541 27279 13599 27285
rect 14182 27276 14188 27288
rect 14240 27276 14246 27328
rect 15194 27276 15200 27328
rect 15252 27316 15258 27328
rect 16209 27319 16267 27325
rect 16209 27316 16221 27319
rect 15252 27288 16221 27316
rect 15252 27276 15258 27288
rect 16209 27285 16221 27288
rect 16255 27285 16267 27319
rect 16209 27279 16267 27285
rect 17678 27276 17684 27328
rect 17736 27316 17742 27328
rect 23198 27316 23204 27328
rect 17736 27288 23204 27316
rect 17736 27276 17742 27288
rect 23198 27276 23204 27288
rect 23256 27316 23262 27328
rect 23845 27319 23903 27325
rect 23845 27316 23857 27319
rect 23256 27288 23857 27316
rect 23256 27276 23262 27288
rect 23845 27285 23857 27288
rect 23891 27285 23903 27319
rect 24670 27316 24676 27328
rect 24631 27288 24676 27316
rect 23845 27279 23903 27285
rect 24670 27276 24676 27288
rect 24728 27276 24734 27328
rect 28626 27276 28632 27328
rect 28684 27316 28690 27328
rect 30929 27319 30987 27325
rect 30929 27316 30941 27319
rect 28684 27288 30941 27316
rect 28684 27276 28690 27288
rect 30929 27285 30941 27288
rect 30975 27285 30987 27319
rect 32324 27316 32352 27415
rect 32398 27449 32456 27455
rect 32398 27442 32410 27449
rect 32444 27442 32456 27449
rect 32398 27390 32404 27442
rect 32456 27390 32462 27442
rect 32514 27421 32526 27455
rect 32560 27452 32572 27455
rect 32600 27452 32628 27492
rect 34054 27480 34060 27492
rect 34112 27480 34118 27532
rect 34514 27480 34520 27532
rect 34572 27520 34578 27532
rect 34572 27492 35296 27520
rect 34572 27480 34578 27492
rect 32560 27424 32628 27452
rect 32677 27455 32735 27461
rect 32560 27421 32572 27424
rect 32514 27415 32572 27421
rect 32677 27421 32689 27455
rect 32723 27452 32735 27455
rect 32766 27452 32772 27464
rect 32723 27424 32772 27452
rect 32723 27421 32735 27424
rect 32677 27415 32735 27421
rect 32766 27412 32772 27424
rect 32824 27412 32830 27464
rect 35268 27461 35296 27492
rect 35253 27455 35311 27461
rect 32876 27424 35020 27452
rect 32876 27316 32904 27424
rect 33137 27387 33195 27393
rect 33137 27353 33149 27387
rect 33183 27353 33195 27387
rect 33137 27347 33195 27353
rect 32324 27288 32904 27316
rect 33152 27316 33180 27347
rect 33318 27344 33324 27396
rect 33376 27384 33382 27396
rect 33376 27356 33421 27384
rect 33376 27344 33382 27356
rect 34698 27316 34704 27328
rect 33152 27288 34704 27316
rect 30929 27279 30987 27285
rect 34698 27276 34704 27288
rect 34756 27276 34762 27328
rect 34992 27316 35020 27424
rect 35253 27421 35265 27455
rect 35299 27421 35311 27455
rect 35253 27415 35311 27421
rect 35342 27412 35348 27464
rect 35400 27452 35406 27464
rect 35897 27455 35955 27461
rect 35897 27452 35909 27455
rect 35400 27424 35909 27452
rect 35400 27412 35406 27424
rect 35897 27421 35909 27424
rect 35943 27421 35955 27455
rect 35897 27415 35955 27421
rect 35986 27412 35992 27464
rect 36044 27452 36050 27464
rect 36153 27455 36211 27461
rect 36153 27452 36165 27455
rect 36044 27424 36165 27452
rect 36044 27412 36050 27424
rect 36153 27421 36165 27424
rect 36199 27421 36211 27455
rect 36924 27452 36952 27560
rect 37277 27557 37289 27560
rect 37323 27588 37335 27591
rect 38102 27588 38108 27600
rect 37323 27560 38108 27588
rect 37323 27557 37335 27560
rect 37277 27551 37335 27557
rect 38102 27548 38108 27560
rect 38160 27548 38166 27600
rect 46293 27523 46351 27529
rect 46293 27489 46305 27523
rect 46339 27520 46351 27523
rect 47026 27520 47032 27532
rect 46339 27492 47032 27520
rect 46339 27489 46351 27492
rect 46293 27483 46351 27489
rect 47026 27480 47032 27492
rect 47084 27480 47090 27532
rect 48133 27523 48191 27529
rect 48133 27489 48145 27523
rect 48179 27520 48191 27523
rect 48222 27520 48228 27532
rect 48179 27492 48228 27520
rect 48179 27489 48191 27492
rect 48133 27483 48191 27489
rect 48222 27480 48228 27492
rect 48280 27480 48286 27532
rect 36153 27415 36211 27421
rect 36740 27424 36952 27452
rect 35069 27387 35127 27393
rect 35069 27353 35081 27387
rect 35115 27384 35127 27387
rect 36740 27384 36768 27424
rect 35115 27356 36768 27384
rect 46477 27387 46535 27393
rect 35115 27353 35127 27356
rect 35069 27347 35127 27353
rect 46477 27353 46489 27387
rect 46523 27384 46535 27387
rect 46658 27384 46664 27396
rect 46523 27356 46664 27384
rect 46523 27353 46535 27356
rect 46477 27347 46535 27353
rect 46658 27344 46664 27356
rect 46716 27344 46722 27396
rect 46934 27316 46940 27328
rect 34992 27288 46940 27316
rect 46934 27276 46940 27288
rect 46992 27276 46998 27328
rect 1104 27226 48852 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 48852 27226
rect 1104 27152 48852 27174
rect 2130 27112 2136 27124
rect 2091 27084 2136 27112
rect 2130 27072 2136 27084
rect 2188 27072 2194 27124
rect 9490 27072 9496 27124
rect 9548 27112 9554 27124
rect 9585 27115 9643 27121
rect 9585 27112 9597 27115
rect 9548 27084 9597 27112
rect 9548 27072 9554 27084
rect 9585 27081 9597 27084
rect 9631 27081 9643 27115
rect 10318 27112 10324 27124
rect 9585 27075 9643 27081
rect 9981 27084 10324 27112
rect 1394 27004 1400 27056
rect 1452 27044 1458 27056
rect 1452 27016 2912 27044
rect 1452 27004 1458 27016
rect 2884 26985 2912 27016
rect 9981 26991 10009 27084
rect 10318 27072 10324 27084
rect 10376 27072 10382 27124
rect 15378 27112 15384 27124
rect 14476 27084 15384 27112
rect 10410 27004 10416 27056
rect 10468 27044 10474 27056
rect 10781 27047 10839 27053
rect 10781 27044 10793 27047
rect 10468 27016 10793 27044
rect 10468 27004 10474 27016
rect 10781 27013 10793 27016
rect 10827 27013 10839 27047
rect 14182 27044 14188 27056
rect 14143 27016 14188 27044
rect 10781 27007 10839 27013
rect 14182 27004 14188 27016
rect 14240 27004 14246 27056
rect 2041 26979 2099 26985
rect 2041 26945 2053 26979
rect 2087 26945 2099 26979
rect 2041 26939 2099 26945
rect 2869 26979 2927 26985
rect 2869 26945 2881 26979
rect 2915 26945 2927 26979
rect 8662 26976 8668 26988
rect 8623 26948 8668 26976
rect 2869 26939 2927 26945
rect 2056 26908 2084 26939
rect 8662 26936 8668 26948
rect 8720 26936 8726 26988
rect 8846 26976 8852 26988
rect 8807 26948 8852 26976
rect 8846 26936 8852 26948
rect 8904 26936 8910 26988
rect 9030 26976 9036 26988
rect 8991 26948 9036 26976
rect 9030 26936 9036 26948
rect 9088 26936 9094 26988
rect 9966 26985 10024 26991
rect 9861 26979 9919 26985
rect 9861 26945 9873 26979
rect 9907 26945 9919 26979
rect 9966 26951 9978 26985
rect 10012 26951 10024 26985
rect 9966 26945 10024 26951
rect 10066 26979 10124 26985
rect 10066 26945 10078 26979
rect 10112 26945 10124 26979
rect 9861 26939 9919 26945
rect 10066 26939 10124 26945
rect 10229 26979 10287 26985
rect 10229 26945 10241 26979
rect 10275 26976 10287 26979
rect 10428 26976 10456 27004
rect 10686 26976 10692 26988
rect 10275 26948 10456 26976
rect 10647 26948 10692 26976
rect 10275 26945 10287 26948
rect 10229 26939 10287 26945
rect 2498 26908 2504 26920
rect 2056 26880 2504 26908
rect 2498 26868 2504 26880
rect 2556 26908 2562 26920
rect 8941 26911 8999 26917
rect 2556 26880 5212 26908
rect 2556 26868 2562 26880
rect 2314 26800 2320 26852
rect 2372 26840 2378 26852
rect 5184 26840 5212 26880
rect 8941 26877 8953 26911
rect 8987 26908 8999 26911
rect 9122 26908 9128 26920
rect 8987 26880 9128 26908
rect 8987 26877 8999 26880
rect 8941 26871 8999 26877
rect 9122 26868 9128 26880
rect 9180 26908 9186 26920
rect 9876 26908 9904 26939
rect 9180 26880 9904 26908
rect 10081 26908 10109 26939
rect 10686 26936 10692 26948
rect 10744 26936 10750 26988
rect 10870 26976 10876 26988
rect 10831 26948 10876 26976
rect 10870 26936 10876 26948
rect 10928 26936 10934 26988
rect 14476 26976 14504 27084
rect 15378 27072 15384 27084
rect 15436 27072 15442 27124
rect 22922 27112 22928 27124
rect 22883 27084 22928 27112
rect 22922 27072 22928 27084
rect 22980 27072 22986 27124
rect 24854 27112 24860 27124
rect 23308 27084 24860 27112
rect 14550 27004 14556 27056
rect 14608 27044 14614 27056
rect 15105 27047 15163 27053
rect 15105 27044 15117 27047
rect 14608 27016 15117 27044
rect 14608 27004 14614 27016
rect 15105 27013 15117 27016
rect 15151 27013 15163 27047
rect 15105 27007 15163 27013
rect 14829 26979 14887 26985
rect 14829 26976 14841 26979
rect 14476 26948 14841 26976
rect 14829 26945 14841 26948
rect 14875 26945 14887 26979
rect 19518 26976 19524 26988
rect 14829 26939 14887 26945
rect 14936 26948 19524 26976
rect 10594 26908 10600 26920
rect 10081 26880 10600 26908
rect 9180 26868 9186 26880
rect 9674 26840 9680 26852
rect 2372 26812 2774 26840
rect 5184 26812 9680 26840
rect 2372 26800 2378 26812
rect 1394 26732 1400 26784
rect 1452 26772 1458 26784
rect 1581 26775 1639 26781
rect 1581 26772 1593 26775
rect 1452 26744 1593 26772
rect 1452 26732 1458 26744
rect 1581 26741 1593 26744
rect 1627 26741 1639 26775
rect 2746 26772 2774 26812
rect 9674 26800 9680 26812
rect 9732 26800 9738 26852
rect 9784 26840 9812 26880
rect 10594 26868 10600 26880
rect 10652 26868 10658 26920
rect 10704 26908 10732 26936
rect 14936 26908 14964 26948
rect 19518 26936 19524 26948
rect 19576 26936 19582 26988
rect 23198 26976 23204 26988
rect 23159 26948 23204 26976
rect 23198 26936 23204 26948
rect 23256 26936 23262 26988
rect 23308 26985 23336 27084
rect 24854 27072 24860 27084
rect 24912 27072 24918 27124
rect 30558 27112 30564 27124
rect 24964 27084 30564 27112
rect 24670 27044 24676 27056
rect 23400 27016 24676 27044
rect 23400 26985 23428 27016
rect 24670 27004 24676 27016
rect 24728 27004 24734 27056
rect 24762 27004 24768 27056
rect 24820 27044 24826 27056
rect 24964 27044 24992 27084
rect 30558 27072 30564 27084
rect 30616 27072 30622 27124
rect 34698 27072 34704 27124
rect 34756 27112 34762 27124
rect 36078 27112 36084 27124
rect 34756 27084 36084 27112
rect 34756 27072 34762 27084
rect 36078 27072 36084 27084
rect 36136 27072 36142 27124
rect 24820 27016 24992 27044
rect 24820 27004 24826 27016
rect 33686 27004 33692 27056
rect 33744 27044 33750 27056
rect 46382 27044 46388 27056
rect 33744 27016 46388 27044
rect 33744 27004 33750 27016
rect 46382 27004 46388 27016
rect 46440 27004 46446 27056
rect 23293 26979 23351 26985
rect 23293 26945 23305 26979
rect 23339 26945 23351 26979
rect 23293 26939 23351 26945
rect 23385 26979 23443 26985
rect 23385 26945 23397 26979
rect 23431 26945 23443 26979
rect 23385 26939 23443 26945
rect 23569 26979 23627 26985
rect 23569 26945 23581 26979
rect 23615 26945 23627 26979
rect 27062 26976 27068 26988
rect 27023 26948 27068 26976
rect 23569 26939 23627 26945
rect 10704 26880 14964 26908
rect 15010 26868 15016 26920
rect 15068 26908 15074 26920
rect 15105 26911 15163 26917
rect 15105 26908 15117 26911
rect 15068 26880 15117 26908
rect 15068 26868 15074 26880
rect 15105 26877 15117 26880
rect 15151 26877 15163 26911
rect 15105 26871 15163 26877
rect 20990 26868 20996 26920
rect 21048 26908 21054 26920
rect 23584 26908 23612 26939
rect 27062 26936 27068 26948
rect 27120 26936 27126 26988
rect 32674 26976 32680 26988
rect 32635 26948 32680 26976
rect 32674 26936 32680 26948
rect 32732 26936 32738 26988
rect 32769 26979 32827 26985
rect 32769 26945 32781 26979
rect 32815 26945 32827 26979
rect 32769 26939 32827 26945
rect 27246 26908 27252 26920
rect 21048 26880 23612 26908
rect 27207 26880 27252 26908
rect 21048 26868 21054 26880
rect 27246 26868 27252 26880
rect 27304 26868 27310 26920
rect 28074 26908 28080 26920
rect 28035 26880 28080 26908
rect 28074 26868 28080 26880
rect 28132 26868 28138 26920
rect 29733 26911 29791 26917
rect 29733 26877 29745 26911
rect 29779 26877 29791 26911
rect 29914 26908 29920 26920
rect 29875 26880 29920 26908
rect 29733 26871 29791 26877
rect 9784 26812 9996 26840
rect 7558 26772 7564 26784
rect 2746 26744 7564 26772
rect 1581 26735 1639 26741
rect 7558 26732 7564 26744
rect 7616 26732 7622 26784
rect 9125 26775 9183 26781
rect 9125 26741 9137 26775
rect 9171 26772 9183 26775
rect 9858 26772 9864 26784
rect 9171 26744 9864 26772
rect 9171 26741 9183 26744
rect 9125 26735 9183 26741
rect 9858 26732 9864 26744
rect 9916 26732 9922 26784
rect 9968 26772 9996 26812
rect 10042 26800 10048 26852
rect 10100 26840 10106 26852
rect 26326 26840 26332 26852
rect 10100 26812 26332 26840
rect 10100 26800 10106 26812
rect 26326 26800 26332 26812
rect 26384 26800 26390 26852
rect 26418 26800 26424 26852
rect 26476 26840 26482 26852
rect 29748 26840 29776 26871
rect 29914 26868 29920 26880
rect 29972 26868 29978 26920
rect 31573 26911 31631 26917
rect 31573 26877 31585 26911
rect 31619 26908 31631 26911
rect 32784 26908 32812 26939
rect 32858 26936 32864 26988
rect 32916 26976 32922 26988
rect 33045 26979 33103 26985
rect 32916 26948 32961 26976
rect 32916 26936 32922 26948
rect 33045 26945 33057 26979
rect 33091 26976 33103 26979
rect 33134 26976 33140 26988
rect 33091 26948 33140 26976
rect 33091 26945 33103 26948
rect 33045 26939 33103 26945
rect 33134 26936 33140 26948
rect 33192 26936 33198 26988
rect 33965 26979 34023 26985
rect 33965 26976 33977 26979
rect 33244 26948 33977 26976
rect 32950 26908 32956 26920
rect 31619 26880 32536 26908
rect 32784 26880 32956 26908
rect 31619 26877 31631 26880
rect 31573 26871 31631 26877
rect 26476 26812 29776 26840
rect 26476 26800 26482 26812
rect 10502 26772 10508 26784
rect 9968 26744 10508 26772
rect 10502 26732 10508 26744
rect 10560 26732 10566 26784
rect 14090 26732 14096 26784
rect 14148 26772 14154 26784
rect 14274 26772 14280 26784
rect 14148 26744 14280 26772
rect 14148 26732 14154 26744
rect 14274 26732 14280 26744
rect 14332 26732 14338 26784
rect 14921 26775 14979 26781
rect 14921 26741 14933 26775
rect 14967 26772 14979 26775
rect 15102 26772 15108 26784
rect 14967 26744 15108 26772
rect 14967 26741 14979 26744
rect 14921 26735 14979 26741
rect 15102 26732 15108 26744
rect 15160 26732 15166 26784
rect 21082 26732 21088 26784
rect 21140 26772 21146 26784
rect 32214 26772 32220 26784
rect 21140 26744 32220 26772
rect 21140 26732 21146 26744
rect 32214 26732 32220 26744
rect 32272 26732 32278 26784
rect 32398 26772 32404 26784
rect 32359 26744 32404 26772
rect 32398 26732 32404 26744
rect 32456 26732 32462 26784
rect 32508 26772 32536 26880
rect 32950 26868 32956 26880
rect 33008 26908 33014 26920
rect 33244 26908 33272 26948
rect 33965 26945 33977 26948
rect 34011 26945 34023 26979
rect 33965 26939 34023 26945
rect 34057 26979 34115 26985
rect 34057 26945 34069 26979
rect 34103 26945 34115 26979
rect 34057 26939 34115 26945
rect 34149 26979 34207 26985
rect 34149 26945 34161 26979
rect 34195 26945 34207 26979
rect 34330 26976 34336 26988
rect 34291 26948 34336 26976
rect 34149 26939 34207 26945
rect 34072 26908 34100 26939
rect 33008 26880 33272 26908
rect 33520 26880 34100 26908
rect 33008 26868 33014 26880
rect 33226 26800 33232 26852
rect 33284 26840 33290 26852
rect 33520 26840 33548 26880
rect 34164 26840 34192 26939
rect 34330 26936 34336 26948
rect 34388 26936 34394 26988
rect 35066 26976 35072 26988
rect 35027 26948 35072 26976
rect 35066 26936 35072 26948
rect 35124 26936 35130 26988
rect 35161 26979 35219 26985
rect 35161 26945 35173 26979
rect 35207 26945 35219 26979
rect 35161 26939 35219 26945
rect 35253 26979 35311 26985
rect 35253 26945 35265 26979
rect 35299 26945 35311 26979
rect 35253 26939 35311 26945
rect 35437 26979 35495 26985
rect 35437 26945 35449 26979
rect 35483 26945 35495 26979
rect 35437 26939 35495 26945
rect 35897 26979 35955 26985
rect 35897 26945 35909 26979
rect 35943 26976 35955 26979
rect 35986 26976 35992 26988
rect 35943 26948 35992 26976
rect 35943 26945 35955 26948
rect 35897 26939 35955 26945
rect 34238 26868 34244 26920
rect 34296 26908 34302 26920
rect 35176 26908 35204 26939
rect 34296 26880 35204 26908
rect 34296 26868 34302 26880
rect 35268 26840 35296 26939
rect 35452 26908 35480 26939
rect 35986 26936 35992 26948
rect 36044 26936 36050 26988
rect 36078 26936 36084 26988
rect 36136 26976 36142 26988
rect 36136 26948 36181 26976
rect 36136 26936 36142 26948
rect 36265 26911 36323 26917
rect 36265 26908 36277 26911
rect 35452 26880 36277 26908
rect 36265 26877 36277 26880
rect 36311 26877 36323 26911
rect 36265 26871 36323 26877
rect 35526 26840 35532 26852
rect 33284 26812 33548 26840
rect 33612 26812 35532 26840
rect 33284 26800 33290 26812
rect 32766 26772 32772 26784
rect 32508 26744 32772 26772
rect 32766 26732 32772 26744
rect 32824 26732 32830 26784
rect 32858 26732 32864 26784
rect 32916 26772 32922 26784
rect 33612 26772 33640 26812
rect 35526 26800 35532 26812
rect 35584 26800 35590 26852
rect 32916 26744 33640 26772
rect 33689 26775 33747 26781
rect 32916 26732 32922 26744
rect 33689 26741 33701 26775
rect 33735 26772 33747 26775
rect 34606 26772 34612 26784
rect 33735 26744 34612 26772
rect 33735 26741 33747 26744
rect 33689 26735 33747 26741
rect 34606 26732 34612 26744
rect 34664 26732 34670 26784
rect 34793 26775 34851 26781
rect 34793 26741 34805 26775
rect 34839 26772 34851 26775
rect 35434 26772 35440 26784
rect 34839 26744 35440 26772
rect 34839 26741 34851 26744
rect 34793 26735 34851 26741
rect 35434 26732 35440 26744
rect 35492 26732 35498 26784
rect 1104 26682 48852 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 48852 26682
rect 1104 26608 48852 26630
rect 6178 26568 6184 26580
rect 6139 26540 6184 26568
rect 6178 26528 6184 26540
rect 6236 26528 6242 26580
rect 9766 26568 9772 26580
rect 8266 26540 9536 26568
rect 9727 26540 9772 26568
rect 6641 26503 6699 26509
rect 6641 26469 6653 26503
rect 6687 26500 6699 26503
rect 8266 26500 8294 26540
rect 6687 26472 8294 26500
rect 6687 26469 6699 26472
rect 6641 26463 6699 26469
rect 9306 26460 9312 26512
rect 9364 26460 9370 26512
rect 9508 26500 9536 26540
rect 9766 26528 9772 26540
rect 9824 26528 9830 26580
rect 10428 26540 19472 26568
rect 10428 26500 10456 26540
rect 10594 26500 10600 26512
rect 9508 26472 10456 26500
rect 10555 26472 10600 26500
rect 10594 26460 10600 26472
rect 10652 26460 10658 26512
rect 12066 26500 12072 26512
rect 12027 26472 12072 26500
rect 12066 26460 12072 26472
rect 12124 26460 12130 26512
rect 14093 26503 14151 26509
rect 14093 26469 14105 26503
rect 14139 26500 14151 26503
rect 14826 26500 14832 26512
rect 14139 26472 14832 26500
rect 14139 26469 14151 26472
rect 14093 26463 14151 26469
rect 14826 26460 14832 26472
rect 14884 26460 14890 26512
rect 18138 26460 18144 26512
rect 18196 26460 18202 26512
rect 1394 26432 1400 26444
rect 1355 26404 1400 26432
rect 1394 26392 1400 26404
rect 1452 26392 1458 26444
rect 2774 26392 2780 26444
rect 2832 26432 2838 26444
rect 6270 26432 6276 26444
rect 2832 26404 2877 26432
rect 6231 26404 6276 26432
rect 2832 26392 2838 26404
rect 6270 26392 6276 26404
rect 6328 26392 6334 26444
rect 7558 26392 7564 26444
rect 7616 26432 7622 26444
rect 9214 26432 9220 26444
rect 7616 26404 9220 26432
rect 7616 26392 7622 26404
rect 9214 26392 9220 26404
rect 9272 26392 9278 26444
rect 9324 26432 9352 26460
rect 9324 26404 9536 26432
rect 6454 26364 6460 26376
rect 6415 26336 6460 26364
rect 6454 26324 6460 26336
rect 6512 26324 6518 26376
rect 9508 26373 9536 26404
rect 9383 26367 9441 26373
rect 9383 26333 9395 26367
rect 9429 26333 9441 26367
rect 9383 26327 9441 26333
rect 9483 26367 9541 26373
rect 9483 26333 9495 26367
rect 9529 26333 9541 26367
rect 9483 26327 9541 26333
rect 9585 26367 9643 26373
rect 9585 26333 9597 26367
rect 9631 26364 9643 26367
rect 10318 26364 10324 26376
rect 9631 26336 10324 26364
rect 9631 26333 9643 26336
rect 9585 26327 9643 26333
rect 1578 26296 1584 26308
rect 1539 26268 1584 26296
rect 1578 26256 1584 26268
rect 1636 26256 1642 26308
rect 5905 26299 5963 26305
rect 5905 26265 5917 26299
rect 5951 26296 5963 26299
rect 6181 26299 6239 26305
rect 6181 26296 6193 26299
rect 5951 26268 6193 26296
rect 5951 26265 5963 26268
rect 5905 26259 5963 26265
rect 6181 26265 6193 26268
rect 6227 26296 6239 26299
rect 6362 26296 6368 26308
rect 6227 26268 6368 26296
rect 6227 26265 6239 26268
rect 6181 26259 6239 26265
rect 6362 26256 6368 26268
rect 6420 26256 6426 26308
rect 9214 26256 9220 26308
rect 9272 26256 9278 26308
rect 9407 26296 9435 26327
rect 10318 26324 10324 26336
rect 10376 26324 10382 26376
rect 10413 26367 10471 26373
rect 10413 26333 10425 26367
rect 10459 26364 10471 26367
rect 10870 26364 10876 26376
rect 10459 26336 10876 26364
rect 10459 26333 10471 26336
rect 10413 26327 10471 26333
rect 10870 26324 10876 26336
rect 10928 26324 10934 26376
rect 12342 26364 12348 26376
rect 12303 26336 12348 26364
rect 12342 26324 12348 26336
rect 12400 26324 12406 26376
rect 14090 26364 14096 26376
rect 14051 26336 14096 26364
rect 14090 26324 14096 26336
rect 14148 26324 14154 26376
rect 14366 26364 14372 26376
rect 14327 26336 14372 26364
rect 14366 26324 14372 26336
rect 14424 26324 14430 26376
rect 14829 26367 14887 26373
rect 14829 26333 14841 26367
rect 14875 26364 14887 26367
rect 15194 26364 15200 26376
rect 14875 26336 15200 26364
rect 14875 26333 14887 26336
rect 14829 26327 14887 26333
rect 15194 26324 15200 26336
rect 15252 26324 15258 26376
rect 15286 26324 15292 26376
rect 15344 26364 15350 26376
rect 15344 26336 15389 26364
rect 15344 26324 15350 26336
rect 17586 26324 17592 26376
rect 17644 26364 17650 26376
rect 17819 26367 17877 26373
rect 18070 26367 18128 26373
rect 17819 26364 17831 26367
rect 17644 26336 17831 26364
rect 17644 26324 17650 26336
rect 17819 26333 17831 26336
rect 17865 26333 17877 26367
rect 17819 26327 17877 26333
rect 17954 26361 18012 26367
rect 17954 26327 17966 26361
rect 18000 26327 18012 26361
rect 18070 26333 18082 26367
rect 18116 26364 18128 26367
rect 18156 26364 18184 26460
rect 19444 26432 19472 26540
rect 19518 26528 19524 26580
rect 19576 26568 19582 26580
rect 21545 26571 21603 26577
rect 21545 26568 21557 26571
rect 19576 26540 21557 26568
rect 19576 26528 19582 26540
rect 21545 26537 21557 26540
rect 21591 26537 21603 26571
rect 21545 26531 21603 26537
rect 27157 26571 27215 26577
rect 27157 26537 27169 26571
rect 27203 26568 27215 26571
rect 27246 26568 27252 26580
rect 27203 26540 27252 26568
rect 27203 26537 27215 26540
rect 27157 26531 27215 26537
rect 27246 26528 27252 26540
rect 27304 26528 27310 26580
rect 29914 26568 29920 26580
rect 29875 26540 29920 26568
rect 29914 26528 29920 26540
rect 29972 26528 29978 26580
rect 34149 26571 34207 26577
rect 34149 26537 34161 26571
rect 34195 26568 34207 26571
rect 34330 26568 34336 26580
rect 34195 26540 34336 26568
rect 34195 26537 34207 26540
rect 34149 26531 34207 26537
rect 34330 26528 34336 26540
rect 34388 26528 34394 26580
rect 35986 26528 35992 26580
rect 36044 26568 36050 26580
rect 38930 26568 38936 26580
rect 36044 26540 36768 26568
rect 38891 26540 38936 26568
rect 36044 26528 36050 26540
rect 36740 26509 36768 26540
rect 38930 26528 38936 26540
rect 38988 26528 38994 26580
rect 36725 26503 36783 26509
rect 36725 26469 36737 26503
rect 36771 26500 36783 26503
rect 37274 26500 37280 26512
rect 36771 26472 37280 26500
rect 36771 26469 36783 26472
rect 36725 26463 36783 26469
rect 37274 26460 37280 26472
rect 37332 26460 37338 26512
rect 19444 26404 20300 26432
rect 18116 26336 18184 26364
rect 18233 26367 18291 26373
rect 18116 26333 18128 26336
rect 18070 26327 18128 26333
rect 18233 26333 18245 26367
rect 18279 26364 18291 26367
rect 19518 26364 19524 26376
rect 18279 26336 19104 26364
rect 19479 26336 19524 26364
rect 18279 26333 18291 26336
rect 18233 26327 18291 26333
rect 17954 26321 18012 26327
rect 10134 26296 10140 26308
rect 9407 26268 10140 26296
rect 10134 26256 10140 26268
rect 10192 26256 10198 26308
rect 10229 26299 10287 26305
rect 10229 26265 10241 26299
rect 10275 26296 10287 26299
rect 10686 26296 10692 26308
rect 10275 26268 10692 26296
rect 10275 26265 10287 26268
rect 10229 26259 10287 26265
rect 1946 26188 1952 26240
rect 2004 26228 2010 26240
rect 5718 26228 5724 26240
rect 2004 26200 5724 26228
rect 2004 26188 2010 26200
rect 5718 26188 5724 26200
rect 5776 26188 5782 26240
rect 9232 26228 9260 26256
rect 10244 26228 10272 26259
rect 10686 26256 10692 26268
rect 10744 26256 10750 26308
rect 12069 26299 12127 26305
rect 12069 26265 12081 26299
rect 12115 26296 12127 26299
rect 12158 26296 12164 26308
rect 12115 26268 12164 26296
rect 12115 26265 12127 26268
rect 12069 26259 12127 26265
rect 12158 26256 12164 26268
rect 12216 26256 12222 26308
rect 15010 26256 15016 26308
rect 15068 26296 15074 26308
rect 15378 26296 15384 26308
rect 15068 26268 15148 26296
rect 15068 26256 15074 26268
rect 12250 26228 12256 26240
rect 9232 26200 10272 26228
rect 12211 26200 12256 26228
rect 12250 26188 12256 26200
rect 12308 26188 12314 26240
rect 14274 26228 14280 26240
rect 14235 26200 14280 26228
rect 14274 26188 14280 26200
rect 14332 26188 14338 26240
rect 15120 26237 15148 26268
rect 15212 26268 15384 26296
rect 15212 26237 15240 26268
rect 15378 26256 15384 26268
rect 15436 26256 15442 26308
rect 15105 26231 15163 26237
rect 15105 26197 15117 26231
rect 15151 26197 15163 26231
rect 15105 26191 15163 26197
rect 15197 26231 15255 26237
rect 15197 26197 15209 26231
rect 15243 26197 15255 26231
rect 15197 26191 15255 26197
rect 16942 26188 16948 26240
rect 17000 26228 17006 26240
rect 17589 26231 17647 26237
rect 17589 26228 17601 26231
rect 17000 26200 17601 26228
rect 17000 26188 17006 26200
rect 17589 26197 17601 26200
rect 17635 26197 17647 26231
rect 17972 26228 18000 26321
rect 18138 26228 18144 26240
rect 17972 26200 18144 26228
rect 17589 26191 17647 26197
rect 18138 26188 18144 26200
rect 18196 26188 18202 26240
rect 19076 26228 19104 26336
rect 19518 26324 19524 26336
rect 19576 26324 19582 26376
rect 20070 26324 20076 26376
rect 20128 26364 20134 26376
rect 20165 26367 20223 26373
rect 20165 26364 20177 26367
rect 20128 26336 20177 26364
rect 20128 26324 20134 26336
rect 20165 26333 20177 26336
rect 20211 26333 20223 26367
rect 20272 26364 20300 26404
rect 23566 26392 23572 26444
rect 23624 26432 23630 26444
rect 31849 26435 31907 26441
rect 31849 26432 31861 26435
rect 23624 26404 31861 26432
rect 23624 26392 23630 26404
rect 31849 26401 31861 26404
rect 31895 26401 31907 26435
rect 31849 26395 31907 26401
rect 32125 26435 32183 26441
rect 32125 26401 32137 26435
rect 32171 26432 32183 26435
rect 32858 26432 32864 26444
rect 32171 26404 32864 26432
rect 32171 26401 32183 26404
rect 32125 26395 32183 26401
rect 32858 26392 32864 26404
rect 32916 26392 32922 26444
rect 24762 26364 24768 26376
rect 20272 26336 24768 26364
rect 20165 26327 20223 26333
rect 24762 26324 24768 26336
rect 24820 26324 24826 26376
rect 27065 26367 27123 26373
rect 27065 26333 27077 26367
rect 27111 26364 27123 26367
rect 27430 26364 27436 26376
rect 27111 26336 27436 26364
rect 27111 26333 27123 26336
rect 27065 26327 27123 26333
rect 27430 26324 27436 26336
rect 27488 26324 27494 26376
rect 29822 26364 29828 26376
rect 29783 26336 29828 26364
rect 29822 26324 29828 26336
rect 29880 26324 29886 26376
rect 30742 26364 30748 26376
rect 30703 26336 30748 26364
rect 30742 26324 30748 26336
rect 30800 26324 30806 26376
rect 33781 26367 33839 26373
rect 33781 26333 33793 26367
rect 33827 26364 33839 26367
rect 33827 26336 34468 26364
rect 33827 26333 33839 26336
rect 33781 26327 33839 26333
rect 19150 26256 19156 26308
rect 19208 26296 19214 26308
rect 19337 26299 19395 26305
rect 19337 26296 19349 26299
rect 19208 26268 19349 26296
rect 19208 26256 19214 26268
rect 19337 26265 19349 26268
rect 19383 26265 19395 26299
rect 19337 26259 19395 26265
rect 20254 26256 20260 26308
rect 20312 26296 20318 26308
rect 20410 26299 20468 26305
rect 20410 26296 20422 26299
rect 20312 26268 20422 26296
rect 20312 26256 20318 26268
rect 20410 26265 20422 26268
rect 20456 26265 20468 26299
rect 20410 26259 20468 26265
rect 26326 26256 26332 26308
rect 26384 26296 26390 26308
rect 31110 26296 31116 26308
rect 26384 26268 31116 26296
rect 26384 26256 26390 26268
rect 31110 26256 31116 26268
rect 31168 26256 31174 26308
rect 31202 26256 31208 26308
rect 31260 26296 31266 26308
rect 33965 26299 34023 26305
rect 33965 26296 33977 26299
rect 31260 26268 33977 26296
rect 31260 26256 31266 26268
rect 33965 26265 33977 26268
rect 34011 26296 34023 26299
rect 34330 26296 34336 26308
rect 34011 26268 34336 26296
rect 34011 26265 34023 26268
rect 33965 26259 34023 26265
rect 34330 26256 34336 26268
rect 34388 26256 34394 26308
rect 34440 26296 34468 26336
rect 34514 26324 34520 26376
rect 34572 26364 34578 26376
rect 35342 26364 35348 26376
rect 34572 26336 35348 26364
rect 34572 26324 34578 26336
rect 35342 26324 35348 26336
rect 35400 26324 35406 26376
rect 35434 26324 35440 26376
rect 35492 26364 35498 26376
rect 35601 26367 35659 26373
rect 35601 26364 35613 26367
rect 35492 26336 35613 26364
rect 35492 26324 35498 26336
rect 35601 26333 35613 26336
rect 35647 26333 35659 26367
rect 35601 26327 35659 26333
rect 37366 26324 37372 26376
rect 37424 26364 37430 26376
rect 38105 26367 38163 26373
rect 38105 26364 38117 26367
rect 37424 26336 38117 26364
rect 37424 26324 37430 26336
rect 38105 26333 38117 26336
rect 38151 26364 38163 26367
rect 38749 26367 38807 26373
rect 38749 26364 38761 26367
rect 38151 26336 38761 26364
rect 38151 26333 38163 26336
rect 38105 26327 38163 26333
rect 38749 26333 38761 26336
rect 38795 26333 38807 26367
rect 38749 26327 38807 26333
rect 35250 26296 35256 26308
rect 34440 26268 35256 26296
rect 35250 26256 35256 26268
rect 35308 26256 35314 26308
rect 47946 26296 47952 26308
rect 47907 26268 47952 26296
rect 47946 26256 47952 26268
rect 48004 26256 48010 26308
rect 48038 26256 48044 26308
rect 48096 26296 48102 26308
rect 48133 26299 48191 26305
rect 48133 26296 48145 26299
rect 48096 26268 48145 26296
rect 48096 26256 48102 26268
rect 48133 26265 48145 26268
rect 48179 26265 48191 26299
rect 48133 26259 48191 26265
rect 19426 26228 19432 26240
rect 19076 26200 19432 26228
rect 19426 26188 19432 26200
rect 19484 26188 19490 26240
rect 19705 26231 19763 26237
rect 19705 26197 19717 26231
rect 19751 26228 19763 26231
rect 20530 26228 20536 26240
rect 19751 26200 20536 26228
rect 19751 26197 19763 26200
rect 19705 26191 19763 26197
rect 20530 26188 20536 26200
rect 20588 26188 20594 26240
rect 20806 26188 20812 26240
rect 20864 26228 20870 26240
rect 30190 26228 30196 26240
rect 20864 26200 30196 26228
rect 20864 26188 20870 26200
rect 30190 26188 30196 26200
rect 30248 26188 30254 26240
rect 30374 26188 30380 26240
rect 30432 26228 30438 26240
rect 36538 26228 36544 26240
rect 30432 26200 36544 26228
rect 30432 26188 30438 26200
rect 36538 26188 36544 26200
rect 36596 26188 36602 26240
rect 38197 26231 38255 26237
rect 38197 26197 38209 26231
rect 38243 26228 38255 26231
rect 38286 26228 38292 26240
rect 38243 26200 38292 26228
rect 38243 26197 38255 26200
rect 38197 26191 38255 26197
rect 38286 26188 38292 26200
rect 38344 26188 38350 26240
rect 1104 26138 48852 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 48852 26138
rect 1104 26064 48852 26086
rect 1578 25984 1584 26036
rect 1636 26024 1642 26036
rect 2225 26027 2283 26033
rect 2225 26024 2237 26027
rect 1636 25996 2237 26024
rect 1636 25984 1642 25996
rect 2225 25993 2237 25996
rect 2271 25993 2283 26027
rect 12621 26027 12679 26033
rect 2225 25987 2283 25993
rect 2516 25996 2774 26024
rect 2516 25900 2544 25996
rect 1578 25888 1584 25900
rect 1539 25860 1584 25888
rect 1578 25848 1584 25860
rect 1636 25848 1642 25900
rect 2133 25891 2191 25897
rect 2133 25857 2145 25891
rect 2179 25888 2191 25891
rect 2498 25888 2504 25900
rect 2179 25860 2504 25888
rect 2179 25857 2191 25860
rect 2133 25851 2191 25857
rect 2498 25848 2504 25860
rect 2556 25848 2562 25900
rect 2746 25888 2774 25996
rect 12621 25993 12633 26027
rect 12667 26024 12679 26027
rect 12894 26024 12900 26036
rect 12667 25996 12900 26024
rect 12667 25993 12679 25996
rect 12621 25987 12679 25993
rect 12894 25984 12900 25996
rect 12952 25984 12958 26036
rect 13262 25984 13268 26036
rect 13320 26024 13326 26036
rect 17954 26024 17960 26036
rect 13320 25996 17960 26024
rect 13320 25984 13326 25996
rect 17954 25984 17960 25996
rect 18012 25984 18018 26036
rect 18046 25984 18052 26036
rect 18104 26024 18110 26036
rect 18417 26027 18475 26033
rect 18417 26024 18429 26027
rect 18104 25996 18429 26024
rect 18104 25984 18110 25996
rect 18417 25993 18429 25996
rect 18463 26024 18475 26027
rect 19058 26024 19064 26036
rect 18463 25996 19064 26024
rect 18463 25993 18475 25996
rect 18417 25987 18475 25993
rect 19058 25984 19064 25996
rect 19116 25984 19122 26036
rect 20073 26027 20131 26033
rect 20073 25993 20085 26027
rect 20119 26024 20131 26027
rect 20254 26024 20260 26036
rect 20119 25996 20260 26024
rect 20119 25993 20131 25996
rect 20073 25987 20131 25993
rect 20254 25984 20260 25996
rect 20312 25984 20318 26036
rect 23385 26027 23443 26033
rect 23385 25993 23397 26027
rect 23431 25993 23443 26027
rect 23385 25987 23443 25993
rect 5718 25916 5724 25968
rect 5776 25956 5782 25968
rect 19886 25956 19892 25968
rect 5776 25928 19892 25956
rect 5776 25916 5782 25928
rect 19886 25916 19892 25928
rect 19944 25916 19950 25968
rect 22922 25956 22928 25968
rect 22883 25928 22928 25956
rect 22922 25916 22928 25928
rect 22980 25916 22986 25968
rect 23400 25956 23428 25987
rect 23934 25984 23940 26036
rect 23992 26024 23998 26036
rect 24394 26024 24400 26036
rect 23992 25996 24400 26024
rect 23992 25984 23998 25996
rect 24394 25984 24400 25996
rect 24452 25984 24458 26036
rect 24670 25984 24676 26036
rect 24728 26024 24734 26036
rect 30374 26024 30380 26036
rect 24728 25996 30380 26024
rect 24728 25984 24734 25996
rect 30374 25984 30380 25996
rect 30432 25984 30438 26036
rect 31754 25984 31760 26036
rect 31812 26024 31818 26036
rect 32122 26024 32128 26036
rect 31812 25996 32128 26024
rect 31812 25984 31818 25996
rect 32122 25984 32128 25996
rect 32180 25984 32186 26036
rect 32582 25984 32588 26036
rect 32640 25984 32646 26036
rect 33318 25984 33324 26036
rect 33376 26024 33382 26036
rect 33689 26027 33747 26033
rect 33689 26024 33701 26027
rect 33376 25996 33701 26024
rect 33376 25984 33382 25996
rect 33689 25993 33701 25996
rect 33735 25993 33747 26027
rect 34514 26024 34520 26036
rect 33689 25987 33747 25993
rect 34256 25996 34520 26024
rect 24765 25959 24823 25965
rect 24765 25956 24777 25959
rect 23400 25928 24777 25956
rect 24765 25925 24777 25928
rect 24811 25925 24823 25959
rect 27982 25956 27988 25968
rect 24765 25919 24823 25925
rect 26160 25928 27988 25956
rect 10229 25891 10287 25897
rect 2746 25860 6316 25888
rect 1397 25755 1455 25761
rect 1397 25721 1409 25755
rect 1443 25752 1455 25755
rect 6178 25752 6184 25764
rect 1443 25724 6184 25752
rect 1443 25721 1455 25724
rect 1397 25715 1455 25721
rect 6178 25712 6184 25724
rect 6236 25712 6242 25764
rect 6288 25684 6316 25860
rect 10229 25857 10241 25891
rect 10275 25888 10287 25891
rect 10318 25888 10324 25900
rect 10275 25860 10324 25888
rect 10275 25857 10287 25860
rect 10229 25851 10287 25857
rect 10318 25848 10324 25860
rect 10376 25848 10382 25900
rect 12161 25891 12219 25897
rect 12161 25857 12173 25891
rect 12207 25888 12219 25891
rect 12437 25891 12495 25897
rect 12207 25860 12388 25888
rect 12207 25857 12219 25860
rect 12161 25851 12219 25857
rect 6825 25823 6883 25829
rect 6825 25789 6837 25823
rect 6871 25789 6883 25823
rect 7006 25820 7012 25832
rect 6967 25792 7012 25820
rect 6825 25783 6883 25789
rect 6840 25752 6868 25783
rect 7006 25780 7012 25792
rect 7064 25780 7070 25832
rect 8662 25820 8668 25832
rect 8623 25792 8668 25820
rect 8662 25780 8668 25792
rect 8720 25780 8726 25832
rect 9953 25823 10011 25829
rect 9953 25789 9965 25823
rect 9999 25820 10011 25823
rect 10134 25820 10140 25832
rect 9999 25792 10140 25820
rect 9999 25789 10011 25792
rect 9953 25783 10011 25789
rect 10134 25780 10140 25792
rect 10192 25780 10198 25832
rect 11054 25780 11060 25832
rect 11112 25820 11118 25832
rect 12253 25823 12311 25829
rect 12253 25820 12265 25823
rect 11112 25792 12265 25820
rect 11112 25780 11118 25792
rect 12253 25789 12265 25792
rect 12299 25789 12311 25823
rect 12360 25820 12388 25860
rect 12437 25857 12449 25891
rect 12483 25888 12495 25891
rect 12526 25888 12532 25900
rect 12483 25860 12532 25888
rect 12483 25857 12495 25860
rect 12437 25851 12495 25857
rect 12526 25848 12532 25860
rect 12584 25848 12590 25900
rect 13538 25848 13544 25900
rect 13596 25888 13602 25900
rect 13725 25891 13783 25897
rect 13725 25888 13737 25891
rect 13596 25860 13737 25888
rect 13596 25848 13602 25860
rect 13725 25857 13737 25860
rect 13771 25857 13783 25891
rect 14550 25888 14556 25900
rect 14511 25860 14556 25888
rect 13725 25851 13783 25857
rect 14550 25848 14556 25860
rect 14608 25848 14614 25900
rect 14826 25888 14832 25900
rect 14787 25860 14832 25888
rect 14826 25848 14832 25860
rect 14884 25848 14890 25900
rect 16942 25897 16948 25900
rect 16936 25888 16948 25897
rect 16903 25860 16948 25888
rect 16936 25851 16948 25860
rect 16942 25848 16948 25851
rect 17000 25848 17006 25900
rect 17954 25848 17960 25900
rect 18012 25888 18018 25900
rect 18874 25888 18880 25900
rect 18012 25860 18880 25888
rect 18012 25848 18018 25860
rect 18874 25848 18880 25860
rect 18932 25848 18938 25900
rect 19058 25888 19064 25900
rect 19019 25860 19064 25888
rect 19058 25848 19064 25860
rect 19116 25848 19122 25900
rect 19153 25891 19211 25897
rect 19153 25857 19165 25891
rect 19199 25857 19211 25891
rect 19153 25851 19211 25857
rect 13630 25820 13636 25832
rect 12360 25792 13400 25820
rect 13591 25792 13636 25820
rect 12253 25783 12311 25789
rect 8386 25752 8392 25764
rect 6840 25724 8392 25752
rect 8386 25712 8392 25724
rect 8444 25712 8450 25764
rect 8496 25724 12434 25752
rect 8496 25684 8524 25724
rect 6288 25656 8524 25684
rect 9582 25644 9588 25696
rect 9640 25684 9646 25696
rect 10870 25684 10876 25696
rect 9640 25656 10876 25684
rect 9640 25644 9646 25656
rect 10870 25644 10876 25656
rect 10928 25644 10934 25696
rect 12066 25644 12072 25696
rect 12124 25684 12130 25696
rect 12161 25687 12219 25693
rect 12161 25684 12173 25687
rect 12124 25656 12173 25684
rect 12124 25644 12130 25656
rect 12161 25653 12173 25656
rect 12207 25653 12219 25687
rect 12406 25684 12434 25724
rect 13262 25684 13268 25696
rect 12406 25656 13268 25684
rect 12161 25647 12219 25653
rect 13262 25644 13268 25656
rect 13320 25644 13326 25696
rect 13372 25684 13400 25792
rect 13630 25780 13636 25792
rect 13688 25780 13694 25832
rect 14645 25823 14703 25829
rect 14645 25820 14657 25823
rect 14108 25792 14657 25820
rect 14108 25761 14136 25792
rect 14645 25789 14657 25792
rect 14691 25789 14703 25823
rect 16666 25820 16672 25832
rect 16627 25792 16672 25820
rect 14645 25783 14703 25789
rect 16666 25780 16672 25792
rect 16724 25780 16730 25832
rect 18138 25780 18144 25832
rect 18196 25820 18202 25832
rect 19168 25820 19196 25851
rect 19242 25848 19248 25900
rect 19300 25888 19306 25900
rect 19300 25860 19345 25888
rect 19300 25848 19306 25860
rect 19426 25848 19432 25900
rect 19484 25888 19490 25900
rect 19484 25860 19529 25888
rect 19484 25848 19490 25860
rect 20254 25848 20260 25900
rect 20312 25897 20318 25900
rect 20312 25891 20361 25897
rect 20312 25857 20315 25891
rect 20349 25857 20361 25891
rect 20312 25851 20361 25857
rect 20441 25891 20499 25897
rect 20441 25857 20453 25891
rect 20487 25857 20499 25891
rect 20441 25851 20499 25857
rect 20312 25848 20318 25851
rect 20456 25820 20484 25851
rect 20530 25848 20536 25900
rect 20588 25888 20594 25900
rect 20588 25860 20633 25888
rect 20588 25848 20594 25860
rect 20714 25848 20720 25900
rect 20772 25888 20778 25900
rect 23201 25891 23259 25897
rect 20772 25860 20817 25888
rect 20772 25848 20778 25860
rect 23201 25857 23213 25891
rect 23247 25857 23259 25891
rect 23842 25888 23848 25900
rect 23803 25860 23848 25888
rect 23201 25851 23259 25857
rect 20806 25820 20812 25832
rect 18196 25792 20812 25820
rect 18196 25780 18202 25792
rect 20806 25780 20812 25792
rect 20864 25780 20870 25832
rect 23106 25820 23112 25832
rect 23067 25792 23112 25820
rect 23106 25780 23112 25792
rect 23164 25780 23170 25832
rect 14093 25755 14151 25761
rect 14093 25721 14105 25755
rect 14139 25721 14151 25755
rect 15013 25755 15071 25761
rect 15013 25752 15025 25755
rect 14093 25715 14151 25721
rect 14200 25724 15025 25752
rect 14200 25684 14228 25724
rect 15013 25721 15025 25724
rect 15059 25721 15071 25755
rect 19978 25752 19984 25764
rect 15013 25715 15071 25721
rect 17604 25724 19984 25752
rect 13372 25656 14228 25684
rect 14458 25644 14464 25696
rect 14516 25684 14522 25696
rect 14553 25687 14611 25693
rect 14553 25684 14565 25687
rect 14516 25656 14565 25684
rect 14516 25644 14522 25656
rect 14553 25653 14565 25656
rect 14599 25653 14611 25687
rect 14553 25647 14611 25653
rect 17034 25644 17040 25696
rect 17092 25684 17098 25696
rect 17604 25684 17632 25724
rect 19978 25712 19984 25724
rect 20036 25712 20042 25764
rect 18046 25684 18052 25696
rect 17092 25656 17632 25684
rect 18007 25656 18052 25684
rect 17092 25644 17098 25656
rect 18046 25644 18052 25656
rect 18104 25644 18110 25696
rect 18782 25684 18788 25696
rect 18743 25656 18788 25684
rect 18782 25644 18788 25656
rect 18840 25644 18846 25696
rect 19886 25644 19892 25696
rect 19944 25684 19950 25696
rect 22557 25687 22615 25693
rect 22557 25684 22569 25687
rect 19944 25656 22569 25684
rect 19944 25644 19950 25656
rect 22557 25653 22569 25656
rect 22603 25684 22615 25687
rect 22925 25687 22983 25693
rect 22925 25684 22937 25687
rect 22603 25656 22937 25684
rect 22603 25653 22615 25656
rect 22557 25647 22615 25653
rect 22925 25653 22937 25656
rect 22971 25653 22983 25687
rect 23216 25684 23244 25851
rect 23842 25848 23848 25860
rect 23900 25848 23906 25900
rect 24026 25848 24032 25900
rect 24084 25888 24090 25900
rect 24121 25891 24179 25897
rect 24121 25888 24133 25891
rect 24084 25860 24133 25888
rect 24084 25848 24090 25860
rect 24121 25857 24133 25860
rect 24167 25857 24179 25891
rect 24121 25851 24179 25857
rect 24302 25848 24308 25900
rect 24360 25848 24366 25900
rect 24949 25891 25007 25897
rect 24949 25888 24961 25891
rect 24510 25860 24961 25888
rect 23937 25823 23995 25829
rect 23937 25789 23949 25823
rect 23983 25820 23995 25823
rect 24320 25820 24348 25848
rect 23983 25792 24348 25820
rect 23983 25789 23995 25792
rect 23937 25783 23995 25789
rect 24305 25755 24363 25761
rect 24305 25721 24317 25755
rect 24351 25752 24363 25755
rect 24510 25752 24538 25860
rect 24949 25857 24961 25860
rect 24995 25857 25007 25891
rect 24949 25851 25007 25857
rect 25041 25891 25099 25897
rect 25041 25857 25053 25891
rect 25087 25888 25099 25891
rect 25958 25888 25964 25900
rect 25087 25860 25964 25888
rect 25087 25857 25099 25860
rect 25041 25851 25099 25857
rect 25958 25848 25964 25860
rect 26016 25848 26022 25900
rect 26160 25897 26188 25928
rect 27982 25916 27988 25928
rect 28040 25916 28046 25968
rect 29822 25916 29828 25968
rect 29880 25956 29886 25968
rect 31297 25959 31355 25965
rect 31297 25956 31309 25959
rect 29880 25928 31309 25956
rect 29880 25916 29886 25928
rect 31297 25925 31309 25928
rect 31343 25925 31355 25959
rect 32600 25956 32628 25984
rect 34256 25956 34284 25996
rect 34514 25984 34520 25996
rect 34572 25984 34578 26036
rect 35250 25984 35256 26036
rect 35308 26024 35314 26036
rect 35618 26024 35624 26036
rect 35308 25996 35624 26024
rect 35308 25984 35314 25996
rect 35618 25984 35624 25996
rect 35676 25984 35682 26036
rect 36538 25984 36544 26036
rect 36596 26024 36602 26036
rect 46842 26024 46848 26036
rect 36596 25996 46848 26024
rect 36596 25984 36602 25996
rect 46842 25984 46848 25996
rect 46900 25984 46906 26036
rect 31297 25919 31355 25925
rect 32324 25928 34284 25956
rect 26145 25891 26203 25897
rect 26145 25857 26157 25891
rect 26191 25857 26203 25891
rect 26145 25851 26203 25857
rect 26329 25891 26387 25897
rect 26329 25857 26341 25891
rect 26375 25857 26387 25891
rect 26329 25851 26387 25857
rect 29917 25891 29975 25897
rect 29917 25857 29929 25891
rect 29963 25888 29975 25891
rect 30742 25888 30748 25900
rect 29963 25860 30748 25888
rect 29963 25857 29975 25860
rect 29917 25851 29975 25857
rect 26145 25755 26203 25761
rect 26145 25752 26157 25755
rect 24351 25724 24538 25752
rect 24964 25724 26157 25752
rect 24351 25721 24363 25724
rect 24305 25715 24363 25721
rect 23753 25687 23811 25693
rect 23753 25684 23765 25687
rect 23216 25656 23765 25684
rect 22925 25647 22983 25653
rect 23753 25653 23765 25656
rect 23799 25684 23811 25687
rect 23934 25684 23940 25696
rect 23799 25656 23940 25684
rect 23799 25653 23811 25656
rect 23753 25647 23811 25653
rect 23934 25644 23940 25656
rect 23992 25644 23998 25696
rect 24118 25684 24124 25696
rect 24079 25656 24124 25684
rect 24118 25644 24124 25656
rect 24176 25644 24182 25696
rect 24762 25684 24768 25696
rect 24723 25656 24768 25684
rect 24762 25644 24768 25656
rect 24820 25644 24826 25696
rect 24854 25644 24860 25696
rect 24912 25684 24918 25696
rect 24964 25684 24992 25724
rect 26145 25721 26157 25724
rect 26191 25721 26203 25755
rect 26145 25715 26203 25721
rect 25222 25684 25228 25696
rect 24912 25656 24992 25684
rect 25183 25656 25228 25684
rect 24912 25644 24918 25656
rect 25222 25644 25228 25656
rect 25280 25644 25286 25696
rect 26344 25684 26372 25851
rect 30742 25848 30748 25860
rect 30800 25888 30806 25900
rect 30929 25891 30987 25897
rect 30929 25888 30941 25891
rect 30800 25860 30941 25888
rect 30800 25848 30806 25860
rect 30929 25857 30941 25860
rect 30975 25857 30987 25891
rect 32214 25888 32220 25900
rect 30929 25851 30987 25857
rect 31036 25860 32220 25888
rect 30098 25820 30104 25832
rect 30059 25792 30104 25820
rect 30098 25780 30104 25792
rect 30156 25820 30162 25832
rect 31036 25820 31064 25860
rect 32214 25848 32220 25860
rect 32272 25848 32278 25900
rect 30156 25792 31064 25820
rect 30156 25780 30162 25792
rect 32122 25780 32128 25832
rect 32180 25820 32186 25832
rect 32324 25829 32352 25928
rect 32398 25848 32404 25900
rect 32456 25888 32462 25900
rect 34256 25897 34284 25928
rect 34606 25916 34612 25968
rect 34664 25916 34670 25968
rect 38286 25956 38292 25968
rect 38247 25928 38292 25956
rect 38286 25916 38292 25928
rect 38344 25916 38350 25968
rect 46474 25956 46480 25968
rect 39500 25928 46480 25956
rect 32565 25891 32623 25897
rect 32565 25888 32577 25891
rect 32456 25860 32577 25888
rect 32456 25848 32462 25860
rect 32565 25857 32577 25860
rect 32611 25857 32623 25891
rect 32565 25851 32623 25857
rect 34241 25891 34299 25897
rect 34241 25857 34253 25891
rect 34287 25857 34299 25891
rect 34241 25851 34299 25857
rect 34508 25891 34566 25897
rect 34508 25857 34520 25891
rect 34554 25888 34566 25891
rect 34624 25888 34652 25916
rect 38102 25888 38108 25900
rect 34554 25860 34652 25888
rect 38063 25860 38108 25888
rect 34554 25857 34566 25860
rect 34508 25851 34566 25857
rect 38102 25848 38108 25860
rect 38160 25848 38166 25900
rect 32309 25823 32367 25829
rect 32309 25820 32321 25823
rect 32180 25792 32321 25820
rect 32180 25780 32186 25792
rect 32309 25789 32321 25792
rect 32355 25789 32367 25823
rect 32309 25783 32367 25789
rect 39500 25752 39528 25928
rect 46474 25916 46480 25928
rect 46532 25956 46538 25968
rect 46937 25959 46995 25965
rect 46937 25956 46949 25959
rect 46532 25928 46949 25956
rect 46532 25916 46538 25928
rect 46937 25925 46949 25928
rect 46983 25925 46995 25959
rect 46937 25919 46995 25925
rect 46842 25888 46848 25900
rect 46803 25860 46848 25888
rect 46842 25848 46848 25860
rect 46900 25848 46906 25900
rect 39945 25823 40003 25829
rect 39945 25789 39957 25823
rect 39991 25820 40003 25823
rect 48498 25820 48504 25832
rect 39991 25792 48504 25820
rect 39991 25789 40003 25792
rect 39945 25783 40003 25789
rect 48498 25780 48504 25792
rect 48556 25780 48562 25832
rect 36464 25724 39528 25752
rect 36464 25684 36492 25724
rect 26344 25656 36492 25684
rect 36538 25644 36544 25696
rect 36596 25684 36602 25696
rect 45186 25684 45192 25696
rect 36596 25656 45192 25684
rect 36596 25644 36602 25656
rect 45186 25644 45192 25656
rect 45244 25644 45250 25696
rect 47762 25684 47768 25696
rect 47723 25656 47768 25684
rect 47762 25644 47768 25656
rect 47820 25644 47826 25696
rect 1104 25594 48852 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 48852 25594
rect 1104 25520 48852 25542
rect 7006 25480 7012 25492
rect 6967 25452 7012 25480
rect 7006 25440 7012 25452
rect 7064 25440 7070 25492
rect 9217 25483 9275 25489
rect 9217 25449 9229 25483
rect 9263 25480 9275 25483
rect 9306 25480 9312 25492
rect 9263 25452 9312 25480
rect 9263 25449 9275 25452
rect 9217 25443 9275 25449
rect 9306 25440 9312 25452
rect 9364 25440 9370 25492
rect 9950 25480 9956 25492
rect 9407 25452 9956 25480
rect 9407 25412 9435 25452
rect 9950 25440 9956 25452
rect 10008 25440 10014 25492
rect 10134 25480 10140 25492
rect 10095 25452 10140 25480
rect 10134 25440 10140 25452
rect 10192 25440 10198 25492
rect 11054 25480 11060 25492
rect 11015 25452 11060 25480
rect 11054 25440 11060 25452
rect 11112 25440 11118 25492
rect 12250 25440 12256 25492
rect 12308 25480 12314 25492
rect 12345 25483 12403 25489
rect 12345 25480 12357 25483
rect 12308 25452 12357 25480
rect 12308 25440 12314 25452
rect 12345 25449 12357 25452
rect 12391 25449 12403 25483
rect 12526 25480 12532 25492
rect 12487 25452 12532 25480
rect 12345 25443 12403 25449
rect 12526 25440 12532 25452
rect 12584 25440 12590 25492
rect 14274 25480 14280 25492
rect 14235 25452 14280 25480
rect 14274 25440 14280 25452
rect 14332 25440 14338 25492
rect 14458 25480 14464 25492
rect 14419 25452 14464 25480
rect 14458 25440 14464 25452
rect 14516 25440 14522 25492
rect 14550 25440 14556 25492
rect 14608 25480 14614 25492
rect 19518 25480 19524 25492
rect 14608 25452 19524 25480
rect 14608 25440 14614 25452
rect 19518 25440 19524 25452
rect 19576 25480 19582 25492
rect 21453 25483 21511 25489
rect 21453 25480 21465 25483
rect 19576 25452 21465 25480
rect 19576 25440 19582 25452
rect 21453 25449 21465 25452
rect 21499 25449 21511 25483
rect 21453 25443 21511 25449
rect 22189 25483 22247 25489
rect 22189 25449 22201 25483
rect 22235 25480 22247 25483
rect 23566 25480 23572 25492
rect 22235 25452 23572 25480
rect 22235 25449 22247 25452
rect 22189 25443 22247 25449
rect 23566 25440 23572 25452
rect 23624 25440 23630 25492
rect 23750 25480 23756 25492
rect 23711 25452 23756 25480
rect 23750 25440 23756 25452
rect 23808 25440 23814 25492
rect 30098 25480 30104 25492
rect 23860 25452 30104 25480
rect 12268 25412 12296 25440
rect 9048 25384 9435 25412
rect 9876 25384 12296 25412
rect 6638 25236 6644 25288
rect 6696 25276 6702 25288
rect 6914 25276 6920 25288
rect 6696 25248 6920 25276
rect 6696 25236 6702 25248
rect 6914 25236 6920 25248
rect 6972 25236 6978 25288
rect 9048 25285 9076 25384
rect 9306 25344 9312 25356
rect 9267 25316 9312 25344
rect 9306 25304 9312 25316
rect 9364 25304 9370 25356
rect 9876 25344 9904 25384
rect 21174 25372 21180 25424
rect 21232 25412 21238 25424
rect 21232 25384 22094 25412
rect 21232 25372 21238 25384
rect 10686 25344 10692 25356
rect 9784 25316 9904 25344
rect 10647 25316 10692 25344
rect 9784 25285 9812 25316
rect 10686 25304 10692 25316
rect 10744 25304 10750 25356
rect 10870 25304 10876 25356
rect 10928 25344 10934 25356
rect 17034 25344 17040 25356
rect 10928 25316 17040 25344
rect 10928 25304 10934 25316
rect 17034 25304 17040 25316
rect 17092 25304 17098 25356
rect 18230 25304 18236 25356
rect 18288 25344 18294 25356
rect 22066 25344 22094 25384
rect 23860 25344 23888 25452
rect 30098 25440 30104 25452
rect 30156 25440 30162 25492
rect 30190 25440 30196 25492
rect 30248 25480 30254 25492
rect 37645 25483 37703 25489
rect 37645 25480 37657 25483
rect 30248 25452 37657 25480
rect 30248 25440 30254 25452
rect 37645 25449 37657 25452
rect 37691 25449 37703 25483
rect 38102 25480 38108 25492
rect 38063 25452 38108 25480
rect 37645 25443 37703 25449
rect 23934 25372 23940 25424
rect 23992 25412 23998 25424
rect 36538 25412 36544 25424
rect 23992 25384 36544 25412
rect 23992 25372 23998 25384
rect 36538 25372 36544 25384
rect 36596 25372 36602 25424
rect 18288 25316 20208 25344
rect 22066 25316 23888 25344
rect 18288 25304 18294 25316
rect 9033 25279 9091 25285
rect 9033 25245 9045 25279
rect 9079 25245 9091 25279
rect 9033 25239 9091 25245
rect 9125 25279 9183 25285
rect 9125 25245 9137 25279
rect 9171 25276 9183 25279
rect 9769 25279 9827 25285
rect 9769 25276 9781 25279
rect 9171 25248 9781 25276
rect 9171 25245 9183 25248
rect 9125 25239 9183 25245
rect 9769 25245 9781 25248
rect 9815 25245 9827 25279
rect 9769 25239 9827 25245
rect 9953 25279 10011 25285
rect 9953 25245 9965 25279
rect 9999 25276 10011 25279
rect 10042 25276 10048 25288
rect 9999 25248 10048 25276
rect 9999 25245 10011 25248
rect 9953 25239 10011 25245
rect 9306 25168 9312 25220
rect 9364 25208 9370 25220
rect 9490 25208 9496 25220
rect 9364 25180 9496 25208
rect 9364 25168 9370 25180
rect 9490 25168 9496 25180
rect 9548 25208 9554 25220
rect 9968 25208 9996 25239
rect 10042 25236 10048 25248
rect 10100 25236 10106 25288
rect 10778 25276 10784 25288
rect 10739 25248 10784 25276
rect 10778 25236 10784 25248
rect 10836 25236 10842 25288
rect 12989 25279 13047 25285
rect 12989 25245 13001 25279
rect 13035 25276 13047 25279
rect 16574 25276 16580 25288
rect 13035 25248 16580 25276
rect 13035 25245 13047 25248
rect 12989 25239 13047 25245
rect 16574 25236 16580 25248
rect 16632 25236 16638 25288
rect 16666 25236 16672 25288
rect 16724 25276 16730 25288
rect 17221 25279 17279 25285
rect 17221 25276 17233 25279
rect 16724 25248 17233 25276
rect 16724 25236 16730 25248
rect 17221 25245 17233 25248
rect 17267 25276 17279 25279
rect 20070 25276 20076 25288
rect 17267 25248 20076 25276
rect 17267 25245 17279 25248
rect 17221 25239 17279 25245
rect 20070 25236 20076 25248
rect 20128 25236 20134 25288
rect 20180 25276 20208 25316
rect 24946 25304 24952 25356
rect 25004 25344 25010 25356
rect 25225 25347 25283 25353
rect 25004 25316 25176 25344
rect 25004 25304 25010 25316
rect 20180 25248 20438 25276
rect 12158 25208 12164 25220
rect 9548 25180 9996 25208
rect 12119 25180 12164 25208
rect 9548 25168 9554 25180
rect 12158 25168 12164 25180
rect 12216 25168 12222 25220
rect 12342 25168 12348 25220
rect 12400 25217 12406 25220
rect 12400 25211 12419 25217
rect 12407 25177 12419 25211
rect 12400 25171 12419 25177
rect 14093 25211 14151 25217
rect 14093 25177 14105 25211
rect 14139 25208 14151 25211
rect 14182 25208 14188 25220
rect 14139 25180 14188 25208
rect 14139 25177 14151 25180
rect 14093 25171 14151 25177
rect 12400 25168 12406 25171
rect 14182 25168 14188 25180
rect 14240 25168 14246 25220
rect 14366 25217 14372 25220
rect 14309 25211 14372 25217
rect 14309 25177 14321 25211
rect 14355 25177 14372 25211
rect 14309 25171 14372 25177
rect 14366 25168 14372 25171
rect 14424 25168 14430 25220
rect 17488 25211 17546 25217
rect 17488 25177 17500 25211
rect 17534 25208 17546 25211
rect 18782 25208 18788 25220
rect 17534 25180 18788 25208
rect 17534 25177 17546 25180
rect 17488 25171 17546 25177
rect 18782 25168 18788 25180
rect 18840 25168 18846 25220
rect 19150 25168 19156 25220
rect 19208 25208 19214 25220
rect 19245 25211 19303 25217
rect 19245 25208 19257 25211
rect 19208 25180 19257 25208
rect 19208 25168 19214 25180
rect 19245 25177 19257 25180
rect 19291 25177 19303 25211
rect 19245 25171 19303 25177
rect 19429 25211 19487 25217
rect 19429 25177 19441 25211
rect 19475 25208 19487 25211
rect 19518 25208 19524 25220
rect 19475 25180 19524 25208
rect 19475 25177 19487 25180
rect 19429 25171 19487 25177
rect 19518 25168 19524 25180
rect 19576 25168 19582 25220
rect 20162 25168 20168 25220
rect 20220 25208 20226 25220
rect 20318 25211 20376 25217
rect 20318 25208 20330 25211
rect 20220 25180 20330 25208
rect 20220 25168 20226 25180
rect 20318 25177 20330 25180
rect 20364 25177 20376 25211
rect 20410 25208 20438 25248
rect 21266 25236 21272 25288
rect 21324 25276 21330 25288
rect 21910 25276 21916 25288
rect 21324 25248 21916 25276
rect 21324 25236 21330 25248
rect 21910 25236 21916 25248
rect 21968 25276 21974 25288
rect 22005 25279 22063 25285
rect 22005 25276 22017 25279
rect 21968 25248 22017 25276
rect 21968 25236 21974 25248
rect 22005 25245 22017 25248
rect 22051 25245 22063 25279
rect 22005 25239 22063 25245
rect 22112 25248 23520 25276
rect 22112 25208 22140 25248
rect 23382 25208 23388 25220
rect 20410 25180 22140 25208
rect 23343 25180 23388 25208
rect 20318 25171 20376 25177
rect 23382 25168 23388 25180
rect 23440 25168 23446 25220
rect 23492 25208 23520 25248
rect 24118 25236 24124 25288
rect 24176 25276 24182 25288
rect 24394 25276 24400 25288
rect 24176 25248 24400 25276
rect 24176 25236 24182 25248
rect 24394 25236 24400 25248
rect 24452 25236 24458 25288
rect 25148 25285 25176 25316
rect 25225 25313 25237 25347
rect 25271 25344 25283 25347
rect 25271 25316 25452 25344
rect 25271 25313 25283 25316
rect 25225 25307 25283 25313
rect 25133 25279 25191 25285
rect 25133 25245 25145 25279
rect 25179 25245 25191 25279
rect 25314 25276 25320 25288
rect 25275 25248 25320 25276
rect 25133 25239 25191 25245
rect 25314 25236 25320 25248
rect 25372 25236 25378 25288
rect 25424 25276 25452 25316
rect 25958 25304 25964 25356
rect 26016 25344 26022 25356
rect 37660 25344 37688 25443
rect 38102 25440 38108 25452
rect 38160 25440 38166 25492
rect 38105 25347 38163 25353
rect 38105 25344 38117 25347
rect 26016 25316 35112 25344
rect 37660 25316 38117 25344
rect 26016 25304 26022 25316
rect 25590 25276 25596 25288
rect 25424 25248 25596 25276
rect 25590 25236 25596 25248
rect 25648 25236 25654 25288
rect 30742 25236 30748 25288
rect 30800 25276 30806 25288
rect 31113 25279 31171 25285
rect 31113 25276 31125 25279
rect 30800 25248 31125 25276
rect 30800 25236 30806 25248
rect 31113 25245 31125 25248
rect 31159 25276 31171 25279
rect 31478 25276 31484 25288
rect 31159 25248 31484 25276
rect 31159 25245 31171 25248
rect 31113 25239 31171 25245
rect 31478 25236 31484 25248
rect 31536 25276 31542 25288
rect 32677 25279 32735 25285
rect 32677 25276 32689 25279
rect 31536 25248 32689 25276
rect 31536 25236 31542 25248
rect 32677 25245 32689 25248
rect 32723 25245 32735 25279
rect 32677 25239 32735 25245
rect 24670 25208 24676 25220
rect 23492 25180 24676 25208
rect 24670 25168 24676 25180
rect 24728 25168 24734 25220
rect 31662 25168 31668 25220
rect 31720 25208 31726 25220
rect 31941 25211 31999 25217
rect 31941 25208 31953 25211
rect 31720 25180 31953 25208
rect 31720 25168 31726 25180
rect 31941 25177 31953 25180
rect 31987 25177 31999 25211
rect 35084 25208 35112 25316
rect 38105 25313 38117 25316
rect 38151 25313 38163 25347
rect 38105 25307 38163 25313
rect 46293 25347 46351 25353
rect 46293 25313 46305 25347
rect 46339 25344 46351 25347
rect 47762 25344 47768 25356
rect 46339 25316 47768 25344
rect 46339 25313 46351 25316
rect 46293 25307 46351 25313
rect 47762 25304 47768 25316
rect 47820 25304 47826 25356
rect 38010 25276 38016 25288
rect 37971 25248 38016 25276
rect 38010 25236 38016 25248
rect 38068 25236 38074 25288
rect 38286 25276 38292 25288
rect 38247 25248 38292 25276
rect 38286 25236 38292 25248
rect 38344 25236 38350 25288
rect 46474 25208 46480 25220
rect 35084 25180 38516 25208
rect 46435 25180 46480 25208
rect 31941 25171 31999 25177
rect 13078 25140 13084 25152
rect 13039 25112 13084 25140
rect 13078 25100 13084 25112
rect 13136 25100 13142 25152
rect 14826 25100 14832 25152
rect 14884 25140 14890 25152
rect 17954 25140 17960 25152
rect 14884 25112 17960 25140
rect 14884 25100 14890 25112
rect 17954 25100 17960 25112
rect 18012 25100 18018 25152
rect 18230 25100 18236 25152
rect 18288 25140 18294 25152
rect 18601 25143 18659 25149
rect 18601 25140 18613 25143
rect 18288 25112 18613 25140
rect 18288 25100 18294 25112
rect 18601 25109 18613 25112
rect 18647 25109 18659 25143
rect 18601 25103 18659 25109
rect 19613 25143 19671 25149
rect 19613 25109 19625 25143
rect 19659 25140 19671 25143
rect 20530 25140 20536 25152
rect 19659 25112 20536 25140
rect 19659 25109 19671 25112
rect 19613 25103 19671 25109
rect 20530 25100 20536 25112
rect 20588 25100 20594 25152
rect 22462 25100 22468 25152
rect 22520 25140 22526 25152
rect 22922 25140 22928 25152
rect 22520 25112 22928 25140
rect 22520 25100 22526 25112
rect 22922 25100 22928 25112
rect 22980 25100 22986 25152
rect 23566 25140 23572 25152
rect 23527 25112 23572 25140
rect 23566 25100 23572 25112
rect 23624 25100 23630 25152
rect 24394 25100 24400 25152
rect 24452 25140 24458 25152
rect 24581 25143 24639 25149
rect 24581 25140 24593 25143
rect 24452 25112 24593 25140
rect 24452 25100 24458 25112
rect 24581 25109 24593 25112
rect 24627 25109 24639 25143
rect 24581 25103 24639 25109
rect 25130 25100 25136 25152
rect 25188 25140 25194 25152
rect 29822 25140 29828 25152
rect 25188 25112 29828 25140
rect 25188 25100 25194 25112
rect 29822 25100 29828 25112
rect 29880 25100 29886 25152
rect 32766 25140 32772 25152
rect 32727 25112 32772 25140
rect 32766 25100 32772 25112
rect 32824 25100 32830 25152
rect 38488 25149 38516 25180
rect 46474 25168 46480 25180
rect 46532 25168 46538 25220
rect 48130 25208 48136 25220
rect 48091 25180 48136 25208
rect 48130 25168 48136 25180
rect 48188 25168 48194 25220
rect 38473 25143 38531 25149
rect 38473 25109 38485 25143
rect 38519 25109 38531 25143
rect 38473 25103 38531 25109
rect 1104 25050 48852 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 48852 25050
rect 1104 24976 48852 24998
rect 11514 24936 11520 24948
rect 8220 24908 11520 24936
rect 7650 24800 7656 24812
rect 7611 24772 7656 24800
rect 7650 24760 7656 24772
rect 7708 24760 7714 24812
rect 2222 24692 2228 24744
rect 2280 24732 2286 24744
rect 8220 24732 8248 24908
rect 11514 24896 11520 24908
rect 11572 24896 11578 24948
rect 14093 24939 14151 24945
rect 14093 24905 14105 24939
rect 14139 24936 14151 24939
rect 14366 24936 14372 24948
rect 14139 24908 14372 24936
rect 14139 24905 14151 24908
rect 14093 24899 14151 24905
rect 14366 24896 14372 24908
rect 14424 24896 14430 24948
rect 16574 24896 16580 24948
rect 16632 24936 16638 24948
rect 18417 24939 18475 24945
rect 16632 24908 18368 24936
rect 16632 24896 16638 24908
rect 8478 24868 8484 24880
rect 8312 24840 8484 24868
rect 8312 24809 8340 24840
rect 8478 24828 8484 24840
rect 8536 24828 8542 24880
rect 10042 24828 10048 24880
rect 10100 24868 10106 24880
rect 18230 24868 18236 24880
rect 10100 24840 18236 24868
rect 10100 24828 10106 24840
rect 18230 24828 18236 24840
rect 18288 24828 18294 24880
rect 18340 24868 18368 24908
rect 18417 24905 18429 24939
rect 18463 24936 18475 24939
rect 19242 24936 19248 24948
rect 18463 24908 19248 24936
rect 18463 24905 18475 24908
rect 18417 24899 18475 24905
rect 19242 24896 19248 24908
rect 19300 24896 19306 24948
rect 20073 24939 20131 24945
rect 20073 24905 20085 24939
rect 20119 24936 20131 24939
rect 20162 24936 20168 24948
rect 20119 24908 20168 24936
rect 20119 24905 20131 24908
rect 20073 24899 20131 24905
rect 20162 24896 20168 24908
rect 20220 24896 20226 24948
rect 23566 24896 23572 24948
rect 23624 24936 23630 24948
rect 23845 24939 23903 24945
rect 23845 24936 23857 24939
rect 23624 24908 23857 24936
rect 23624 24896 23630 24908
rect 23845 24905 23857 24908
rect 23891 24936 23903 24939
rect 24670 24936 24676 24948
rect 23891 24908 24676 24936
rect 23891 24905 23903 24908
rect 23845 24899 23903 24905
rect 24670 24896 24676 24908
rect 24728 24936 24734 24948
rect 24765 24939 24823 24945
rect 24765 24936 24777 24939
rect 24728 24908 24777 24936
rect 24728 24896 24734 24908
rect 24765 24905 24777 24908
rect 24811 24905 24823 24939
rect 24765 24899 24823 24905
rect 24949 24939 25007 24945
rect 24949 24905 24961 24939
rect 24995 24936 25007 24939
rect 25498 24936 25504 24948
rect 24995 24908 25504 24936
rect 24995 24905 25007 24908
rect 24949 24899 25007 24905
rect 25498 24896 25504 24908
rect 25556 24896 25562 24948
rect 25682 24896 25688 24948
rect 25740 24936 25746 24948
rect 47486 24936 47492 24948
rect 25740 24908 47492 24936
rect 25740 24896 25746 24908
rect 47486 24896 47492 24908
rect 47544 24896 47550 24948
rect 19886 24868 19892 24880
rect 18340 24840 19892 24868
rect 19886 24828 19892 24840
rect 19944 24828 19950 24880
rect 24581 24871 24639 24877
rect 20272 24840 22508 24868
rect 8297 24803 8355 24809
rect 8297 24769 8309 24803
rect 8343 24769 8355 24803
rect 8297 24763 8355 24769
rect 13262 24760 13268 24812
rect 13320 24800 13326 24812
rect 13320 24772 13492 24800
rect 13320 24760 13326 24772
rect 2280 24704 8248 24732
rect 8481 24735 8539 24741
rect 2280 24692 2286 24704
rect 8481 24701 8493 24735
rect 8527 24701 8539 24735
rect 8481 24695 8539 24701
rect 7745 24667 7803 24673
rect 7745 24633 7757 24667
rect 7791 24664 7803 24667
rect 8496 24664 8524 24695
rect 8754 24692 8760 24744
rect 8812 24732 8818 24744
rect 11514 24732 11520 24744
rect 8812 24704 8857 24732
rect 11475 24704 11520 24732
rect 8812 24692 8818 24704
rect 11514 24692 11520 24704
rect 11572 24692 11578 24744
rect 11701 24735 11759 24741
rect 11701 24701 11713 24735
rect 11747 24732 11759 24735
rect 13078 24732 13084 24744
rect 11747 24704 13084 24732
rect 11747 24701 11759 24704
rect 11701 24695 11759 24701
rect 13078 24692 13084 24704
rect 13136 24692 13142 24744
rect 13354 24732 13360 24744
rect 13315 24704 13360 24732
rect 13354 24692 13360 24704
rect 13412 24692 13418 24744
rect 13464 24732 13492 24772
rect 13722 24760 13728 24812
rect 13780 24800 13786 24812
rect 13817 24803 13875 24809
rect 13817 24800 13829 24803
rect 13780 24772 13829 24800
rect 13780 24760 13786 24772
rect 13817 24769 13829 24772
rect 13863 24769 13875 24803
rect 13817 24763 13875 24769
rect 17221 24803 17279 24809
rect 17221 24769 17233 24803
rect 17267 24769 17279 24803
rect 17402 24800 17408 24812
rect 17363 24772 17408 24800
rect 17221 24763 17279 24769
rect 14093 24735 14151 24741
rect 14093 24732 14105 24735
rect 13464 24704 14105 24732
rect 14093 24701 14105 24704
rect 14139 24732 14151 24735
rect 14182 24732 14188 24744
rect 14139 24704 14188 24732
rect 14139 24701 14151 24704
rect 14093 24695 14151 24701
rect 14182 24692 14188 24704
rect 14240 24692 14246 24744
rect 17236 24732 17264 24763
rect 17402 24760 17408 24772
rect 17460 24760 17466 24812
rect 17589 24803 17647 24809
rect 17589 24769 17601 24803
rect 17635 24800 17647 24803
rect 17678 24800 17684 24812
rect 17635 24772 17684 24800
rect 17635 24769 17647 24772
rect 17589 24763 17647 24769
rect 17678 24760 17684 24772
rect 17736 24760 17742 24812
rect 18049 24803 18107 24809
rect 18049 24769 18061 24803
rect 18095 24800 18107 24803
rect 19150 24800 19156 24812
rect 18095 24772 19156 24800
rect 18095 24769 18107 24772
rect 18049 24763 18107 24769
rect 18064 24732 18092 24763
rect 19150 24760 19156 24772
rect 19208 24760 19214 24812
rect 19426 24760 19432 24812
rect 19484 24800 19490 24812
rect 20272 24800 20300 24840
rect 19484 24772 20300 24800
rect 20349 24803 20407 24809
rect 19484 24760 19490 24772
rect 20349 24769 20361 24803
rect 20395 24769 20407 24803
rect 20349 24763 20407 24769
rect 20441 24803 20499 24809
rect 20441 24769 20453 24803
rect 20487 24769 20499 24803
rect 20441 24763 20499 24769
rect 17236 24704 18092 24732
rect 18414 24692 18420 24744
rect 18472 24732 18478 24744
rect 18782 24732 18788 24744
rect 18472 24704 18788 24732
rect 18472 24692 18478 24704
rect 18782 24692 18788 24704
rect 18840 24692 18846 24744
rect 7791 24636 8524 24664
rect 8588 24636 17264 24664
rect 7791 24633 7803 24636
rect 7745 24627 7803 24633
rect 1578 24556 1584 24608
rect 1636 24596 1642 24608
rect 8588 24596 8616 24636
rect 1636 24568 8616 24596
rect 1636 24556 1642 24568
rect 12250 24556 12256 24608
rect 12308 24596 12314 24608
rect 13446 24596 13452 24608
rect 12308 24568 13452 24596
rect 12308 24556 12314 24568
rect 13446 24556 13452 24568
rect 13504 24556 13510 24608
rect 13538 24556 13544 24608
rect 13596 24596 13602 24608
rect 13909 24599 13967 24605
rect 13909 24596 13921 24599
rect 13596 24568 13921 24596
rect 13596 24556 13602 24568
rect 13909 24565 13921 24568
rect 13955 24596 13967 24599
rect 15102 24596 15108 24608
rect 13955 24568 15108 24596
rect 13955 24565 13967 24568
rect 13909 24559 13967 24565
rect 15102 24556 15108 24568
rect 15160 24556 15166 24608
rect 17236 24596 17264 24636
rect 17402 24624 17408 24676
rect 17460 24664 17466 24676
rect 18046 24664 18052 24676
rect 17460 24636 18052 24664
rect 17460 24624 17466 24636
rect 18046 24624 18052 24636
rect 18104 24624 18110 24676
rect 20364 24664 20392 24763
rect 20456 24732 20484 24763
rect 20530 24760 20536 24812
rect 20588 24800 20594 24812
rect 20588 24772 20633 24800
rect 20588 24760 20594 24772
rect 20714 24760 20720 24812
rect 20772 24800 20778 24812
rect 20824 24800 20852 24840
rect 20772 24772 20865 24800
rect 20772 24760 20778 24772
rect 21818 24760 21824 24812
rect 21876 24800 21882 24812
rect 22051 24803 22109 24809
rect 22051 24800 22063 24803
rect 21876 24772 22063 24800
rect 21876 24760 21882 24772
rect 22051 24769 22063 24772
rect 22097 24769 22109 24803
rect 22051 24763 22109 24769
rect 22189 24806 22247 24812
rect 22480 24809 22508 24840
rect 24581 24837 24593 24871
rect 24627 24868 24639 24871
rect 24854 24868 24860 24880
rect 24627 24840 24860 24868
rect 24627 24837 24639 24840
rect 24581 24831 24639 24837
rect 24854 24828 24860 24840
rect 24912 24828 24918 24880
rect 25516 24840 29224 24868
rect 22189 24772 22201 24806
rect 22235 24772 22247 24806
rect 22189 24766 22247 24772
rect 22281 24803 22339 24809
rect 22281 24769 22293 24803
rect 22327 24769 22339 24803
rect 20806 24732 20812 24744
rect 20456 24704 20812 24732
rect 20806 24692 20812 24704
rect 20864 24732 20870 24744
rect 20864 24704 22048 24732
rect 20864 24692 20870 24704
rect 21910 24664 21916 24676
rect 20364 24636 21916 24664
rect 21910 24624 21916 24636
rect 21968 24624 21974 24676
rect 22020 24664 22048 24704
rect 22204 24664 22232 24766
rect 22281 24763 22339 24769
rect 22465 24803 22523 24809
rect 22465 24769 22477 24803
rect 22511 24769 22523 24803
rect 22465 24763 22523 24769
rect 23753 24803 23811 24809
rect 23753 24769 23765 24803
rect 23799 24769 23811 24803
rect 23934 24800 23940 24812
rect 23895 24772 23940 24800
rect 23753 24763 23811 24769
rect 22296 24732 22324 24763
rect 22738 24732 22744 24744
rect 22296 24704 22744 24732
rect 22738 24692 22744 24704
rect 22796 24692 22802 24744
rect 23774 24732 23802 24763
rect 23934 24760 23940 24772
rect 23992 24760 23998 24812
rect 24673 24803 24731 24809
rect 24673 24769 24685 24803
rect 24719 24800 24731 24803
rect 24946 24800 24952 24812
rect 24719 24772 24952 24800
rect 24719 24769 24731 24772
rect 24673 24763 24731 24769
rect 24946 24760 24952 24772
rect 25004 24800 25010 24812
rect 25516 24809 25544 24840
rect 25501 24803 25559 24809
rect 25501 24800 25513 24803
rect 25004 24772 25513 24800
rect 25004 24760 25010 24772
rect 25501 24769 25513 24772
rect 25547 24769 25559 24803
rect 25501 24763 25559 24769
rect 27154 24760 27160 24812
rect 27212 24800 27218 24812
rect 27249 24803 27307 24809
rect 27249 24800 27261 24803
rect 27212 24772 27261 24800
rect 27212 24760 27218 24772
rect 27249 24769 27261 24772
rect 27295 24769 27307 24803
rect 27249 24763 27307 24769
rect 27341 24803 27399 24809
rect 27341 24769 27353 24803
rect 27387 24769 27399 24803
rect 27341 24763 27399 24769
rect 25222 24732 25228 24744
rect 23774 24704 25228 24732
rect 25222 24692 25228 24704
rect 25280 24692 25286 24744
rect 22020 24636 22232 24664
rect 24397 24667 24455 24673
rect 24397 24633 24409 24667
rect 24443 24633 24455 24667
rect 24397 24627 24455 24633
rect 21542 24596 21548 24608
rect 17236 24568 21548 24596
rect 21542 24556 21548 24568
rect 21600 24556 21606 24608
rect 21818 24596 21824 24608
rect 21779 24568 21824 24596
rect 21818 24556 21824 24568
rect 21876 24556 21882 24608
rect 23474 24556 23480 24608
rect 23532 24596 23538 24608
rect 24412 24596 24440 24627
rect 24578 24624 24584 24676
rect 24636 24664 24642 24676
rect 25593 24667 25651 24673
rect 25593 24664 25605 24667
rect 24636 24636 25605 24664
rect 24636 24624 24642 24636
rect 25593 24633 25605 24636
rect 25639 24633 25651 24667
rect 25593 24627 25651 24633
rect 26694 24624 26700 24676
rect 26752 24664 26758 24676
rect 27356 24664 27384 24763
rect 27430 24760 27436 24812
rect 27488 24800 27494 24812
rect 27488 24772 27533 24800
rect 27488 24760 27494 24772
rect 27614 24760 27620 24812
rect 27672 24800 27678 24812
rect 28902 24800 28908 24812
rect 27672 24772 28908 24800
rect 27672 24760 27678 24772
rect 28902 24760 28908 24772
rect 28960 24760 28966 24812
rect 29196 24732 29224 24840
rect 29270 24828 29276 24880
rect 29328 24868 29334 24880
rect 31478 24868 31484 24880
rect 29328 24840 29705 24868
rect 31439 24840 31484 24868
rect 29328 24828 29334 24840
rect 29677 24812 29705 24840
rect 31478 24828 31484 24840
rect 31536 24828 31542 24880
rect 37461 24871 37519 24877
rect 37461 24868 37473 24871
rect 37292 24840 37473 24868
rect 29362 24760 29368 24812
rect 29420 24809 29426 24812
rect 29420 24803 29469 24809
rect 29420 24769 29423 24803
rect 29457 24769 29469 24803
rect 29420 24763 29469 24769
rect 29530 24803 29588 24809
rect 29530 24769 29542 24803
rect 29576 24769 29588 24803
rect 29530 24766 29588 24769
rect 29662 24806 29720 24812
rect 29662 24772 29674 24806
rect 29708 24772 29720 24806
rect 29662 24766 29720 24772
rect 29825 24803 29883 24809
rect 29825 24769 29837 24803
rect 29871 24800 29883 24803
rect 30190 24800 30196 24812
rect 29871 24772 30196 24800
rect 29871 24769 29883 24772
rect 29530 24763 29592 24766
rect 29825 24763 29883 24769
rect 29420 24760 29426 24763
rect 29544 24744 29592 24763
rect 30190 24760 30196 24772
rect 30248 24760 30254 24812
rect 30374 24760 30380 24812
rect 30432 24800 30438 24812
rect 30837 24803 30895 24809
rect 30837 24800 30849 24803
rect 30432 24772 30849 24800
rect 30432 24760 30438 24772
rect 30837 24769 30849 24772
rect 30883 24800 30895 24803
rect 31297 24803 31355 24809
rect 31297 24800 31309 24803
rect 30883 24772 31309 24800
rect 30883 24769 30895 24772
rect 30837 24763 30895 24769
rect 31297 24769 31309 24772
rect 31343 24769 31355 24803
rect 31297 24763 31355 24769
rect 32214 24760 32220 24812
rect 32272 24800 32278 24812
rect 32585 24803 32643 24809
rect 32585 24800 32597 24803
rect 32272 24772 32597 24800
rect 32272 24760 32278 24772
rect 32585 24769 32597 24772
rect 32631 24800 32643 24803
rect 33134 24800 33140 24812
rect 32631 24772 33140 24800
rect 32631 24769 32643 24772
rect 32585 24763 32643 24769
rect 33134 24760 33140 24772
rect 33192 24760 33198 24812
rect 33318 24760 33324 24812
rect 33376 24800 33382 24812
rect 33597 24803 33655 24809
rect 33597 24800 33609 24803
rect 33376 24772 33609 24800
rect 33376 24760 33382 24772
rect 33597 24769 33609 24772
rect 33643 24769 33655 24803
rect 36538 24800 36544 24812
rect 36499 24772 36544 24800
rect 33597 24763 33655 24769
rect 36538 24760 36544 24772
rect 36596 24760 36602 24812
rect 36633 24803 36691 24809
rect 36633 24769 36645 24803
rect 36679 24800 36691 24803
rect 37292 24800 37320 24840
rect 37461 24837 37473 24840
rect 37507 24837 37519 24871
rect 37461 24831 37519 24837
rect 39114 24800 39120 24812
rect 36679 24772 37320 24800
rect 39075 24772 39120 24800
rect 36679 24769 36691 24772
rect 36633 24763 36691 24769
rect 39114 24760 39120 24772
rect 39172 24760 39178 24812
rect 47946 24800 47952 24812
rect 47907 24772 47952 24800
rect 47946 24760 47952 24772
rect 48004 24760 48010 24812
rect 29544 24738 29552 24744
rect 29196 24704 29408 24732
rect 29270 24664 29276 24676
rect 26752 24636 29276 24664
rect 26752 24624 26758 24636
rect 29270 24624 29276 24636
rect 29328 24624 29334 24676
rect 29380 24664 29408 24704
rect 29546 24692 29552 24738
rect 29604 24692 29610 24744
rect 33781 24735 33839 24741
rect 33781 24701 33793 24735
rect 33827 24732 33839 24735
rect 34790 24732 34796 24744
rect 33827 24704 34796 24732
rect 33827 24701 33839 24704
rect 33781 24695 33839 24701
rect 34790 24692 34796 24704
rect 34848 24692 34854 24744
rect 35434 24732 35440 24744
rect 35395 24704 35440 24732
rect 35434 24692 35440 24704
rect 35492 24692 35498 24744
rect 35618 24692 35624 24744
rect 35676 24732 35682 24744
rect 37277 24735 37335 24741
rect 37277 24732 37289 24735
rect 35676 24704 37289 24732
rect 35676 24692 35682 24704
rect 37277 24701 37289 24704
rect 37323 24701 37335 24735
rect 37277 24695 37335 24701
rect 37384 24704 38654 24732
rect 37384 24664 37412 24704
rect 29380 24636 37412 24664
rect 38626 24664 38654 24704
rect 48133 24667 48191 24673
rect 48133 24664 48145 24667
rect 38626 24636 48145 24664
rect 48133 24633 48145 24636
rect 48179 24633 48191 24667
rect 48133 24627 48191 24633
rect 25314 24596 25320 24608
rect 23532 24568 25320 24596
rect 23532 24556 23538 24568
rect 25314 24556 25320 24568
rect 25372 24556 25378 24608
rect 26973 24599 27031 24605
rect 26973 24565 26985 24599
rect 27019 24596 27031 24599
rect 27062 24596 27068 24608
rect 27019 24568 27068 24596
rect 27019 24565 27031 24568
rect 26973 24559 27031 24565
rect 27062 24556 27068 24568
rect 27120 24556 27126 24608
rect 29181 24599 29239 24605
rect 29181 24565 29193 24599
rect 29227 24596 29239 24599
rect 29822 24596 29828 24608
rect 29227 24568 29828 24596
rect 29227 24565 29239 24568
rect 29181 24559 29239 24565
rect 29822 24556 29828 24568
rect 29880 24556 29886 24608
rect 32490 24556 32496 24608
rect 32548 24596 32554 24608
rect 32677 24599 32735 24605
rect 32677 24596 32689 24599
rect 32548 24568 32689 24596
rect 32548 24556 32554 24568
rect 32677 24565 32689 24568
rect 32723 24565 32735 24599
rect 32677 24559 32735 24565
rect 32766 24556 32772 24608
rect 32824 24596 32830 24608
rect 36538 24596 36544 24608
rect 32824 24568 36544 24596
rect 32824 24556 32830 24568
rect 36538 24556 36544 24568
rect 36596 24596 36602 24608
rect 37366 24596 37372 24608
rect 36596 24568 37372 24596
rect 36596 24556 36602 24568
rect 37366 24556 37372 24568
rect 37424 24556 37430 24608
rect 38562 24556 38568 24608
rect 38620 24596 38626 24608
rect 39114 24596 39120 24608
rect 38620 24568 39120 24596
rect 38620 24556 38626 24568
rect 39114 24556 39120 24568
rect 39172 24556 39178 24608
rect 1104 24506 48852 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 48852 24506
rect 1104 24432 48852 24454
rect 1578 24392 1584 24404
rect 1539 24364 1584 24392
rect 1578 24352 1584 24364
rect 1636 24352 1642 24404
rect 1762 24352 1768 24404
rect 1820 24392 1826 24404
rect 10413 24395 10471 24401
rect 1820 24364 2774 24392
rect 1820 24352 1826 24364
rect 2746 24324 2774 24364
rect 10413 24361 10425 24395
rect 10459 24392 10471 24395
rect 10686 24392 10692 24404
rect 10459 24364 10692 24392
rect 10459 24361 10471 24364
rect 10413 24355 10471 24361
rect 10686 24352 10692 24364
rect 10744 24352 10750 24404
rect 12342 24352 12348 24404
rect 12400 24392 12406 24404
rect 12437 24395 12495 24401
rect 12437 24392 12449 24395
rect 12400 24364 12449 24392
rect 12400 24352 12406 24364
rect 12437 24361 12449 24364
rect 12483 24361 12495 24395
rect 13262 24392 13268 24404
rect 13223 24364 13268 24392
rect 12437 24355 12495 24361
rect 13262 24352 13268 24364
rect 13320 24352 13326 24404
rect 13446 24392 13452 24404
rect 13407 24364 13452 24392
rect 13446 24352 13452 24364
rect 13504 24352 13510 24404
rect 13722 24352 13728 24404
rect 13780 24392 13786 24404
rect 14093 24395 14151 24401
rect 14093 24392 14105 24395
rect 13780 24364 14105 24392
rect 13780 24352 13786 24364
rect 14093 24361 14105 24364
rect 14139 24361 14151 24395
rect 14093 24355 14151 24361
rect 14642 24352 14648 24404
rect 14700 24392 14706 24404
rect 22646 24392 22652 24404
rect 14700 24364 22508 24392
rect 22607 24364 22652 24392
rect 14700 24352 14706 24364
rect 22480 24324 22508 24364
rect 22646 24352 22652 24364
rect 22704 24352 22710 24404
rect 32766 24392 32772 24404
rect 22756 24364 32772 24392
rect 22756 24324 22784 24364
rect 32766 24352 32772 24364
rect 32824 24352 32830 24404
rect 34790 24392 34796 24404
rect 34751 24364 34796 24392
rect 34790 24352 34796 24364
rect 34848 24352 34854 24404
rect 2746 24296 22416 24324
rect 22480 24296 22784 24324
rect 3789 24259 3847 24265
rect 3789 24225 3801 24259
rect 3835 24256 3847 24259
rect 8202 24256 8208 24268
rect 3835 24228 8208 24256
rect 3835 24225 3847 24228
rect 3789 24219 3847 24225
rect 8202 24216 8208 24228
rect 8260 24216 8266 24268
rect 10137 24259 10195 24265
rect 10137 24225 10149 24259
rect 10183 24256 10195 24259
rect 12250 24256 12256 24268
rect 10183 24228 12256 24256
rect 10183 24225 10195 24228
rect 10137 24219 10195 24225
rect 12250 24216 12256 24228
rect 12308 24216 12314 24268
rect 13081 24259 13139 24265
rect 13081 24225 13093 24259
rect 13127 24256 13139 24259
rect 13906 24256 13912 24268
rect 13127 24228 13912 24256
rect 13127 24225 13139 24228
rect 13081 24219 13139 24225
rect 13906 24216 13912 24228
rect 13964 24216 13970 24268
rect 18138 24256 18144 24268
rect 18099 24228 18144 24256
rect 18138 24216 18144 24228
rect 18196 24216 18202 24268
rect 20257 24259 20315 24265
rect 20257 24225 20269 24259
rect 20303 24256 20315 24259
rect 22388 24256 22416 24296
rect 23290 24284 23296 24336
rect 23348 24324 23354 24336
rect 23934 24324 23940 24336
rect 23348 24296 23940 24324
rect 23348 24284 23354 24296
rect 23934 24284 23940 24296
rect 23992 24284 23998 24336
rect 28997 24327 29055 24333
rect 28997 24293 29009 24327
rect 29043 24324 29055 24327
rect 29178 24324 29184 24336
rect 29043 24296 29184 24324
rect 29043 24293 29055 24296
rect 28997 24287 29055 24293
rect 29178 24284 29184 24296
rect 29236 24284 29242 24336
rect 32674 24284 32680 24336
rect 32732 24324 32738 24336
rect 43990 24324 43996 24336
rect 32732 24296 43996 24324
rect 32732 24284 32738 24296
rect 43990 24284 43996 24296
rect 44048 24284 44054 24336
rect 26602 24256 26608 24268
rect 20303 24228 22324 24256
rect 22388 24228 25728 24256
rect 20303 24225 20315 24228
rect 20257 24219 20315 24225
rect 1394 24188 1400 24200
rect 1355 24160 1400 24188
rect 1394 24148 1400 24160
rect 1452 24148 1458 24200
rect 3053 24191 3111 24197
rect 3053 24157 3065 24191
rect 3099 24157 3111 24191
rect 3053 24151 3111 24157
rect 3068 24064 3096 24151
rect 8846 24148 8852 24200
rect 8904 24188 8910 24200
rect 9950 24188 9956 24200
rect 8904 24160 9956 24188
rect 8904 24148 8910 24160
rect 9950 24148 9956 24160
rect 10008 24188 10014 24200
rect 10045 24191 10103 24197
rect 10045 24188 10057 24191
rect 10008 24160 10057 24188
rect 10008 24148 10014 24160
rect 10045 24157 10057 24160
rect 10091 24157 10103 24191
rect 10045 24151 10103 24157
rect 12345 24191 12403 24197
rect 12345 24157 12357 24191
rect 12391 24157 12403 24191
rect 12345 24151 12403 24157
rect 12529 24191 12587 24197
rect 12529 24157 12541 24191
rect 12575 24188 12587 24191
rect 12894 24188 12900 24200
rect 12575 24160 12900 24188
rect 12575 24157 12587 24160
rect 12529 24151 12587 24157
rect 3145 24123 3203 24129
rect 3145 24089 3157 24123
rect 3191 24120 3203 24123
rect 3973 24123 4031 24129
rect 3973 24120 3985 24123
rect 3191 24092 3985 24120
rect 3191 24089 3203 24092
rect 3145 24083 3203 24089
rect 3973 24089 3985 24092
rect 4019 24089 4031 24123
rect 3973 24083 4031 24089
rect 4062 24080 4068 24132
rect 4120 24120 4126 24132
rect 5629 24123 5687 24129
rect 5629 24120 5641 24123
rect 4120 24092 5641 24120
rect 4120 24080 4126 24092
rect 5629 24089 5641 24092
rect 5675 24089 5687 24123
rect 12250 24120 12256 24132
rect 5629 24083 5687 24089
rect 5736 24092 12256 24120
rect 3050 24052 3056 24064
rect 2963 24024 3056 24052
rect 3050 24012 3056 24024
rect 3108 24052 3114 24064
rect 5736 24052 5764 24092
rect 12250 24080 12256 24092
rect 12308 24080 12314 24132
rect 3108 24024 5764 24052
rect 12360 24052 12388 24151
rect 12894 24148 12900 24160
rect 12952 24188 12958 24200
rect 13265 24191 13323 24197
rect 13265 24188 13277 24191
rect 12952 24160 13277 24188
rect 12952 24148 12958 24160
rect 13265 24157 13277 24160
rect 13311 24157 13323 24191
rect 13265 24151 13323 24157
rect 14093 24191 14151 24197
rect 14093 24157 14105 24191
rect 14139 24157 14151 24191
rect 14093 24151 14151 24157
rect 12986 24120 12992 24132
rect 12947 24092 12992 24120
rect 12986 24080 12992 24092
rect 13044 24120 13050 24132
rect 14108 24120 14136 24151
rect 14182 24148 14188 24200
rect 14240 24188 14246 24200
rect 14277 24191 14335 24197
rect 14277 24188 14289 24191
rect 14240 24160 14289 24188
rect 14240 24148 14246 24160
rect 14277 24157 14289 24160
rect 14323 24188 14335 24191
rect 16942 24188 16948 24200
rect 14323 24160 16948 24188
rect 14323 24157 14335 24160
rect 14277 24151 14335 24157
rect 16942 24148 16948 24160
rect 17000 24148 17006 24200
rect 17862 24188 17868 24200
rect 17823 24160 17868 24188
rect 17862 24148 17868 24160
rect 17920 24148 17926 24200
rect 19150 24148 19156 24200
rect 19208 24188 19214 24200
rect 19889 24191 19947 24197
rect 19889 24188 19901 24191
rect 19208 24160 19901 24188
rect 19208 24148 19214 24160
rect 19889 24157 19901 24160
rect 19935 24157 19947 24191
rect 19889 24151 19947 24157
rect 20073 24191 20131 24197
rect 20073 24157 20085 24191
rect 20119 24188 20131 24191
rect 22186 24188 22192 24200
rect 20119 24160 22192 24188
rect 20119 24157 20131 24160
rect 20073 24151 20131 24157
rect 22186 24148 22192 24160
rect 22244 24148 22250 24200
rect 22296 24188 22324 24228
rect 22738 24188 22744 24200
rect 22296 24160 22744 24188
rect 22738 24148 22744 24160
rect 22796 24148 22802 24200
rect 23658 24148 23664 24200
rect 23716 24188 23722 24200
rect 24578 24188 24584 24200
rect 23716 24160 24584 24188
rect 23716 24148 23722 24160
rect 24578 24148 24584 24160
rect 24636 24148 24642 24200
rect 24670 24148 24676 24200
rect 24728 24188 24734 24200
rect 25130 24188 25136 24200
rect 24728 24160 24773 24188
rect 25043 24160 25136 24188
rect 24728 24148 24734 24160
rect 25130 24148 25136 24160
rect 25188 24188 25194 24200
rect 25590 24188 25596 24200
rect 25188 24160 25596 24188
rect 25188 24148 25194 24160
rect 25590 24148 25596 24160
rect 25648 24148 25654 24200
rect 25700 24188 25728 24228
rect 26068 24228 26608 24256
rect 26068 24197 26096 24228
rect 26602 24216 26608 24228
rect 26660 24216 26666 24268
rect 26786 24256 26792 24268
rect 26747 24228 26792 24256
rect 26786 24216 26792 24228
rect 26844 24216 26850 24268
rect 32490 24256 32496 24268
rect 32451 24228 32496 24256
rect 32490 24216 32496 24228
rect 32548 24216 32554 24268
rect 33134 24216 33140 24268
rect 33192 24256 33198 24268
rect 37274 24256 37280 24268
rect 33192 24228 34744 24256
rect 37235 24228 37280 24256
rect 33192 24216 33198 24228
rect 25961 24191 26019 24197
rect 25961 24188 25973 24191
rect 25700 24160 25973 24188
rect 25961 24157 25973 24160
rect 26007 24157 26019 24191
rect 25961 24151 26019 24157
rect 26053 24191 26111 24197
rect 26053 24157 26065 24191
rect 26099 24157 26111 24191
rect 26053 24151 26111 24157
rect 26145 24191 26203 24197
rect 26145 24157 26157 24191
rect 26191 24188 26203 24191
rect 26234 24188 26240 24200
rect 26191 24160 26240 24188
rect 26191 24157 26203 24160
rect 26145 24151 26203 24157
rect 26234 24148 26240 24160
rect 26292 24148 26298 24200
rect 26326 24148 26332 24200
rect 26384 24188 26390 24200
rect 29546 24188 29552 24200
rect 26384 24160 26429 24188
rect 29507 24160 29552 24188
rect 26384 24148 26390 24160
rect 29546 24148 29552 24160
rect 29604 24148 29610 24200
rect 29822 24197 29828 24200
rect 29816 24151 29828 24197
rect 29880 24188 29886 24200
rect 32306 24188 32312 24200
rect 29880 24160 29916 24188
rect 32267 24160 32312 24188
rect 29822 24148 29828 24151
rect 29880 24148 29886 24160
rect 32306 24148 32312 24160
rect 32364 24148 32370 24200
rect 34716 24197 34744 24228
rect 37274 24216 37280 24228
rect 37332 24216 37338 24268
rect 46934 24216 46940 24268
rect 46992 24256 46998 24268
rect 47581 24259 47639 24265
rect 47581 24256 47593 24259
rect 46992 24228 47593 24256
rect 46992 24216 46998 24228
rect 47581 24225 47593 24228
rect 47627 24225 47639 24259
rect 47581 24219 47639 24225
rect 34701 24191 34759 24197
rect 34701 24157 34713 24191
rect 34747 24157 34759 24191
rect 47302 24188 47308 24200
rect 47263 24160 47308 24188
rect 34701 24151 34759 24157
rect 47302 24148 47308 24160
rect 47360 24148 47366 24200
rect 21358 24120 21364 24132
rect 13044 24092 14136 24120
rect 21319 24092 21364 24120
rect 13044 24080 13050 24092
rect 21358 24080 21364 24092
rect 21416 24080 21422 24132
rect 21542 24080 21548 24132
rect 21600 24120 21606 24132
rect 23842 24120 23848 24132
rect 21600 24092 23848 24120
rect 21600 24080 21606 24092
rect 23842 24080 23848 24092
rect 23900 24080 23906 24132
rect 25041 24123 25099 24129
rect 25041 24089 25053 24123
rect 25087 24089 25099 24123
rect 25041 24083 25099 24089
rect 25685 24123 25743 24129
rect 25685 24089 25697 24123
rect 25731 24120 25743 24123
rect 27034 24123 27092 24129
rect 27034 24120 27046 24123
rect 25731 24092 27046 24120
rect 25731 24089 25743 24092
rect 25685 24083 25743 24089
rect 27034 24089 27046 24092
rect 27080 24089 27092 24123
rect 27034 24083 27092 24089
rect 14274 24052 14280 24064
rect 12360 24024 14280 24052
rect 3108 24012 3114 24024
rect 14274 24012 14280 24024
rect 14332 24052 14338 24064
rect 14461 24055 14519 24061
rect 14461 24052 14473 24055
rect 14332 24024 14473 24052
rect 14332 24012 14338 24024
rect 14461 24021 14473 24024
rect 14507 24021 14519 24055
rect 14461 24015 14519 24021
rect 17586 24012 17592 24064
rect 17644 24052 17650 24064
rect 20162 24052 20168 24064
rect 17644 24024 20168 24052
rect 17644 24012 17650 24024
rect 20162 24012 20168 24024
rect 20220 24012 20226 24064
rect 25056 24052 25084 24083
rect 28442 24080 28448 24132
rect 28500 24120 28506 24132
rect 28629 24123 28687 24129
rect 28629 24120 28641 24123
rect 28500 24092 28641 24120
rect 28500 24080 28506 24092
rect 28629 24089 28641 24092
rect 28675 24089 28687 24123
rect 28629 24083 28687 24089
rect 28813 24123 28871 24129
rect 28813 24089 28825 24123
rect 28859 24089 28871 24123
rect 28813 24083 28871 24089
rect 34149 24123 34207 24129
rect 34149 24089 34161 24123
rect 34195 24089 34207 24123
rect 37458 24120 37464 24132
rect 37419 24092 37464 24120
rect 34149 24083 34207 24089
rect 27982 24052 27988 24064
rect 25056 24024 27988 24052
rect 27982 24012 27988 24024
rect 28040 24012 28046 24064
rect 28166 24052 28172 24064
rect 28127 24024 28172 24052
rect 28166 24012 28172 24024
rect 28224 24012 28230 24064
rect 28534 24012 28540 24064
rect 28592 24052 28598 24064
rect 28828 24052 28856 24083
rect 30929 24055 30987 24061
rect 30929 24052 30941 24055
rect 28592 24024 30941 24052
rect 28592 24012 28598 24024
rect 30929 24021 30941 24024
rect 30975 24021 30987 24055
rect 34164 24052 34192 24083
rect 37458 24080 37464 24092
rect 37516 24080 37522 24132
rect 39114 24120 39120 24132
rect 39075 24092 39120 24120
rect 39114 24080 39120 24092
rect 39172 24080 39178 24132
rect 38654 24052 38660 24064
rect 34164 24024 38660 24052
rect 30929 24015 30987 24021
rect 38654 24012 38660 24024
rect 38712 24012 38718 24064
rect 1104 23962 48852 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 48852 23962
rect 1104 23888 48852 23910
rect 4706 23808 4712 23860
rect 4764 23848 4770 23860
rect 4764 23820 17954 23848
rect 4764 23808 4770 23820
rect 8294 23780 8300 23792
rect 7852 23752 8300 23780
rect 7852 23721 7880 23752
rect 8294 23740 8300 23752
rect 8352 23740 8358 23792
rect 17221 23783 17279 23789
rect 17221 23749 17233 23783
rect 17267 23780 17279 23783
rect 17586 23780 17592 23792
rect 17267 23752 17592 23780
rect 17267 23749 17279 23752
rect 17221 23743 17279 23749
rect 17586 23740 17592 23752
rect 17644 23740 17650 23792
rect 17926 23780 17954 23820
rect 19150 23808 19156 23860
rect 19208 23848 19214 23860
rect 19337 23851 19395 23857
rect 19337 23848 19349 23851
rect 19208 23820 19349 23848
rect 19208 23808 19214 23820
rect 19337 23817 19349 23820
rect 19383 23817 19395 23851
rect 27154 23848 27160 23860
rect 19337 23811 19395 23817
rect 23124 23820 27160 23848
rect 23124 23780 23152 23820
rect 27154 23808 27160 23820
rect 27212 23808 27218 23860
rect 27982 23808 27988 23860
rect 28040 23848 28046 23860
rect 30466 23848 30472 23860
rect 28040 23820 30472 23848
rect 28040 23808 28046 23820
rect 30466 23808 30472 23820
rect 30524 23808 30530 23860
rect 31113 23851 31171 23857
rect 31113 23817 31125 23851
rect 31159 23817 31171 23851
rect 37458 23848 37464 23860
rect 37419 23820 37464 23848
rect 31113 23811 31171 23817
rect 23474 23780 23480 23792
rect 17926 23752 23152 23780
rect 23216 23752 23480 23780
rect 7837 23715 7895 23721
rect 7837 23681 7849 23715
rect 7883 23681 7895 23715
rect 7837 23675 7895 23681
rect 8104 23715 8162 23721
rect 8104 23681 8116 23715
rect 8150 23712 8162 23715
rect 8938 23712 8944 23724
rect 8150 23684 8944 23712
rect 8150 23681 8162 23684
rect 8104 23675 8162 23681
rect 8938 23672 8944 23684
rect 8996 23672 9002 23724
rect 12986 23672 12992 23724
rect 13044 23712 13050 23724
rect 13173 23715 13231 23721
rect 13173 23712 13185 23715
rect 13044 23684 13185 23712
rect 13044 23672 13050 23684
rect 13173 23681 13185 23684
rect 13219 23681 13231 23715
rect 13173 23675 13231 23681
rect 13906 23672 13912 23724
rect 13964 23712 13970 23724
rect 14642 23712 14648 23724
rect 13964 23684 14057 23712
rect 14603 23684 14648 23712
rect 13964 23672 13970 23684
rect 14642 23672 14648 23684
rect 14700 23672 14706 23724
rect 17328 23702 18184 23712
rect 17297 23684 18184 23702
rect 17297 23674 17356 23684
rect 13924 23644 13952 23672
rect 15102 23644 15108 23656
rect 13924 23616 15108 23644
rect 15102 23604 15108 23616
rect 15160 23604 15166 23656
rect 11514 23536 11520 23588
rect 11572 23576 11578 23588
rect 17297 23576 17325 23674
rect 17586 23604 17592 23656
rect 17644 23644 17650 23656
rect 18049 23647 18107 23653
rect 18049 23644 18061 23647
rect 17644 23616 18061 23644
rect 17644 23604 17650 23616
rect 18049 23613 18061 23616
rect 18095 23613 18107 23647
rect 18049 23607 18107 23613
rect 11572 23548 17325 23576
rect 17405 23579 17463 23585
rect 11572 23536 11578 23548
rect 17405 23545 17417 23579
rect 17451 23576 17463 23579
rect 17954 23576 17960 23588
rect 17451 23548 17960 23576
rect 17451 23545 17463 23548
rect 17405 23539 17463 23545
rect 17954 23536 17960 23548
rect 18012 23536 18018 23588
rect 18156 23576 18184 23684
rect 19242 23672 19248 23724
rect 19300 23712 19306 23724
rect 19521 23715 19579 23721
rect 19521 23712 19533 23715
rect 19300 23684 19533 23712
rect 19300 23672 19306 23684
rect 19521 23681 19533 23684
rect 19567 23681 19579 23715
rect 19521 23675 19579 23681
rect 18325 23647 18383 23653
rect 18325 23613 18337 23647
rect 18371 23644 18383 23647
rect 19426 23644 19432 23656
rect 18371 23616 19432 23644
rect 18371 23613 18383 23616
rect 18325 23607 18383 23613
rect 19426 23604 19432 23616
rect 19484 23604 19490 23656
rect 18156 23548 19196 23576
rect 2038 23508 2044 23520
rect 1999 23480 2044 23508
rect 2038 23468 2044 23480
rect 2096 23468 2102 23520
rect 8202 23468 8208 23520
rect 8260 23508 8266 23520
rect 9217 23511 9275 23517
rect 9217 23508 9229 23511
rect 8260 23480 9229 23508
rect 8260 23468 8266 23480
rect 9217 23477 9229 23480
rect 9263 23477 9275 23511
rect 9217 23471 9275 23477
rect 13265 23511 13323 23517
rect 13265 23477 13277 23511
rect 13311 23508 13323 23511
rect 13538 23508 13544 23520
rect 13311 23480 13544 23508
rect 13311 23477 13323 23480
rect 13265 23471 13323 23477
rect 13538 23468 13544 23480
rect 13596 23468 13602 23520
rect 13722 23468 13728 23520
rect 13780 23508 13786 23520
rect 14001 23511 14059 23517
rect 14001 23508 14013 23511
rect 13780 23480 14013 23508
rect 13780 23468 13786 23480
rect 14001 23477 14013 23480
rect 14047 23477 14059 23511
rect 14734 23508 14740 23520
rect 14695 23480 14740 23508
rect 14001 23471 14059 23477
rect 14734 23468 14740 23480
rect 14792 23468 14798 23520
rect 16850 23468 16856 23520
rect 16908 23508 16914 23520
rect 17678 23508 17684 23520
rect 16908 23480 17684 23508
rect 16908 23468 16914 23480
rect 17678 23468 17684 23480
rect 17736 23468 17742 23520
rect 19168 23508 19196 23548
rect 20162 23536 20168 23588
rect 20220 23576 20226 23588
rect 23106 23576 23112 23588
rect 20220 23548 23112 23576
rect 20220 23536 20226 23548
rect 23106 23536 23112 23548
rect 23164 23536 23170 23588
rect 23216 23508 23244 23752
rect 23474 23740 23480 23752
rect 23532 23740 23538 23792
rect 25958 23740 25964 23792
rect 26016 23780 26022 23792
rect 28994 23780 29000 23792
rect 26016 23752 29000 23780
rect 26016 23740 26022 23752
rect 28994 23740 29000 23752
rect 29052 23740 29058 23792
rect 29089 23783 29147 23789
rect 29089 23749 29101 23783
rect 29135 23780 29147 23783
rect 31018 23780 31024 23792
rect 29135 23752 31024 23780
rect 29135 23749 29147 23752
rect 29089 23743 29147 23749
rect 31018 23740 31024 23752
rect 31076 23780 31082 23792
rect 31128 23780 31156 23811
rect 37458 23808 37464 23820
rect 37516 23808 37522 23860
rect 31076 23752 31156 23780
rect 31076 23740 31082 23752
rect 32398 23740 32404 23792
rect 32456 23780 32462 23792
rect 48038 23780 48044 23792
rect 32456 23752 48044 23780
rect 32456 23740 32462 23752
rect 48038 23740 48044 23752
rect 48096 23740 48102 23792
rect 23385 23715 23443 23721
rect 23385 23681 23397 23715
rect 23431 23712 23443 23715
rect 23431 23684 23612 23712
rect 23431 23681 23443 23684
rect 23385 23675 23443 23681
rect 23477 23647 23535 23653
rect 23477 23613 23489 23647
rect 23523 23613 23535 23647
rect 23584 23644 23612 23684
rect 23658 23672 23664 23724
rect 23716 23712 23722 23724
rect 24397 23715 24455 23721
rect 23716 23684 23761 23712
rect 23716 23672 23722 23684
rect 24397 23681 24409 23715
rect 24443 23712 24455 23715
rect 24673 23715 24731 23721
rect 24443 23684 24624 23712
rect 24443 23681 24455 23684
rect 24397 23675 24455 23681
rect 24412 23644 24440 23675
rect 23584 23616 24440 23644
rect 24489 23647 24547 23653
rect 23477 23607 23535 23613
rect 24489 23613 24501 23647
rect 24535 23613 24547 23647
rect 24596 23644 24624 23684
rect 24673 23681 24685 23715
rect 24719 23712 24731 23715
rect 24946 23712 24952 23724
rect 24719 23684 24952 23712
rect 24719 23681 24731 23684
rect 24673 23675 24731 23681
rect 24946 23672 24952 23684
rect 25004 23672 25010 23724
rect 25593 23715 25651 23721
rect 25593 23681 25605 23715
rect 25639 23712 25651 23715
rect 26694 23712 26700 23724
rect 25639 23684 26700 23712
rect 25639 23681 25651 23684
rect 25593 23675 25651 23681
rect 26694 23672 26700 23684
rect 26752 23672 26758 23724
rect 26786 23672 26792 23724
rect 26844 23712 26850 23724
rect 26973 23715 27031 23721
rect 26973 23712 26985 23715
rect 26844 23684 26985 23712
rect 26844 23672 26850 23684
rect 26973 23681 26985 23684
rect 27019 23681 27031 23715
rect 26973 23675 27031 23681
rect 27062 23672 27068 23724
rect 27120 23712 27126 23724
rect 27229 23715 27287 23721
rect 27229 23712 27241 23715
rect 27120 23684 27241 23712
rect 27120 23672 27126 23684
rect 27229 23681 27241 23684
rect 27275 23681 27287 23715
rect 27229 23675 27287 23681
rect 28442 23672 28448 23724
rect 28500 23712 28506 23724
rect 28905 23715 28963 23721
rect 28905 23712 28917 23715
rect 28500 23684 28917 23712
rect 28500 23672 28506 23684
rect 28905 23681 28917 23684
rect 28951 23681 28963 23715
rect 28905 23675 28963 23681
rect 29546 23672 29552 23724
rect 29604 23712 29610 23724
rect 29989 23715 30047 23721
rect 29989 23712 30001 23715
rect 29604 23684 30001 23712
rect 29604 23672 29610 23684
rect 29989 23681 30001 23684
rect 30035 23681 30047 23715
rect 37366 23712 37372 23724
rect 37327 23684 37372 23712
rect 29989 23675 30047 23681
rect 37366 23672 37372 23684
rect 37424 23672 37430 23724
rect 25130 23644 25136 23656
rect 24596 23616 25136 23644
rect 24489 23607 24547 23613
rect 23492 23576 23520 23607
rect 24504 23576 24532 23607
rect 25130 23604 25136 23616
rect 25188 23604 25194 23656
rect 25317 23647 25375 23653
rect 25317 23613 25329 23647
rect 25363 23613 25375 23647
rect 25317 23607 25375 23613
rect 25222 23576 25228 23588
rect 23492 23548 25228 23576
rect 25222 23536 25228 23548
rect 25280 23536 25286 23588
rect 23382 23508 23388 23520
rect 19168 23480 23244 23508
rect 23343 23480 23388 23508
rect 23382 23468 23388 23480
rect 23440 23468 23446 23520
rect 23474 23468 23480 23520
rect 23532 23508 23538 23520
rect 23845 23511 23903 23517
rect 23845 23508 23857 23511
rect 23532 23480 23857 23508
rect 23532 23468 23538 23480
rect 23845 23477 23857 23480
rect 23891 23477 23903 23511
rect 24670 23508 24676 23520
rect 24631 23480 24676 23508
rect 23845 23471 23903 23477
rect 24670 23468 24676 23480
rect 24728 23468 24734 23520
rect 24854 23508 24860 23520
rect 24815 23480 24860 23508
rect 24854 23468 24860 23480
rect 24912 23468 24918 23520
rect 25038 23468 25044 23520
rect 25096 23508 25102 23520
rect 25332 23508 25360 23607
rect 27982 23604 27988 23656
rect 28040 23644 28046 23656
rect 29086 23644 29092 23656
rect 28040 23616 29092 23644
rect 28040 23604 28046 23616
rect 29086 23604 29092 23616
rect 29144 23604 29150 23656
rect 29730 23644 29736 23656
rect 29691 23616 29736 23644
rect 29730 23604 29736 23616
rect 29788 23604 29794 23656
rect 33226 23644 33232 23656
rect 33187 23616 33232 23644
rect 33226 23604 33232 23616
rect 33284 23604 33290 23656
rect 33410 23644 33416 23656
rect 33371 23616 33416 23644
rect 33410 23604 33416 23616
rect 33468 23604 33474 23656
rect 35069 23647 35127 23653
rect 35069 23613 35081 23647
rect 35115 23644 35127 23647
rect 40034 23644 40040 23656
rect 35115 23616 40040 23644
rect 35115 23613 35127 23616
rect 35069 23607 35127 23613
rect 40034 23604 40040 23616
rect 40092 23604 40098 23656
rect 28626 23536 28632 23588
rect 28684 23576 28690 23588
rect 28684 23548 29776 23576
rect 28684 23536 28690 23548
rect 25096 23480 25360 23508
rect 25096 23468 25102 23480
rect 27890 23468 27896 23520
rect 27948 23508 27954 23520
rect 28353 23511 28411 23517
rect 28353 23508 28365 23511
rect 27948 23480 28365 23508
rect 27948 23468 27954 23480
rect 28353 23477 28365 23480
rect 28399 23477 28411 23511
rect 28353 23471 28411 23477
rect 29273 23511 29331 23517
rect 29273 23477 29285 23511
rect 29319 23508 29331 23511
rect 29638 23508 29644 23520
rect 29319 23480 29644 23508
rect 29319 23477 29331 23480
rect 29273 23471 29331 23477
rect 29638 23468 29644 23480
rect 29696 23468 29702 23520
rect 29748 23508 29776 23548
rect 47670 23508 47676 23520
rect 29748 23480 47676 23508
rect 47670 23468 47676 23480
rect 47728 23468 47734 23520
rect 1104 23418 48852 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 48852 23418
rect 1104 23344 48852 23366
rect 23014 23304 23020 23316
rect 2746 23276 23020 23304
rect 1578 23196 1584 23248
rect 1636 23236 1642 23248
rect 2746 23236 2774 23276
rect 23014 23264 23020 23276
rect 23072 23264 23078 23316
rect 23106 23264 23112 23316
rect 23164 23304 23170 23316
rect 23164 23276 23520 23304
rect 23164 23264 23170 23276
rect 8938 23236 8944 23248
rect 1636 23208 2774 23236
rect 8899 23208 8944 23236
rect 1636 23196 1642 23208
rect 8938 23196 8944 23208
rect 8996 23196 9002 23248
rect 9306 23196 9312 23248
rect 9364 23196 9370 23248
rect 12066 23196 12072 23248
rect 12124 23236 12130 23248
rect 12124 23208 13124 23236
rect 12124 23196 12130 23208
rect 1397 23171 1455 23177
rect 1397 23137 1409 23171
rect 1443 23168 1455 23171
rect 2038 23168 2044 23180
rect 1443 23140 2044 23168
rect 1443 23137 1455 23140
rect 1397 23131 1455 23137
rect 2038 23128 2044 23140
rect 2096 23128 2102 23180
rect 2774 23128 2780 23180
rect 2832 23168 2838 23180
rect 9324 23168 9352 23196
rect 13096 23177 13124 23208
rect 15102 23196 15108 23248
rect 15160 23236 15166 23248
rect 15473 23239 15531 23245
rect 15473 23236 15485 23239
rect 15160 23208 15485 23236
rect 15160 23196 15166 23208
rect 15473 23205 15485 23208
rect 15519 23205 15531 23239
rect 15473 23199 15531 23205
rect 16942 23196 16948 23248
rect 17000 23236 17006 23248
rect 17313 23239 17371 23245
rect 17313 23236 17325 23239
rect 17000 23208 17325 23236
rect 17000 23196 17006 23208
rect 17313 23205 17325 23208
rect 17359 23205 17371 23239
rect 17313 23199 17371 23205
rect 19978 23196 19984 23248
rect 20036 23236 20042 23248
rect 20254 23236 20260 23248
rect 20036 23208 20260 23236
rect 20036 23196 20042 23208
rect 20254 23196 20260 23208
rect 20312 23196 20318 23248
rect 22186 23236 22192 23248
rect 22099 23208 22192 23236
rect 22186 23196 22192 23208
rect 22244 23236 22250 23248
rect 23198 23236 23204 23248
rect 22244 23208 23204 23236
rect 22244 23196 22250 23208
rect 23198 23196 23204 23208
rect 23256 23196 23262 23248
rect 23492 23236 23520 23276
rect 23566 23264 23572 23316
rect 23624 23304 23630 23316
rect 23753 23307 23811 23313
rect 23753 23304 23765 23307
rect 23624 23276 23765 23304
rect 23624 23264 23630 23276
rect 23753 23273 23765 23276
rect 23799 23304 23811 23307
rect 25038 23304 25044 23316
rect 23799 23276 25044 23304
rect 23799 23273 23811 23276
rect 23753 23267 23811 23273
rect 25038 23264 25044 23276
rect 25096 23264 25102 23316
rect 26234 23264 26240 23316
rect 26292 23304 26298 23316
rect 27525 23307 27583 23313
rect 27525 23304 27537 23307
rect 26292 23276 27537 23304
rect 26292 23264 26298 23276
rect 27525 23273 27537 23276
rect 27571 23273 27583 23307
rect 27525 23267 27583 23273
rect 27706 23264 27712 23316
rect 27764 23304 27770 23316
rect 28258 23304 28264 23316
rect 27764 23276 28264 23304
rect 27764 23264 27770 23276
rect 28258 23264 28264 23276
rect 28316 23264 28322 23316
rect 29546 23304 29552 23316
rect 29507 23276 29552 23304
rect 29546 23264 29552 23276
rect 29604 23264 29610 23316
rect 29730 23264 29736 23316
rect 29788 23304 29794 23316
rect 32122 23304 32128 23316
rect 29788 23276 32128 23304
rect 29788 23264 29794 23276
rect 32122 23264 32128 23276
rect 32180 23264 32186 23316
rect 33229 23307 33287 23313
rect 33229 23273 33241 23307
rect 33275 23304 33287 23307
rect 33410 23304 33416 23316
rect 33275 23276 33416 23304
rect 33275 23273 33287 23276
rect 33229 23267 33287 23273
rect 33410 23264 33416 23276
rect 33468 23264 33474 23316
rect 47854 23304 47860 23316
rect 47815 23276 47860 23304
rect 47854 23264 47860 23276
rect 47912 23264 47918 23316
rect 24762 23236 24768 23248
rect 23492 23208 24768 23236
rect 24762 23196 24768 23208
rect 24820 23236 24826 23248
rect 24820 23208 25820 23236
rect 24820 23196 24826 23208
rect 2832 23140 2877 23168
rect 9321 23140 9352 23168
rect 13081 23171 13139 23177
rect 2832 23128 2838 23140
rect 8202 23100 8208 23112
rect 8163 23072 8208 23100
rect 8202 23060 8208 23072
rect 8260 23060 8266 23112
rect 8846 23060 8852 23112
rect 8904 23100 8910 23112
rect 9217 23103 9275 23109
rect 8904 23097 9168 23100
rect 9217 23097 9229 23103
rect 8904 23072 9229 23097
rect 8904 23060 8910 23072
rect 9140 23069 9229 23072
rect 9263 23069 9275 23103
rect 9321 23106 9349 23140
rect 13081 23137 13093 23171
rect 13127 23137 13139 23171
rect 19150 23168 19156 23180
rect 13081 23131 13139 23137
rect 18156 23140 19156 23168
rect 9321 23100 9380 23106
rect 9597 23103 9655 23109
rect 9321 23069 9334 23100
rect 9217 23063 9275 23069
rect 9322 23066 9334 23069
rect 9368 23066 9380 23100
rect 9322 23060 9380 23066
rect 9422 23097 9480 23103
rect 9422 23063 9434 23097
rect 9468 23094 9480 23097
rect 9468 23066 9536 23094
rect 9468 23063 9480 23066
rect 9422 23057 9480 23063
rect 1581 23035 1639 23041
rect 1581 23001 1593 23035
rect 1627 23032 1639 23035
rect 2314 23032 2320 23044
rect 1627 23004 2320 23032
rect 1627 23001 1639 23004
rect 1581 22995 1639 23001
rect 2314 22992 2320 23004
rect 2372 22992 2378 23044
rect 8018 23032 8024 23044
rect 7979 23004 8024 23032
rect 8018 22992 8024 23004
rect 8076 22992 8082 23044
rect 8386 23032 8392 23044
rect 8347 23004 8392 23032
rect 8386 22992 8392 23004
rect 8444 22992 8450 23044
rect 9508 23032 9536 23066
rect 9597 23069 9609 23103
rect 9643 23100 9655 23103
rect 9766 23100 9772 23112
rect 9643 23072 9772 23100
rect 9643 23069 9655 23072
rect 9597 23063 9655 23069
rect 9766 23060 9772 23072
rect 9824 23060 9830 23112
rect 11790 23060 11796 23112
rect 11848 23109 11854 23112
rect 11848 23103 11897 23109
rect 11848 23069 11851 23103
rect 11885 23069 11897 23103
rect 11974 23100 11980 23112
rect 11935 23072 11980 23100
rect 11848 23063 11897 23069
rect 11848 23060 11854 23063
rect 11974 23060 11980 23072
rect 12032 23060 12038 23112
rect 12066 23060 12072 23112
rect 12124 23100 12130 23112
rect 12253 23103 12311 23109
rect 12124 23072 12169 23100
rect 12124 23060 12130 23072
rect 12253 23069 12265 23103
rect 12299 23100 12311 23103
rect 12342 23100 12348 23112
rect 12299 23072 12348 23100
rect 12299 23069 12311 23072
rect 12253 23063 12311 23069
rect 12342 23060 12348 23072
rect 12400 23060 12406 23112
rect 12713 23103 12771 23109
rect 12713 23069 12725 23103
rect 12759 23100 12771 23103
rect 13446 23100 13452 23112
rect 12759 23072 13452 23100
rect 12759 23069 12771 23072
rect 12713 23063 12771 23069
rect 13446 23060 13452 23072
rect 13504 23060 13510 23112
rect 14093 23103 14151 23109
rect 14093 23069 14105 23103
rect 14139 23100 14151 23103
rect 15933 23103 15991 23109
rect 15933 23100 15945 23103
rect 14139 23072 15945 23100
rect 14139 23069 14151 23072
rect 14093 23063 14151 23069
rect 15933 23069 15945 23072
rect 15979 23100 15991 23103
rect 17034 23100 17040 23112
rect 15979 23072 17040 23100
rect 15979 23069 15991 23072
rect 15933 23063 15991 23069
rect 17034 23060 17040 23072
rect 17092 23060 17098 23112
rect 18156 23109 18184 23140
rect 19150 23128 19156 23140
rect 19208 23168 19214 23180
rect 19208 23140 19334 23168
rect 19208 23128 19214 23140
rect 18049 23103 18107 23109
rect 18049 23100 18061 23103
rect 17144 23072 18061 23100
rect 9858 23032 9864 23044
rect 9508 23004 9864 23032
rect 9858 22992 9864 23004
rect 9916 22992 9922 23044
rect 12894 23032 12900 23044
rect 10060 23004 11744 23032
rect 12855 23004 12900 23032
rect 4614 22924 4620 22976
rect 4672 22964 4678 22976
rect 10060 22964 10088 23004
rect 11606 22964 11612 22976
rect 4672 22936 10088 22964
rect 11567 22936 11612 22964
rect 4672 22924 4678 22936
rect 11606 22924 11612 22936
rect 11664 22924 11670 22976
rect 11716 22964 11744 23004
rect 12894 22992 12900 23004
rect 12952 22992 12958 23044
rect 14182 22992 14188 23044
rect 14240 23032 14246 23044
rect 14338 23035 14396 23041
rect 14338 23032 14350 23035
rect 14240 23004 14350 23032
rect 14240 22992 14246 23004
rect 14338 23001 14350 23004
rect 14384 23001 14396 23035
rect 14338 22995 14396 23001
rect 15562 22992 15568 23044
rect 15620 23032 15626 23044
rect 16178 23035 16236 23041
rect 16178 23032 16190 23035
rect 15620 23004 16190 23032
rect 15620 22992 15626 23004
rect 16178 23001 16190 23004
rect 16224 23001 16236 23035
rect 16178 22995 16236 23001
rect 17144 22964 17172 23072
rect 18049 23069 18061 23072
rect 18095 23069 18107 23103
rect 18049 23063 18107 23069
rect 18141 23103 18199 23109
rect 18141 23069 18153 23103
rect 18187 23069 18199 23103
rect 18141 23063 18199 23069
rect 18230 23060 18236 23112
rect 18288 23100 18294 23112
rect 18417 23103 18475 23109
rect 18288 23072 18333 23100
rect 18288 23060 18294 23072
rect 18417 23069 18429 23103
rect 18463 23100 18475 23103
rect 18690 23100 18696 23112
rect 18463 23072 18696 23100
rect 18463 23069 18475 23072
rect 18417 23063 18475 23069
rect 17954 22992 17960 23044
rect 18012 23032 18018 23044
rect 18432 23032 18460 23063
rect 18690 23060 18696 23072
rect 18748 23060 18754 23112
rect 18012 23004 18460 23032
rect 19306 23032 19334 23140
rect 19886 23128 19892 23180
rect 19944 23168 19950 23180
rect 20809 23171 20867 23177
rect 20809 23168 20821 23171
rect 19944 23140 20821 23168
rect 19944 23128 19950 23140
rect 20809 23137 20821 23140
rect 20855 23137 20867 23171
rect 20809 23131 20867 23137
rect 19426 23100 19432 23112
rect 19484 23109 19490 23112
rect 19395 23072 19432 23100
rect 19426 23060 19432 23072
rect 19484 23063 19495 23109
rect 19484 23060 19490 23063
rect 20162 23060 20168 23112
rect 20220 23100 20226 23112
rect 20898 23100 20904 23112
rect 20220 23072 20904 23100
rect 20220 23060 20226 23072
rect 20898 23060 20904 23072
rect 20956 23060 20962 23112
rect 21076 23103 21134 23109
rect 21076 23069 21088 23103
rect 21122 23100 21134 23103
rect 21818 23100 21824 23112
rect 21122 23072 21824 23100
rect 21122 23069 21134 23072
rect 21076 23063 21134 23069
rect 21818 23060 21824 23072
rect 21876 23060 21882 23112
rect 22741 23103 22799 23109
rect 22741 23069 22753 23103
rect 22787 23100 22799 23103
rect 23474 23100 23480 23112
rect 22787 23072 23480 23100
rect 22787 23069 22799 23072
rect 22741 23063 22799 23069
rect 23474 23060 23480 23072
rect 23532 23060 23538 23112
rect 24673 23103 24731 23109
rect 24673 23069 24685 23103
rect 24719 23100 24731 23103
rect 24854 23100 24860 23112
rect 24719 23072 24860 23100
rect 24719 23069 24731 23072
rect 24673 23063 24731 23069
rect 24854 23060 24860 23072
rect 24912 23060 24918 23112
rect 25593 23103 25651 23109
rect 25593 23069 25605 23103
rect 25639 23100 25651 23103
rect 25792 23100 25820 23208
rect 26418 23196 26424 23248
rect 26476 23236 26482 23248
rect 27982 23236 27988 23248
rect 26476 23208 27988 23236
rect 26476 23196 26482 23208
rect 27982 23196 27988 23208
rect 28040 23196 28046 23248
rect 48222 23236 48228 23248
rect 29820 23208 48228 23236
rect 25869 23171 25927 23177
rect 25869 23137 25881 23171
rect 25915 23168 25927 23171
rect 26326 23168 26332 23180
rect 25915 23140 26332 23168
rect 25915 23137 25927 23140
rect 25869 23131 25927 23137
rect 26326 23128 26332 23140
rect 26384 23128 26390 23180
rect 25639 23072 25820 23100
rect 27341 23103 27399 23109
rect 25639 23069 25651 23072
rect 25593 23063 25651 23069
rect 27341 23069 27353 23103
rect 27387 23100 27399 23103
rect 28166 23100 28172 23112
rect 27387 23072 28172 23100
rect 27387 23069 27399 23072
rect 27341 23063 27399 23069
rect 28166 23060 28172 23072
rect 28224 23060 28230 23112
rect 28626 23109 28632 23112
rect 28583 23103 28632 23109
rect 28583 23069 28595 23103
rect 28629 23069 28632 23103
rect 28583 23063 28632 23069
rect 28626 23060 28632 23063
rect 28684 23060 28690 23112
rect 28721 23103 28779 23109
rect 28721 23069 28733 23103
rect 28767 23069 28779 23103
rect 28721 23063 28779 23069
rect 24949 23035 25007 23041
rect 19306 23004 22876 23032
rect 18012 22992 18018 23004
rect 17770 22964 17776 22976
rect 11716 22936 17172 22964
rect 17731 22936 17776 22964
rect 17770 22924 17776 22936
rect 17828 22924 17834 22976
rect 19242 22964 19248 22976
rect 19203 22936 19248 22964
rect 19242 22924 19248 22936
rect 19300 22924 19306 22976
rect 20070 22924 20076 22976
rect 20128 22964 20134 22976
rect 20438 22964 20444 22976
rect 20128 22936 20444 22964
rect 20128 22924 20134 22936
rect 20438 22924 20444 22936
rect 20496 22924 20502 22976
rect 22848 22973 22876 23004
rect 24949 23001 24961 23035
rect 24995 23032 25007 23035
rect 25682 23032 25688 23044
rect 24995 23004 25688 23032
rect 24995 23001 25007 23004
rect 24949 22995 25007 23001
rect 25682 22992 25688 23004
rect 25740 22992 25746 23044
rect 26970 22992 26976 23044
rect 27028 23032 27034 23044
rect 27157 23035 27215 23041
rect 27157 23032 27169 23035
rect 27028 23004 27169 23032
rect 27028 22992 27034 23004
rect 27157 23001 27169 23004
rect 27203 23001 27215 23035
rect 28736 23032 28764 23063
rect 28810 23060 28816 23112
rect 28868 23097 28874 23112
rect 28868 23069 28910 23097
rect 28868 23060 28874 23069
rect 28994 23060 29000 23112
rect 29052 23100 29058 23112
rect 29820 23109 29848 23208
rect 48222 23196 48228 23208
rect 48280 23196 48286 23248
rect 45738 23128 45744 23180
rect 45796 23168 45802 23180
rect 47397 23171 47455 23177
rect 47397 23168 47409 23171
rect 45796 23140 47409 23168
rect 45796 23128 45802 23140
rect 47397 23137 47409 23140
rect 47443 23137 47455 23171
rect 47397 23131 47455 23137
rect 29805 23103 29863 23109
rect 29052 23072 29097 23100
rect 29052 23060 29058 23072
rect 29805 23069 29817 23103
rect 29851 23069 29863 23103
rect 29805 23063 29863 23069
rect 29917 23103 29975 23109
rect 29917 23069 29929 23103
rect 29963 23069 29975 23103
rect 29917 23063 29975 23069
rect 30009 23103 30067 23109
rect 30009 23069 30021 23103
rect 30055 23069 30067 23103
rect 30009 23063 30067 23069
rect 29454 23032 29460 23044
rect 28736 23004 29460 23032
rect 27157 22995 27215 23001
rect 29454 22992 29460 23004
rect 29512 23032 29518 23044
rect 29932 23032 29960 23063
rect 29512 23004 29960 23032
rect 29512 22992 29518 23004
rect 22833 22967 22891 22973
rect 22833 22933 22845 22967
rect 22879 22933 22891 22967
rect 22833 22927 22891 22933
rect 28353 22967 28411 22973
rect 28353 22933 28365 22967
rect 28399 22964 28411 22967
rect 29362 22964 29368 22976
rect 28399 22936 29368 22964
rect 28399 22933 28411 22936
rect 28353 22927 28411 22933
rect 29362 22924 29368 22936
rect 29420 22924 29426 22976
rect 29638 22924 29644 22976
rect 29696 22964 29702 22976
rect 30024 22964 30052 23063
rect 30190 23060 30196 23112
rect 30248 23100 30254 23112
rect 33134 23100 33140 23112
rect 30248 23072 30293 23100
rect 33095 23072 33140 23100
rect 30248 23060 30254 23072
rect 33134 23060 33140 23072
rect 33192 23060 33198 23112
rect 47486 23060 47492 23112
rect 47544 23100 47550 23112
rect 47857 23103 47915 23109
rect 47544 23072 47589 23100
rect 47544 23060 47550 23072
rect 47857 23069 47869 23103
rect 47903 23069 47915 23103
rect 47857 23063 47915 23069
rect 46658 22992 46664 23044
rect 46716 23032 46722 23044
rect 47872 23032 47900 23063
rect 46716 23004 47900 23032
rect 46716 22992 46722 23004
rect 48038 22964 48044 22976
rect 29696 22936 30052 22964
rect 47999 22936 48044 22964
rect 29696 22924 29702 22936
rect 48038 22924 48044 22936
rect 48096 22924 48102 22976
rect 1104 22874 48852 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 48852 22874
rect 1104 22800 48852 22822
rect 1578 22760 1584 22772
rect 1539 22732 1584 22760
rect 1578 22720 1584 22732
rect 1636 22720 1642 22772
rect 2314 22760 2320 22772
rect 2275 22732 2320 22760
rect 2314 22720 2320 22732
rect 2372 22720 2378 22772
rect 8018 22720 8024 22772
rect 8076 22760 8082 22772
rect 8076 22732 9076 22760
rect 8076 22720 8082 22732
rect 8294 22692 8300 22704
rect 7208 22664 8300 22692
rect 1394 22624 1400 22636
rect 1355 22596 1400 22624
rect 1394 22584 1400 22596
rect 1452 22584 1458 22636
rect 2130 22584 2136 22636
rect 2188 22624 2194 22636
rect 7208 22633 7236 22664
rect 8294 22652 8300 22664
rect 8352 22692 8358 22704
rect 8938 22692 8944 22704
rect 8352 22664 8944 22692
rect 8352 22652 8358 22664
rect 8938 22652 8944 22664
rect 8996 22652 9002 22704
rect 9048 22701 9076 22732
rect 11974 22720 11980 22772
rect 12032 22760 12038 22772
rect 14182 22760 14188 22772
rect 12032 22732 14044 22760
rect 14143 22732 14188 22760
rect 12032 22720 12038 22732
rect 9033 22695 9091 22701
rect 9033 22661 9045 22695
rect 9079 22692 9091 22695
rect 9079 22664 10364 22692
rect 9079 22661 9091 22664
rect 9033 22655 9091 22661
rect 2225 22627 2283 22633
rect 2225 22624 2237 22627
rect 2188 22596 2237 22624
rect 2188 22584 2194 22596
rect 2225 22593 2237 22596
rect 2271 22593 2283 22627
rect 2225 22587 2283 22593
rect 7193 22627 7251 22633
rect 7193 22593 7205 22627
rect 7239 22593 7251 22627
rect 7193 22587 7251 22593
rect 7460 22627 7518 22633
rect 7460 22593 7472 22627
rect 7506 22624 7518 22627
rect 8846 22624 8852 22636
rect 7506 22596 8852 22624
rect 7506 22593 7518 22596
rect 7460 22587 7518 22593
rect 8846 22584 8852 22596
rect 8904 22584 8910 22636
rect 9217 22627 9275 22633
rect 9217 22593 9229 22627
rect 9263 22593 9275 22627
rect 9217 22587 9275 22593
rect 9232 22556 9260 22587
rect 10336 22565 10364 22664
rect 11606 22652 11612 22704
rect 11664 22692 11670 22704
rect 11762 22695 11820 22701
rect 11762 22692 11774 22695
rect 11664 22664 11774 22692
rect 11664 22652 11670 22664
rect 11762 22661 11774 22664
rect 11808 22661 11820 22695
rect 11762 22655 11820 22661
rect 13541 22695 13599 22701
rect 13541 22661 13553 22695
rect 13587 22692 13599 22695
rect 13722 22692 13728 22704
rect 13587 22664 13728 22692
rect 13587 22661 13599 22664
rect 13541 22655 13599 22661
rect 13722 22652 13728 22664
rect 13780 22652 13786 22704
rect 14016 22692 14044 22732
rect 14182 22720 14188 22732
rect 14240 22720 14246 22772
rect 14458 22720 14464 22772
rect 14516 22760 14522 22772
rect 15473 22763 15531 22769
rect 14516 22732 15424 22760
rect 14516 22720 14522 22732
rect 14274 22692 14280 22704
rect 14016 22664 14280 22692
rect 14274 22652 14280 22664
rect 14332 22692 14338 22704
rect 15396 22692 15424 22732
rect 15473 22729 15485 22763
rect 15519 22760 15531 22763
rect 15562 22760 15568 22772
rect 15519 22732 15568 22760
rect 15519 22729 15531 22732
rect 15473 22723 15531 22729
rect 15562 22720 15568 22732
rect 15620 22720 15626 22772
rect 15746 22720 15752 22772
rect 15804 22760 15810 22772
rect 16206 22760 16212 22772
rect 15804 22732 16212 22760
rect 15804 22720 15810 22732
rect 16206 22720 16212 22732
rect 16264 22720 16270 22772
rect 27341 22763 27399 22769
rect 16316 22732 26924 22760
rect 16316 22692 16344 22732
rect 14332 22664 15148 22692
rect 15396 22664 16344 22692
rect 17512 22664 21864 22692
rect 14332 22652 14338 22664
rect 11514 22624 11520 22636
rect 11475 22596 11520 22624
rect 11514 22584 11520 22596
rect 11572 22584 11578 22636
rect 13357 22627 13415 22633
rect 13357 22593 13369 22627
rect 13403 22624 13415 22627
rect 13446 22624 13452 22636
rect 13403 22596 13452 22624
rect 13403 22593 13415 22596
rect 13357 22587 13415 22593
rect 13446 22584 13452 22596
rect 13504 22584 13510 22636
rect 14458 22624 14464 22636
rect 14419 22596 14464 22624
rect 14458 22584 14464 22596
rect 14516 22584 14522 22636
rect 14568 22633 14596 22664
rect 14553 22627 14611 22633
rect 14553 22593 14565 22627
rect 14599 22593 14611 22627
rect 14553 22587 14611 22593
rect 14645 22627 14703 22633
rect 14645 22593 14657 22627
rect 14691 22624 14703 22627
rect 14829 22627 14887 22633
rect 14691 22596 14780 22624
rect 14691 22593 14703 22596
rect 14645 22587 14703 22593
rect 8588 22528 9260 22556
rect 10045 22559 10103 22565
rect 8202 22380 8208 22432
rect 8260 22420 8266 22432
rect 8588 22429 8616 22528
rect 10045 22525 10057 22559
rect 10091 22525 10103 22559
rect 10045 22519 10103 22525
rect 10321 22559 10379 22565
rect 10321 22525 10333 22559
rect 10367 22556 10379 22559
rect 10778 22556 10784 22568
rect 10367 22528 10784 22556
rect 10367 22525 10379 22528
rect 10321 22519 10379 22525
rect 8573 22423 8631 22429
rect 8573 22420 8585 22423
rect 8260 22392 8585 22420
rect 8260 22380 8266 22392
rect 8573 22389 8585 22392
rect 8619 22389 8631 22423
rect 9398 22420 9404 22432
rect 9359 22392 9404 22420
rect 8573 22383 8631 22389
rect 9398 22380 9404 22392
rect 9456 22380 9462 22432
rect 10060 22420 10088 22519
rect 10778 22516 10784 22528
rect 10836 22516 10842 22568
rect 13725 22559 13783 22565
rect 13725 22525 13737 22559
rect 13771 22556 13783 22559
rect 14752 22556 14780 22596
rect 14829 22593 14841 22627
rect 14875 22624 14955 22627
rect 15010 22624 15016 22636
rect 14875 22599 15016 22624
rect 14875 22593 14887 22599
rect 14927 22596 15016 22599
rect 14829 22587 14887 22593
rect 15010 22584 15016 22596
rect 15068 22584 15074 22636
rect 13771 22528 14780 22556
rect 15120 22556 15148 22664
rect 15197 22627 15255 22633
rect 15197 22593 15209 22627
rect 15243 22624 15255 22627
rect 15746 22624 15752 22636
rect 15243 22596 15752 22624
rect 15243 22593 15255 22596
rect 15197 22587 15255 22593
rect 15746 22584 15752 22596
rect 15804 22584 15810 22636
rect 15841 22627 15899 22633
rect 15841 22593 15853 22627
rect 15887 22593 15899 22627
rect 15841 22587 15899 22593
rect 15856 22556 15884 22587
rect 15930 22584 15936 22636
rect 15988 22624 15994 22636
rect 16117 22627 16175 22633
rect 15988 22596 16033 22624
rect 15988 22584 15994 22596
rect 16117 22593 16129 22627
rect 16163 22624 16175 22627
rect 16206 22624 16212 22636
rect 16163 22596 16212 22624
rect 16163 22593 16175 22596
rect 16117 22587 16175 22593
rect 16206 22584 16212 22596
rect 16264 22584 16270 22636
rect 16853 22627 16911 22633
rect 16853 22593 16865 22627
rect 16899 22593 16911 22627
rect 16853 22587 16911 22593
rect 15120 22528 15884 22556
rect 16868 22556 16896 22587
rect 17034 22584 17040 22636
rect 17092 22624 17098 22636
rect 17512 22633 17540 22664
rect 17770 22633 17776 22636
rect 17497 22627 17555 22633
rect 17497 22624 17509 22627
rect 17092 22596 17509 22624
rect 17092 22584 17098 22596
rect 17497 22593 17509 22596
rect 17543 22593 17555 22627
rect 17764 22624 17776 22633
rect 17731 22596 17776 22624
rect 17497 22587 17555 22593
rect 17764 22587 17776 22596
rect 17770 22584 17776 22587
rect 17828 22584 17834 22636
rect 19352 22633 19380 22664
rect 19337 22627 19395 22633
rect 19337 22593 19349 22627
rect 19383 22593 19395 22627
rect 19337 22587 19395 22593
rect 19426 22584 19432 22636
rect 19484 22624 19490 22636
rect 21836 22633 21864 22664
rect 21910 22652 21916 22704
rect 21968 22692 21974 22704
rect 22066 22695 22124 22701
rect 22066 22692 22078 22695
rect 21968 22664 22078 22692
rect 21968 22652 21974 22664
rect 22066 22661 22078 22664
rect 22112 22661 22124 22695
rect 26418 22692 26424 22704
rect 22066 22655 22124 22661
rect 24320 22664 26424 22692
rect 19593 22627 19651 22633
rect 19593 22624 19605 22627
rect 19484 22596 19605 22624
rect 19484 22584 19490 22596
rect 19593 22593 19605 22596
rect 19639 22593 19651 22627
rect 19593 22587 19651 22593
rect 21821 22627 21879 22633
rect 21821 22593 21833 22627
rect 21867 22593 21879 22627
rect 23474 22624 23480 22636
rect 21821 22587 21879 22593
rect 21928 22596 23480 22624
rect 21928 22556 21956 22596
rect 23474 22584 23480 22596
rect 23532 22584 23538 22636
rect 24118 22624 24124 22636
rect 24079 22596 24124 22624
rect 24118 22584 24124 22596
rect 24176 22584 24182 22636
rect 24320 22633 24348 22664
rect 26418 22652 26424 22664
rect 26476 22652 26482 22704
rect 26896 22692 26924 22732
rect 27341 22729 27353 22763
rect 27387 22760 27399 22763
rect 27430 22760 27436 22772
rect 27387 22732 27436 22760
rect 27387 22729 27399 22732
rect 27341 22723 27399 22729
rect 27430 22720 27436 22732
rect 27488 22720 27494 22772
rect 28810 22760 28816 22772
rect 28771 22732 28816 22760
rect 28810 22720 28816 22732
rect 28868 22720 28874 22772
rect 41874 22760 41880 22772
rect 28920 22732 41880 22760
rect 28920 22692 28948 22732
rect 41874 22720 41880 22732
rect 41932 22720 41938 22772
rect 47486 22720 47492 22772
rect 47544 22760 47550 22772
rect 47949 22763 48007 22769
rect 47949 22760 47961 22763
rect 47544 22732 47961 22760
rect 47544 22720 47550 22732
rect 47949 22729 47961 22732
rect 47995 22729 48007 22763
rect 47949 22723 48007 22729
rect 29730 22692 29736 22704
rect 26896 22664 28948 22692
rect 29288 22664 29736 22692
rect 24305 22627 24363 22633
rect 24305 22593 24317 22627
rect 24351 22593 24363 22627
rect 24305 22587 24363 22593
rect 24397 22627 24455 22633
rect 24397 22593 24409 22627
rect 24443 22593 24455 22627
rect 25038 22624 25044 22636
rect 24999 22596 25044 22624
rect 24397 22587 24455 22593
rect 16868 22528 17080 22556
rect 13771 22525 13783 22528
rect 13725 22519 13783 22525
rect 15856 22488 15884 22528
rect 15856 22460 16988 22488
rect 12710 22420 12716 22432
rect 10060 22392 12716 22420
rect 12710 22380 12716 22392
rect 12768 22380 12774 22432
rect 12894 22420 12900 22432
rect 12855 22392 12900 22420
rect 12894 22380 12900 22392
rect 12952 22380 12958 22432
rect 16960 22429 16988 22460
rect 16945 22423 17003 22429
rect 16945 22389 16957 22423
rect 16991 22389 17003 22423
rect 17052 22420 17080 22528
rect 20364 22528 21956 22556
rect 18432 22460 19012 22488
rect 17862 22420 17868 22432
rect 17052 22392 17868 22420
rect 16945 22383 17003 22389
rect 17862 22380 17868 22392
rect 17920 22420 17926 22432
rect 18432 22420 18460 22460
rect 18874 22420 18880 22432
rect 17920 22392 18460 22420
rect 18835 22392 18880 22420
rect 17920 22380 17926 22392
rect 18874 22380 18880 22392
rect 18932 22380 18938 22432
rect 18984 22420 19012 22460
rect 20364 22420 20392 22528
rect 23566 22448 23572 22500
rect 23624 22488 23630 22500
rect 24412 22488 24440 22587
rect 25038 22584 25044 22596
rect 25096 22584 25102 22636
rect 25317 22627 25375 22633
rect 25317 22624 25329 22627
rect 25148 22596 25329 22624
rect 25148 22556 25176 22596
rect 25317 22593 25329 22596
rect 25363 22593 25375 22627
rect 26142 22624 26148 22636
rect 26103 22596 26148 22624
rect 25317 22587 25375 22593
rect 26142 22584 26148 22596
rect 26200 22584 26206 22636
rect 26970 22624 26976 22636
rect 26883 22596 26976 22624
rect 26970 22584 26976 22596
rect 27028 22584 27034 22636
rect 27157 22627 27215 22633
rect 27157 22593 27169 22627
rect 27203 22624 27215 22627
rect 27798 22624 27804 22636
rect 27203 22596 27804 22624
rect 27203 22593 27215 22596
rect 27157 22587 27215 22593
rect 27798 22584 27804 22596
rect 27856 22584 27862 22636
rect 28442 22584 28448 22636
rect 28500 22624 28506 22636
rect 29288 22633 29316 22664
rect 29730 22652 29736 22664
rect 29788 22652 29794 22704
rect 30374 22652 30380 22704
rect 30432 22692 30438 22704
rect 32370 22695 32428 22701
rect 32370 22692 32382 22695
rect 30432 22664 32382 22692
rect 30432 22652 30438 22664
rect 32370 22661 32382 22664
rect 32416 22661 32428 22695
rect 32370 22655 32428 22661
rect 28629 22627 28687 22633
rect 28500 22596 28593 22624
rect 28500 22584 28506 22596
rect 28629 22593 28641 22627
rect 28675 22593 28687 22627
rect 28629 22587 28687 22593
rect 29273 22627 29331 22633
rect 29273 22593 29285 22627
rect 29319 22593 29331 22627
rect 29273 22587 29331 22593
rect 24596 22528 25176 22556
rect 25225 22559 25283 22565
rect 24596 22497 24624 22528
rect 25225 22525 25237 22559
rect 25271 22556 25283 22559
rect 25498 22556 25504 22568
rect 25271 22528 25504 22556
rect 25271 22525 25283 22528
rect 25225 22519 25283 22525
rect 25498 22516 25504 22528
rect 25556 22516 25562 22568
rect 26988 22556 27016 22584
rect 28460 22556 28488 22584
rect 25976 22528 28488 22556
rect 23624 22460 24440 22488
rect 24581 22491 24639 22497
rect 23624 22448 23630 22460
rect 24581 22457 24593 22491
rect 24627 22457 24639 22491
rect 24581 22451 24639 22457
rect 24670 22448 24676 22500
rect 24728 22488 24734 22500
rect 25976 22497 26004 22528
rect 25961 22491 26019 22497
rect 24728 22460 25544 22488
rect 24728 22448 24734 22460
rect 20714 22420 20720 22432
rect 18984 22392 20392 22420
rect 20675 22392 20720 22420
rect 20714 22380 20720 22392
rect 20772 22380 20778 22432
rect 22186 22380 22192 22432
rect 22244 22420 22250 22432
rect 23201 22423 23259 22429
rect 23201 22420 23213 22423
rect 22244 22392 23213 22420
rect 22244 22380 22250 22392
rect 23201 22389 23213 22392
rect 23247 22389 23259 22423
rect 24210 22420 24216 22432
rect 24171 22392 24216 22420
rect 23201 22383 23259 22389
rect 24210 22380 24216 22392
rect 24268 22380 24274 22432
rect 25314 22420 25320 22432
rect 25275 22392 25320 22420
rect 25314 22380 25320 22392
rect 25372 22380 25378 22432
rect 25516 22429 25544 22460
rect 25961 22457 25973 22491
rect 26007 22457 26019 22491
rect 25961 22451 26019 22457
rect 25501 22423 25559 22429
rect 25501 22389 25513 22423
rect 25547 22389 25559 22423
rect 25501 22383 25559 22389
rect 28074 22380 28080 22432
rect 28132 22420 28138 22432
rect 28644 22420 28672 22587
rect 29362 22584 29368 22636
rect 29420 22624 29426 22636
rect 29529 22627 29587 22633
rect 29529 22624 29541 22627
rect 29420 22596 29541 22624
rect 29420 22584 29426 22596
rect 29529 22593 29541 22596
rect 29575 22593 29587 22627
rect 32122 22624 32128 22636
rect 32083 22596 32128 22624
rect 29529 22587 29587 22593
rect 32122 22584 32128 22596
rect 32180 22584 32186 22636
rect 48130 22624 48136 22636
rect 48091 22596 48136 22624
rect 48130 22584 48136 22596
rect 48188 22584 48194 22636
rect 33226 22448 33232 22500
rect 33284 22488 33290 22500
rect 33502 22488 33508 22500
rect 33284 22460 33508 22488
rect 33284 22448 33290 22460
rect 33502 22448 33508 22460
rect 33560 22448 33566 22500
rect 30653 22423 30711 22429
rect 30653 22420 30665 22423
rect 28132 22392 30665 22420
rect 28132 22380 28138 22392
rect 30653 22389 30665 22392
rect 30699 22389 30711 22423
rect 30653 22383 30711 22389
rect 1104 22330 48852 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 48852 22330
rect 1104 22256 48852 22278
rect 12986 22216 12992 22228
rect 2746 22188 12848 22216
rect 12947 22188 12992 22216
rect 2130 22108 2136 22160
rect 2188 22148 2194 22160
rect 2746 22148 2774 22188
rect 2188 22120 2774 22148
rect 2188 22108 2194 22120
rect 9030 22108 9036 22160
rect 9088 22148 9094 22160
rect 11514 22148 11520 22160
rect 9088 22120 11520 22148
rect 9088 22108 9094 22120
rect 11514 22108 11520 22120
rect 11572 22148 11578 22160
rect 12820 22148 12848 22188
rect 12986 22176 12992 22188
rect 13044 22176 13050 22228
rect 15930 22216 15936 22228
rect 15891 22188 15936 22216
rect 15930 22176 15936 22188
rect 15988 22176 15994 22228
rect 16206 22176 16212 22228
rect 16264 22216 16270 22228
rect 16577 22219 16635 22225
rect 16577 22216 16589 22219
rect 16264 22188 16589 22216
rect 16264 22176 16270 22188
rect 16577 22185 16589 22188
rect 16623 22185 16635 22219
rect 16577 22179 16635 22185
rect 18230 22176 18236 22228
rect 18288 22216 18294 22228
rect 18325 22219 18383 22225
rect 18325 22216 18337 22219
rect 18288 22188 18337 22216
rect 18288 22176 18294 22188
rect 18325 22185 18337 22188
rect 18371 22185 18383 22219
rect 19794 22216 19800 22228
rect 18325 22179 18383 22185
rect 18616 22188 19800 22216
rect 18616 22148 18644 22188
rect 19794 22176 19800 22188
rect 19852 22176 19858 22228
rect 20809 22219 20867 22225
rect 20809 22185 20821 22219
rect 20855 22216 20867 22219
rect 21910 22216 21916 22228
rect 20855 22188 21916 22216
rect 20855 22185 20867 22188
rect 20809 22179 20867 22185
rect 21910 22176 21916 22188
rect 21968 22176 21974 22228
rect 23014 22176 23020 22228
rect 23072 22216 23078 22228
rect 27706 22216 27712 22228
rect 23072 22188 27712 22216
rect 23072 22176 23078 22188
rect 27706 22176 27712 22188
rect 27764 22176 27770 22228
rect 30374 22216 30380 22228
rect 30335 22188 30380 22216
rect 30374 22176 30380 22188
rect 30432 22176 30438 22228
rect 33781 22219 33839 22225
rect 33781 22216 33793 22219
rect 30944 22188 33793 22216
rect 11572 22120 11652 22148
rect 12820 22120 18644 22148
rect 11572 22108 11578 22120
rect 6457 22083 6515 22089
rect 6457 22049 6469 22083
rect 6503 22080 6515 22083
rect 8202 22080 8208 22092
rect 6503 22052 8208 22080
rect 6503 22049 6515 22052
rect 6457 22043 6515 22049
rect 8202 22040 8208 22052
rect 8260 22040 8266 22092
rect 8846 22040 8852 22092
rect 8904 22080 8910 22092
rect 11624 22089 11652 22120
rect 18690 22108 18696 22160
rect 18748 22148 18754 22160
rect 19886 22148 19892 22160
rect 18748 22120 19892 22148
rect 18748 22108 18754 22120
rect 19886 22108 19892 22120
rect 19944 22108 19950 22160
rect 21174 22108 21180 22160
rect 21232 22148 21238 22160
rect 21232 22120 22048 22148
rect 21232 22108 21238 22120
rect 8941 22083 8999 22089
rect 8941 22080 8953 22083
rect 8904 22052 8953 22080
rect 8904 22040 8910 22052
rect 8941 22049 8953 22052
rect 8987 22049 8999 22083
rect 8941 22043 8999 22049
rect 11609 22083 11667 22089
rect 11609 22049 11621 22083
rect 11655 22049 11667 22083
rect 11609 22043 11667 22049
rect 19245 22083 19303 22089
rect 19245 22049 19257 22083
rect 19291 22080 19303 22083
rect 19426 22080 19432 22092
rect 19291 22052 19432 22080
rect 19291 22049 19303 22052
rect 19245 22043 19303 22049
rect 19426 22040 19432 22052
rect 19484 22040 19490 22092
rect 22020 22089 22048 22120
rect 25314 22108 25320 22160
rect 25372 22148 25378 22160
rect 30650 22148 30656 22160
rect 25372 22120 30656 22148
rect 25372 22108 25378 22120
rect 30650 22108 30656 22120
rect 30708 22108 30714 22160
rect 22005 22083 22063 22089
rect 19536 22052 21128 22080
rect 9214 22012 9220 22024
rect 9175 21984 9220 22012
rect 9214 21972 9220 21984
rect 9272 21972 9278 22024
rect 9422 22015 9480 22021
rect 9306 22009 9364 22015
rect 9306 21975 9318 22009
rect 9352 21975 9364 22009
rect 9422 21981 9434 22015
rect 9468 22012 9480 22015
rect 9585 22015 9643 22021
rect 9468 21984 9536 22012
rect 9468 21981 9480 21984
rect 9422 21975 9480 21981
rect 9306 21969 9364 21975
rect 6641 21947 6699 21953
rect 6641 21913 6653 21947
rect 6687 21944 6699 21947
rect 6730 21944 6736 21956
rect 6687 21916 6736 21944
rect 6687 21913 6699 21916
rect 6641 21907 6699 21913
rect 6730 21904 6736 21916
rect 6788 21904 6794 21956
rect 8297 21947 8355 21953
rect 8297 21944 8309 21947
rect 6840 21916 8309 21944
rect 4062 21836 4068 21888
rect 4120 21876 4126 21888
rect 6840 21876 6868 21916
rect 8297 21913 8309 21916
rect 8343 21913 8355 21947
rect 8297 21907 8355 21913
rect 9324 21888 9352 21969
rect 4120 21848 6868 21876
rect 4120 21836 4126 21848
rect 9306 21836 9312 21888
rect 9364 21836 9370 21888
rect 9398 21836 9404 21888
rect 9456 21876 9462 21888
rect 9508 21876 9536 21984
rect 9585 21981 9597 22015
rect 9631 22012 9643 22015
rect 9766 22012 9772 22024
rect 9631 21984 9772 22012
rect 9631 21981 9643 21984
rect 9585 21975 9643 21981
rect 9766 21972 9772 21984
rect 9824 21972 9830 22024
rect 16485 22015 16543 22021
rect 16485 21981 16497 22015
rect 16531 22012 16543 22015
rect 17586 22012 17592 22024
rect 16531 21984 17592 22012
rect 16531 21981 16543 21984
rect 16485 21975 16543 21981
rect 17586 21972 17592 21984
rect 17644 21972 17650 22024
rect 19536 22021 19564 22052
rect 19521 22015 19579 22021
rect 19521 21981 19533 22015
rect 19567 21981 19579 22015
rect 19521 21975 19579 21981
rect 19613 22015 19671 22021
rect 19613 21981 19625 22015
rect 19659 21981 19671 22015
rect 19613 21975 19671 21981
rect 19705 22015 19763 22021
rect 19705 21981 19717 22015
rect 19751 22012 19763 22015
rect 19751 21984 19840 22012
rect 19751 21981 19763 21984
rect 19705 21975 19763 21981
rect 10413 21947 10471 21953
rect 10413 21913 10425 21947
rect 10459 21944 10471 21947
rect 10459 21916 11468 21944
rect 10459 21913 10471 21916
rect 10413 21907 10471 21913
rect 9456 21848 9536 21876
rect 9456 21836 9462 21848
rect 10134 21836 10140 21888
rect 10192 21876 10198 21888
rect 10505 21879 10563 21885
rect 10505 21876 10517 21879
rect 10192 21848 10517 21876
rect 10192 21836 10198 21848
rect 10505 21845 10517 21848
rect 10551 21845 10563 21879
rect 11440 21876 11468 21916
rect 11606 21904 11612 21956
rect 11664 21944 11670 21956
rect 11854 21947 11912 21953
rect 11854 21944 11866 21947
rect 11664 21916 11866 21944
rect 11664 21904 11670 21916
rect 11854 21913 11866 21916
rect 11900 21913 11912 21947
rect 11854 21907 11912 21913
rect 13446 21904 13452 21956
rect 13504 21944 13510 21956
rect 15565 21947 15623 21953
rect 15565 21944 15577 21947
rect 13504 21916 15577 21944
rect 13504 21904 13510 21916
rect 15565 21913 15577 21916
rect 15611 21913 15623 21947
rect 15565 21907 15623 21913
rect 15749 21947 15807 21953
rect 15749 21913 15761 21947
rect 15795 21944 15807 21947
rect 16942 21944 16948 21956
rect 15795 21916 16948 21944
rect 15795 21913 15807 21916
rect 15749 21907 15807 21913
rect 12802 21876 12808 21888
rect 11440 21848 12808 21876
rect 10505 21839 10563 21845
rect 12802 21836 12808 21848
rect 12860 21836 12866 21888
rect 15580 21876 15608 21907
rect 16942 21904 16948 21916
rect 17000 21904 17006 21956
rect 17957 21947 18015 21953
rect 17957 21913 17969 21947
rect 18003 21944 18015 21947
rect 18046 21944 18052 21956
rect 18003 21916 18052 21944
rect 18003 21913 18015 21916
rect 17957 21907 18015 21913
rect 18046 21904 18052 21916
rect 18104 21904 18110 21956
rect 18141 21947 18199 21953
rect 18141 21913 18153 21947
rect 18187 21944 18199 21947
rect 18874 21944 18880 21956
rect 18187 21916 18880 21944
rect 18187 21913 18199 21916
rect 18141 21907 18199 21913
rect 18874 21904 18880 21916
rect 18932 21904 18938 21956
rect 17494 21876 17500 21888
rect 15580 21848 17500 21876
rect 17494 21836 17500 21848
rect 17552 21836 17558 21888
rect 19150 21836 19156 21888
rect 19208 21876 19214 21888
rect 19628 21876 19656 21975
rect 19812 21944 19840 21984
rect 19886 21972 19892 22024
rect 19944 22012 19950 22024
rect 20898 22012 20904 22024
rect 19944 21984 20904 22012
rect 19944 21972 19950 21984
rect 20898 21972 20904 21984
rect 20956 21972 20962 22024
rect 20993 22015 21051 22021
rect 20993 21981 21005 22015
rect 21039 21981 21051 22015
rect 21100 22012 21128 22052
rect 22005 22049 22017 22083
rect 22051 22049 22063 22083
rect 22005 22043 22063 22049
rect 23290 22040 23296 22092
rect 23348 22080 23354 22092
rect 23348 22052 24716 22080
rect 23348 22040 23354 22052
rect 24688 22021 24716 22052
rect 24673 22015 24731 22021
rect 21100 21984 24624 22012
rect 20993 21975 21051 21981
rect 20346 21944 20352 21956
rect 19812 21916 20352 21944
rect 20346 21904 20352 21916
rect 20404 21904 20410 21956
rect 19208 21848 19656 21876
rect 21008 21876 21036 21975
rect 21821 21947 21879 21953
rect 21821 21913 21833 21947
rect 21867 21944 21879 21947
rect 22186 21944 22192 21956
rect 21867 21916 22192 21944
rect 21867 21913 21879 21916
rect 21821 21907 21879 21913
rect 22186 21904 22192 21916
rect 22244 21944 22250 21956
rect 22738 21944 22744 21956
rect 22244 21916 22744 21944
rect 22244 21904 22250 21916
rect 22738 21904 22744 21916
rect 22796 21904 22802 21956
rect 24118 21904 24124 21956
rect 24176 21944 24182 21956
rect 24397 21947 24455 21953
rect 24397 21944 24409 21947
rect 24176 21916 24409 21944
rect 24176 21904 24182 21916
rect 24397 21913 24409 21916
rect 24443 21913 24455 21947
rect 24596 21944 24624 21984
rect 24673 21981 24685 22015
rect 24719 21981 24731 22015
rect 24673 21975 24731 21981
rect 25130 21972 25136 22024
rect 25188 22012 25194 22024
rect 30739 22021 30745 22024
rect 30607 22015 30665 22021
rect 30607 22012 30619 22015
rect 25188 21984 30619 22012
rect 25188 21972 25194 21984
rect 30607 21981 30619 21984
rect 30653 21981 30665 22015
rect 30607 21975 30665 21981
rect 30726 22015 30745 22021
rect 30726 21981 30738 22015
rect 30726 21975 30745 21981
rect 30739 21972 30745 21975
rect 30797 21972 30803 22024
rect 30842 22015 30900 22021
rect 30842 21981 30854 22015
rect 30888 22012 30900 22015
rect 30944 22012 30972 22188
rect 33781 22185 33793 22188
rect 33827 22185 33839 22219
rect 33781 22179 33839 22185
rect 31478 22148 31484 22160
rect 31036 22120 31484 22148
rect 31036 22021 31064 22120
rect 31478 22108 31484 22120
rect 31536 22108 31542 22160
rect 31570 22108 31576 22160
rect 31628 22148 31634 22160
rect 48038 22148 48044 22160
rect 31628 22120 48044 22148
rect 31628 22108 31634 22120
rect 48038 22108 48044 22120
rect 48096 22108 48102 22160
rect 31220 22052 31889 22080
rect 30888 21984 30972 22012
rect 31021 22015 31079 22021
rect 30888 21981 30900 21984
rect 30842 21975 30900 21981
rect 31021 21981 31033 22015
rect 31067 21981 31079 22015
rect 31021 21975 31079 21981
rect 30374 21944 30380 21956
rect 24596 21916 30380 21944
rect 24397 21907 24455 21913
rect 30374 21904 30380 21916
rect 30432 21904 30438 21956
rect 30760 21944 30788 21972
rect 31220 21944 31248 22052
rect 31861 22021 31889 22052
rect 32030 22040 32036 22092
rect 32088 22080 32094 22092
rect 48133 22083 48191 22089
rect 48133 22080 48145 22083
rect 32088 22052 48145 22080
rect 32088 22040 32094 22052
rect 48133 22049 48145 22052
rect 48179 22049 48191 22083
rect 48133 22043 48191 22049
rect 31757 22015 31815 22021
rect 31757 21981 31769 22015
rect 31803 21981 31815 22015
rect 31757 21975 31815 21981
rect 31846 22015 31904 22021
rect 31846 21981 31858 22015
rect 31892 21981 31904 22015
rect 31846 21975 31904 21981
rect 31941 22009 31999 22015
rect 32122 22012 32128 22024
rect 31941 21975 31953 22009
rect 31987 21975 31999 22009
rect 32083 21984 32128 22012
rect 31772 21944 31800 21975
rect 31941 21969 31999 21975
rect 32122 21972 32128 21984
rect 32180 21972 32186 22024
rect 32582 22012 32588 22024
rect 32495 21984 32588 22012
rect 32582 21972 32588 21984
rect 32640 22012 32646 22024
rect 33413 22015 33471 22021
rect 33413 22012 33425 22015
rect 32640 21984 33425 22012
rect 32640 21972 32646 21984
rect 33413 21981 33425 21984
rect 33459 21981 33471 22015
rect 33413 21975 33471 21981
rect 33502 21972 33508 22024
rect 33560 22012 33566 22024
rect 33597 22015 33655 22021
rect 33597 22012 33609 22015
rect 33560 21984 33609 22012
rect 33560 21972 33566 21984
rect 33597 21981 33609 21984
rect 33643 21981 33655 22015
rect 33597 21975 33655 21981
rect 34701 22015 34759 22021
rect 34701 21981 34713 22015
rect 34747 21981 34759 22015
rect 34701 21975 34759 21981
rect 36541 22015 36599 22021
rect 36541 21981 36553 22015
rect 36587 22012 36599 22015
rect 45462 22012 45468 22024
rect 36587 21984 45468 22012
rect 36587 21981 36599 21984
rect 36541 21975 36599 21981
rect 30760 21916 31248 21944
rect 31312 21916 31800 21944
rect 21453 21879 21511 21885
rect 21453 21876 21465 21879
rect 21008 21848 21465 21876
rect 19208 21836 19214 21848
rect 21453 21845 21465 21848
rect 21499 21845 21511 21879
rect 21453 21839 21511 21845
rect 21542 21836 21548 21888
rect 21600 21876 21606 21888
rect 21913 21879 21971 21885
rect 21913 21876 21925 21879
rect 21600 21848 21925 21876
rect 21600 21836 21606 21848
rect 21913 21845 21925 21848
rect 21959 21845 21971 21879
rect 21913 21839 21971 21845
rect 23382 21836 23388 21888
rect 23440 21876 23446 21888
rect 24495 21879 24553 21885
rect 24495 21876 24507 21879
rect 23440 21848 24507 21876
rect 23440 21836 23446 21848
rect 24495 21845 24507 21848
rect 24541 21845 24553 21879
rect 24495 21839 24553 21845
rect 24581 21879 24639 21885
rect 24581 21845 24593 21879
rect 24627 21876 24639 21879
rect 24670 21876 24676 21888
rect 24627 21848 24676 21876
rect 24627 21845 24639 21848
rect 24581 21839 24639 21845
rect 24670 21836 24676 21848
rect 24728 21836 24734 21888
rect 24854 21836 24860 21888
rect 24912 21876 24918 21888
rect 25958 21876 25964 21888
rect 24912 21848 25964 21876
rect 24912 21836 24918 21848
rect 25958 21836 25964 21848
rect 26016 21836 26022 21888
rect 28258 21836 28264 21888
rect 28316 21876 28322 21888
rect 31312 21876 31340 21916
rect 31478 21876 31484 21888
rect 28316 21848 31340 21876
rect 31439 21848 31484 21876
rect 28316 21836 28322 21848
rect 31478 21836 31484 21848
rect 31536 21836 31542 21888
rect 31956 21876 31984 21969
rect 32769 21947 32827 21953
rect 32769 21913 32781 21947
rect 32815 21944 32827 21947
rect 33318 21944 33324 21956
rect 32815 21916 33324 21944
rect 32815 21913 32827 21916
rect 32769 21907 32827 21913
rect 33318 21904 33324 21916
rect 33376 21944 33382 21956
rect 34716 21944 34744 21975
rect 45462 21972 45468 21984
rect 45520 21972 45526 22024
rect 33376 21916 34744 21944
rect 34885 21947 34943 21953
rect 33376 21904 33382 21916
rect 34885 21913 34897 21947
rect 34931 21913 34943 21947
rect 47946 21944 47952 21956
rect 47907 21916 47952 21944
rect 34885 21907 34943 21913
rect 32953 21879 33011 21885
rect 32953 21876 32965 21879
rect 31956 21848 32965 21876
rect 32953 21845 32965 21848
rect 32999 21845 33011 21879
rect 32953 21839 33011 21845
rect 34790 21836 34796 21888
rect 34848 21876 34854 21888
rect 34900 21876 34928 21907
rect 47946 21904 47952 21916
rect 48004 21904 48010 21956
rect 34848 21848 34928 21876
rect 34848 21836 34854 21848
rect 1104 21786 48852 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 48852 21786
rect 1104 21712 48852 21734
rect 6730 21672 6736 21684
rect 6691 21644 6736 21672
rect 6730 21632 6736 21644
rect 6788 21632 6794 21684
rect 8478 21632 8484 21684
rect 8536 21672 8542 21684
rect 11606 21672 11612 21684
rect 8536 21644 10272 21672
rect 11567 21644 11612 21672
rect 8536 21632 8542 21644
rect 9306 21564 9312 21616
rect 9364 21604 9370 21616
rect 10134 21604 10140 21616
rect 9364 21576 10140 21604
rect 9364 21564 9370 21576
rect 9597 21548 9625 21576
rect 10134 21564 10140 21576
rect 10192 21564 10198 21616
rect 6638 21536 6644 21548
rect 6599 21508 6644 21536
rect 6638 21496 6644 21508
rect 6696 21496 6702 21548
rect 9398 21496 9404 21548
rect 9456 21502 9462 21548
rect 9493 21539 9551 21545
rect 9493 21505 9505 21539
rect 9539 21505 9551 21539
rect 9493 21502 9551 21505
rect 9582 21542 9640 21548
rect 9582 21508 9594 21542
rect 9628 21508 9640 21542
rect 9582 21502 9640 21508
rect 9677 21539 9735 21545
rect 9677 21505 9689 21539
rect 9723 21505 9735 21539
rect 9456 21499 9551 21502
rect 9677 21499 9735 21505
rect 9456 21496 9536 21499
rect 9416 21474 9536 21496
rect 9692 21468 9720 21499
rect 9858 21496 9864 21548
rect 9916 21536 9922 21548
rect 10244 21536 10272 21644
rect 11606 21632 11612 21644
rect 11664 21632 11670 21684
rect 11974 21632 11980 21684
rect 12032 21632 12038 21684
rect 18969 21675 19027 21681
rect 18969 21641 18981 21675
rect 19015 21672 19027 21675
rect 20346 21672 20352 21684
rect 19015 21644 20352 21672
rect 19015 21641 19027 21644
rect 18969 21635 19027 21641
rect 20346 21632 20352 21644
rect 20404 21632 20410 21684
rect 24029 21675 24087 21681
rect 24029 21672 24041 21675
rect 22204 21644 24041 21672
rect 12005 21551 12033 21632
rect 12713 21607 12771 21613
rect 12713 21573 12725 21607
rect 12759 21604 12771 21607
rect 13446 21604 13452 21616
rect 12759 21576 13452 21604
rect 12759 21573 12771 21576
rect 12713 21567 12771 21573
rect 13446 21564 13452 21576
rect 13504 21564 13510 21616
rect 14001 21607 14059 21613
rect 14001 21573 14013 21607
rect 14047 21604 14059 21607
rect 14734 21604 14740 21616
rect 14047 21576 14740 21604
rect 14047 21573 14059 21576
rect 14001 21567 14059 21573
rect 14734 21564 14740 21576
rect 14792 21564 14798 21616
rect 17773 21607 17831 21613
rect 17773 21573 17785 21607
rect 17819 21604 17831 21607
rect 18046 21604 18052 21616
rect 17819 21576 18052 21604
rect 17819 21573 17831 21576
rect 17773 21567 17831 21573
rect 18046 21564 18052 21576
rect 18104 21604 18110 21616
rect 18601 21607 18659 21613
rect 18601 21604 18613 21607
rect 18104 21576 18613 21604
rect 18104 21564 18110 21576
rect 18601 21573 18613 21576
rect 18647 21604 18659 21607
rect 19058 21604 19064 21616
rect 18647 21576 19064 21604
rect 18647 21573 18659 21576
rect 18601 21567 18659 21573
rect 19058 21564 19064 21576
rect 19116 21604 19122 21616
rect 19242 21604 19248 21616
rect 19116 21576 19248 21604
rect 19116 21564 19122 21576
rect 19242 21564 19248 21576
rect 19300 21564 19306 21616
rect 11990 21545 12048 21551
rect 11839 21539 11897 21545
rect 11839 21536 11851 21539
rect 9916 21508 9961 21536
rect 10244 21508 11851 21536
rect 9916 21496 9922 21508
rect 11839 21505 11851 21508
rect 11885 21505 11897 21539
rect 11990 21511 12002 21545
rect 12036 21511 12048 21545
rect 11990 21505 12048 21511
rect 12090 21539 12148 21545
rect 12090 21505 12102 21539
rect 12136 21536 12148 21539
rect 12253 21539 12311 21545
rect 12136 21508 12204 21536
rect 12136 21505 12148 21508
rect 11839 21499 11897 21505
rect 12090 21499 12148 21505
rect 11146 21468 11152 21480
rect 9692 21440 11152 21468
rect 11146 21428 11152 21440
rect 11204 21428 11210 21480
rect 12176 21468 12204 21508
rect 12253 21505 12265 21539
rect 12299 21536 12311 21539
rect 12342 21536 12348 21548
rect 12299 21508 12348 21536
rect 12299 21505 12311 21508
rect 12253 21499 12311 21505
rect 12342 21496 12348 21508
rect 12400 21496 12406 21548
rect 12897 21539 12955 21545
rect 12897 21505 12909 21539
rect 12943 21536 12955 21539
rect 13538 21536 13544 21548
rect 12943 21508 13544 21536
rect 12943 21505 12955 21508
rect 12897 21499 12955 21505
rect 13538 21496 13544 21508
rect 13596 21496 13602 21548
rect 17957 21539 18015 21545
rect 17957 21505 17969 21539
rect 18003 21536 18015 21539
rect 18414 21536 18420 21548
rect 18003 21508 18420 21536
rect 18003 21505 18015 21508
rect 17957 21499 18015 21505
rect 18414 21496 18420 21508
rect 18472 21496 18478 21548
rect 18785 21539 18843 21545
rect 18785 21505 18797 21539
rect 18831 21505 18843 21539
rect 18785 21499 18843 21505
rect 13081 21471 13139 21477
rect 13081 21468 13093 21471
rect 12176 21440 13093 21468
rect 13081 21437 13093 21440
rect 13127 21437 13139 21471
rect 13814 21468 13820 21480
rect 13775 21440 13820 21468
rect 13081 21431 13139 21437
rect 13814 21428 13820 21440
rect 13872 21428 13878 21480
rect 14277 21471 14335 21477
rect 14277 21437 14289 21471
rect 14323 21437 14335 21471
rect 18800 21468 18828 21499
rect 18874 21496 18880 21548
rect 18932 21536 18938 21548
rect 22204 21536 22232 21644
rect 24029 21641 24041 21644
rect 24075 21672 24087 21675
rect 25590 21672 25596 21684
rect 24075 21644 25596 21672
rect 24075 21641 24087 21644
rect 24029 21635 24087 21641
rect 25590 21632 25596 21644
rect 25648 21632 25654 21684
rect 33318 21632 33324 21684
rect 33376 21672 33382 21684
rect 33873 21675 33931 21681
rect 33873 21672 33885 21675
rect 33376 21644 33885 21672
rect 33376 21632 33382 21644
rect 33873 21641 33885 21644
rect 33919 21641 33931 21675
rect 33873 21635 33931 21641
rect 22738 21604 22744 21616
rect 22699 21576 22744 21604
rect 22738 21564 22744 21576
rect 22796 21564 22802 21616
rect 23106 21564 23112 21616
rect 23164 21604 23170 21616
rect 24121 21607 24179 21613
rect 24121 21604 24133 21607
rect 23164 21576 24133 21604
rect 23164 21564 23170 21576
rect 24121 21573 24133 21576
rect 24167 21573 24179 21607
rect 27614 21604 27620 21616
rect 24121 21567 24179 21573
rect 24964 21576 27620 21604
rect 18932 21508 22232 21536
rect 18932 21496 18938 21508
rect 22370 21496 22376 21548
rect 22428 21536 22434 21548
rect 22649 21539 22707 21545
rect 22649 21536 22661 21539
rect 22428 21508 22661 21536
rect 22428 21496 22434 21508
rect 22649 21505 22661 21508
rect 22695 21505 22707 21539
rect 24854 21536 24860 21548
rect 22649 21499 22707 21505
rect 22848 21508 24860 21536
rect 18800 21440 18920 21468
rect 14277 21431 14335 21437
rect 3970 21360 3976 21412
rect 4028 21400 4034 21412
rect 14292 21400 14320 21431
rect 18892 21400 18920 21440
rect 18966 21428 18972 21480
rect 19024 21468 19030 21480
rect 22848 21468 22876 21508
rect 24854 21496 24860 21508
rect 24912 21496 24918 21548
rect 24964 21545 24992 21576
rect 27614 21564 27620 21576
rect 27672 21564 27678 21616
rect 31478 21564 31484 21616
rect 31536 21604 31542 21616
rect 32738 21607 32796 21613
rect 32738 21604 32750 21607
rect 31536 21576 32750 21604
rect 31536 21564 31542 21576
rect 32738 21573 32750 21576
rect 32784 21573 32796 21607
rect 32738 21567 32796 21573
rect 25222 21545 25228 21548
rect 24949 21539 25007 21545
rect 24949 21505 24961 21539
rect 24995 21505 25007 21539
rect 24949 21499 25007 21505
rect 25216 21499 25228 21545
rect 25280 21536 25286 21548
rect 25280 21508 25316 21536
rect 25222 21496 25228 21499
rect 25280 21496 25286 21508
rect 25590 21496 25596 21548
rect 25648 21536 25654 21548
rect 31205 21539 31263 21545
rect 31205 21536 31217 21539
rect 25648 21508 31217 21536
rect 25648 21496 25654 21508
rect 31205 21505 31217 21508
rect 31251 21505 31263 21539
rect 31205 21499 31263 21505
rect 31297 21539 31355 21545
rect 31297 21505 31309 21539
rect 31343 21505 31355 21539
rect 31297 21499 31355 21505
rect 19024 21440 22876 21468
rect 22925 21471 22983 21477
rect 19024 21428 19030 21440
rect 22925 21437 22937 21471
rect 22971 21468 22983 21471
rect 24210 21468 24216 21480
rect 22971 21440 24216 21468
rect 22971 21437 22983 21440
rect 22925 21431 22983 21437
rect 24210 21428 24216 21440
rect 24268 21428 24274 21480
rect 30742 21428 30748 21480
rect 30800 21468 30806 21480
rect 31312 21468 31340 21499
rect 31386 21496 31392 21548
rect 31444 21536 31450 21548
rect 31444 21508 31489 21536
rect 31444 21496 31450 21508
rect 31570 21496 31576 21548
rect 31628 21536 31634 21548
rect 32122 21536 32128 21548
rect 31628 21508 32128 21536
rect 31628 21496 31634 21508
rect 32122 21496 32128 21508
rect 32180 21496 32186 21548
rect 30800 21440 31340 21468
rect 30800 21428 30806 21440
rect 31478 21428 31484 21480
rect 31536 21468 31542 21480
rect 32493 21471 32551 21477
rect 32493 21468 32505 21471
rect 31536 21440 32505 21468
rect 31536 21428 31542 21440
rect 32493 21437 32505 21440
rect 32539 21437 32551 21471
rect 34514 21468 34520 21480
rect 34475 21440 34520 21468
rect 32493 21431 32551 21437
rect 34514 21428 34520 21440
rect 34572 21428 34578 21480
rect 34698 21468 34704 21480
rect 34659 21440 34704 21468
rect 34698 21428 34704 21440
rect 34756 21428 34762 21480
rect 36357 21471 36415 21477
rect 36357 21437 36369 21471
rect 36403 21468 36415 21471
rect 46566 21468 46572 21480
rect 36403 21440 46572 21468
rect 36403 21437 36415 21440
rect 36357 21431 36415 21437
rect 46566 21428 46572 21440
rect 46624 21428 46630 21480
rect 20714 21400 20720 21412
rect 4028 21372 14320 21400
rect 17972 21372 18828 21400
rect 18892 21372 20720 21400
rect 4028 21360 4034 21372
rect 9214 21332 9220 21344
rect 9175 21304 9220 21332
rect 9214 21292 9220 21304
rect 9272 21292 9278 21344
rect 12802 21292 12808 21344
rect 12860 21332 12866 21344
rect 17972 21332 18000 21372
rect 18138 21332 18144 21344
rect 12860 21304 18000 21332
rect 18099 21304 18144 21332
rect 12860 21292 12866 21304
rect 18138 21292 18144 21304
rect 18196 21292 18202 21344
rect 18800 21332 18828 21372
rect 20714 21360 20720 21372
rect 20772 21360 20778 21412
rect 21818 21360 21824 21412
rect 21876 21400 21882 21412
rect 23106 21400 23112 21412
rect 21876 21372 23112 21400
rect 21876 21360 21882 21372
rect 23106 21360 23112 21372
rect 23164 21400 23170 21412
rect 24946 21400 24952 21412
rect 23164 21372 24952 21400
rect 23164 21360 23170 21372
rect 24946 21360 24952 21372
rect 25004 21360 25010 21412
rect 22094 21332 22100 21344
rect 18800 21304 22100 21332
rect 22094 21292 22100 21304
rect 22152 21292 22158 21344
rect 22278 21332 22284 21344
rect 22239 21304 22284 21332
rect 22278 21292 22284 21304
rect 22336 21292 22342 21344
rect 23290 21292 23296 21344
rect 23348 21332 23354 21344
rect 23661 21335 23719 21341
rect 23661 21332 23673 21335
rect 23348 21304 23673 21332
rect 23348 21292 23354 21304
rect 23661 21301 23673 21304
rect 23707 21301 23719 21335
rect 23661 21295 23719 21301
rect 24670 21292 24676 21344
rect 24728 21332 24734 21344
rect 24854 21332 24860 21344
rect 24728 21304 24860 21332
rect 24728 21292 24734 21304
rect 24854 21292 24860 21304
rect 24912 21292 24918 21344
rect 24964 21332 24992 21360
rect 26329 21335 26387 21341
rect 26329 21332 26341 21335
rect 24964 21304 26341 21332
rect 26329 21301 26341 21304
rect 26375 21301 26387 21335
rect 26329 21295 26387 21301
rect 30929 21335 30987 21341
rect 30929 21301 30941 21335
rect 30975 21332 30987 21335
rect 32766 21332 32772 21344
rect 30975 21304 32772 21332
rect 30975 21301 30987 21304
rect 30929 21295 30987 21301
rect 32766 21292 32772 21304
rect 32824 21292 32830 21344
rect 1104 21242 48852 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 48852 21242
rect 1104 21168 48852 21190
rect 11146 21128 11152 21140
rect 11107 21100 11152 21128
rect 11146 21088 11152 21100
rect 11204 21088 11210 21140
rect 15562 21088 15568 21140
rect 15620 21128 15626 21140
rect 18966 21128 18972 21140
rect 15620 21100 18972 21128
rect 15620 21088 15626 21100
rect 18966 21088 18972 21100
rect 19024 21088 19030 21140
rect 21542 21088 21548 21140
rect 21600 21128 21606 21140
rect 21729 21131 21787 21137
rect 21729 21128 21741 21131
rect 21600 21100 21741 21128
rect 21600 21088 21606 21100
rect 21729 21097 21741 21100
rect 21775 21097 21787 21131
rect 22370 21128 22376 21140
rect 21729 21091 21787 21097
rect 21836 21100 22376 21128
rect 18414 21060 18420 21072
rect 18327 21032 18420 21060
rect 18414 21020 18420 21032
rect 18472 21060 18478 21072
rect 21836 21060 21864 21100
rect 22370 21088 22376 21100
rect 22428 21128 22434 21140
rect 23109 21131 23167 21137
rect 22428 21100 22876 21128
rect 22428 21088 22434 21100
rect 22741 21063 22799 21069
rect 22741 21060 22753 21063
rect 18472 21032 21864 21060
rect 22020 21032 22753 21060
rect 18472 21020 18478 21032
rect 17034 20992 17040 21004
rect 16995 20964 17040 20992
rect 17034 20952 17040 20964
rect 17092 20952 17098 21004
rect 21269 20995 21327 21001
rect 21269 20961 21281 20995
rect 21315 20992 21327 20995
rect 21542 20992 21548 21004
rect 21315 20964 21548 20992
rect 21315 20961 21327 20964
rect 21269 20955 21327 20961
rect 21542 20952 21548 20964
rect 21600 20952 21606 21004
rect 22020 20992 22048 21032
rect 22741 21029 22753 21032
rect 22787 21029 22799 21063
rect 22848 21060 22876 21100
rect 23109 21097 23121 21131
rect 23155 21128 23167 21131
rect 23290 21128 23296 21140
rect 23155 21100 23296 21128
rect 23155 21097 23167 21100
rect 23109 21091 23167 21097
rect 23290 21088 23296 21100
rect 23348 21088 23354 21140
rect 25222 21088 25228 21140
rect 25280 21128 25286 21140
rect 25409 21131 25467 21137
rect 25409 21128 25421 21131
rect 25280 21100 25421 21128
rect 25280 21088 25286 21100
rect 25409 21097 25421 21100
rect 25455 21097 25467 21131
rect 25409 21091 25467 21097
rect 25682 21088 25688 21140
rect 25740 21128 25746 21140
rect 25740 21100 30512 21128
rect 25740 21088 25746 21100
rect 25130 21060 25136 21072
rect 22848 21032 25136 21060
rect 22741 21023 22799 21029
rect 21928 20964 22048 20992
rect 5626 20884 5632 20936
rect 5684 20924 5690 20936
rect 6638 20924 6644 20936
rect 5684 20896 6644 20924
rect 5684 20884 5690 20896
rect 6638 20884 6644 20896
rect 6696 20884 6702 20936
rect 8018 20924 8024 20936
rect 7979 20896 8024 20924
rect 8018 20884 8024 20896
rect 8076 20884 8082 20936
rect 8938 20924 8944 20936
rect 8851 20896 8944 20924
rect 8938 20884 8944 20896
rect 8996 20884 9002 20936
rect 9214 20933 9220 20936
rect 9208 20924 9220 20933
rect 9175 20896 9220 20924
rect 9208 20887 9220 20896
rect 9214 20884 9220 20887
rect 9272 20884 9278 20936
rect 10778 20924 10784 20936
rect 10739 20896 10784 20924
rect 10778 20884 10784 20896
rect 10836 20884 10842 20936
rect 12986 20884 12992 20936
rect 13044 20924 13050 20936
rect 14185 20927 14243 20933
rect 14185 20924 14197 20927
rect 13044 20896 14197 20924
rect 13044 20884 13050 20896
rect 14185 20893 14197 20896
rect 14231 20924 14243 20927
rect 15930 20924 15936 20936
rect 14231 20896 15936 20924
rect 14231 20893 14243 20896
rect 14185 20887 14243 20893
rect 15930 20884 15936 20896
rect 15988 20884 15994 20936
rect 20990 20924 20996 20936
rect 20951 20896 20996 20924
rect 20990 20884 20996 20896
rect 21048 20884 21054 20936
rect 21082 20884 21088 20936
rect 21140 20924 21146 20936
rect 21928 20933 21956 20964
rect 22186 20952 22192 21004
rect 22244 20992 22250 21004
rect 22244 20964 22289 20992
rect 22244 20952 22250 20964
rect 21913 20927 21971 20933
rect 21140 20896 21185 20924
rect 21140 20884 21146 20896
rect 21913 20893 21925 20927
rect 21959 20893 21971 20927
rect 21913 20887 21971 20893
rect 22005 20927 22063 20933
rect 22005 20893 22017 20927
rect 22051 20893 22063 20927
rect 22005 20887 22063 20893
rect 22281 20927 22339 20933
rect 22281 20893 22293 20927
rect 22327 20893 22339 20927
rect 22281 20887 22339 20893
rect 8202 20856 8208 20868
rect 8163 20828 8208 20856
rect 8202 20816 8208 20828
rect 8260 20816 8266 20868
rect 8956 20856 8984 20884
rect 9122 20856 9128 20868
rect 8956 20828 9128 20856
rect 9122 20816 9128 20828
rect 9180 20816 9186 20868
rect 10965 20859 11023 20865
rect 10965 20825 10977 20859
rect 11011 20825 11023 20859
rect 10965 20819 11023 20825
rect 6638 20748 6644 20800
rect 6696 20788 6702 20800
rect 6733 20791 6791 20797
rect 6733 20788 6745 20791
rect 6696 20760 6745 20788
rect 6696 20748 6702 20760
rect 6733 20757 6745 20760
rect 6779 20757 6791 20791
rect 6733 20751 6791 20757
rect 8389 20791 8447 20797
rect 8389 20757 8401 20791
rect 8435 20788 8447 20791
rect 9398 20788 9404 20800
rect 8435 20760 9404 20788
rect 8435 20757 8447 20760
rect 8389 20751 8447 20757
rect 9398 20748 9404 20760
rect 9456 20748 9462 20800
rect 10318 20788 10324 20800
rect 10279 20760 10324 20788
rect 10318 20748 10324 20760
rect 10376 20788 10382 20800
rect 10980 20788 11008 20819
rect 13906 20816 13912 20868
rect 13964 20856 13970 20868
rect 14430 20859 14488 20865
rect 14430 20856 14442 20859
rect 13964 20828 14442 20856
rect 13964 20816 13970 20828
rect 14430 20825 14442 20828
rect 14476 20825 14488 20859
rect 14430 20819 14488 20825
rect 16850 20816 16856 20868
rect 16908 20856 16914 20868
rect 17282 20859 17340 20865
rect 17282 20856 17294 20859
rect 16908 20828 17294 20856
rect 16908 20816 16914 20828
rect 17282 20825 17294 20828
rect 17328 20825 17340 20859
rect 17282 20819 17340 20825
rect 21269 20859 21327 20865
rect 21269 20825 21281 20859
rect 21315 20856 21327 20859
rect 22020 20856 22048 20887
rect 21315 20828 22048 20856
rect 22296 20856 22324 20887
rect 22370 20884 22376 20936
rect 22428 20924 22434 20936
rect 22925 20927 22983 20933
rect 22925 20924 22937 20927
rect 22428 20896 22937 20924
rect 22428 20884 22434 20896
rect 22925 20893 22937 20896
rect 22971 20893 22983 20927
rect 22925 20887 22983 20893
rect 23032 20856 23060 21032
rect 25130 21020 25136 21032
rect 25188 21020 25194 21072
rect 25700 21032 26648 21060
rect 23474 20952 23480 21004
rect 23532 20992 23538 21004
rect 24394 20992 24400 21004
rect 23532 20964 24400 20992
rect 23532 20952 23538 20964
rect 24394 20952 24400 20964
rect 24452 20952 24458 21004
rect 24946 20992 24952 21004
rect 24907 20964 24952 20992
rect 24946 20952 24952 20964
rect 25004 20952 25010 21004
rect 25041 20995 25099 21001
rect 25041 20961 25053 20995
rect 25087 20992 25099 20995
rect 25314 20992 25320 21004
rect 25087 20964 25320 20992
rect 25087 20961 25099 20964
rect 25041 20955 25099 20961
rect 25314 20952 25320 20964
rect 25372 20952 25378 21004
rect 23106 20884 23112 20936
rect 23164 20924 23170 20936
rect 23201 20927 23259 20933
rect 23201 20924 23213 20927
rect 23164 20896 23213 20924
rect 23164 20884 23170 20896
rect 23201 20893 23213 20896
rect 23247 20893 23259 20927
rect 23845 20927 23903 20933
rect 23845 20924 23857 20927
rect 23201 20887 23259 20893
rect 23492 20896 23857 20924
rect 22296 20828 23060 20856
rect 21315 20825 21327 20828
rect 21269 20819 21327 20825
rect 23492 20800 23520 20896
rect 23845 20893 23857 20896
rect 23891 20893 23903 20927
rect 24670 20924 24676 20936
rect 24631 20896 24676 20924
rect 23845 20887 23903 20893
rect 24670 20884 24676 20896
rect 24728 20884 24734 20936
rect 24857 20927 24915 20933
rect 24857 20893 24869 20927
rect 24903 20924 24915 20927
rect 25130 20924 25136 20936
rect 24903 20896 25136 20924
rect 24903 20893 24915 20896
rect 24857 20887 24915 20893
rect 25130 20884 25136 20896
rect 25188 20884 25194 20936
rect 25225 20927 25283 20933
rect 25225 20893 25237 20927
rect 25271 20924 25283 20927
rect 25590 20924 25596 20936
rect 25271 20896 25596 20924
rect 25271 20893 25283 20896
rect 25225 20887 25283 20893
rect 25590 20884 25596 20896
rect 25648 20884 25654 20936
rect 24946 20816 24952 20868
rect 25004 20856 25010 20868
rect 25700 20856 25728 21032
rect 26142 20992 26148 21004
rect 26103 20964 26148 20992
rect 26142 20952 26148 20964
rect 26200 20952 26206 21004
rect 25866 20924 25872 20936
rect 25827 20896 25872 20924
rect 25866 20884 25872 20896
rect 25924 20884 25930 20936
rect 25958 20884 25964 20936
rect 26016 20924 26022 20936
rect 26620 20933 26648 21032
rect 30484 21001 30512 21100
rect 31386 21088 31392 21140
rect 31444 21128 31450 21140
rect 32217 21131 32275 21137
rect 32217 21128 32229 21131
rect 31444 21100 32229 21128
rect 31444 21088 31450 21100
rect 32217 21097 32229 21100
rect 32263 21097 32275 21131
rect 34790 21128 34796 21140
rect 34751 21100 34796 21128
rect 32217 21091 32275 21097
rect 34790 21088 34796 21100
rect 34848 21088 34854 21140
rect 30469 20995 30527 21001
rect 30469 20961 30481 20995
rect 30515 20961 30527 20995
rect 30742 20992 30748 21004
rect 30703 20964 30748 20992
rect 30469 20955 30527 20961
rect 30742 20952 30748 20964
rect 30800 20952 30806 21004
rect 26605 20927 26663 20933
rect 26016 20896 26061 20924
rect 26016 20884 26022 20896
rect 26605 20893 26617 20927
rect 26651 20893 26663 20927
rect 26605 20887 26663 20893
rect 26789 20927 26847 20933
rect 26789 20893 26801 20927
rect 26835 20893 26847 20927
rect 27614 20924 27620 20936
rect 27527 20896 27620 20924
rect 26789 20887 26847 20893
rect 25004 20828 25728 20856
rect 25976 20856 26004 20884
rect 26804 20856 26832 20887
rect 27614 20884 27620 20896
rect 27672 20924 27678 20936
rect 28626 20924 28632 20936
rect 27672 20896 28632 20924
rect 27672 20884 27678 20896
rect 28626 20884 28632 20896
rect 28684 20924 28690 20936
rect 31478 20924 31484 20936
rect 28684 20896 31484 20924
rect 28684 20884 28690 20896
rect 31478 20884 31484 20896
rect 31536 20884 31542 20936
rect 32122 20884 32128 20936
rect 32180 20924 32186 20936
rect 32677 20927 32735 20933
rect 32677 20924 32689 20927
rect 32180 20896 32689 20924
rect 32180 20884 32186 20896
rect 32677 20893 32689 20896
rect 32723 20893 32735 20927
rect 32677 20887 32735 20893
rect 32766 20884 32772 20936
rect 32824 20924 32830 20936
rect 32933 20927 32991 20933
rect 32933 20924 32945 20927
rect 32824 20896 32945 20924
rect 32824 20884 32830 20896
rect 32933 20893 32945 20896
rect 32979 20893 32991 20927
rect 32933 20887 32991 20893
rect 34238 20884 34244 20936
rect 34296 20924 34302 20936
rect 34701 20927 34759 20933
rect 34701 20924 34713 20927
rect 34296 20896 34713 20924
rect 34296 20884 34302 20896
rect 34701 20893 34713 20896
rect 34747 20893 34759 20927
rect 34701 20887 34759 20893
rect 25976 20828 26832 20856
rect 25004 20816 25010 20828
rect 27706 20816 27712 20868
rect 27764 20856 27770 20868
rect 27862 20859 27920 20865
rect 27862 20856 27874 20859
rect 27764 20828 27874 20856
rect 27764 20816 27770 20828
rect 27862 20825 27874 20828
rect 27908 20825 27920 20859
rect 27862 20819 27920 20825
rect 31849 20859 31907 20865
rect 31849 20825 31861 20859
rect 31895 20825 31907 20859
rect 31849 20819 31907 20825
rect 32033 20859 32091 20865
rect 32033 20825 32045 20859
rect 32079 20856 32091 20859
rect 34514 20856 34520 20868
rect 32079 20828 34520 20856
rect 32079 20825 32091 20828
rect 32033 20819 32091 20825
rect 15562 20788 15568 20800
rect 10376 20760 11008 20788
rect 15523 20760 15568 20788
rect 10376 20748 10382 20760
rect 15562 20748 15568 20760
rect 15620 20748 15626 20800
rect 21542 20748 21548 20800
rect 21600 20788 21606 20800
rect 23474 20788 23480 20800
rect 21600 20760 23480 20788
rect 21600 20748 21606 20760
rect 23474 20748 23480 20760
rect 23532 20748 23538 20800
rect 23658 20788 23664 20800
rect 23619 20760 23664 20788
rect 23658 20748 23664 20760
rect 23716 20748 23722 20800
rect 23750 20748 23756 20800
rect 23808 20788 23814 20800
rect 26145 20791 26203 20797
rect 26145 20788 26157 20791
rect 23808 20760 26157 20788
rect 23808 20748 23814 20760
rect 26145 20757 26157 20760
rect 26191 20757 26203 20791
rect 26145 20751 26203 20757
rect 26418 20748 26424 20800
rect 26476 20788 26482 20800
rect 26697 20791 26755 20797
rect 26697 20788 26709 20791
rect 26476 20760 26709 20788
rect 26476 20748 26482 20760
rect 26697 20757 26709 20760
rect 26743 20757 26755 20791
rect 28994 20788 29000 20800
rect 28955 20760 29000 20788
rect 26697 20751 26755 20757
rect 28994 20748 29000 20760
rect 29052 20748 29058 20800
rect 31864 20788 31892 20819
rect 32214 20788 32220 20800
rect 31864 20760 32220 20788
rect 32214 20748 32220 20760
rect 32272 20788 32278 20800
rect 32582 20788 32588 20800
rect 32272 20760 32588 20788
rect 32272 20748 32278 20760
rect 32582 20748 32588 20760
rect 32640 20748 32646 20800
rect 34072 20797 34100 20828
rect 34514 20816 34520 20828
rect 34572 20816 34578 20868
rect 34057 20791 34115 20797
rect 34057 20757 34069 20791
rect 34103 20757 34115 20791
rect 34057 20751 34115 20757
rect 1104 20698 48852 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 48852 20698
rect 1104 20624 48852 20646
rect 10318 20584 10324 20596
rect 7852 20556 10324 20584
rect 5721 20519 5779 20525
rect 5721 20485 5733 20519
rect 5767 20516 5779 20519
rect 6549 20519 6607 20525
rect 6549 20516 6561 20519
rect 5767 20488 6561 20516
rect 5767 20485 5779 20488
rect 5721 20479 5779 20485
rect 6549 20485 6561 20488
rect 6595 20485 6607 20519
rect 6549 20479 6607 20485
rect 5626 20448 5632 20460
rect 5587 20420 5632 20448
rect 5626 20408 5632 20420
rect 5684 20408 5690 20460
rect 6365 20383 6423 20389
rect 6365 20349 6377 20383
rect 6411 20380 6423 20383
rect 7852 20380 7880 20556
rect 10318 20544 10324 20556
rect 10376 20544 10382 20596
rect 13906 20584 13912 20596
rect 13867 20556 13912 20584
rect 13906 20544 13912 20556
rect 13964 20544 13970 20596
rect 14826 20584 14832 20596
rect 14200 20556 14832 20584
rect 9122 20516 9128 20528
rect 8680 20488 9128 20516
rect 8680 20457 8708 20488
rect 9122 20476 9128 20488
rect 9180 20476 9186 20528
rect 10505 20519 10563 20525
rect 10505 20485 10517 20519
rect 10551 20516 10563 20519
rect 10778 20516 10784 20528
rect 10551 20488 10784 20516
rect 10551 20485 10563 20488
rect 10505 20479 10563 20485
rect 10778 20476 10784 20488
rect 10836 20476 10842 20528
rect 14200 20516 14228 20556
rect 14826 20544 14832 20556
rect 14884 20544 14890 20596
rect 16850 20584 16856 20596
rect 16811 20556 16856 20584
rect 16850 20544 16856 20556
rect 16908 20544 16914 20596
rect 19150 20584 19156 20596
rect 17236 20556 19156 20584
rect 17236 20516 17264 20556
rect 18138 20516 18144 20528
rect 13280 20488 14228 20516
rect 15948 20488 17264 20516
rect 8938 20457 8944 20460
rect 8665 20451 8723 20457
rect 8665 20417 8677 20451
rect 8711 20417 8723 20451
rect 8665 20411 8723 20417
rect 8932 20411 8944 20457
rect 8996 20448 9002 20460
rect 10686 20448 10692 20460
rect 8996 20420 9032 20448
rect 10647 20420 10692 20448
rect 8938 20408 8944 20411
rect 8996 20408 9002 20420
rect 10686 20408 10692 20420
rect 10744 20408 10750 20460
rect 13280 20457 13308 20488
rect 14182 20457 14188 20460
rect 13265 20451 13323 20457
rect 13265 20417 13277 20451
rect 13311 20417 13323 20451
rect 13265 20411 13323 20417
rect 14165 20451 14188 20457
rect 14165 20417 14177 20451
rect 14165 20411 14188 20417
rect 14182 20408 14188 20411
rect 14240 20408 14246 20460
rect 14277 20451 14335 20457
rect 14277 20417 14289 20451
rect 14323 20417 14335 20451
rect 14277 20411 14335 20417
rect 14390 20451 14448 20457
rect 14390 20417 14402 20451
rect 14436 20417 14448 20451
rect 14390 20411 14448 20417
rect 8018 20380 8024 20392
rect 6411 20352 7880 20380
rect 7979 20352 8024 20380
rect 6411 20349 6423 20352
rect 6365 20343 6423 20349
rect 8018 20340 8024 20352
rect 8076 20340 8082 20392
rect 14292 20324 14320 20411
rect 14405 20380 14433 20411
rect 14550 20408 14556 20460
rect 14608 20448 14614 20460
rect 15948 20457 15976 20488
rect 15933 20451 15991 20457
rect 14608 20420 14653 20448
rect 14608 20408 14614 20420
rect 15933 20417 15945 20451
rect 15979 20417 15991 20451
rect 15933 20411 15991 20417
rect 16117 20451 16175 20457
rect 16117 20417 16129 20451
rect 16163 20448 16175 20451
rect 16574 20448 16580 20460
rect 16163 20420 16580 20448
rect 16163 20417 16175 20420
rect 16117 20411 16175 20417
rect 16574 20408 16580 20420
rect 16632 20408 16638 20460
rect 17126 20448 17132 20460
rect 17087 20420 17132 20448
rect 17126 20408 17132 20420
rect 17184 20408 17190 20460
rect 17236 20457 17264 20488
rect 17328 20488 18144 20516
rect 17328 20457 17356 20488
rect 18138 20476 18144 20488
rect 18196 20476 18202 20528
rect 17221 20451 17279 20457
rect 17221 20417 17233 20451
rect 17267 20417 17279 20451
rect 17221 20411 17279 20417
rect 17313 20451 17371 20457
rect 17313 20417 17325 20451
rect 17359 20417 17371 20451
rect 17313 20411 17371 20417
rect 17497 20451 17555 20457
rect 17497 20417 17509 20451
rect 17543 20417 17555 20451
rect 18230 20448 18236 20460
rect 18191 20420 18236 20448
rect 17497 20411 17555 20417
rect 16025 20383 16083 20389
rect 16025 20380 16037 20383
rect 14405 20352 16037 20380
rect 16025 20349 16037 20352
rect 16071 20349 16083 20383
rect 17512 20380 17540 20411
rect 18230 20408 18236 20420
rect 18288 20408 18294 20460
rect 18340 20457 18368 20556
rect 19150 20544 19156 20556
rect 19208 20544 19214 20596
rect 20070 20544 20076 20596
rect 20128 20544 20134 20596
rect 23290 20544 23296 20596
rect 23348 20544 23354 20596
rect 23477 20587 23535 20593
rect 23477 20553 23489 20587
rect 23523 20584 23535 20587
rect 24118 20584 24124 20596
rect 23523 20556 24124 20584
rect 23523 20553 23535 20556
rect 23477 20547 23535 20553
rect 24118 20544 24124 20556
rect 24176 20584 24182 20596
rect 24486 20584 24492 20596
rect 24176 20556 24492 20584
rect 24176 20544 24182 20556
rect 24486 20544 24492 20556
rect 24544 20544 24550 20596
rect 25866 20544 25872 20596
rect 25924 20584 25930 20596
rect 32858 20584 32864 20596
rect 25924 20556 32864 20584
rect 25924 20544 25930 20556
rect 32858 20544 32864 20556
rect 32916 20544 32922 20596
rect 34425 20587 34483 20593
rect 34425 20553 34437 20587
rect 34471 20584 34483 20587
rect 34698 20584 34704 20596
rect 34471 20556 34704 20584
rect 34471 20553 34483 20556
rect 34425 20547 34483 20553
rect 34698 20544 34704 20556
rect 34756 20544 34762 20596
rect 19429 20519 19487 20525
rect 19429 20516 19441 20519
rect 18432 20488 19441 20516
rect 18432 20457 18460 20488
rect 19429 20485 19441 20488
rect 19475 20485 19487 20519
rect 20088 20516 20116 20544
rect 19429 20479 19487 20485
rect 19536 20488 20116 20516
rect 22189 20519 22247 20525
rect 18325 20451 18383 20457
rect 18325 20417 18337 20451
rect 18371 20417 18383 20451
rect 18325 20411 18383 20417
rect 18417 20451 18475 20457
rect 18417 20417 18429 20451
rect 18463 20417 18475 20451
rect 18417 20411 18475 20417
rect 18601 20451 18659 20457
rect 18601 20417 18613 20451
rect 18647 20448 18659 20451
rect 18690 20448 18696 20460
rect 18647 20420 18696 20448
rect 18647 20417 18659 20420
rect 18601 20411 18659 20417
rect 18616 20380 18644 20411
rect 18690 20408 18696 20420
rect 18748 20408 18754 20460
rect 19058 20448 19064 20460
rect 19019 20420 19064 20448
rect 19058 20408 19064 20420
rect 19116 20408 19122 20460
rect 19242 20448 19248 20460
rect 19203 20420 19248 20448
rect 19242 20408 19248 20420
rect 19300 20408 19306 20460
rect 17512 20352 18644 20380
rect 16025 20343 16083 20349
rect 19150 20340 19156 20392
rect 19208 20380 19214 20392
rect 19536 20380 19564 20488
rect 22189 20485 22201 20519
rect 22235 20516 22247 20519
rect 22278 20516 22284 20528
rect 22235 20488 22284 20516
rect 22235 20485 22247 20488
rect 22189 20479 22247 20485
rect 22278 20476 22284 20488
rect 22336 20476 22342 20528
rect 22373 20519 22431 20525
rect 22373 20485 22385 20519
rect 22419 20516 22431 20519
rect 23308 20516 23336 20544
rect 24210 20516 24216 20528
rect 22419 20488 23336 20516
rect 23584 20488 24216 20516
rect 22419 20485 22431 20488
rect 22373 20479 22431 20485
rect 20070 20408 20076 20460
rect 20128 20448 20134 20460
rect 20165 20451 20223 20457
rect 20165 20448 20177 20451
rect 20128 20420 20177 20448
rect 20128 20408 20134 20420
rect 20165 20417 20177 20420
rect 20211 20417 20223 20451
rect 20530 20448 20536 20460
rect 20165 20411 20223 20417
rect 20456 20420 20536 20448
rect 20456 20389 20484 20420
rect 20530 20408 20536 20420
rect 20588 20448 20594 20460
rect 20901 20451 20959 20457
rect 20901 20448 20913 20451
rect 20588 20420 20913 20448
rect 20588 20408 20594 20420
rect 20901 20417 20913 20420
rect 20947 20417 20959 20451
rect 20901 20411 20959 20417
rect 20990 20408 20996 20460
rect 21048 20448 21054 20460
rect 21085 20451 21143 20457
rect 21085 20448 21097 20451
rect 21048 20420 21097 20448
rect 21048 20408 21054 20420
rect 21085 20417 21097 20420
rect 21131 20448 21143 20451
rect 21542 20448 21548 20460
rect 21131 20420 21548 20448
rect 21131 20417 21143 20420
rect 21085 20411 21143 20417
rect 21542 20408 21548 20420
rect 21600 20408 21606 20460
rect 23293 20451 23351 20457
rect 23293 20417 23305 20451
rect 23339 20448 23351 20451
rect 23584 20448 23612 20488
rect 24210 20476 24216 20488
rect 24268 20516 24274 20528
rect 27893 20519 27951 20525
rect 24268 20488 26096 20516
rect 24268 20476 24274 20488
rect 23339 20420 23612 20448
rect 23339 20417 23351 20420
rect 23293 20411 23351 20417
rect 23658 20408 23664 20460
rect 23716 20448 23722 20460
rect 24305 20451 24363 20457
rect 24305 20448 24317 20451
rect 23716 20420 24317 20448
rect 23716 20408 23722 20420
rect 24305 20417 24317 20420
rect 24351 20448 24363 20451
rect 25133 20451 25191 20457
rect 25133 20448 25145 20451
rect 24351 20420 25145 20448
rect 24351 20417 24363 20420
rect 24305 20411 24363 20417
rect 25133 20417 25145 20420
rect 25179 20448 25191 20451
rect 25958 20448 25964 20460
rect 25179 20420 25964 20448
rect 25179 20417 25191 20420
rect 25133 20411 25191 20417
rect 25958 20408 25964 20420
rect 26016 20408 26022 20460
rect 19208 20352 19564 20380
rect 20441 20383 20499 20389
rect 19208 20340 19214 20352
rect 20441 20349 20453 20383
rect 20487 20349 20499 20383
rect 20441 20343 20499 20349
rect 21266 20340 21272 20392
rect 21324 20380 21330 20392
rect 21634 20380 21640 20392
rect 21324 20352 21640 20380
rect 21324 20340 21330 20352
rect 21634 20340 21640 20352
rect 21692 20340 21698 20392
rect 26068 20380 26096 20488
rect 27893 20485 27905 20519
rect 27939 20516 27951 20519
rect 28994 20516 29000 20528
rect 27939 20488 29000 20516
rect 27939 20485 27951 20488
rect 27893 20479 27951 20485
rect 28994 20476 29000 20488
rect 29052 20476 29058 20528
rect 27798 20448 27804 20460
rect 27711 20420 27804 20448
rect 27798 20408 27804 20420
rect 27856 20448 27862 20460
rect 28813 20451 28871 20457
rect 27856 20420 28764 20448
rect 27856 20408 27862 20420
rect 27982 20380 27988 20392
rect 26068 20352 27988 20380
rect 27982 20340 27988 20352
rect 28040 20340 28046 20392
rect 28736 20380 28764 20420
rect 28813 20417 28825 20451
rect 28859 20448 28871 20451
rect 29178 20448 29184 20460
rect 28859 20420 29184 20448
rect 28859 20417 28871 20420
rect 28813 20411 28871 20417
rect 29178 20408 29184 20420
rect 29236 20408 29242 20460
rect 30466 20408 30472 20460
rect 30524 20448 30530 20460
rect 30837 20451 30895 20457
rect 30837 20448 30849 20451
rect 30524 20420 30849 20448
rect 30524 20408 30530 20420
rect 30837 20417 30849 20420
rect 30883 20417 30895 20451
rect 32125 20451 32183 20457
rect 32125 20448 32137 20451
rect 30837 20411 30895 20417
rect 31726 20420 32137 20448
rect 29089 20383 29147 20389
rect 29089 20380 29101 20383
rect 28736 20352 29101 20380
rect 29089 20349 29101 20352
rect 29135 20380 29147 20383
rect 30374 20380 30380 20392
rect 29135 20352 30380 20380
rect 29135 20349 29147 20352
rect 29089 20343 29147 20349
rect 30374 20340 30380 20352
rect 30432 20340 30438 20392
rect 31726 20324 31754 20420
rect 32125 20417 32137 20420
rect 32171 20448 32183 20451
rect 32214 20448 32220 20460
rect 32171 20420 32220 20448
rect 32171 20417 32183 20420
rect 32125 20411 32183 20417
rect 32214 20408 32220 20420
rect 32272 20408 32278 20460
rect 32309 20451 32367 20457
rect 32309 20417 32321 20451
rect 32355 20448 32367 20451
rect 32582 20448 32588 20460
rect 32355 20420 32588 20448
rect 32355 20417 32367 20420
rect 32309 20411 32367 20417
rect 32582 20408 32588 20420
rect 32640 20408 32646 20460
rect 34238 20408 34244 20460
rect 34296 20448 34302 20460
rect 34333 20451 34391 20457
rect 34333 20448 34345 20451
rect 34296 20420 34345 20448
rect 34296 20408 34302 20420
rect 34333 20417 34345 20420
rect 34379 20417 34391 20451
rect 34333 20411 34391 20417
rect 14274 20272 14280 20324
rect 14332 20272 14338 20324
rect 20257 20315 20315 20321
rect 20257 20281 20269 20315
rect 20303 20312 20315 20315
rect 22557 20315 22615 20321
rect 22557 20312 22569 20315
rect 20303 20284 22569 20312
rect 20303 20281 20315 20284
rect 20257 20275 20315 20281
rect 21008 20256 21036 20284
rect 22557 20281 22569 20284
rect 22603 20281 22615 20315
rect 22557 20275 22615 20281
rect 25409 20315 25467 20321
rect 25409 20281 25421 20315
rect 25455 20312 25467 20315
rect 27798 20312 27804 20324
rect 25455 20284 27804 20312
rect 25455 20281 25467 20284
rect 25409 20275 25467 20281
rect 27798 20272 27804 20284
rect 27856 20312 27862 20324
rect 28718 20312 28724 20324
rect 27856 20284 28724 20312
rect 27856 20272 27862 20284
rect 28718 20272 28724 20284
rect 28776 20272 28782 20324
rect 30653 20315 30711 20321
rect 30653 20281 30665 20315
rect 30699 20312 30711 20315
rect 31726 20312 31760 20324
rect 30699 20284 31760 20312
rect 30699 20281 30711 20284
rect 30653 20275 30711 20281
rect 31754 20272 31760 20284
rect 31812 20272 31818 20324
rect 8202 20204 8208 20256
rect 8260 20244 8266 20256
rect 10045 20247 10103 20253
rect 10045 20244 10057 20247
rect 8260 20216 10057 20244
rect 8260 20204 8266 20216
rect 10045 20213 10057 20216
rect 10091 20213 10103 20247
rect 10045 20207 10103 20213
rect 10134 20204 10140 20256
rect 10192 20244 10198 20256
rect 10873 20247 10931 20253
rect 10873 20244 10885 20247
rect 10192 20216 10885 20244
rect 10192 20204 10198 20216
rect 10873 20213 10885 20216
rect 10919 20213 10931 20247
rect 10873 20207 10931 20213
rect 12526 20204 12532 20256
rect 12584 20244 12590 20256
rect 13357 20247 13415 20253
rect 13357 20244 13369 20247
rect 12584 20216 13369 20244
rect 12584 20204 12590 20216
rect 13357 20213 13369 20216
rect 13403 20213 13415 20247
rect 13357 20207 13415 20213
rect 17586 20204 17592 20256
rect 17644 20244 17650 20256
rect 17957 20247 18015 20253
rect 17957 20244 17969 20247
rect 17644 20216 17969 20244
rect 17644 20204 17650 20216
rect 17957 20213 17969 20216
rect 18003 20213 18015 20247
rect 17957 20207 18015 20213
rect 20346 20204 20352 20256
rect 20404 20244 20410 20256
rect 20990 20244 20996 20256
rect 20404 20216 20449 20244
rect 20951 20216 20996 20244
rect 20404 20204 20410 20216
rect 20990 20204 20996 20216
rect 21048 20204 21054 20256
rect 21269 20247 21327 20253
rect 21269 20213 21281 20247
rect 21315 20244 21327 20247
rect 22278 20244 22284 20256
rect 21315 20216 22284 20244
rect 21315 20213 21327 20216
rect 21269 20207 21327 20213
rect 22278 20204 22284 20216
rect 22336 20204 22342 20256
rect 24486 20244 24492 20256
rect 24447 20216 24492 20244
rect 24486 20204 24492 20216
rect 24544 20244 24550 20256
rect 24762 20244 24768 20256
rect 24544 20216 24768 20244
rect 24544 20204 24550 20216
rect 24762 20204 24768 20216
rect 24820 20204 24826 20256
rect 25314 20204 25320 20256
rect 25372 20244 25378 20256
rect 25682 20244 25688 20256
rect 25372 20216 25688 20244
rect 25372 20204 25378 20216
rect 25682 20204 25688 20216
rect 25740 20244 25746 20256
rect 26145 20247 26203 20253
rect 26145 20244 26157 20247
rect 25740 20216 26157 20244
rect 25740 20204 25746 20216
rect 26145 20213 26157 20216
rect 26191 20213 26203 20247
rect 26145 20207 26203 20213
rect 26694 20204 26700 20256
rect 26752 20244 26758 20256
rect 27433 20247 27491 20253
rect 27433 20244 27445 20247
rect 26752 20216 27445 20244
rect 26752 20204 26758 20216
rect 27433 20213 27445 20216
rect 27479 20213 27491 20247
rect 27433 20207 27491 20213
rect 27522 20204 27528 20256
rect 27580 20244 27586 20256
rect 28629 20247 28687 20253
rect 28629 20244 28641 20247
rect 27580 20216 28641 20244
rect 27580 20204 27586 20216
rect 28629 20213 28641 20216
rect 28675 20213 28687 20247
rect 28629 20207 28687 20213
rect 28997 20247 29055 20253
rect 28997 20213 29009 20247
rect 29043 20244 29055 20247
rect 29086 20244 29092 20256
rect 29043 20216 29092 20244
rect 29043 20213 29055 20216
rect 28997 20207 29055 20213
rect 29086 20204 29092 20216
rect 29144 20204 29150 20256
rect 32493 20247 32551 20253
rect 32493 20213 32505 20247
rect 32539 20244 32551 20247
rect 33134 20244 33140 20256
rect 32539 20216 33140 20244
rect 32539 20213 32551 20216
rect 32493 20207 32551 20213
rect 33134 20204 33140 20216
rect 33192 20204 33198 20256
rect 46290 20204 46296 20256
rect 46348 20244 46354 20256
rect 47765 20247 47823 20253
rect 47765 20244 47777 20247
rect 46348 20216 47777 20244
rect 46348 20204 46354 20216
rect 47765 20213 47777 20216
rect 47811 20213 47823 20247
rect 47765 20207 47823 20213
rect 1104 20154 48852 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 48852 20154
rect 1104 20080 48852 20102
rect 8938 20040 8944 20052
rect 8899 20012 8944 20040
rect 8938 20000 8944 20012
rect 8996 20000 9002 20052
rect 18598 20040 18604 20052
rect 12406 20012 18604 20040
rect 8202 19972 8208 19984
rect 6472 19944 8208 19972
rect 6472 19913 6500 19944
rect 8202 19932 8208 19944
rect 8260 19932 8266 19984
rect 12406 19972 12434 20012
rect 18598 20000 18604 20012
rect 18656 20000 18662 20052
rect 18693 20043 18751 20049
rect 18693 20009 18705 20043
rect 18739 20040 18751 20043
rect 19242 20040 19248 20052
rect 18739 20012 19248 20040
rect 18739 20009 18751 20012
rect 18693 20003 18751 20009
rect 19242 20000 19248 20012
rect 19300 20040 19306 20052
rect 21450 20040 21456 20052
rect 19300 20012 21456 20040
rect 19300 20000 19306 20012
rect 21450 20000 21456 20012
rect 21508 20000 21514 20052
rect 27706 20040 27712 20052
rect 27667 20012 27712 20040
rect 27706 20000 27712 20012
rect 27764 20000 27770 20052
rect 8312 19944 12434 19972
rect 6457 19907 6515 19913
rect 6457 19873 6469 19907
rect 6503 19873 6515 19907
rect 6638 19904 6644 19916
rect 6599 19876 6644 19904
rect 6457 19867 6515 19873
rect 6638 19864 6644 19876
rect 6696 19864 6702 19916
rect 6914 19904 6920 19916
rect 6875 19876 6920 19904
rect 6914 19864 6920 19876
rect 6972 19864 6978 19916
rect 8312 19836 8340 19944
rect 20530 19932 20536 19984
rect 20588 19972 20594 19984
rect 21085 19975 21143 19981
rect 21085 19972 21097 19975
rect 20588 19944 21097 19972
rect 20588 19932 20594 19944
rect 21085 19941 21097 19944
rect 21131 19941 21143 19975
rect 21085 19935 21143 19941
rect 21174 19932 21180 19984
rect 21232 19972 21238 19984
rect 22186 19972 22192 19984
rect 21232 19944 22192 19972
rect 21232 19932 21238 19944
rect 22186 19932 22192 19944
rect 22244 19972 22250 19984
rect 23569 19975 23627 19981
rect 23569 19972 23581 19975
rect 22244 19944 23581 19972
rect 22244 19932 22250 19944
rect 23569 19941 23581 19944
rect 23615 19941 23627 19975
rect 23569 19935 23627 19941
rect 30742 19932 30748 19984
rect 30800 19972 30806 19984
rect 30800 19944 33088 19972
rect 30800 19932 30806 19944
rect 10137 19907 10195 19913
rect 10137 19873 10149 19907
rect 10183 19904 10195 19907
rect 21634 19904 21640 19916
rect 10183 19876 12434 19904
rect 21595 19876 21640 19904
rect 10183 19873 10195 19876
rect 10137 19867 10195 19873
rect 7852 19808 8340 19836
rect 3970 19728 3976 19780
rect 4028 19768 4034 19780
rect 7852 19768 7880 19808
rect 9030 19796 9036 19848
rect 9088 19836 9094 19848
rect 9171 19839 9229 19845
rect 9171 19836 9183 19839
rect 9088 19808 9183 19836
rect 9088 19796 9094 19808
rect 9171 19805 9183 19808
rect 9217 19805 9229 19839
rect 9306 19836 9312 19848
rect 9267 19808 9312 19836
rect 9171 19799 9229 19805
rect 9306 19796 9312 19808
rect 9364 19796 9370 19848
rect 9398 19796 9404 19848
rect 9456 19833 9462 19848
rect 9585 19839 9643 19845
rect 9456 19805 9498 19833
rect 9585 19805 9597 19839
rect 9631 19836 9643 19839
rect 9766 19836 9772 19848
rect 9631 19808 9772 19836
rect 9631 19805 9643 19808
rect 9456 19796 9462 19805
rect 9585 19799 9643 19805
rect 9766 19796 9772 19808
rect 9824 19836 9830 19848
rect 10226 19836 10232 19848
rect 9824 19808 10232 19836
rect 9824 19796 9830 19808
rect 10226 19796 10232 19808
rect 10284 19836 10290 19848
rect 10413 19839 10471 19845
rect 10413 19836 10425 19839
rect 10284 19808 10425 19836
rect 10284 19796 10290 19808
rect 10413 19805 10425 19808
rect 10459 19805 10471 19839
rect 12406 19836 12434 19876
rect 21634 19864 21640 19876
rect 21692 19864 21698 19916
rect 22278 19864 22284 19916
rect 22336 19904 22342 19916
rect 22557 19907 22615 19913
rect 22557 19904 22569 19907
rect 22336 19876 22569 19904
rect 22336 19864 22342 19876
rect 22557 19873 22569 19876
rect 22603 19873 22615 19907
rect 22557 19867 22615 19873
rect 22741 19907 22799 19913
rect 22741 19873 22753 19907
rect 22787 19904 22799 19907
rect 23750 19904 23756 19916
rect 22787 19876 23756 19904
rect 22787 19873 22799 19876
rect 22741 19867 22799 19873
rect 23750 19864 23756 19876
rect 23808 19864 23814 19916
rect 24578 19864 24584 19916
rect 24636 19904 24642 19916
rect 24765 19907 24823 19913
rect 24765 19904 24777 19907
rect 24636 19876 24777 19904
rect 24636 19864 24642 19876
rect 24765 19873 24777 19876
rect 24811 19873 24823 19907
rect 24765 19867 24823 19873
rect 27430 19864 27436 19916
rect 27488 19864 27494 19916
rect 13630 19836 13636 19848
rect 12406 19808 13636 19836
rect 10413 19799 10471 19805
rect 13630 19796 13636 19808
rect 13688 19796 13694 19848
rect 13814 19796 13820 19848
rect 13872 19836 13878 19848
rect 14277 19839 14335 19845
rect 14277 19836 14289 19839
rect 13872 19808 14289 19836
rect 13872 19796 13878 19808
rect 14277 19805 14289 19808
rect 14323 19805 14335 19839
rect 17310 19836 17316 19848
rect 17271 19808 17316 19836
rect 14277 19799 14335 19805
rect 17310 19796 17316 19808
rect 17368 19796 17374 19848
rect 17586 19845 17592 19848
rect 17580 19836 17592 19845
rect 17547 19808 17592 19836
rect 17580 19799 17592 19808
rect 17586 19796 17592 19799
rect 17644 19796 17650 19848
rect 17862 19796 17868 19848
rect 17920 19836 17926 19848
rect 19245 19839 19303 19845
rect 19245 19836 19257 19839
rect 17920 19808 19257 19836
rect 17920 19796 17926 19808
rect 19245 19805 19257 19808
rect 19291 19805 19303 19839
rect 19245 19799 19303 19805
rect 20346 19796 20352 19848
rect 20404 19836 20410 19848
rect 22465 19839 22523 19845
rect 22465 19836 22477 19839
rect 20404 19808 22477 19836
rect 20404 19796 20410 19808
rect 22465 19805 22477 19808
rect 22511 19805 22523 19839
rect 22465 19799 22523 19805
rect 22649 19839 22707 19845
rect 22649 19805 22661 19839
rect 22695 19836 22707 19839
rect 23014 19836 23020 19848
rect 22695 19808 23020 19836
rect 22695 19805 22707 19808
rect 22649 19799 22707 19805
rect 23014 19796 23020 19808
rect 23072 19796 23078 19848
rect 23385 19839 23443 19845
rect 23385 19805 23397 19839
rect 23431 19836 23443 19839
rect 23474 19836 23480 19848
rect 23431 19808 23480 19836
rect 23431 19805 23443 19808
rect 23385 19799 23443 19805
rect 23474 19796 23480 19808
rect 23532 19836 23538 19848
rect 25041 19839 25099 19845
rect 25041 19836 25053 19839
rect 23532 19808 25053 19836
rect 23532 19796 23538 19808
rect 25041 19805 25053 19808
rect 25087 19805 25099 19839
rect 26418 19836 26424 19848
rect 26379 19808 26424 19836
rect 25041 19799 25099 19805
rect 26418 19796 26424 19808
rect 26476 19796 26482 19848
rect 26694 19836 26700 19848
rect 26655 19808 26700 19836
rect 26694 19796 26700 19808
rect 26752 19796 26758 19848
rect 27157 19839 27215 19845
rect 27157 19805 27169 19839
rect 27203 19836 27215 19839
rect 27448 19836 27476 19864
rect 27203 19808 27476 19836
rect 27525 19839 27583 19845
rect 27203 19805 27215 19808
rect 27157 19799 27215 19805
rect 27525 19805 27537 19839
rect 27571 19836 27583 19839
rect 27614 19836 27620 19848
rect 27571 19808 27620 19836
rect 27571 19805 27583 19808
rect 27525 19799 27583 19805
rect 27614 19796 27620 19808
rect 27672 19796 27678 19848
rect 28718 19796 28724 19848
rect 28776 19836 28782 19848
rect 30285 19839 30343 19845
rect 30285 19836 30297 19839
rect 28776 19808 30297 19836
rect 28776 19796 28782 19808
rect 30285 19805 30297 19808
rect 30331 19805 30343 19839
rect 30285 19799 30343 19805
rect 30374 19796 30380 19848
rect 30432 19836 30438 19848
rect 31956 19845 31984 19944
rect 32306 19904 32312 19916
rect 32140 19876 32312 19904
rect 31803 19839 31861 19845
rect 31803 19836 31815 19839
rect 30432 19808 31815 19836
rect 30432 19796 30438 19808
rect 31803 19805 31815 19808
rect 31849 19805 31861 19839
rect 31803 19799 31861 19805
rect 31941 19839 31999 19845
rect 31941 19805 31953 19839
rect 31987 19805 31999 19839
rect 31941 19799 31999 19805
rect 32033 19839 32091 19845
rect 32033 19805 32045 19839
rect 32079 19836 32091 19839
rect 32140 19836 32168 19876
rect 32306 19864 32312 19876
rect 32364 19864 32370 19916
rect 33060 19845 33088 19944
rect 46290 19904 46296 19916
rect 46251 19876 46296 19904
rect 46290 19864 46296 19876
rect 46348 19864 46354 19916
rect 32079 19808 32168 19836
rect 32217 19839 32275 19845
rect 32079 19805 32091 19808
rect 32033 19799 32091 19805
rect 32217 19805 32229 19839
rect 32263 19805 32275 19839
rect 32217 19799 32275 19805
rect 32953 19839 33011 19845
rect 32953 19805 32965 19839
rect 32999 19805 33011 19839
rect 32953 19799 33011 19805
rect 33045 19839 33103 19845
rect 33045 19805 33057 19839
rect 33091 19805 33103 19839
rect 33045 19799 33103 19805
rect 4028 19740 7880 19768
rect 14093 19771 14151 19777
rect 4028 19728 4034 19740
rect 14093 19737 14105 19771
rect 14139 19768 14151 19771
rect 14366 19768 14372 19780
rect 14139 19740 14372 19768
rect 14139 19737 14151 19740
rect 14093 19731 14151 19737
rect 14366 19728 14372 19740
rect 14424 19728 14430 19780
rect 19512 19771 19570 19777
rect 19512 19737 19524 19771
rect 19558 19768 19570 19771
rect 20898 19768 20904 19780
rect 19558 19740 20904 19768
rect 19558 19737 19570 19740
rect 19512 19731 19570 19737
rect 20898 19728 20904 19740
rect 20956 19728 20962 19780
rect 21545 19771 21603 19777
rect 21545 19768 21557 19771
rect 21008 19740 21557 19768
rect 14461 19703 14519 19709
rect 14461 19669 14473 19703
rect 14507 19700 14519 19703
rect 15102 19700 15108 19712
rect 14507 19672 15108 19700
rect 14507 19669 14519 19672
rect 14461 19663 14519 19669
rect 15102 19660 15108 19672
rect 15160 19660 15166 19712
rect 20622 19700 20628 19712
rect 20583 19672 20628 19700
rect 20622 19660 20628 19672
rect 20680 19700 20686 19712
rect 21008 19700 21036 19740
rect 21545 19737 21557 19740
rect 21591 19737 21603 19771
rect 25866 19768 25872 19780
rect 21545 19731 21603 19737
rect 22066 19740 25872 19768
rect 21450 19700 21456 19712
rect 20680 19672 21036 19700
rect 21363 19672 21456 19700
rect 20680 19660 20686 19672
rect 21450 19660 21456 19672
rect 21508 19700 21514 19712
rect 22066 19700 22094 19740
rect 25866 19728 25872 19740
rect 25924 19728 25930 19780
rect 26237 19771 26295 19777
rect 26237 19737 26249 19771
rect 26283 19768 26295 19771
rect 27341 19771 27399 19777
rect 27341 19768 27353 19771
rect 26283 19740 27353 19768
rect 26283 19737 26295 19740
rect 26237 19731 26295 19737
rect 27341 19737 27353 19740
rect 27387 19737 27399 19771
rect 27341 19731 27399 19737
rect 27433 19771 27491 19777
rect 27433 19737 27445 19771
rect 27479 19768 27491 19771
rect 28994 19768 29000 19780
rect 27479 19740 29000 19768
rect 27479 19737 27491 19740
rect 27433 19731 27491 19737
rect 28994 19728 29000 19740
rect 29052 19728 29058 19780
rect 31478 19768 31484 19780
rect 30622 19740 31484 19768
rect 22278 19700 22284 19712
rect 21508 19672 22094 19700
rect 22239 19672 22284 19700
rect 21508 19660 21514 19672
rect 22278 19660 22284 19672
rect 22336 19660 22342 19712
rect 26605 19703 26663 19709
rect 26605 19669 26617 19703
rect 26651 19700 26663 19703
rect 27522 19700 27528 19712
rect 26651 19672 27528 19700
rect 26651 19669 26663 19672
rect 26605 19663 26663 19669
rect 27522 19660 27528 19672
rect 27580 19660 27586 19712
rect 30515 19703 30573 19709
rect 30515 19669 30527 19703
rect 30561 19700 30573 19703
rect 30622 19700 30650 19740
rect 31478 19728 31484 19740
rect 31536 19768 31542 19780
rect 32232 19768 32260 19799
rect 31536 19740 32812 19768
rect 31536 19728 31542 19740
rect 31570 19700 31576 19712
rect 30561 19672 30650 19700
rect 31531 19672 31576 19700
rect 30561 19669 30573 19672
rect 30515 19663 30573 19669
rect 31570 19660 31576 19672
rect 31628 19660 31634 19712
rect 32674 19700 32680 19712
rect 32635 19672 32680 19700
rect 32674 19660 32680 19672
rect 32732 19660 32738 19712
rect 32784 19700 32812 19740
rect 32858 19728 32864 19780
rect 32916 19768 32922 19780
rect 32968 19768 32996 19799
rect 33134 19796 33140 19848
rect 33192 19836 33198 19848
rect 33321 19839 33379 19845
rect 33192 19808 33237 19836
rect 33192 19796 33198 19808
rect 33321 19805 33333 19839
rect 33367 19805 33379 19839
rect 48130 19836 48136 19848
rect 48091 19808 48136 19836
rect 33321 19799 33379 19805
rect 32916 19740 32996 19768
rect 32916 19728 32922 19740
rect 33336 19700 33364 19799
rect 48130 19796 48136 19808
rect 48188 19796 48194 19848
rect 46477 19771 46535 19777
rect 46477 19737 46489 19771
rect 46523 19768 46535 19771
rect 46934 19768 46940 19780
rect 46523 19740 46940 19768
rect 46523 19737 46535 19740
rect 46477 19731 46535 19737
rect 46934 19728 46940 19740
rect 46992 19728 46998 19780
rect 32784 19672 33364 19700
rect 1104 19610 48852 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 48852 19610
rect 1104 19536 48852 19558
rect 2314 19496 2320 19508
rect 2148 19468 2320 19496
rect 2148 19369 2176 19468
rect 2314 19456 2320 19468
rect 2372 19496 2378 19508
rect 3970 19496 3976 19508
rect 2372 19468 3976 19496
rect 2372 19456 2378 19468
rect 3970 19456 3976 19468
rect 4028 19456 4034 19508
rect 4062 19456 4068 19508
rect 4120 19496 4126 19508
rect 15930 19496 15936 19508
rect 4120 19468 14228 19496
rect 15891 19468 15936 19496
rect 4120 19456 4126 19468
rect 12526 19428 12532 19440
rect 12487 19400 12532 19428
rect 12526 19388 12532 19400
rect 12584 19388 12590 19440
rect 14200 19437 14228 19468
rect 15930 19456 15936 19468
rect 15988 19456 15994 19508
rect 17034 19456 17040 19508
rect 17092 19496 17098 19508
rect 17681 19499 17739 19505
rect 17681 19496 17693 19499
rect 17092 19468 17693 19496
rect 17092 19456 17098 19468
rect 17681 19465 17693 19468
rect 17727 19496 17739 19499
rect 17862 19496 17868 19508
rect 17727 19468 17868 19496
rect 17727 19465 17739 19468
rect 17681 19459 17739 19465
rect 17862 19456 17868 19468
rect 17920 19456 17926 19508
rect 20257 19499 20315 19505
rect 20257 19465 20269 19499
rect 20303 19496 20315 19499
rect 22278 19496 22284 19508
rect 20303 19468 22284 19496
rect 20303 19465 20315 19468
rect 20257 19459 20315 19465
rect 22278 19456 22284 19468
rect 22336 19456 22342 19508
rect 23385 19499 23443 19505
rect 23385 19465 23397 19499
rect 23431 19496 23443 19499
rect 24670 19496 24676 19508
rect 23431 19468 24676 19496
rect 23431 19465 23443 19468
rect 23385 19459 23443 19465
rect 24670 19456 24676 19468
rect 24728 19456 24734 19508
rect 25590 19456 25596 19508
rect 25648 19496 25654 19508
rect 27893 19499 27951 19505
rect 25648 19468 26832 19496
rect 25648 19456 25654 19468
rect 14185 19431 14243 19437
rect 14185 19397 14197 19431
rect 14231 19397 14243 19431
rect 14185 19391 14243 19397
rect 15841 19431 15899 19437
rect 15841 19397 15853 19431
rect 15887 19428 15899 19431
rect 16758 19428 16764 19440
rect 15887 19400 16764 19428
rect 15887 19397 15899 19400
rect 15841 19391 15899 19397
rect 16758 19388 16764 19400
rect 16816 19428 16822 19440
rect 17589 19431 17647 19437
rect 17589 19428 17601 19431
rect 16816 19400 17601 19428
rect 16816 19388 16822 19400
rect 17589 19397 17601 19400
rect 17635 19397 17647 19431
rect 21913 19431 21971 19437
rect 21913 19428 21925 19431
rect 17589 19391 17647 19397
rect 20640 19400 21925 19428
rect 20640 19372 20668 19400
rect 21913 19397 21925 19400
rect 21959 19397 21971 19431
rect 21913 19391 21971 19397
rect 22066 19400 23428 19428
rect 9398 19369 9404 19372
rect 2133 19363 2191 19369
rect 2133 19329 2145 19363
rect 2179 19329 2191 19363
rect 2133 19323 2191 19329
rect 9392 19323 9404 19369
rect 9456 19360 9462 19372
rect 9456 19332 9492 19360
rect 9398 19320 9404 19323
rect 9456 19320 9462 19332
rect 9858 19320 9864 19372
rect 9916 19360 9922 19372
rect 10686 19360 10692 19372
rect 9916 19332 10692 19360
rect 9916 19320 9922 19332
rect 9122 19292 9128 19304
rect 9083 19264 9128 19292
rect 9122 19252 9128 19264
rect 9180 19252 9186 19304
rect 10520 19233 10548 19332
rect 10686 19320 10692 19332
rect 10744 19320 10750 19372
rect 13722 19320 13728 19372
rect 13780 19360 13786 19372
rect 14921 19363 14979 19369
rect 14921 19360 14933 19363
rect 13780 19332 14933 19360
rect 13780 19320 13786 19332
rect 14921 19329 14933 19332
rect 14967 19329 14979 19363
rect 14921 19323 14979 19329
rect 15013 19363 15071 19369
rect 15013 19329 15025 19363
rect 15059 19329 15071 19363
rect 15013 19323 15071 19329
rect 12345 19295 12403 19301
rect 12345 19261 12357 19295
rect 12391 19292 12403 19295
rect 12618 19292 12624 19304
rect 12391 19264 12624 19292
rect 12391 19261 12403 19264
rect 12345 19255 12403 19261
rect 12618 19252 12624 19264
rect 12676 19252 12682 19304
rect 14458 19252 14464 19304
rect 14516 19292 14522 19304
rect 15028 19292 15056 19323
rect 15102 19320 15108 19372
rect 15160 19360 15166 19372
rect 15160 19332 15205 19360
rect 15160 19320 15166 19332
rect 15286 19320 15292 19372
rect 15344 19360 15350 19372
rect 16666 19360 16672 19372
rect 15344 19332 15389 19360
rect 16132 19332 16672 19360
rect 15344 19320 15350 19332
rect 14516 19264 15056 19292
rect 14516 19252 14522 19264
rect 10505 19227 10563 19233
rect 10505 19193 10517 19227
rect 10551 19193 10563 19227
rect 15562 19224 15568 19236
rect 10505 19187 10563 19193
rect 14476 19196 15568 19224
rect 1394 19116 1400 19168
rect 1452 19156 1458 19168
rect 1673 19159 1731 19165
rect 1673 19156 1685 19159
rect 1452 19128 1685 19156
rect 1452 19116 1458 19128
rect 1673 19125 1685 19128
rect 1719 19125 1731 19159
rect 2222 19156 2228 19168
rect 2183 19128 2228 19156
rect 1673 19119 1731 19125
rect 2222 19116 2228 19128
rect 2280 19116 2286 19168
rect 9766 19116 9772 19168
rect 9824 19156 9830 19168
rect 14476 19156 14504 19196
rect 15562 19184 15568 19196
rect 15620 19224 15626 19236
rect 16132 19224 16160 19332
rect 16666 19320 16672 19332
rect 16724 19320 16730 19372
rect 20622 19360 20628 19372
rect 20583 19332 20628 19360
rect 20622 19320 20628 19332
rect 20680 19320 20686 19372
rect 20717 19363 20775 19369
rect 20717 19329 20729 19363
rect 20763 19360 20775 19363
rect 22066 19360 22094 19400
rect 20763 19332 21404 19360
rect 20763 19329 20775 19332
rect 20717 19323 20775 19329
rect 16574 19252 16580 19304
rect 16632 19292 16638 19304
rect 16761 19295 16819 19301
rect 16761 19292 16773 19295
rect 16632 19264 16773 19292
rect 16632 19252 16638 19264
rect 16761 19261 16773 19264
rect 16807 19261 16819 19295
rect 20898 19292 20904 19304
rect 20859 19264 20904 19292
rect 16761 19255 16819 19261
rect 20898 19252 20904 19264
rect 20956 19252 20962 19304
rect 15620 19196 16160 19224
rect 15620 19184 15626 19196
rect 21082 19184 21088 19236
rect 21140 19224 21146 19236
rect 21376 19224 21404 19332
rect 21468 19332 22094 19360
rect 22189 19363 22247 19369
rect 21468 19303 21496 19332
rect 22189 19329 22201 19363
rect 22235 19360 22247 19363
rect 22738 19360 22744 19372
rect 22235 19332 22744 19360
rect 22235 19329 22247 19332
rect 22189 19323 22247 19329
rect 22738 19320 22744 19332
rect 22796 19320 22802 19372
rect 23124 19369 23152 19400
rect 23109 19363 23167 19369
rect 23109 19329 23121 19363
rect 23155 19329 23167 19363
rect 23109 19323 23167 19329
rect 23201 19363 23259 19369
rect 23201 19329 23213 19363
rect 23247 19360 23259 19363
rect 23290 19360 23296 19372
rect 23247 19332 23296 19360
rect 23247 19329 23259 19332
rect 23201 19323 23259 19329
rect 23290 19320 23296 19332
rect 23348 19320 23354 19372
rect 23400 19360 23428 19400
rect 23474 19388 23480 19440
rect 23532 19428 23538 19440
rect 23937 19431 23995 19437
rect 23937 19428 23949 19431
rect 23532 19400 23949 19428
rect 23532 19388 23538 19400
rect 23937 19397 23949 19400
rect 23983 19397 23995 19431
rect 23937 19391 23995 19397
rect 24210 19388 24216 19440
rect 24268 19428 24274 19440
rect 24762 19428 24768 19440
rect 24268 19400 24768 19428
rect 24268 19388 24274 19400
rect 24762 19388 24768 19400
rect 24820 19388 24826 19440
rect 26053 19431 26111 19437
rect 26053 19397 26065 19431
rect 26099 19428 26111 19431
rect 26694 19428 26700 19440
rect 26099 19400 26700 19428
rect 26099 19397 26111 19400
rect 26053 19391 26111 19397
rect 26694 19388 26700 19400
rect 26752 19388 26758 19440
rect 26804 19428 26832 19468
rect 27893 19465 27905 19499
rect 27939 19496 27951 19499
rect 28350 19496 28356 19508
rect 27939 19468 28356 19496
rect 27939 19465 27951 19468
rect 27893 19459 27951 19465
rect 28350 19456 28356 19468
rect 28408 19496 28414 19508
rect 30009 19499 30067 19505
rect 30009 19496 30021 19499
rect 28408 19468 30021 19496
rect 28408 19456 28414 19468
rect 30009 19465 30021 19468
rect 30055 19465 30067 19499
rect 31754 19496 31760 19508
rect 30009 19459 30067 19465
rect 31220 19468 31760 19496
rect 29178 19428 29184 19440
rect 26804 19400 29184 19428
rect 29178 19388 29184 19400
rect 29236 19388 29242 19440
rect 31220 19437 31248 19468
rect 31754 19456 31760 19468
rect 31812 19456 31818 19508
rect 32306 19456 32312 19508
rect 32364 19456 32370 19508
rect 32582 19456 32588 19508
rect 32640 19496 32646 19508
rect 33505 19499 33563 19505
rect 33505 19496 33517 19499
rect 32640 19468 33517 19496
rect 32640 19456 32646 19468
rect 33505 19465 33517 19468
rect 33551 19465 33563 19499
rect 46934 19496 46940 19508
rect 46895 19468 46940 19496
rect 33505 19459 33563 19465
rect 46934 19456 46940 19468
rect 46992 19456 46998 19508
rect 31205 19431 31263 19437
rect 31205 19397 31217 19431
rect 31251 19397 31263 19431
rect 31205 19391 31263 19397
rect 31573 19431 31631 19437
rect 31573 19397 31585 19431
rect 31619 19428 31631 19431
rect 32324 19428 32352 19456
rect 31619 19400 32352 19428
rect 32392 19431 32450 19437
rect 31619 19397 31631 19400
rect 31573 19391 31631 19397
rect 32392 19397 32404 19431
rect 32438 19428 32450 19431
rect 32674 19428 32680 19440
rect 32438 19400 32680 19428
rect 32438 19397 32450 19400
rect 32392 19391 32450 19397
rect 32674 19388 32680 19400
rect 32732 19388 32738 19440
rect 24854 19360 24860 19372
rect 23400 19332 24860 19360
rect 24854 19320 24860 19332
rect 24912 19320 24918 19372
rect 26237 19363 26295 19369
rect 26237 19329 26249 19363
rect 26283 19360 26295 19363
rect 27338 19360 27344 19372
rect 26283 19332 27344 19360
rect 26283 19329 26295 19332
rect 26237 19323 26295 19329
rect 27338 19320 27344 19332
rect 27396 19320 27402 19372
rect 27801 19363 27859 19369
rect 27801 19329 27813 19363
rect 27847 19360 27859 19363
rect 28258 19360 28264 19372
rect 27847 19332 28264 19360
rect 27847 19329 27859 19332
rect 27801 19323 27859 19329
rect 28258 19320 28264 19332
rect 28316 19320 28322 19372
rect 28626 19360 28632 19372
rect 28587 19332 28632 19360
rect 28626 19320 28632 19332
rect 28684 19320 28690 19372
rect 28902 19369 28908 19372
rect 28896 19323 28908 19369
rect 28960 19360 28966 19372
rect 31389 19363 31447 19369
rect 28960 19332 28996 19360
rect 28902 19320 28908 19323
rect 28960 19320 28966 19332
rect 31389 19329 31401 19363
rect 31435 19360 31447 19363
rect 31754 19360 31760 19372
rect 31435 19332 31760 19360
rect 31435 19329 31447 19332
rect 31389 19323 31447 19329
rect 31754 19320 31760 19332
rect 31812 19320 31818 19372
rect 32122 19360 32128 19372
rect 32083 19332 32128 19360
rect 32122 19320 32128 19332
rect 32180 19320 32186 19372
rect 46750 19320 46756 19372
rect 46808 19360 46814 19372
rect 46845 19363 46903 19369
rect 46845 19360 46857 19363
rect 46808 19332 46857 19360
rect 46808 19320 46814 19332
rect 46845 19329 46857 19332
rect 46891 19329 46903 19363
rect 47946 19360 47952 19372
rect 47907 19332 47952 19360
rect 46845 19323 46903 19329
rect 47946 19320 47952 19332
rect 48004 19320 48010 19372
rect 21140 19196 21404 19224
rect 21459 19275 21496 19303
rect 21140 19184 21146 19196
rect 14642 19156 14648 19168
rect 9824 19128 14504 19156
rect 14603 19128 14648 19156
rect 9824 19116 9830 19128
rect 14642 19116 14648 19128
rect 14700 19116 14706 19168
rect 20070 19116 20076 19168
rect 20128 19156 20134 19168
rect 21459 19156 21487 19275
rect 21910 19252 21916 19304
rect 21968 19292 21974 19304
rect 22005 19295 22063 19301
rect 22005 19292 22017 19295
rect 21968 19264 22017 19292
rect 21968 19252 21974 19264
rect 22005 19261 22017 19264
rect 22051 19261 22063 19295
rect 23382 19292 23388 19304
rect 23343 19264 23388 19292
rect 22005 19255 22063 19261
rect 23382 19252 23388 19264
rect 23440 19252 23446 19304
rect 24581 19295 24639 19301
rect 24581 19261 24593 19295
rect 24627 19292 24639 19295
rect 26418 19292 26424 19304
rect 24627 19264 26424 19292
rect 24627 19261 24639 19264
rect 24581 19255 24639 19261
rect 26418 19252 26424 19264
rect 26476 19252 26482 19304
rect 27982 19292 27988 19304
rect 27943 19264 27988 19292
rect 27982 19252 27988 19264
rect 28040 19252 28046 19304
rect 23014 19184 23020 19236
rect 23072 19224 23078 19236
rect 24121 19227 24179 19233
rect 24121 19224 24133 19227
rect 23072 19196 24133 19224
rect 23072 19184 23078 19196
rect 24121 19193 24133 19196
rect 24167 19224 24179 19227
rect 24854 19224 24860 19236
rect 24167 19196 24860 19224
rect 24167 19193 24179 19196
rect 24121 19187 24179 19193
rect 24854 19184 24860 19196
rect 24912 19184 24918 19236
rect 20128 19128 21487 19156
rect 20128 19116 20134 19128
rect 21818 19116 21824 19168
rect 21876 19156 21882 19168
rect 21913 19159 21971 19165
rect 21913 19156 21925 19159
rect 21876 19128 21925 19156
rect 21876 19116 21882 19128
rect 21913 19125 21925 19128
rect 21959 19125 21971 19159
rect 22370 19156 22376 19168
rect 22331 19128 22376 19156
rect 21913 19119 21971 19125
rect 22370 19116 22376 19128
rect 22428 19116 22434 19168
rect 25958 19116 25964 19168
rect 26016 19156 26022 19168
rect 26421 19159 26479 19165
rect 26421 19156 26433 19159
rect 26016 19128 26433 19156
rect 26016 19116 26022 19128
rect 26421 19125 26433 19128
rect 26467 19125 26479 19159
rect 26421 19119 26479 19125
rect 27338 19116 27344 19168
rect 27396 19156 27402 19168
rect 27433 19159 27491 19165
rect 27433 19156 27445 19159
rect 27396 19128 27445 19156
rect 27396 19116 27402 19128
rect 27433 19125 27445 19128
rect 27479 19125 27491 19159
rect 48038 19156 48044 19168
rect 47999 19128 48044 19156
rect 27433 19119 27491 19125
rect 48038 19116 48044 19128
rect 48096 19116 48102 19168
rect 1104 19066 48852 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 48852 19066
rect 1104 18992 48852 19014
rect 9398 18912 9404 18964
rect 9456 18952 9462 18964
rect 9585 18955 9643 18961
rect 9585 18952 9597 18955
rect 9456 18924 9597 18952
rect 9456 18912 9462 18924
rect 9585 18921 9597 18924
rect 9631 18921 9643 18955
rect 12618 18952 12624 18964
rect 12579 18924 12624 18952
rect 9585 18915 9643 18921
rect 12618 18912 12624 18924
rect 12676 18912 12682 18964
rect 20395 18955 20453 18961
rect 20395 18921 20407 18955
rect 20441 18952 20453 18955
rect 20990 18952 20996 18964
rect 20441 18924 20996 18952
rect 20441 18921 20453 18924
rect 20395 18915 20453 18921
rect 20990 18912 20996 18924
rect 21048 18952 21054 18964
rect 21177 18955 21235 18961
rect 21177 18952 21189 18955
rect 21048 18924 21189 18952
rect 21048 18912 21054 18924
rect 21177 18921 21189 18924
rect 21223 18921 21235 18955
rect 25409 18955 25467 18961
rect 25409 18952 25421 18955
rect 21177 18915 21235 18921
rect 21560 18924 25421 18952
rect 14366 18844 14372 18896
rect 14424 18844 14430 18896
rect 20806 18844 20812 18896
rect 20864 18884 20870 18896
rect 21450 18884 21456 18896
rect 20864 18856 21456 18884
rect 20864 18844 20870 18856
rect 21450 18844 21456 18856
rect 21508 18884 21514 18896
rect 21560 18884 21588 18924
rect 25409 18921 25421 18924
rect 25455 18952 25467 18955
rect 25590 18952 25596 18964
rect 25455 18924 25596 18952
rect 25455 18921 25467 18924
rect 25409 18915 25467 18921
rect 25590 18912 25596 18924
rect 25648 18952 25654 18964
rect 25866 18952 25872 18964
rect 25648 18924 25872 18952
rect 25648 18912 25654 18924
rect 25866 18912 25872 18924
rect 25924 18912 25930 18964
rect 26237 18955 26295 18961
rect 26237 18921 26249 18955
rect 26283 18952 26295 18955
rect 26694 18952 26700 18964
rect 26283 18924 26700 18952
rect 26283 18921 26295 18924
rect 26237 18915 26295 18921
rect 26694 18912 26700 18924
rect 26752 18912 26758 18964
rect 26786 18912 26792 18964
rect 26844 18952 26850 18964
rect 27065 18955 27123 18961
rect 27065 18952 27077 18955
rect 26844 18924 27077 18952
rect 26844 18912 26850 18924
rect 27065 18921 27077 18924
rect 27111 18921 27123 18955
rect 27522 18952 27528 18964
rect 27483 18924 27528 18952
rect 27065 18915 27123 18921
rect 27522 18912 27528 18924
rect 27580 18912 27586 18964
rect 28258 18912 28264 18964
rect 28316 18952 28322 18964
rect 28813 18955 28871 18961
rect 28316 18924 28672 18952
rect 28316 18912 28322 18924
rect 21508 18856 21588 18884
rect 21508 18844 21514 18856
rect 21634 18844 21640 18896
rect 21692 18884 21698 18896
rect 21818 18884 21824 18896
rect 21692 18856 21824 18884
rect 21692 18844 21698 18856
rect 21818 18844 21824 18856
rect 21876 18844 21882 18896
rect 23106 18884 23112 18896
rect 22066 18856 23112 18884
rect 1394 18816 1400 18828
rect 1355 18788 1400 18816
rect 1394 18776 1400 18788
rect 1452 18776 1458 18828
rect 1581 18819 1639 18825
rect 1581 18785 1593 18819
rect 1627 18816 1639 18819
rect 2222 18816 2228 18828
rect 1627 18788 2228 18816
rect 1627 18785 1639 18788
rect 1581 18779 1639 18785
rect 2222 18776 2228 18788
rect 2280 18776 2286 18828
rect 2774 18776 2780 18828
rect 2832 18816 2838 18828
rect 2832 18788 2877 18816
rect 2832 18776 2838 18788
rect 9306 18776 9312 18828
rect 9364 18816 9370 18828
rect 12986 18816 12992 18828
rect 9364 18788 9996 18816
rect 9364 18776 9370 18788
rect 9766 18708 9772 18760
rect 9824 18757 9830 18760
rect 9968 18757 9996 18788
rect 12544 18788 12992 18816
rect 9824 18751 9873 18757
rect 9824 18717 9827 18751
rect 9861 18717 9873 18751
rect 9824 18711 9873 18717
rect 9953 18751 10011 18757
rect 9953 18717 9965 18751
rect 9999 18717 10011 18751
rect 9953 18711 10011 18717
rect 10045 18748 10103 18754
rect 10134 18748 10140 18760
rect 10045 18714 10057 18748
rect 10091 18720 10140 18748
rect 10091 18714 10103 18720
rect 9824 18708 9830 18711
rect 10045 18708 10103 18714
rect 10134 18708 10140 18720
rect 10192 18708 10198 18760
rect 10226 18708 10232 18760
rect 10284 18748 10290 18760
rect 11238 18748 11244 18760
rect 10284 18720 10329 18748
rect 11151 18720 11244 18748
rect 10284 18708 10290 18720
rect 11238 18708 11244 18720
rect 11296 18748 11302 18760
rect 12544 18748 12572 18788
rect 12986 18776 12992 18788
rect 13044 18776 13050 18828
rect 14384 18816 14412 18844
rect 13372 18788 14412 18816
rect 11296 18720 12572 18748
rect 11296 18708 11302 18720
rect 12618 18708 12624 18760
rect 12676 18748 12682 18760
rect 13265 18751 13323 18757
rect 13265 18748 13277 18751
rect 12676 18720 13277 18748
rect 12676 18708 12682 18720
rect 13265 18717 13277 18720
rect 13311 18717 13323 18751
rect 13265 18711 13323 18717
rect 11508 18683 11566 18689
rect 11508 18649 11520 18683
rect 11554 18680 11566 18683
rect 13081 18683 13139 18689
rect 11554 18652 13032 18680
rect 11554 18649 11566 18652
rect 11508 18643 11566 18649
rect 13004 18612 13032 18652
rect 13081 18649 13093 18683
rect 13127 18680 13139 18683
rect 13372 18680 13400 18788
rect 16666 18776 16672 18828
rect 16724 18816 16730 18828
rect 20530 18816 20536 18828
rect 16724 18788 17724 18816
rect 20443 18788 20536 18816
rect 16724 18776 16730 18788
rect 13538 18708 13544 18760
rect 13596 18748 13602 18760
rect 14323 18751 14381 18757
rect 14323 18748 14335 18751
rect 13596 18720 14335 18748
rect 13596 18708 13602 18720
rect 14323 18717 14335 18720
rect 14369 18717 14381 18751
rect 14458 18748 14464 18760
rect 14419 18720 14464 18748
rect 14323 18711 14381 18717
rect 14458 18708 14464 18720
rect 14516 18708 14522 18760
rect 14553 18751 14611 18757
rect 14553 18717 14565 18751
rect 14599 18717 14611 18751
rect 14553 18711 14611 18717
rect 14737 18751 14795 18757
rect 14737 18717 14749 18751
rect 14783 18748 14795 18751
rect 15286 18748 15292 18760
rect 14783 18720 15292 18748
rect 14783 18717 14795 18720
rect 14737 18711 14795 18717
rect 13127 18652 13400 18680
rect 13449 18683 13507 18689
rect 13127 18649 13139 18652
rect 13081 18643 13139 18649
rect 13449 18649 13461 18683
rect 13495 18680 13507 18683
rect 14568 18680 14596 18711
rect 15286 18708 15292 18720
rect 15344 18708 15350 18760
rect 15657 18751 15715 18757
rect 15657 18717 15669 18751
rect 15703 18748 15715 18751
rect 17310 18748 17316 18760
rect 15703 18720 17316 18748
rect 15703 18717 15715 18720
rect 15657 18711 15715 18717
rect 17310 18708 17316 18720
rect 17368 18708 17374 18760
rect 17696 18757 17724 18788
rect 20530 18776 20536 18788
rect 20588 18816 20594 18828
rect 21269 18819 21327 18825
rect 21269 18816 21281 18819
rect 20588 18788 21281 18816
rect 20588 18776 20594 18788
rect 21269 18785 21281 18788
rect 21315 18785 21327 18819
rect 21542 18816 21548 18828
rect 21455 18788 21548 18816
rect 21269 18779 21327 18785
rect 17497 18751 17555 18757
rect 17497 18717 17509 18751
rect 17543 18717 17555 18751
rect 17497 18711 17555 18717
rect 17681 18751 17739 18757
rect 17681 18717 17693 18751
rect 17727 18717 17739 18751
rect 17681 18711 17739 18717
rect 13495 18652 14596 18680
rect 15924 18683 15982 18689
rect 13495 18649 13507 18652
rect 13449 18643 13507 18649
rect 15924 18649 15936 18683
rect 15970 18680 15982 18683
rect 16666 18680 16672 18692
rect 15970 18652 16672 18680
rect 15970 18649 15982 18652
rect 15924 18643 15982 18649
rect 16666 18640 16672 18652
rect 16724 18640 16730 18692
rect 17218 18680 17224 18692
rect 17052 18652 17224 18680
rect 17052 18621 17080 18652
rect 17218 18640 17224 18652
rect 17276 18680 17282 18692
rect 17512 18680 17540 18711
rect 20070 18708 20076 18760
rect 20128 18748 20134 18760
rect 21468 18757 21496 18788
rect 21542 18776 21548 18788
rect 21600 18816 21606 18828
rect 22066 18816 22094 18856
rect 23106 18844 23112 18856
rect 23164 18884 23170 18896
rect 26418 18884 26424 18896
rect 23164 18856 26424 18884
rect 23164 18844 23170 18856
rect 26418 18844 26424 18856
rect 26476 18844 26482 18896
rect 27172 18856 28488 18884
rect 26145 18819 26203 18825
rect 21600 18788 22094 18816
rect 23400 18788 24440 18816
rect 21600 18776 21606 18788
rect 23400 18760 23428 18788
rect 20257 18751 20315 18757
rect 20257 18748 20269 18751
rect 20128 18720 20269 18748
rect 20128 18708 20134 18720
rect 20257 18717 20269 18720
rect 20303 18717 20315 18751
rect 20257 18711 20315 18717
rect 20717 18751 20775 18757
rect 20717 18717 20729 18751
rect 20763 18748 20775 18751
rect 21453 18751 21511 18757
rect 20763 18720 21220 18748
rect 20763 18717 20775 18720
rect 20717 18711 20775 18717
rect 21192 18689 21220 18720
rect 21453 18717 21465 18751
rect 21499 18717 21511 18751
rect 21453 18711 21511 18717
rect 21634 18708 21640 18760
rect 21692 18748 21698 18760
rect 22097 18751 22155 18757
rect 22097 18748 22109 18751
rect 21692 18720 22109 18748
rect 21692 18708 21698 18720
rect 22097 18717 22109 18720
rect 22143 18717 22155 18751
rect 23382 18748 23388 18760
rect 23343 18720 23388 18748
rect 22097 18711 22155 18717
rect 23382 18708 23388 18720
rect 23440 18708 23446 18760
rect 23474 18708 23480 18760
rect 23532 18748 23538 18760
rect 24412 18757 24440 18788
rect 26145 18785 26157 18819
rect 26191 18816 26203 18819
rect 26786 18816 26792 18828
rect 26191 18788 26792 18816
rect 26191 18785 26203 18788
rect 26145 18779 26203 18785
rect 26786 18776 26792 18788
rect 26844 18776 26850 18828
rect 24397 18751 24455 18757
rect 23532 18720 23577 18748
rect 23532 18708 23538 18720
rect 24397 18717 24409 18751
rect 24443 18717 24455 18751
rect 24397 18711 24455 18717
rect 24765 18751 24823 18757
rect 24765 18717 24777 18751
rect 24811 18748 24823 18751
rect 25225 18751 25283 18757
rect 25225 18748 25237 18751
rect 24811 18720 25237 18748
rect 24811 18717 24823 18720
rect 24765 18711 24823 18717
rect 25225 18717 25237 18720
rect 25271 18748 25283 18751
rect 25958 18748 25964 18760
rect 25271 18720 25452 18748
rect 25919 18720 25964 18748
rect 25271 18717 25283 18720
rect 25225 18711 25283 18717
rect 17276 18652 17540 18680
rect 21177 18683 21235 18689
rect 17276 18640 17282 18652
rect 21177 18649 21189 18683
rect 21223 18680 21235 18683
rect 22189 18683 22247 18689
rect 22189 18680 22201 18683
rect 21223 18652 22201 18680
rect 21223 18649 21235 18652
rect 21177 18643 21235 18649
rect 22189 18649 22201 18652
rect 22235 18649 22247 18683
rect 22189 18643 22247 18649
rect 23661 18683 23719 18689
rect 23661 18649 23673 18683
rect 23707 18649 23719 18683
rect 23661 18643 23719 18649
rect 24581 18683 24639 18689
rect 24581 18649 24593 18683
rect 24627 18680 24639 18683
rect 25314 18680 25320 18692
rect 24627 18652 25320 18680
rect 24627 18649 24639 18652
rect 24581 18643 24639 18649
rect 14093 18615 14151 18621
rect 14093 18612 14105 18615
rect 13004 18584 14105 18612
rect 14093 18581 14105 18584
rect 14139 18581 14151 18615
rect 14093 18575 14151 18581
rect 17037 18615 17095 18621
rect 17037 18581 17049 18615
rect 17083 18581 17095 18615
rect 17037 18575 17095 18581
rect 17681 18615 17739 18621
rect 17681 18581 17693 18615
rect 17727 18612 17739 18615
rect 17770 18612 17776 18624
rect 17727 18584 17776 18612
rect 17727 18581 17739 18584
rect 17681 18575 17739 18581
rect 17770 18572 17776 18584
rect 17828 18572 17834 18624
rect 20717 18615 20775 18621
rect 20717 18581 20729 18615
rect 20763 18612 20775 18615
rect 21542 18612 21548 18624
rect 20763 18584 21548 18612
rect 20763 18581 20775 18584
rect 20717 18575 20775 18581
rect 21542 18572 21548 18584
rect 21600 18572 21606 18624
rect 21637 18615 21695 18621
rect 21637 18581 21649 18615
rect 21683 18612 21695 18615
rect 22094 18612 22100 18624
rect 21683 18584 22100 18612
rect 21683 18581 21695 18584
rect 21637 18575 21695 18581
rect 22094 18572 22100 18584
rect 22152 18572 22158 18624
rect 23676 18612 23704 18643
rect 25314 18640 25320 18652
rect 25372 18640 25378 18692
rect 25424 18680 25452 18720
rect 25958 18708 25964 18720
rect 26016 18708 26022 18760
rect 26237 18751 26295 18757
rect 26237 18717 26249 18751
rect 26283 18748 26295 18751
rect 26878 18748 26884 18760
rect 26283 18720 26884 18748
rect 26283 18717 26295 18720
rect 26237 18711 26295 18717
rect 26878 18708 26884 18720
rect 26936 18708 26942 18760
rect 26973 18751 27031 18757
rect 26973 18717 26985 18751
rect 27019 18748 27031 18751
rect 27062 18748 27068 18760
rect 27019 18720 27068 18748
rect 27019 18717 27031 18720
rect 26973 18711 27031 18717
rect 27062 18708 27068 18720
rect 27120 18708 27126 18760
rect 26142 18680 26148 18692
rect 25424 18652 26148 18680
rect 26142 18640 26148 18652
rect 26200 18640 26206 18692
rect 24670 18612 24676 18624
rect 23676 18584 24676 18612
rect 24670 18572 24676 18584
rect 24728 18572 24734 18624
rect 25682 18572 25688 18624
rect 25740 18612 25746 18624
rect 27172 18612 27200 18856
rect 28350 18816 28356 18828
rect 28311 18788 28356 18816
rect 28350 18776 28356 18788
rect 28408 18776 28414 18828
rect 28460 18825 28488 18856
rect 28445 18819 28503 18825
rect 28445 18785 28457 18819
rect 28491 18785 28503 18819
rect 28445 18779 28503 18785
rect 27338 18748 27344 18760
rect 27299 18720 27344 18748
rect 27338 18708 27344 18720
rect 27396 18708 27402 18760
rect 27798 18708 27804 18760
rect 27856 18748 27862 18760
rect 28077 18751 28135 18757
rect 28077 18748 28089 18751
rect 27856 18720 28089 18748
rect 27856 18708 27862 18720
rect 28077 18717 28089 18720
rect 28123 18717 28135 18751
rect 28258 18748 28264 18760
rect 28219 18720 28264 18748
rect 28077 18711 28135 18717
rect 28258 18708 28264 18720
rect 28316 18708 28322 18760
rect 28644 18757 28672 18924
rect 28813 18921 28825 18955
rect 28859 18952 28871 18955
rect 28902 18952 28908 18964
rect 28859 18924 28908 18952
rect 28859 18921 28871 18924
rect 28813 18915 28871 18921
rect 28902 18912 28908 18924
rect 28960 18912 28966 18964
rect 28629 18751 28687 18757
rect 28629 18717 28641 18751
rect 28675 18717 28687 18751
rect 28629 18711 28687 18717
rect 28718 18708 28724 18760
rect 28776 18748 28782 18760
rect 30837 18751 30895 18757
rect 30837 18748 30849 18751
rect 28776 18720 30849 18748
rect 28776 18708 28782 18720
rect 30837 18717 30849 18720
rect 30883 18717 30895 18751
rect 30837 18711 30895 18717
rect 31104 18751 31162 18757
rect 31104 18717 31116 18751
rect 31150 18748 31162 18751
rect 31570 18748 31576 18760
rect 31150 18720 31576 18748
rect 31150 18717 31162 18720
rect 31104 18711 31162 18717
rect 31570 18708 31576 18720
rect 31628 18708 31634 18760
rect 25740 18584 27200 18612
rect 25740 18572 25746 18584
rect 31754 18572 31760 18624
rect 31812 18612 31818 18624
rect 32217 18615 32275 18621
rect 32217 18612 32229 18615
rect 31812 18584 32229 18612
rect 31812 18572 31818 18584
rect 32217 18581 32229 18584
rect 32263 18581 32275 18615
rect 32217 18575 32275 18581
rect 1104 18522 48852 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 48852 18522
rect 1104 18448 48852 18470
rect 13814 18368 13820 18420
rect 13872 18408 13878 18420
rect 14185 18411 14243 18417
rect 14185 18408 14197 18411
rect 13872 18380 14197 18408
rect 13872 18368 13878 18380
rect 14185 18377 14197 18380
rect 14231 18377 14243 18411
rect 16666 18408 16672 18420
rect 16627 18380 16672 18408
rect 14185 18371 14243 18377
rect 16666 18368 16672 18380
rect 16724 18368 16730 18420
rect 17770 18408 17776 18420
rect 17731 18380 17776 18408
rect 17770 18368 17776 18380
rect 17828 18368 17834 18420
rect 20533 18411 20591 18417
rect 20533 18377 20545 18411
rect 20579 18408 20591 18411
rect 21634 18408 21640 18420
rect 20579 18380 21640 18408
rect 20579 18377 20591 18380
rect 20533 18371 20591 18377
rect 21634 18368 21640 18380
rect 21692 18368 21698 18420
rect 21818 18368 21824 18420
rect 21876 18408 21882 18420
rect 21876 18380 22968 18408
rect 21876 18368 21882 18380
rect 12986 18300 12992 18352
rect 13044 18300 13050 18352
rect 14366 18300 14372 18352
rect 14424 18340 14430 18352
rect 15749 18343 15807 18349
rect 15749 18340 15761 18343
rect 14424 18312 15761 18340
rect 14424 18300 14430 18312
rect 15749 18309 15761 18312
rect 15795 18309 15807 18343
rect 15749 18303 15807 18309
rect 15933 18343 15991 18349
rect 15933 18309 15945 18343
rect 15979 18340 15991 18343
rect 16022 18340 16028 18352
rect 15979 18312 16028 18340
rect 15979 18309 15991 18312
rect 15933 18303 15991 18309
rect 16022 18300 16028 18312
rect 16080 18300 16086 18352
rect 16574 18300 16580 18352
rect 16632 18340 16638 18352
rect 17037 18343 17095 18349
rect 17037 18340 17049 18343
rect 16632 18312 17049 18340
rect 16632 18300 16638 18312
rect 17037 18309 17049 18312
rect 17083 18309 17095 18343
rect 17037 18303 17095 18309
rect 17589 18343 17647 18349
rect 17589 18309 17601 18343
rect 17635 18340 17647 18343
rect 20346 18340 20352 18352
rect 17635 18312 20352 18340
rect 17635 18309 17647 18312
rect 17589 18303 17647 18309
rect 20346 18300 20352 18312
rect 20404 18300 20410 18352
rect 20990 18340 20996 18352
rect 20903 18312 20996 18340
rect 20990 18300 20996 18312
rect 21048 18340 21054 18352
rect 21910 18340 21916 18352
rect 21048 18312 21916 18340
rect 21048 18300 21054 18312
rect 21910 18300 21916 18312
rect 21968 18300 21974 18352
rect 12805 18275 12863 18281
rect 12805 18241 12817 18275
rect 12851 18272 12863 18275
rect 13004 18272 13032 18300
rect 12851 18244 13032 18272
rect 13072 18275 13130 18281
rect 12851 18241 12863 18244
rect 12805 18235 12863 18241
rect 13072 18241 13084 18275
rect 13118 18272 13130 18275
rect 14642 18272 14648 18284
rect 13118 18244 14648 18272
rect 13118 18241 13130 18244
rect 13072 18235 13130 18241
rect 14642 18232 14648 18244
rect 14700 18232 14706 18284
rect 14918 18281 14924 18284
rect 14901 18275 14924 18281
rect 14901 18241 14913 18275
rect 14901 18235 14924 18241
rect 14918 18232 14924 18235
rect 14976 18232 14982 18284
rect 15013 18275 15071 18281
rect 15013 18241 15025 18275
rect 15059 18241 15071 18275
rect 15013 18235 15071 18241
rect 15105 18275 15163 18281
rect 15105 18241 15117 18275
rect 15151 18241 15163 18275
rect 15286 18272 15292 18284
rect 15247 18244 15292 18272
rect 15105 18235 15163 18241
rect 1765 18207 1823 18213
rect 1765 18173 1777 18207
rect 1811 18173 1823 18207
rect 1946 18204 1952 18216
rect 1907 18176 1952 18204
rect 1765 18167 1823 18173
rect 1780 18068 1808 18167
rect 1946 18164 1952 18176
rect 2004 18164 2010 18216
rect 2774 18164 2780 18216
rect 2832 18204 2838 18216
rect 2832 18176 2877 18204
rect 2832 18164 2838 18176
rect 14458 18164 14464 18216
rect 14516 18204 14522 18216
rect 15028 18204 15056 18235
rect 14516 18176 15056 18204
rect 15120 18204 15148 18235
rect 15286 18232 15292 18244
rect 15344 18232 15350 18284
rect 15838 18232 15844 18284
rect 15896 18272 15902 18284
rect 16853 18275 16911 18281
rect 16853 18272 16865 18275
rect 15896 18244 16865 18272
rect 15896 18232 15902 18244
rect 16853 18241 16865 18244
rect 16899 18241 16911 18275
rect 16853 18235 16911 18241
rect 17129 18275 17187 18281
rect 17129 18241 17141 18275
rect 17175 18272 17187 18275
rect 17218 18272 17224 18284
rect 17175 18244 17224 18272
rect 17175 18241 17187 18244
rect 17129 18235 17187 18241
rect 16117 18207 16175 18213
rect 16117 18204 16129 18207
rect 15120 18176 16129 18204
rect 14516 18164 14522 18176
rect 16117 18173 16129 18176
rect 16163 18173 16175 18207
rect 16868 18204 16896 18235
rect 17218 18232 17224 18244
rect 17276 18232 17282 18284
rect 17865 18275 17923 18281
rect 17865 18241 17877 18275
rect 17911 18272 17923 18275
rect 18506 18272 18512 18284
rect 17911 18244 18512 18272
rect 17911 18241 17923 18244
rect 17865 18235 17923 18241
rect 18506 18232 18512 18244
rect 18564 18232 18570 18284
rect 18598 18232 18604 18284
rect 18656 18272 18662 18284
rect 20714 18272 20720 18284
rect 18656 18244 18701 18272
rect 19444 18244 20720 18272
rect 18656 18232 18662 18244
rect 16868 18176 17264 18204
rect 16117 18167 16175 18173
rect 17236 18148 17264 18176
rect 17402 18164 17408 18216
rect 17460 18204 17466 18216
rect 19444 18204 19472 18244
rect 20714 18232 20720 18244
rect 20772 18272 20778 18284
rect 20898 18272 20904 18284
rect 20772 18244 20904 18272
rect 20772 18232 20778 18244
rect 20898 18232 20904 18244
rect 20956 18232 20962 18284
rect 21818 18272 21824 18284
rect 21192 18244 21824 18272
rect 21192 18213 21220 18244
rect 21818 18232 21824 18244
rect 21876 18232 21882 18284
rect 22094 18232 22100 18284
rect 22152 18272 22158 18284
rect 22940 18272 22968 18380
rect 23658 18368 23664 18420
rect 23716 18408 23722 18420
rect 24210 18408 24216 18420
rect 23716 18380 24216 18408
rect 23716 18368 23722 18380
rect 24210 18368 24216 18380
rect 24268 18368 24274 18420
rect 25130 18368 25136 18420
rect 25188 18408 25194 18420
rect 25777 18411 25835 18417
rect 25777 18408 25789 18411
rect 25188 18380 25789 18408
rect 25188 18368 25194 18380
rect 25777 18377 25789 18380
rect 25823 18408 25835 18411
rect 27798 18408 27804 18420
rect 25823 18380 27660 18408
rect 27759 18380 27804 18408
rect 25823 18377 25835 18380
rect 25777 18371 25835 18377
rect 23014 18300 23020 18352
rect 23072 18340 23078 18352
rect 23293 18343 23351 18349
rect 23293 18340 23305 18343
rect 23072 18312 23305 18340
rect 23072 18300 23078 18312
rect 23293 18309 23305 18312
rect 23339 18340 23351 18343
rect 24026 18340 24032 18352
rect 23339 18312 24032 18340
rect 23339 18309 23351 18312
rect 23293 18303 23351 18309
rect 24026 18300 24032 18312
rect 24084 18300 24090 18352
rect 25685 18343 25743 18349
rect 25685 18309 25697 18343
rect 25731 18340 25743 18343
rect 26142 18340 26148 18352
rect 25731 18312 26148 18340
rect 25731 18309 25743 18312
rect 25685 18303 25743 18309
rect 26142 18300 26148 18312
rect 26200 18300 26206 18352
rect 27522 18340 27528 18352
rect 27264 18312 27528 18340
rect 23109 18275 23167 18281
rect 23109 18272 23121 18275
rect 22152 18244 22197 18272
rect 22940 18244 23121 18272
rect 22152 18232 22158 18244
rect 23109 18241 23121 18244
rect 23155 18272 23167 18275
rect 24118 18272 24124 18284
rect 23155 18244 24124 18272
rect 23155 18241 23167 18244
rect 23109 18235 23167 18241
rect 24118 18232 24124 18244
rect 24176 18232 24182 18284
rect 24949 18275 25007 18281
rect 24949 18241 24961 18275
rect 24995 18272 25007 18275
rect 25314 18272 25320 18284
rect 24995 18244 25320 18272
rect 24995 18241 25007 18244
rect 24949 18235 25007 18241
rect 25314 18232 25320 18244
rect 25372 18232 25378 18284
rect 27264 18281 27292 18312
rect 27522 18300 27528 18312
rect 27580 18300 27586 18352
rect 27632 18340 27660 18380
rect 27798 18368 27804 18380
rect 27856 18368 27862 18420
rect 28258 18340 28264 18352
rect 27632 18312 28264 18340
rect 28258 18300 28264 18312
rect 28316 18300 28322 18352
rect 28350 18300 28356 18352
rect 28408 18340 28414 18352
rect 28629 18343 28687 18349
rect 28629 18340 28641 18343
rect 28408 18312 28641 18340
rect 28408 18300 28414 18312
rect 28629 18309 28641 18312
rect 28675 18309 28687 18343
rect 28629 18303 28687 18309
rect 27249 18275 27307 18281
rect 27249 18241 27261 18275
rect 27295 18241 27307 18275
rect 27249 18235 27307 18241
rect 28534 18232 28540 18284
rect 28592 18272 28598 18284
rect 28905 18275 28963 18281
rect 28905 18272 28917 18275
rect 28592 18244 28917 18272
rect 28592 18232 28598 18244
rect 28905 18241 28917 18244
rect 28951 18241 28963 18275
rect 28905 18235 28963 18241
rect 34330 18232 34336 18284
rect 34388 18272 34394 18284
rect 34388 18244 34560 18272
rect 34388 18232 34394 18244
rect 17460 18176 19472 18204
rect 21177 18207 21235 18213
rect 17460 18164 17466 18176
rect 21177 18173 21189 18207
rect 21223 18173 21235 18207
rect 21177 18167 21235 18173
rect 21542 18164 21548 18216
rect 21600 18204 21606 18216
rect 22005 18207 22063 18213
rect 22005 18204 22017 18207
rect 21600 18176 22017 18204
rect 21600 18164 21606 18176
rect 22005 18173 22017 18176
rect 22051 18173 22063 18207
rect 22005 18167 22063 18173
rect 22189 18207 22247 18213
rect 22189 18173 22201 18207
rect 22235 18173 22247 18207
rect 22189 18167 22247 18173
rect 4062 18096 4068 18148
rect 4120 18136 4126 18148
rect 8294 18136 8300 18148
rect 4120 18108 8300 18136
rect 4120 18096 4126 18108
rect 8294 18096 8300 18108
rect 8352 18096 8358 18148
rect 17218 18096 17224 18148
rect 17276 18096 17282 18148
rect 22204 18136 22232 18167
rect 22278 18164 22284 18216
rect 22336 18204 22342 18216
rect 24210 18204 24216 18216
rect 22336 18176 22381 18204
rect 22480 18176 24216 18204
rect 22336 18164 22342 18176
rect 22480 18136 22508 18176
rect 24210 18164 24216 18176
rect 24268 18164 24274 18216
rect 24670 18164 24676 18216
rect 24728 18204 24734 18216
rect 26142 18204 26148 18216
rect 24728 18176 26148 18204
rect 24728 18164 24734 18176
rect 26142 18164 26148 18176
rect 26200 18204 26206 18216
rect 27525 18207 27583 18213
rect 27525 18204 27537 18207
rect 26200 18176 27537 18204
rect 26200 18164 26206 18176
rect 27525 18173 27537 18176
rect 27571 18173 27583 18207
rect 27525 18167 27583 18173
rect 28813 18207 28871 18213
rect 28813 18173 28825 18207
rect 28859 18204 28871 18207
rect 28994 18204 29000 18216
rect 28859 18176 29000 18204
rect 28859 18173 28871 18176
rect 28813 18167 28871 18173
rect 28994 18164 29000 18176
rect 29052 18164 29058 18216
rect 32858 18204 32864 18216
rect 32819 18176 32864 18204
rect 32858 18164 32864 18176
rect 32916 18164 32922 18216
rect 33045 18207 33103 18213
rect 33045 18173 33057 18207
rect 33091 18204 33103 18207
rect 34422 18204 34428 18216
rect 33091 18176 34428 18204
rect 33091 18173 33103 18176
rect 33045 18167 33103 18173
rect 34422 18164 34428 18176
rect 34480 18164 34486 18216
rect 34532 18213 34560 18244
rect 34517 18207 34575 18213
rect 34517 18173 34529 18207
rect 34563 18173 34575 18207
rect 34517 18167 34575 18173
rect 22204 18108 22508 18136
rect 23290 18096 23296 18148
rect 23348 18136 23354 18148
rect 25133 18139 25191 18145
rect 25133 18136 25145 18139
rect 23348 18108 25145 18136
rect 23348 18096 23354 18108
rect 25133 18105 25145 18108
rect 25179 18136 25191 18139
rect 25590 18136 25596 18148
rect 25179 18108 25596 18136
rect 25179 18105 25191 18108
rect 25133 18099 25191 18105
rect 25590 18096 25596 18108
rect 25648 18096 25654 18148
rect 29089 18139 29147 18145
rect 29089 18136 29101 18139
rect 25700 18108 29101 18136
rect 4249 18071 4307 18077
rect 4249 18068 4261 18071
rect 1780 18040 4261 18068
rect 4249 18037 4261 18040
rect 4295 18037 4307 18071
rect 4249 18031 4307 18037
rect 14645 18071 14703 18077
rect 14645 18037 14657 18071
rect 14691 18068 14703 18071
rect 14918 18068 14924 18080
rect 14691 18040 14924 18068
rect 14691 18037 14703 18040
rect 14645 18031 14703 18037
rect 14918 18028 14924 18040
rect 14976 18028 14982 18080
rect 17494 18028 17500 18080
rect 17552 18068 17558 18080
rect 17589 18071 17647 18077
rect 17589 18068 17601 18071
rect 17552 18040 17601 18068
rect 17552 18028 17558 18040
rect 17589 18037 17601 18040
rect 17635 18037 17647 18071
rect 18690 18068 18696 18080
rect 18651 18040 18696 18068
rect 17589 18031 17647 18037
rect 18690 18028 18696 18040
rect 18748 18028 18754 18080
rect 20714 18028 20720 18080
rect 20772 18068 20778 18080
rect 21821 18071 21879 18077
rect 21821 18068 21833 18071
rect 20772 18040 21833 18068
rect 20772 18028 20778 18040
rect 21821 18037 21833 18040
rect 21867 18037 21879 18071
rect 21821 18031 21879 18037
rect 22186 18028 22192 18080
rect 22244 18068 22250 18080
rect 23106 18068 23112 18080
rect 22244 18040 23112 18068
rect 22244 18028 22250 18040
rect 23106 18028 23112 18040
rect 23164 18068 23170 18080
rect 23382 18068 23388 18080
rect 23164 18040 23388 18068
rect 23164 18028 23170 18040
rect 23382 18028 23388 18040
rect 23440 18068 23446 18080
rect 23477 18071 23535 18077
rect 23477 18068 23489 18071
rect 23440 18040 23489 18068
rect 23440 18028 23446 18040
rect 23477 18037 23489 18040
rect 23523 18037 23535 18071
rect 23477 18031 23535 18037
rect 23566 18028 23572 18080
rect 23624 18068 23630 18080
rect 23937 18071 23995 18077
rect 23937 18068 23949 18071
rect 23624 18040 23949 18068
rect 23624 18028 23630 18040
rect 23937 18037 23949 18040
rect 23983 18037 23995 18071
rect 23937 18031 23995 18037
rect 24026 18028 24032 18080
rect 24084 18068 24090 18080
rect 25700 18068 25728 18108
rect 29089 18105 29101 18108
rect 29135 18105 29147 18139
rect 29089 18099 29147 18105
rect 27614 18068 27620 18080
rect 24084 18040 25728 18068
rect 27575 18040 27620 18068
rect 24084 18028 24090 18040
rect 27614 18028 27620 18040
rect 27672 18028 27678 18080
rect 28718 18068 28724 18080
rect 28679 18040 28724 18068
rect 28718 18028 28724 18040
rect 28776 18028 28782 18080
rect 1104 17978 48852 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 48852 17978
rect 1104 17904 48852 17926
rect 1946 17824 1952 17876
rect 2004 17864 2010 17876
rect 2133 17867 2191 17873
rect 2133 17864 2145 17867
rect 2004 17836 2145 17864
rect 2004 17824 2010 17836
rect 2133 17833 2145 17836
rect 2179 17833 2191 17867
rect 2133 17827 2191 17833
rect 2746 17836 12434 17864
rect 2746 17728 2774 17836
rect 8294 17796 8300 17808
rect 8255 17768 8300 17796
rect 8294 17756 8300 17768
rect 8352 17756 8358 17808
rect 12406 17796 12434 17836
rect 13722 17824 13728 17876
rect 13780 17864 13786 17876
rect 16022 17864 16028 17876
rect 13780 17836 15700 17864
rect 15983 17836 16028 17864
rect 13780 17824 13786 17836
rect 14642 17796 14648 17808
rect 12406 17768 14648 17796
rect 14642 17756 14648 17768
rect 14700 17756 14706 17808
rect 2056 17700 2774 17728
rect 7745 17731 7803 17737
rect 2056 17672 2084 17700
rect 7745 17697 7757 17731
rect 7791 17728 7803 17731
rect 9122 17728 9128 17740
rect 7791 17700 9128 17728
rect 7791 17697 7803 17700
rect 7745 17691 7803 17697
rect 9122 17688 9128 17700
rect 9180 17728 9186 17740
rect 11238 17728 11244 17740
rect 9180 17700 11244 17728
rect 9180 17688 9186 17700
rect 11238 17688 11244 17700
rect 11296 17688 11302 17740
rect 11330 17688 11336 17740
rect 11388 17728 11394 17740
rect 12713 17731 12771 17737
rect 11388 17700 11433 17728
rect 11388 17688 11394 17700
rect 12713 17697 12725 17731
rect 12759 17728 12771 17731
rect 12802 17728 12808 17740
rect 12759 17700 12808 17728
rect 12759 17697 12771 17700
rect 12713 17691 12771 17697
rect 12802 17688 12808 17700
rect 12860 17688 12866 17740
rect 14458 17728 14464 17740
rect 13004 17700 14464 17728
rect 1581 17663 1639 17669
rect 1581 17629 1593 17663
rect 1627 17660 1639 17663
rect 1762 17660 1768 17672
rect 1627 17632 1768 17660
rect 1627 17629 1639 17632
rect 1581 17623 1639 17629
rect 1762 17620 1768 17632
rect 1820 17620 1826 17672
rect 2038 17660 2044 17672
rect 1951 17632 2044 17660
rect 2038 17620 2044 17632
rect 2096 17620 2102 17672
rect 2590 17620 2596 17672
rect 2648 17660 2654 17672
rect 2685 17663 2743 17669
rect 2685 17660 2697 17663
rect 2648 17632 2697 17660
rect 2648 17620 2654 17632
rect 2685 17629 2697 17632
rect 2731 17629 2743 17663
rect 9858 17660 9864 17672
rect 9819 17632 9864 17660
rect 2685 17623 2743 17629
rect 9858 17620 9864 17632
rect 9916 17620 9922 17672
rect 11974 17620 11980 17672
rect 12032 17660 12038 17672
rect 13004 17669 13032 17700
rect 14458 17688 14464 17700
rect 14516 17688 14522 17740
rect 15672 17728 15700 17836
rect 16022 17824 16028 17836
rect 16080 17824 16086 17876
rect 16114 17824 16120 17876
rect 16172 17864 16178 17876
rect 19429 17867 19487 17873
rect 19429 17864 19441 17867
rect 16172 17836 19441 17864
rect 16172 17824 16178 17836
rect 19429 17833 19441 17836
rect 19475 17833 19487 17867
rect 19429 17827 19487 17833
rect 21177 17867 21235 17873
rect 21177 17833 21189 17867
rect 21223 17864 21235 17867
rect 22278 17864 22284 17876
rect 21223 17836 22284 17864
rect 21223 17833 21235 17836
rect 21177 17827 21235 17833
rect 22278 17824 22284 17836
rect 22336 17824 22342 17876
rect 23385 17867 23443 17873
rect 23385 17833 23397 17867
rect 23431 17864 23443 17867
rect 23474 17864 23480 17876
rect 23431 17836 23480 17864
rect 23431 17833 23443 17836
rect 23385 17827 23443 17833
rect 23474 17824 23480 17836
rect 23532 17824 23538 17876
rect 24581 17867 24639 17873
rect 24581 17864 24593 17867
rect 23584 17836 24593 17864
rect 16758 17796 16764 17808
rect 16719 17768 16764 17796
rect 16758 17756 16764 17768
rect 16816 17756 16822 17808
rect 18601 17799 18659 17805
rect 18601 17765 18613 17799
rect 18647 17796 18659 17799
rect 23014 17796 23020 17808
rect 18647 17768 23020 17796
rect 18647 17765 18659 17768
rect 18601 17759 18659 17765
rect 17034 17728 17040 17740
rect 15672 17700 17040 17728
rect 17034 17688 17040 17700
rect 17092 17688 17098 17740
rect 12989 17663 13047 17669
rect 12989 17660 13001 17663
rect 12032 17632 13001 17660
rect 12032 17620 12038 17632
rect 12989 17629 13001 17632
rect 13035 17629 13047 17663
rect 12989 17623 13047 17629
rect 14366 17620 14372 17672
rect 14424 17660 14430 17672
rect 14645 17663 14703 17669
rect 14645 17660 14657 17663
rect 14424 17632 14657 17660
rect 14424 17620 14430 17632
rect 14645 17629 14657 17632
rect 14691 17660 14703 17663
rect 17221 17663 17279 17669
rect 17221 17660 17233 17663
rect 14691 17632 17233 17660
rect 14691 17629 14703 17632
rect 14645 17623 14703 17629
rect 17221 17629 17233 17632
rect 17267 17660 17279 17663
rect 17310 17660 17316 17672
rect 17267 17632 17316 17660
rect 17267 17629 17279 17632
rect 17221 17623 17279 17629
rect 17310 17620 17316 17632
rect 17368 17620 17374 17672
rect 17494 17669 17500 17672
rect 17488 17660 17500 17669
rect 17455 17632 17500 17660
rect 17488 17623 17500 17632
rect 17494 17620 17500 17623
rect 17552 17620 17558 17672
rect 19352 17669 19380 17768
rect 23014 17756 23020 17768
rect 23072 17756 23078 17808
rect 23106 17756 23112 17808
rect 23164 17796 23170 17808
rect 23584 17796 23612 17836
rect 24581 17833 24593 17836
rect 24627 17833 24639 17867
rect 24581 17827 24639 17833
rect 24762 17824 24768 17876
rect 24820 17864 24826 17876
rect 25130 17864 25136 17876
rect 24820 17836 25136 17864
rect 24820 17824 24826 17836
rect 25130 17824 25136 17836
rect 25188 17824 25194 17876
rect 25314 17864 25320 17876
rect 25275 17836 25320 17864
rect 25314 17824 25320 17836
rect 25372 17824 25378 17876
rect 26694 17824 26700 17876
rect 26752 17864 26758 17876
rect 26789 17867 26847 17873
rect 26789 17864 26801 17867
rect 26752 17836 26801 17864
rect 26752 17824 26758 17836
rect 26789 17833 26801 17836
rect 26835 17833 26847 17867
rect 26789 17827 26847 17833
rect 27614 17824 27620 17876
rect 27672 17864 27678 17876
rect 27985 17867 28043 17873
rect 27985 17864 27997 17867
rect 27672 17836 27997 17864
rect 27672 17824 27678 17836
rect 27985 17833 27997 17836
rect 28031 17833 28043 17867
rect 27985 17827 28043 17833
rect 34422 17824 34428 17876
rect 34480 17864 34486 17876
rect 34793 17867 34851 17873
rect 34793 17864 34805 17867
rect 34480 17836 34805 17864
rect 34480 17824 34486 17836
rect 34793 17833 34805 17836
rect 34839 17833 34851 17867
rect 34793 17827 34851 17833
rect 27157 17799 27215 17805
rect 23164 17768 23612 17796
rect 24044 17768 27108 17796
rect 23164 17756 23170 17768
rect 20070 17688 20076 17740
rect 20128 17728 20134 17740
rect 24044 17728 24072 17768
rect 20128 17700 24072 17728
rect 20128 17688 20134 17700
rect 24118 17688 24124 17740
rect 24176 17728 24182 17740
rect 24176 17700 24521 17728
rect 24176 17688 24182 17700
rect 19337 17663 19395 17669
rect 19337 17629 19349 17663
rect 19383 17629 19395 17663
rect 19337 17623 19395 17629
rect 21361 17663 21419 17669
rect 21361 17629 21373 17663
rect 21407 17629 21419 17663
rect 21634 17660 21640 17672
rect 21595 17632 21640 17660
rect 21361 17623 21419 17629
rect 7837 17595 7895 17601
rect 7837 17561 7849 17595
rect 7883 17592 7895 17595
rect 8846 17592 8852 17604
rect 7883 17564 8852 17592
rect 7883 17561 7895 17564
rect 7837 17555 7895 17561
rect 8846 17552 8852 17564
rect 8904 17552 8910 17604
rect 10042 17592 10048 17604
rect 10003 17564 10048 17592
rect 10042 17552 10048 17564
rect 10100 17552 10106 17604
rect 14918 17601 14924 17604
rect 14912 17592 14924 17601
rect 14879 17564 14924 17592
rect 14912 17555 14924 17564
rect 14918 17552 14924 17555
rect 14976 17552 14982 17604
rect 15010 17552 15016 17604
rect 15068 17592 15074 17604
rect 16114 17592 16120 17604
rect 15068 17564 16120 17592
rect 15068 17552 15074 17564
rect 16114 17552 16120 17564
rect 16172 17552 16178 17604
rect 16574 17592 16580 17604
rect 16535 17564 16580 17592
rect 16574 17552 16580 17564
rect 16632 17552 16638 17604
rect 20622 17592 20628 17604
rect 17236 17564 20628 17592
rect 1946 17484 1952 17536
rect 2004 17524 2010 17536
rect 2777 17527 2835 17533
rect 2777 17524 2789 17527
rect 2004 17496 2789 17524
rect 2004 17484 2010 17496
rect 2777 17493 2789 17496
rect 2823 17493 2835 17527
rect 2777 17487 2835 17493
rect 7558 17484 7564 17536
rect 7616 17524 7622 17536
rect 10410 17524 10416 17536
rect 7616 17496 10416 17524
rect 7616 17484 7622 17496
rect 10410 17484 10416 17496
rect 10468 17484 10474 17536
rect 10502 17484 10508 17536
rect 10560 17524 10566 17536
rect 17236 17524 17264 17564
rect 20622 17552 20628 17564
rect 20680 17552 20686 17604
rect 21376 17592 21404 17623
rect 21634 17620 21640 17632
rect 21692 17620 21698 17672
rect 22094 17660 22100 17672
rect 22066 17620 22100 17660
rect 22152 17660 22158 17672
rect 22152 17632 22197 17660
rect 22152 17620 22158 17632
rect 22370 17620 22376 17672
rect 22428 17660 22434 17672
rect 22922 17660 22928 17672
rect 22428 17632 22928 17660
rect 22428 17620 22434 17632
rect 22922 17620 22928 17632
rect 22980 17660 22986 17672
rect 23201 17663 23259 17669
rect 23201 17660 23213 17663
rect 22980 17632 23213 17660
rect 22980 17620 22986 17632
rect 23201 17629 23213 17632
rect 23247 17629 23259 17663
rect 23201 17623 23259 17629
rect 23385 17663 23443 17669
rect 23385 17629 23397 17663
rect 23431 17629 23443 17663
rect 23385 17623 23443 17629
rect 23477 17663 23535 17669
rect 23477 17629 23489 17663
rect 23523 17660 23535 17663
rect 24210 17660 24216 17672
rect 23523 17632 24216 17660
rect 23523 17629 23535 17632
rect 23477 17623 23535 17629
rect 22066 17592 22094 17620
rect 21376 17564 22094 17592
rect 23106 17552 23112 17604
rect 23164 17592 23170 17604
rect 23400 17592 23428 17623
rect 24210 17620 24216 17632
rect 24268 17620 24274 17672
rect 24026 17592 24032 17604
rect 23164 17564 24032 17592
rect 23164 17552 23170 17564
rect 24026 17552 24032 17564
rect 24084 17552 24090 17604
rect 24397 17595 24455 17601
rect 24397 17561 24409 17595
rect 24443 17592 24455 17595
rect 24493 17592 24521 17700
rect 24578 17688 24584 17740
rect 24636 17688 24642 17740
rect 24946 17688 24952 17740
rect 25004 17728 25010 17740
rect 25004 17700 26372 17728
rect 25004 17688 25010 17700
rect 24596 17660 24624 17688
rect 25225 17663 25283 17669
rect 25225 17660 25237 17663
rect 24596 17632 25237 17660
rect 25225 17629 25237 17632
rect 25271 17629 25283 17663
rect 25225 17623 25283 17629
rect 26142 17592 26148 17604
rect 24443 17564 24521 17592
rect 26103 17564 26148 17592
rect 24443 17561 24455 17564
rect 24397 17555 24455 17561
rect 26142 17552 26148 17564
rect 26200 17552 26206 17604
rect 10560 17496 17264 17524
rect 10560 17484 10566 17496
rect 20898 17484 20904 17536
rect 20956 17524 20962 17536
rect 21545 17527 21603 17533
rect 21545 17524 21557 17527
rect 20956 17496 21557 17524
rect 20956 17484 20962 17496
rect 21545 17493 21557 17496
rect 21591 17493 21603 17527
rect 22278 17524 22284 17536
rect 22239 17496 22284 17524
rect 21545 17487 21603 17493
rect 22278 17484 22284 17496
rect 22336 17484 22342 17536
rect 23661 17527 23719 17533
rect 23661 17493 23673 17527
rect 23707 17524 23719 17527
rect 24597 17527 24655 17533
rect 24597 17524 24609 17527
rect 23707 17496 24609 17524
rect 23707 17493 23719 17496
rect 23661 17487 23719 17493
rect 24597 17493 24609 17496
rect 24643 17493 24655 17527
rect 24762 17524 24768 17536
rect 24723 17496 24768 17524
rect 24597 17487 24655 17493
rect 24762 17484 24768 17496
rect 24820 17484 24826 17536
rect 26237 17527 26295 17533
rect 26237 17493 26249 17527
rect 26283 17524 26295 17527
rect 26344 17524 26372 17700
rect 26786 17660 26792 17672
rect 26747 17632 26792 17660
rect 26786 17620 26792 17632
rect 26844 17620 26850 17672
rect 26970 17660 26976 17672
rect 26931 17632 26976 17660
rect 26970 17620 26976 17632
rect 27028 17620 27034 17672
rect 27080 17592 27108 17768
rect 27157 17765 27169 17799
rect 27203 17796 27215 17799
rect 27203 17768 27660 17796
rect 27203 17765 27215 17768
rect 27157 17759 27215 17765
rect 27632 17737 27660 17768
rect 30760 17768 33732 17796
rect 27617 17731 27675 17737
rect 27617 17697 27629 17731
rect 27663 17697 27675 17731
rect 27617 17691 27675 17697
rect 28350 17688 28356 17740
rect 28408 17728 28414 17740
rect 28626 17728 28632 17740
rect 28408 17700 28632 17728
rect 28408 17688 28414 17700
rect 28626 17688 28632 17700
rect 28684 17728 28690 17740
rect 28721 17731 28779 17737
rect 28721 17728 28733 17731
rect 28684 17700 28733 17728
rect 28684 17688 28690 17700
rect 28721 17697 28733 17700
rect 28767 17697 28779 17731
rect 28721 17691 28779 17697
rect 27338 17620 27344 17672
rect 27396 17660 27402 17672
rect 30760 17669 30788 17768
rect 31389 17731 31447 17737
rect 31389 17697 31401 17731
rect 31435 17728 31447 17731
rect 31754 17728 31760 17740
rect 31435 17700 31760 17728
rect 31435 17697 31447 17700
rect 31389 17691 31447 17697
rect 31754 17688 31760 17700
rect 31812 17688 31818 17740
rect 33042 17728 33048 17740
rect 33003 17700 33048 17728
rect 33042 17688 33048 17700
rect 33100 17688 33106 17740
rect 33704 17669 33732 17768
rect 27801 17663 27859 17669
rect 27801 17660 27813 17663
rect 27396 17632 27813 17660
rect 27396 17620 27402 17632
rect 27801 17629 27813 17632
rect 27847 17629 27859 17663
rect 30745 17663 30803 17669
rect 30745 17660 30757 17663
rect 27801 17623 27859 17629
rect 28184 17632 30757 17660
rect 28184 17592 28212 17632
rect 30745 17629 30757 17632
rect 30791 17629 30803 17663
rect 30745 17623 30803 17629
rect 33689 17663 33747 17669
rect 33689 17629 33701 17663
rect 33735 17660 33747 17663
rect 34238 17660 34244 17672
rect 33735 17632 34244 17660
rect 33735 17629 33747 17632
rect 33689 17623 33747 17629
rect 34238 17620 34244 17632
rect 34296 17660 34302 17672
rect 34701 17663 34759 17669
rect 34701 17660 34713 17663
rect 34296 17632 34713 17660
rect 34296 17620 34302 17632
rect 34701 17629 34713 17632
rect 34747 17629 34759 17663
rect 34701 17623 34759 17629
rect 46290 17620 46296 17672
rect 46348 17660 46354 17672
rect 47673 17663 47731 17669
rect 47673 17660 47685 17663
rect 46348 17632 47685 17660
rect 46348 17620 46354 17632
rect 47673 17629 47685 17632
rect 47719 17629 47731 17663
rect 47673 17623 47731 17629
rect 27080 17564 28212 17592
rect 28537 17595 28595 17601
rect 28537 17561 28549 17595
rect 28583 17592 28595 17595
rect 29638 17592 29644 17604
rect 28583 17564 29644 17592
rect 28583 17561 28595 17564
rect 28537 17555 28595 17561
rect 29638 17552 29644 17564
rect 29696 17552 29702 17604
rect 30837 17595 30895 17601
rect 30837 17561 30849 17595
rect 30883 17592 30895 17595
rect 31573 17595 31631 17601
rect 31573 17592 31585 17595
rect 30883 17564 31585 17592
rect 30883 17561 30895 17564
rect 30837 17555 30895 17561
rect 31573 17561 31585 17564
rect 31619 17561 31631 17595
rect 31573 17555 31631 17561
rect 29822 17524 29828 17536
rect 26283 17496 29828 17524
rect 26283 17493 26295 17496
rect 26237 17487 26295 17493
rect 29822 17484 29828 17496
rect 29880 17484 29886 17536
rect 33502 17484 33508 17536
rect 33560 17524 33566 17536
rect 33781 17527 33839 17533
rect 33781 17524 33793 17527
rect 33560 17496 33793 17524
rect 33560 17484 33566 17496
rect 33781 17493 33793 17496
rect 33827 17493 33839 17527
rect 33781 17487 33839 17493
rect 1104 17434 48852 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 48852 17434
rect 1104 17360 48852 17382
rect 1670 17280 1676 17332
rect 1728 17320 1734 17332
rect 7558 17320 7564 17332
rect 1728 17292 7564 17320
rect 1728 17280 1734 17292
rect 7558 17280 7564 17292
rect 7616 17280 7622 17332
rect 8846 17320 8852 17332
rect 8807 17292 8852 17320
rect 8846 17280 8852 17292
rect 8904 17280 8910 17332
rect 10042 17320 10048 17332
rect 10003 17292 10048 17320
rect 10042 17280 10048 17292
rect 10100 17280 10106 17332
rect 15286 17320 15292 17332
rect 14292 17292 15292 17320
rect 1946 17252 1952 17264
rect 1907 17224 1952 17252
rect 1946 17212 1952 17224
rect 2004 17212 2010 17264
rect 12894 17252 12900 17264
rect 11854 17224 12900 17252
rect 1762 17184 1768 17196
rect 1723 17156 1768 17184
rect 1762 17144 1768 17156
rect 1820 17144 1826 17196
rect 8757 17187 8815 17193
rect 8757 17153 8769 17187
rect 8803 17184 8815 17187
rect 9766 17184 9772 17196
rect 8803 17156 9772 17184
rect 8803 17153 8815 17156
rect 8757 17147 8815 17153
rect 9766 17144 9772 17156
rect 9824 17144 9830 17196
rect 9950 17184 9956 17196
rect 9911 17156 9956 17184
rect 9950 17144 9956 17156
rect 10008 17184 10014 17196
rect 10502 17184 10508 17196
rect 10008 17156 10508 17184
rect 10008 17144 10014 17156
rect 10502 17144 10508 17156
rect 10560 17144 10566 17196
rect 10597 17187 10655 17193
rect 10597 17153 10609 17187
rect 10643 17153 10655 17187
rect 10597 17147 10655 17153
rect 10781 17187 10839 17193
rect 10781 17153 10793 17187
rect 10827 17184 10839 17187
rect 11514 17184 11520 17196
rect 10827 17156 11520 17184
rect 10827 17153 10839 17156
rect 10781 17147 10839 17153
rect 2774 17076 2780 17128
rect 2832 17116 2838 17128
rect 2832 17088 2877 17116
rect 2832 17076 2838 17088
rect 10612 17048 10640 17147
rect 11514 17144 11520 17156
rect 11572 17144 11578 17196
rect 11854 17193 11882 17224
rect 12894 17212 12900 17224
rect 12952 17212 12958 17264
rect 11839 17187 11897 17193
rect 11839 17153 11851 17187
rect 11885 17153 11897 17187
rect 11974 17184 11980 17196
rect 11935 17156 11980 17184
rect 11839 17147 11897 17153
rect 11974 17144 11980 17156
rect 12032 17144 12038 17196
rect 12069 17187 12127 17193
rect 12069 17153 12081 17187
rect 12115 17184 12127 17187
rect 12253 17187 12311 17193
rect 12115 17156 12204 17184
rect 12115 17153 12127 17156
rect 12069 17147 12127 17153
rect 10965 17119 11023 17125
rect 10965 17085 10977 17119
rect 11011 17116 11023 17119
rect 12176 17116 12204 17156
rect 12253 17153 12265 17187
rect 12299 17184 12311 17187
rect 12710 17184 12716 17196
rect 12299 17156 12434 17184
rect 12671 17156 12716 17184
rect 12299 17153 12311 17156
rect 12253 17147 12311 17153
rect 11011 17088 12204 17116
rect 12406 17116 12434 17156
rect 12710 17144 12716 17156
rect 12768 17144 12774 17196
rect 14292 17193 14320 17292
rect 15286 17280 15292 17292
rect 15344 17320 15350 17332
rect 15930 17320 15936 17332
rect 15344 17292 15936 17320
rect 15344 17280 15350 17292
rect 15930 17280 15936 17292
rect 15988 17280 15994 17332
rect 18506 17280 18512 17332
rect 18564 17320 18570 17332
rect 20806 17320 20812 17332
rect 18564 17292 20812 17320
rect 18564 17280 18570 17292
rect 20806 17280 20812 17292
rect 20864 17280 20870 17332
rect 20901 17323 20959 17329
rect 20901 17289 20913 17323
rect 20947 17320 20959 17323
rect 20990 17320 20996 17332
rect 20947 17292 20996 17320
rect 20947 17289 20959 17292
rect 20901 17283 20959 17289
rect 20990 17280 20996 17292
rect 21048 17280 21054 17332
rect 21266 17280 21272 17332
rect 21324 17320 21330 17332
rect 21818 17320 21824 17332
rect 21324 17292 21824 17320
rect 21324 17280 21330 17292
rect 21818 17280 21824 17292
rect 21876 17280 21882 17332
rect 22094 17280 22100 17332
rect 22152 17320 22158 17332
rect 22281 17323 22339 17329
rect 22281 17320 22293 17323
rect 22152 17292 22293 17320
rect 22152 17280 22158 17292
rect 22281 17289 22293 17292
rect 22327 17289 22339 17323
rect 24121 17323 24179 17329
rect 24121 17320 24133 17323
rect 22281 17283 22339 17289
rect 22756 17292 24133 17320
rect 14458 17212 14464 17264
rect 14516 17252 14522 17264
rect 14516 17224 15700 17252
rect 14516 17212 14522 17224
rect 14277 17187 14335 17193
rect 14277 17184 14289 17187
rect 12912 17156 14289 17184
rect 12912 17116 12940 17156
rect 14277 17153 14289 17156
rect 14323 17153 14335 17187
rect 14277 17147 14335 17153
rect 15378 17144 15384 17196
rect 15436 17190 15442 17196
rect 15672 17193 15700 17224
rect 16022 17212 16028 17264
rect 16080 17252 16086 17264
rect 22756 17252 22784 17292
rect 24121 17289 24133 17292
rect 24167 17320 24179 17323
rect 24949 17323 25007 17329
rect 24167 17292 24808 17320
rect 24167 17289 24179 17292
rect 24121 17283 24179 17289
rect 22922 17252 22928 17264
rect 16080 17224 22784 17252
rect 22883 17224 22928 17252
rect 16080 17212 16086 17224
rect 22922 17212 22928 17224
rect 22980 17212 22986 17264
rect 23014 17212 23020 17264
rect 23072 17252 23078 17264
rect 24489 17255 24547 17261
rect 24489 17252 24501 17255
rect 23072 17224 24501 17252
rect 23072 17212 23078 17224
rect 24489 17221 24501 17224
rect 24535 17221 24547 17255
rect 24489 17215 24547 17221
rect 15545 17190 15603 17193
rect 15436 17187 15603 17190
rect 15436 17162 15557 17187
rect 15436 17144 15442 17162
rect 15545 17153 15557 17162
rect 15591 17153 15603 17187
rect 15545 17147 15603 17153
rect 15657 17187 15715 17193
rect 15657 17153 15669 17187
rect 15703 17153 15715 17187
rect 15657 17147 15715 17153
rect 15770 17187 15828 17193
rect 15770 17153 15782 17187
rect 15816 17184 15828 17187
rect 15816 17156 15884 17184
rect 15816 17153 15828 17156
rect 15770 17147 15828 17153
rect 12406 17088 12940 17116
rect 11011 17085 11023 17088
rect 10965 17079 11023 17085
rect 13722 17076 13728 17128
rect 13780 17116 13786 17128
rect 14001 17119 14059 17125
rect 14001 17116 14013 17119
rect 13780 17088 14013 17116
rect 13780 17076 13786 17088
rect 14001 17085 14013 17088
rect 14047 17085 14059 17119
rect 14001 17079 14059 17085
rect 15856 17060 15884 17156
rect 15930 17144 15936 17196
rect 15988 17184 15994 17196
rect 17865 17187 17923 17193
rect 15988 17156 16033 17184
rect 15988 17144 15994 17156
rect 17865 17153 17877 17187
rect 17911 17184 17923 17187
rect 18322 17184 18328 17196
rect 17911 17156 18328 17184
rect 17911 17153 17923 17156
rect 17865 17147 17923 17153
rect 18322 17144 18328 17156
rect 18380 17184 18386 17196
rect 18693 17187 18751 17193
rect 18693 17184 18705 17187
rect 18380 17156 18705 17184
rect 18380 17144 18386 17156
rect 18693 17153 18705 17156
rect 18739 17153 18751 17187
rect 18693 17147 18751 17153
rect 19788 17187 19846 17193
rect 19788 17153 19800 17187
rect 19834 17184 19846 17187
rect 20530 17184 20536 17196
rect 19834 17156 20536 17184
rect 19834 17153 19846 17156
rect 19788 17147 19846 17153
rect 20530 17144 20536 17156
rect 20588 17144 20594 17196
rect 22186 17184 22192 17196
rect 22147 17156 22192 17184
rect 22186 17144 22192 17156
rect 22244 17144 22250 17196
rect 22373 17187 22431 17193
rect 22373 17153 22385 17187
rect 22419 17153 22431 17187
rect 23106 17184 23112 17196
rect 23067 17156 23112 17184
rect 22373 17147 22431 17153
rect 17402 17076 17408 17128
rect 17460 17116 17466 17128
rect 19521 17119 19579 17125
rect 19521 17116 19533 17119
rect 17460 17088 19533 17116
rect 17460 17076 17466 17088
rect 19521 17085 19533 17088
rect 19567 17085 19579 17119
rect 19521 17079 19579 17085
rect 20898 17076 20904 17128
rect 20956 17116 20962 17128
rect 21634 17116 21640 17128
rect 20956 17088 21640 17116
rect 20956 17076 20962 17088
rect 21634 17076 21640 17088
rect 21692 17116 21698 17128
rect 22388 17116 22416 17147
rect 23106 17144 23112 17156
rect 23164 17144 23170 17196
rect 23201 17187 23259 17193
rect 23201 17153 23213 17187
rect 23247 17184 23259 17187
rect 23566 17184 23572 17196
rect 23247 17156 23572 17184
rect 23247 17153 23259 17156
rect 23201 17147 23259 17153
rect 23566 17144 23572 17156
rect 23624 17144 23630 17196
rect 24780 17193 24808 17292
rect 24949 17289 24961 17323
rect 24995 17320 25007 17323
rect 25038 17320 25044 17332
rect 24995 17292 25044 17320
rect 24995 17289 25007 17292
rect 24949 17283 25007 17289
rect 25038 17280 25044 17292
rect 25096 17280 25102 17332
rect 25130 17280 25136 17332
rect 25188 17320 25194 17332
rect 25593 17323 25651 17329
rect 25593 17320 25605 17323
rect 25188 17292 25605 17320
rect 25188 17280 25194 17292
rect 25593 17289 25605 17292
rect 25639 17289 25651 17323
rect 25593 17283 25651 17289
rect 26786 17280 26792 17332
rect 26844 17320 26850 17332
rect 27433 17323 27491 17329
rect 27433 17320 27445 17323
rect 26844 17292 27445 17320
rect 26844 17280 26850 17292
rect 27433 17289 27445 17292
rect 27479 17289 27491 17323
rect 29086 17320 29092 17332
rect 27433 17283 27491 17289
rect 27908 17292 29092 17320
rect 24854 17212 24860 17264
rect 24912 17252 24918 17264
rect 27908 17261 27936 17292
rect 29086 17280 29092 17292
rect 29144 17280 29150 17332
rect 27893 17255 27951 17261
rect 27893 17252 27905 17255
rect 24912 17224 27905 17252
rect 24912 17212 24918 17224
rect 27893 17221 27905 17224
rect 27939 17221 27951 17255
rect 28074 17252 28080 17264
rect 28035 17224 28080 17252
rect 27893 17215 27951 17221
rect 28074 17212 28080 17224
rect 28132 17212 28138 17264
rect 28261 17255 28319 17261
rect 28261 17221 28273 17255
rect 28307 17252 28319 17255
rect 29454 17252 29460 17264
rect 28307 17224 29460 17252
rect 28307 17221 28319 17224
rect 28261 17215 28319 17221
rect 29454 17212 29460 17224
rect 29512 17212 29518 17264
rect 33502 17252 33508 17264
rect 33463 17224 33508 17252
rect 33502 17212 33508 17224
rect 33560 17212 33566 17264
rect 23845 17187 23903 17193
rect 23845 17153 23857 17187
rect 23891 17153 23903 17187
rect 23845 17147 23903 17153
rect 24765 17187 24823 17193
rect 24765 17153 24777 17187
rect 24811 17153 24823 17187
rect 24765 17147 24823 17153
rect 23290 17116 23296 17128
rect 21692 17088 23296 17116
rect 21692 17076 21698 17088
rect 23290 17076 23296 17088
rect 23348 17076 23354 17128
rect 23860 17116 23888 17147
rect 25130 17144 25136 17196
rect 25188 17184 25194 17196
rect 25501 17187 25559 17193
rect 25501 17184 25513 17187
rect 25188 17156 25513 17184
rect 25188 17144 25194 17156
rect 25501 17153 25513 17156
rect 25547 17153 25559 17187
rect 25501 17147 25559 17153
rect 27065 17187 27123 17193
rect 27065 17153 27077 17187
rect 27111 17184 27123 17187
rect 27154 17184 27160 17196
rect 27111 17156 27160 17184
rect 27111 17153 27123 17156
rect 27065 17147 27123 17153
rect 27154 17144 27160 17156
rect 27212 17144 27218 17196
rect 27249 17187 27307 17193
rect 27249 17153 27261 17187
rect 27295 17184 27307 17187
rect 27338 17184 27344 17196
rect 27295 17156 27344 17184
rect 27295 17153 27307 17156
rect 27249 17147 27307 17153
rect 27338 17144 27344 17156
rect 27396 17144 27402 17196
rect 29080 17187 29138 17193
rect 29080 17153 29092 17187
rect 29126 17184 29138 17187
rect 30282 17184 30288 17196
rect 29126 17156 30288 17184
rect 29126 17153 29138 17156
rect 29080 17147 29138 17153
rect 30282 17144 30288 17156
rect 30340 17144 30346 17196
rect 47394 17144 47400 17196
rect 47452 17184 47458 17196
rect 47581 17187 47639 17193
rect 47581 17184 47593 17187
rect 47452 17156 47593 17184
rect 47452 17144 47458 17156
rect 47581 17153 47593 17156
rect 47627 17153 47639 17187
rect 47581 17147 47639 17153
rect 24118 17116 24124 17128
rect 23860 17088 24124 17116
rect 24118 17076 24124 17088
rect 24176 17076 24182 17128
rect 24302 17076 24308 17128
rect 24360 17116 24366 17128
rect 24581 17119 24639 17125
rect 24581 17116 24593 17119
rect 24360 17088 24593 17116
rect 24360 17076 24366 17088
rect 24581 17085 24593 17088
rect 24627 17085 24639 17119
rect 24581 17079 24639 17085
rect 28813 17119 28871 17125
rect 28813 17085 28825 17119
rect 28859 17085 28871 17119
rect 28813 17079 28871 17085
rect 33321 17119 33379 17125
rect 33321 17085 33333 17119
rect 33367 17116 33379 17119
rect 33502 17116 33508 17128
rect 33367 17088 33508 17116
rect 33367 17085 33379 17088
rect 33321 17079 33379 17085
rect 10612 17020 11836 17048
rect 11609 16983 11667 16989
rect 11609 16949 11621 16983
rect 11655 16980 11667 16983
rect 11698 16980 11704 16992
rect 11655 16952 11704 16980
rect 11655 16949 11667 16952
rect 11609 16943 11667 16949
rect 11698 16940 11704 16952
rect 11756 16940 11762 16992
rect 11808 16980 11836 17020
rect 11882 17008 11888 17060
rect 11940 17048 11946 17060
rect 15378 17048 15384 17060
rect 11940 17020 15384 17048
rect 11940 17008 11946 17020
rect 15378 17008 15384 17020
rect 15436 17008 15442 17060
rect 15838 17008 15844 17060
rect 15896 17008 15902 17060
rect 20622 17008 20628 17060
rect 20680 17048 20686 17060
rect 22554 17048 22560 17060
rect 20680 17020 22560 17048
rect 20680 17008 20686 17020
rect 22554 17008 22560 17020
rect 22612 17008 22618 17060
rect 23385 17051 23443 17057
rect 23385 17048 23397 17051
rect 22756 17020 23397 17048
rect 12943 16983 13001 16989
rect 12943 16980 12955 16983
rect 11808 16952 12955 16980
rect 12943 16949 12955 16952
rect 12989 16980 13001 16983
rect 14274 16980 14280 16992
rect 12989 16952 14280 16980
rect 12989 16949 13001 16952
rect 12943 16943 13001 16949
rect 14274 16940 14280 16952
rect 14332 16940 14338 16992
rect 15194 16940 15200 16992
rect 15252 16980 15258 16992
rect 15289 16983 15347 16989
rect 15289 16980 15301 16983
rect 15252 16952 15301 16980
rect 15252 16940 15258 16952
rect 15289 16949 15301 16952
rect 15335 16949 15347 16983
rect 15289 16943 15347 16949
rect 15470 16940 15476 16992
rect 15528 16980 15534 16992
rect 17957 16983 18015 16989
rect 17957 16980 17969 16983
rect 15528 16952 17969 16980
rect 15528 16940 15534 16952
rect 17957 16949 17969 16952
rect 18003 16980 18015 16983
rect 18598 16980 18604 16992
rect 18003 16952 18604 16980
rect 18003 16949 18015 16952
rect 17957 16943 18015 16949
rect 18598 16940 18604 16952
rect 18656 16940 18662 16992
rect 18877 16983 18935 16989
rect 18877 16949 18889 16983
rect 18923 16980 18935 16983
rect 18966 16980 18972 16992
rect 18923 16952 18972 16980
rect 18923 16949 18935 16952
rect 18877 16943 18935 16949
rect 18966 16940 18972 16952
rect 19024 16940 19030 16992
rect 20162 16940 20168 16992
rect 20220 16980 20226 16992
rect 20438 16980 20444 16992
rect 20220 16952 20444 16980
rect 20220 16940 20226 16952
rect 20438 16940 20444 16952
rect 20496 16940 20502 16992
rect 20806 16940 20812 16992
rect 20864 16980 20870 16992
rect 22756 16980 22784 17020
rect 23385 17017 23397 17020
rect 23431 17017 23443 17051
rect 23385 17011 23443 17017
rect 23842 17008 23848 17060
rect 23900 17048 23906 17060
rect 24762 17048 24768 17060
rect 23900 17020 24768 17048
rect 23900 17008 23906 17020
rect 24762 17008 24768 17020
rect 24820 17008 24826 17060
rect 27246 17048 27252 17060
rect 25516 17020 27252 17048
rect 20864 16952 22784 16980
rect 23201 16983 23259 16989
rect 20864 16940 20870 16952
rect 23201 16949 23213 16983
rect 23247 16980 23259 16983
rect 23474 16980 23480 16992
rect 23247 16952 23480 16980
rect 23247 16949 23259 16952
rect 23201 16943 23259 16949
rect 23474 16940 23480 16952
rect 23532 16940 23538 16992
rect 23658 16980 23664 16992
rect 23619 16952 23664 16980
rect 23658 16940 23664 16952
rect 23716 16940 23722 16992
rect 24673 16983 24731 16989
rect 24673 16949 24685 16983
rect 24719 16980 24731 16983
rect 25516 16980 25544 17020
rect 27246 17008 27252 17020
rect 27304 17008 27310 17060
rect 24719 16952 25544 16980
rect 28828 16980 28856 17079
rect 33502 17076 33508 17088
rect 33560 17076 33566 17128
rect 33594 17076 33600 17128
rect 33652 17116 33658 17128
rect 33781 17119 33839 17125
rect 33781 17116 33793 17119
rect 33652 17088 33793 17116
rect 33652 17076 33658 17088
rect 33781 17085 33793 17088
rect 33827 17085 33839 17119
rect 33781 17079 33839 17085
rect 29546 16980 29552 16992
rect 28828 16952 29552 16980
rect 24719 16949 24731 16952
rect 24673 16943 24731 16949
rect 29546 16940 29552 16952
rect 29604 16940 29610 16992
rect 30190 16980 30196 16992
rect 30151 16952 30196 16980
rect 30190 16940 30196 16952
rect 30248 16940 30254 16992
rect 47670 16980 47676 16992
rect 47631 16952 47676 16980
rect 47670 16940 47676 16952
rect 47728 16940 47734 16992
rect 1104 16890 48852 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 48852 16890
rect 1104 16816 48852 16838
rect 1949 16779 2007 16785
rect 1949 16745 1961 16779
rect 1995 16776 2007 16779
rect 1995 16748 16528 16776
rect 1995 16745 2007 16748
rect 1949 16739 2007 16745
rect 2682 16668 2688 16720
rect 2740 16708 2746 16720
rect 2740 16668 2774 16708
rect 2746 16640 2774 16668
rect 2746 16612 11192 16640
rect 1854 16572 1860 16584
rect 1815 16544 1860 16572
rect 1854 16532 1860 16544
rect 1912 16532 1918 16584
rect 10796 16581 10824 16612
rect 10781 16575 10839 16581
rect 10781 16541 10793 16575
rect 10827 16541 10839 16575
rect 10781 16535 10839 16541
rect 11164 16504 11192 16612
rect 11238 16600 11244 16652
rect 11296 16640 11302 16652
rect 11425 16643 11483 16649
rect 11425 16640 11437 16643
rect 11296 16612 11437 16640
rect 11296 16600 11302 16612
rect 11425 16609 11437 16612
rect 11471 16609 11483 16643
rect 14366 16640 14372 16652
rect 14327 16612 14372 16640
rect 11425 16603 11483 16609
rect 14366 16600 14372 16612
rect 14424 16600 14430 16652
rect 16500 16640 16528 16748
rect 16574 16736 16580 16788
rect 16632 16776 16638 16788
rect 17678 16776 17684 16788
rect 16632 16748 17684 16776
rect 16632 16736 16638 16748
rect 17678 16736 17684 16748
rect 17736 16776 17742 16788
rect 18417 16779 18475 16785
rect 18417 16776 18429 16779
rect 17736 16748 18429 16776
rect 17736 16736 17742 16748
rect 18417 16745 18429 16748
rect 18463 16745 18475 16779
rect 18417 16739 18475 16745
rect 19981 16779 20039 16785
rect 19981 16745 19993 16779
rect 20027 16776 20039 16779
rect 20070 16776 20076 16788
rect 20027 16748 20076 16776
rect 20027 16745 20039 16748
rect 19981 16739 20039 16745
rect 20070 16736 20076 16748
rect 20128 16736 20134 16788
rect 20530 16776 20536 16788
rect 20491 16748 20536 16776
rect 20530 16736 20536 16748
rect 20588 16736 20594 16788
rect 28350 16776 28356 16788
rect 24412 16748 28356 16776
rect 17402 16708 17408 16720
rect 17363 16680 17408 16708
rect 17402 16668 17408 16680
rect 17460 16668 17466 16720
rect 23014 16640 23020 16652
rect 16500 16612 23020 16640
rect 23014 16600 23020 16612
rect 23072 16600 23078 16652
rect 24412 16649 24440 16748
rect 28350 16736 28356 16748
rect 28408 16736 28414 16788
rect 28902 16736 28908 16788
rect 28960 16776 28966 16788
rect 30282 16776 30288 16788
rect 28960 16748 29868 16776
rect 30243 16748 30288 16776
rect 28960 16736 28966 16748
rect 27617 16711 27675 16717
rect 27617 16677 27629 16711
rect 27663 16708 27675 16711
rect 27663 16680 29776 16708
rect 27663 16677 27675 16680
rect 27617 16671 27675 16677
rect 24397 16643 24455 16649
rect 24397 16609 24409 16643
rect 24443 16609 24455 16643
rect 27154 16640 27160 16652
rect 27115 16612 27160 16640
rect 24397 16603 24455 16609
rect 27154 16600 27160 16612
rect 27212 16640 27218 16652
rect 28534 16640 28540 16652
rect 27212 16612 27660 16640
rect 28495 16612 28540 16640
rect 27212 16600 27218 16612
rect 11698 16581 11704 16584
rect 11692 16572 11704 16581
rect 11659 16544 11704 16572
rect 11692 16535 11704 16544
rect 11698 16532 11704 16535
rect 11756 16532 11762 16584
rect 14636 16575 14694 16581
rect 14636 16541 14648 16575
rect 14682 16572 14694 16575
rect 15194 16572 15200 16584
rect 14682 16544 15200 16572
rect 14682 16541 14694 16544
rect 14636 16535 14694 16541
rect 15194 16532 15200 16544
rect 15252 16532 15258 16584
rect 18325 16575 18383 16581
rect 18325 16541 18337 16575
rect 18371 16572 18383 16575
rect 18371 16544 20668 16572
rect 18371 16541 18383 16544
rect 18325 16535 18383 16541
rect 11882 16504 11888 16516
rect 11164 16476 11888 16504
rect 11882 16464 11888 16476
rect 11940 16464 11946 16516
rect 17221 16507 17279 16513
rect 17221 16473 17233 16507
rect 17267 16504 17279 16507
rect 17862 16504 17868 16516
rect 17267 16476 17868 16504
rect 17267 16473 17279 16476
rect 17221 16467 17279 16473
rect 17862 16464 17868 16476
rect 17920 16464 17926 16516
rect 18966 16464 18972 16516
rect 19024 16504 19030 16516
rect 19705 16507 19763 16513
rect 19705 16504 19717 16507
rect 19024 16476 19717 16504
rect 19024 16464 19030 16476
rect 19705 16473 19717 16476
rect 19751 16473 19763 16507
rect 20640 16504 20668 16544
rect 20714 16532 20720 16584
rect 20772 16572 20778 16584
rect 20901 16575 20959 16581
rect 20772 16544 20817 16572
rect 20772 16532 20778 16544
rect 20901 16541 20913 16575
rect 20947 16541 20959 16575
rect 20901 16535 20959 16541
rect 20806 16504 20812 16516
rect 20640 16476 20812 16504
rect 19705 16467 19763 16473
rect 20806 16464 20812 16476
rect 20864 16464 20870 16516
rect 20916 16504 20944 16535
rect 20990 16532 20996 16584
rect 21048 16572 21054 16584
rect 21048 16544 21093 16572
rect 21048 16532 21054 16544
rect 21450 16532 21456 16584
rect 21508 16572 21514 16584
rect 21545 16575 21603 16581
rect 21545 16572 21557 16575
rect 21508 16544 21557 16572
rect 21508 16532 21514 16544
rect 21545 16541 21557 16544
rect 21591 16541 21603 16575
rect 21545 16535 21603 16541
rect 23658 16532 23664 16584
rect 23716 16572 23722 16584
rect 24653 16575 24711 16581
rect 24653 16572 24665 16575
rect 23716 16544 24665 16572
rect 23716 16532 23722 16544
rect 24653 16541 24665 16544
rect 24699 16541 24711 16575
rect 24653 16535 24711 16541
rect 27249 16575 27307 16581
rect 27249 16541 27261 16575
rect 27295 16572 27307 16575
rect 27430 16572 27436 16584
rect 27295 16544 27436 16572
rect 27295 16541 27307 16544
rect 27249 16535 27307 16541
rect 27430 16532 27436 16544
rect 27488 16532 27494 16584
rect 20916 16476 21036 16504
rect 21008 16448 21036 16476
rect 10873 16439 10931 16445
rect 10873 16405 10885 16439
rect 10919 16436 10931 16439
rect 11698 16436 11704 16448
rect 10919 16408 11704 16436
rect 10919 16405 10931 16408
rect 10873 16399 10931 16405
rect 11698 16396 11704 16408
rect 11756 16396 11762 16448
rect 11790 16396 11796 16448
rect 11848 16436 11854 16448
rect 12805 16439 12863 16445
rect 12805 16436 12817 16439
rect 11848 16408 12817 16436
rect 11848 16396 11854 16408
rect 12805 16405 12817 16408
rect 12851 16405 12863 16439
rect 12805 16399 12863 16405
rect 15749 16439 15807 16445
rect 15749 16405 15761 16439
rect 15795 16436 15807 16439
rect 16666 16436 16672 16448
rect 15795 16408 16672 16436
rect 15795 16405 15807 16408
rect 15749 16399 15807 16405
rect 16666 16396 16672 16408
rect 16724 16396 16730 16448
rect 20990 16396 20996 16448
rect 21048 16436 21054 16448
rect 21637 16439 21695 16445
rect 21637 16436 21649 16439
rect 21048 16408 21649 16436
rect 21048 16396 21054 16408
rect 21637 16405 21649 16408
rect 21683 16405 21695 16439
rect 21637 16399 21695 16405
rect 25130 16396 25136 16448
rect 25188 16436 25194 16448
rect 25777 16439 25835 16445
rect 25777 16436 25789 16439
rect 25188 16408 25789 16436
rect 25188 16396 25194 16408
rect 25777 16405 25789 16408
rect 25823 16405 25835 16439
rect 27632 16436 27660 16612
rect 28534 16600 28540 16612
rect 28592 16600 28598 16652
rect 28626 16600 28632 16652
rect 28684 16640 28690 16652
rect 28684 16612 28729 16640
rect 28684 16600 28690 16612
rect 28074 16532 28080 16584
rect 28132 16572 28138 16584
rect 28445 16575 28503 16581
rect 28445 16572 28457 16575
rect 28132 16544 28457 16572
rect 28132 16532 28138 16544
rect 28445 16541 28457 16544
rect 28491 16541 28503 16575
rect 28552 16572 28580 16600
rect 28552 16544 29408 16572
rect 28445 16535 28503 16541
rect 28077 16439 28135 16445
rect 28077 16436 28089 16439
rect 27632 16408 28089 16436
rect 25777 16399 25835 16405
rect 28077 16405 28089 16408
rect 28123 16405 28135 16439
rect 28460 16436 28488 16535
rect 29380 16504 29408 16544
rect 29454 16532 29460 16584
rect 29512 16572 29518 16584
rect 29748 16581 29776 16680
rect 29840 16640 29868 16748
rect 30282 16736 30288 16748
rect 30340 16736 30346 16788
rect 29917 16643 29975 16649
rect 29917 16640 29929 16643
rect 29840 16612 29929 16640
rect 29917 16609 29929 16612
rect 29963 16609 29975 16643
rect 46290 16640 46296 16652
rect 46251 16612 46296 16640
rect 29917 16603 29975 16609
rect 46290 16600 46296 16612
rect 46348 16600 46354 16652
rect 48130 16640 48136 16652
rect 48091 16612 48136 16640
rect 48130 16600 48136 16612
rect 48188 16600 48194 16652
rect 29549 16575 29607 16581
rect 29549 16572 29561 16575
rect 29512 16544 29561 16572
rect 29512 16532 29518 16544
rect 29549 16541 29561 16544
rect 29595 16541 29607 16575
rect 29549 16535 29607 16541
rect 29733 16575 29791 16581
rect 29733 16541 29745 16575
rect 29779 16541 29791 16575
rect 29733 16535 29791 16541
rect 29822 16532 29828 16584
rect 29880 16572 29886 16584
rect 30101 16575 30159 16581
rect 29880 16544 29925 16572
rect 29880 16532 29886 16544
rect 30101 16541 30113 16575
rect 30147 16572 30159 16575
rect 30190 16572 30196 16584
rect 30147 16544 30196 16572
rect 30147 16541 30159 16544
rect 30101 16535 30159 16541
rect 30116 16504 30144 16535
rect 30190 16532 30196 16544
rect 30248 16532 30254 16584
rect 31757 16575 31815 16581
rect 31757 16541 31769 16575
rect 31803 16572 31815 16575
rect 32858 16572 32864 16584
rect 31803 16544 32864 16572
rect 31803 16541 31815 16544
rect 31757 16535 31815 16541
rect 32858 16532 32864 16544
rect 32916 16532 32922 16584
rect 29380 16476 30144 16504
rect 30374 16464 30380 16516
rect 30432 16504 30438 16516
rect 31478 16504 31484 16516
rect 30432 16476 31484 16504
rect 30432 16464 30438 16476
rect 31478 16464 31484 16476
rect 31536 16464 31542 16516
rect 31573 16507 31631 16513
rect 31573 16473 31585 16507
rect 31619 16504 31631 16507
rect 31662 16504 31668 16516
rect 31619 16476 31668 16504
rect 31619 16473 31631 16476
rect 31573 16467 31631 16473
rect 31662 16464 31668 16476
rect 31720 16464 31726 16516
rect 46477 16507 46535 16513
rect 46477 16473 46489 16507
rect 46523 16504 46535 16507
rect 47670 16504 47676 16516
rect 46523 16476 47676 16504
rect 46523 16473 46535 16476
rect 46477 16467 46535 16473
rect 47670 16464 47676 16476
rect 47728 16464 47734 16516
rect 30742 16436 30748 16448
rect 28460 16408 30748 16436
rect 28077 16399 28135 16405
rect 30742 16396 30748 16408
rect 30800 16396 30806 16448
rect 31938 16436 31944 16448
rect 31899 16408 31944 16436
rect 31938 16396 31944 16408
rect 31996 16396 32002 16448
rect 36538 16396 36544 16448
rect 36596 16436 36602 16448
rect 47486 16436 47492 16448
rect 36596 16408 47492 16436
rect 36596 16396 36602 16408
rect 47486 16396 47492 16408
rect 47544 16396 47550 16448
rect 1104 16346 48852 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 48852 16346
rect 1104 16272 48852 16294
rect 11514 16192 11520 16244
rect 11572 16232 11578 16244
rect 11790 16232 11796 16244
rect 11572 16204 11796 16232
rect 11572 16192 11578 16204
rect 11790 16192 11796 16204
rect 11848 16192 11854 16244
rect 14829 16235 14887 16241
rect 14829 16201 14841 16235
rect 14875 16232 14887 16235
rect 15838 16232 15844 16244
rect 14875 16204 15844 16232
rect 14875 16201 14887 16204
rect 14829 16195 14887 16201
rect 15838 16192 15844 16204
rect 15896 16192 15902 16244
rect 27154 16232 27160 16244
rect 15948 16204 27160 16232
rect 11698 16164 11704 16176
rect 11659 16136 11704 16164
rect 11698 16124 11704 16136
rect 11756 16124 11762 16176
rect 14274 16124 14280 16176
rect 14332 16164 14338 16176
rect 14461 16167 14519 16173
rect 14461 16164 14473 16167
rect 14332 16136 14473 16164
rect 14332 16124 14338 16136
rect 14461 16133 14473 16136
rect 14507 16133 14519 16167
rect 14461 16127 14519 16133
rect 15378 16124 15384 16176
rect 15436 16164 15442 16176
rect 15948 16164 15976 16204
rect 27154 16192 27160 16204
rect 27212 16192 27218 16244
rect 27430 16232 27436 16244
rect 27391 16204 27436 16232
rect 27430 16192 27436 16204
rect 27488 16192 27494 16244
rect 28258 16192 28264 16244
rect 28316 16232 28322 16244
rect 28902 16232 28908 16244
rect 28316 16204 28908 16232
rect 28316 16192 28322 16204
rect 28902 16192 28908 16204
rect 28960 16192 28966 16244
rect 29638 16232 29644 16244
rect 29599 16204 29644 16232
rect 29638 16192 29644 16204
rect 29696 16232 29702 16244
rect 36538 16232 36544 16244
rect 29696 16204 30328 16232
rect 29696 16192 29702 16204
rect 30300 16173 30328 16204
rect 30392 16204 36544 16232
rect 15436 16136 15976 16164
rect 15436 16124 15442 16136
rect 11514 16096 11520 16108
rect 11475 16068 11520 16096
rect 11514 16056 11520 16068
rect 11572 16056 11578 16108
rect 15948 16105 15976 16136
rect 16025 16167 16083 16173
rect 16025 16133 16037 16167
rect 16071 16164 16083 16167
rect 16853 16167 16911 16173
rect 16853 16164 16865 16167
rect 16071 16136 16865 16164
rect 16071 16133 16083 16136
rect 16025 16127 16083 16133
rect 16853 16133 16865 16136
rect 16899 16133 16911 16167
rect 30285 16167 30343 16173
rect 16853 16127 16911 16133
rect 22066 16136 29684 16164
rect 14645 16099 14703 16105
rect 14645 16065 14657 16099
rect 14691 16065 14703 16099
rect 14645 16059 14703 16065
rect 15933 16099 15991 16105
rect 15933 16065 15945 16099
rect 15979 16065 15991 16099
rect 16666 16096 16672 16108
rect 16627 16068 16672 16096
rect 15933 16059 15991 16065
rect 11977 16031 12035 16037
rect 11977 15997 11989 16031
rect 12023 15997 12035 16031
rect 14660 16028 14688 16059
rect 16666 16056 16672 16068
rect 16724 16056 16730 16108
rect 18322 16056 18328 16108
rect 18380 16096 18386 16108
rect 18966 16096 18972 16108
rect 18380 16068 18972 16096
rect 18380 16056 18386 16068
rect 18966 16056 18972 16068
rect 19024 16056 19030 16108
rect 20714 16056 20720 16108
rect 20772 16096 20778 16108
rect 20898 16096 20904 16108
rect 20772 16068 20904 16096
rect 20772 16056 20778 16068
rect 20898 16056 20904 16068
rect 20956 16056 20962 16108
rect 16684 16028 16712 16056
rect 18506 16028 18512 16040
rect 14660 16000 16712 16028
rect 18467 16000 18512 16028
rect 11977 15991 12035 15997
rect 14 15920 20 15972
rect 72 15960 78 15972
rect 11992 15960 12020 15991
rect 18506 15988 18512 16000
rect 18564 15988 18570 16040
rect 19518 16028 19524 16040
rect 19479 16000 19524 16028
rect 19518 15988 19524 16000
rect 19576 16028 19582 16040
rect 20070 16028 20076 16040
rect 19576 16000 20076 16028
rect 19576 15988 19582 16000
rect 20070 15988 20076 16000
rect 20128 16028 20134 16040
rect 22066 16028 22094 16136
rect 25130 16096 25136 16108
rect 25091 16068 25136 16096
rect 25130 16056 25136 16068
rect 25188 16056 25194 16108
rect 25682 16056 25688 16108
rect 25740 16096 25746 16108
rect 28074 16096 28080 16108
rect 25740 16068 28080 16096
rect 25740 16056 25746 16068
rect 28074 16056 28080 16068
rect 28132 16056 28138 16108
rect 28629 16099 28687 16105
rect 28629 16096 28641 16099
rect 28460 16068 28641 16096
rect 20128 16000 22094 16028
rect 20128 15988 20134 16000
rect 26602 15988 26608 16040
rect 26660 16028 26666 16040
rect 26973 16031 27031 16037
rect 26973 16028 26985 16031
rect 26660 16000 26985 16028
rect 26660 15988 26666 16000
rect 26973 15997 26985 16000
rect 27019 15997 27031 16031
rect 26973 15991 27031 15997
rect 72 15932 12020 15960
rect 72 15920 78 15932
rect 20162 15920 20168 15972
rect 20220 15960 20226 15972
rect 20622 15960 20628 15972
rect 20220 15932 20628 15960
rect 20220 15920 20226 15932
rect 20622 15920 20628 15932
rect 20680 15960 20686 15972
rect 21085 15963 21143 15969
rect 21085 15960 21097 15963
rect 20680 15932 21097 15960
rect 20680 15920 20686 15932
rect 21085 15929 21097 15932
rect 21131 15929 21143 15963
rect 21085 15923 21143 15929
rect 13170 15852 13176 15904
rect 13228 15892 13234 15904
rect 23014 15892 23020 15904
rect 13228 15864 23020 15892
rect 13228 15852 13234 15864
rect 23014 15852 23020 15864
rect 23072 15892 23078 15904
rect 25038 15892 25044 15904
rect 23072 15864 25044 15892
rect 23072 15852 23078 15864
rect 25038 15852 25044 15864
rect 25096 15852 25102 15904
rect 25314 15892 25320 15904
rect 25275 15864 25320 15892
rect 25314 15852 25320 15864
rect 25372 15852 25378 15904
rect 26988 15892 27016 15991
rect 27062 15920 27068 15972
rect 27120 15960 27126 15972
rect 27249 15963 27307 15969
rect 27249 15960 27261 15963
rect 27120 15932 27261 15960
rect 27120 15920 27126 15932
rect 27249 15929 27261 15932
rect 27295 15929 27307 15963
rect 27249 15923 27307 15929
rect 27338 15892 27344 15904
rect 26988 15864 27344 15892
rect 27338 15852 27344 15864
rect 27396 15892 27402 15904
rect 28261 15895 28319 15901
rect 28261 15892 28273 15895
rect 27396 15864 28273 15892
rect 27396 15852 27402 15864
rect 28261 15861 28273 15864
rect 28307 15861 28319 15895
rect 28460 15892 28488 16068
rect 28629 16065 28641 16068
rect 28675 16065 28687 16099
rect 28629 16059 28687 16065
rect 28994 16056 29000 16108
rect 29052 16096 29058 16108
rect 29549 16099 29607 16105
rect 29549 16096 29561 16099
rect 29052 16068 29561 16096
rect 29052 16056 29058 16068
rect 29549 16065 29561 16068
rect 29595 16065 29607 16099
rect 29656 16096 29684 16136
rect 30285 16133 30297 16167
rect 30331 16133 30343 16167
rect 30285 16127 30343 16133
rect 30392 16096 30420 16204
rect 36538 16192 36544 16204
rect 36596 16192 36602 16244
rect 30834 16124 30840 16176
rect 30892 16164 30898 16176
rect 31018 16164 31024 16176
rect 30892 16136 31024 16164
rect 30892 16124 30898 16136
rect 31018 16124 31024 16136
rect 31076 16124 31082 16176
rect 31938 16164 31944 16176
rect 31404 16136 31944 16164
rect 29656 16068 30420 16096
rect 29549 16059 29607 16065
rect 30742 16056 30748 16108
rect 30800 16096 30806 16108
rect 31404 16105 31432 16136
rect 31938 16124 31944 16136
rect 31996 16124 32002 16176
rect 31205 16099 31263 16105
rect 31205 16096 31217 16099
rect 30800 16068 31217 16096
rect 30800 16056 30806 16068
rect 31205 16065 31217 16068
rect 31251 16065 31263 16099
rect 31205 16059 31263 16065
rect 31297 16099 31355 16105
rect 31297 16065 31309 16099
rect 31343 16065 31355 16099
rect 31297 16059 31355 16065
rect 31389 16099 31447 16105
rect 31389 16065 31401 16099
rect 31435 16065 31447 16099
rect 31570 16096 31576 16108
rect 31531 16068 31576 16096
rect 31389 16059 31447 16065
rect 28718 16028 28724 16040
rect 28679 16000 28724 16028
rect 28718 15988 28724 16000
rect 28776 15988 28782 16040
rect 28813 16031 28871 16037
rect 28813 15997 28825 16031
rect 28859 15997 28871 16031
rect 28813 15991 28871 15997
rect 28534 15920 28540 15972
rect 28592 15960 28598 15972
rect 28828 15960 28856 15991
rect 29178 15988 29184 16040
rect 29236 16028 29242 16040
rect 30834 16028 30840 16040
rect 29236 16000 30840 16028
rect 29236 15988 29242 16000
rect 30834 15988 30840 16000
rect 30892 15988 30898 16040
rect 31018 15988 31024 16040
rect 31076 16028 31082 16040
rect 31312 16028 31340 16059
rect 31570 16056 31576 16068
rect 31628 16056 31634 16108
rect 32122 16096 32128 16108
rect 32083 16068 32128 16096
rect 32122 16056 32128 16068
rect 32180 16056 32186 16108
rect 32214 16056 32220 16108
rect 32272 16096 32278 16108
rect 32381 16099 32439 16105
rect 32381 16096 32393 16099
rect 32272 16068 32393 16096
rect 32272 16056 32278 16068
rect 32381 16065 32393 16068
rect 32427 16065 32439 16099
rect 32381 16059 32439 16065
rect 31076 16000 31340 16028
rect 31076 15988 31082 16000
rect 31478 15988 31484 16040
rect 31536 16028 31542 16040
rect 32140 16028 32168 16056
rect 31536 16000 32168 16028
rect 31536 15988 31542 16000
rect 28592 15932 28856 15960
rect 28592 15920 28598 15932
rect 29086 15920 29092 15972
rect 29144 15960 29150 15972
rect 46750 15960 46756 15972
rect 29144 15932 32168 15960
rect 29144 15920 29150 15932
rect 29178 15892 29184 15904
rect 28460 15864 29184 15892
rect 28261 15855 28319 15861
rect 29178 15852 29184 15864
rect 29236 15852 29242 15904
rect 29546 15852 29552 15904
rect 29604 15892 29610 15904
rect 30377 15895 30435 15901
rect 30377 15892 30389 15895
rect 29604 15864 30389 15892
rect 29604 15852 29610 15864
rect 30377 15861 30389 15864
rect 30423 15861 30435 15895
rect 30377 15855 30435 15861
rect 30929 15895 30987 15901
rect 30929 15861 30941 15895
rect 30975 15892 30987 15895
rect 31754 15892 31760 15904
rect 30975 15864 31760 15892
rect 30975 15861 30987 15864
rect 30929 15855 30987 15861
rect 31754 15852 31760 15864
rect 31812 15852 31818 15904
rect 32140 15892 32168 15932
rect 33060 15932 46756 15960
rect 33060 15892 33088 15932
rect 46750 15920 46756 15932
rect 46808 15920 46814 15972
rect 33502 15892 33508 15904
rect 32140 15864 33088 15892
rect 33463 15864 33508 15892
rect 33502 15852 33508 15864
rect 33560 15852 33566 15904
rect 46290 15852 46296 15904
rect 46348 15892 46354 15904
rect 47765 15895 47823 15901
rect 47765 15892 47777 15895
rect 46348 15864 47777 15892
rect 46348 15852 46354 15864
rect 47765 15861 47777 15864
rect 47811 15861 47823 15895
rect 47765 15855 47823 15861
rect 1104 15802 48852 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 48852 15802
rect 1104 15728 48852 15750
rect 19518 15688 19524 15700
rect 2746 15660 19524 15688
rect 2406 15580 2412 15632
rect 2464 15620 2470 15632
rect 2746 15620 2774 15660
rect 19518 15648 19524 15660
rect 19576 15648 19582 15700
rect 20993 15691 21051 15697
rect 20993 15657 21005 15691
rect 21039 15688 21051 15691
rect 21174 15688 21180 15700
rect 21039 15660 21180 15688
rect 21039 15657 21051 15660
rect 20993 15651 21051 15657
rect 21174 15648 21180 15660
rect 21232 15648 21238 15700
rect 22554 15688 22560 15700
rect 22515 15660 22560 15688
rect 22554 15648 22560 15660
rect 22612 15648 22618 15700
rect 25038 15648 25044 15700
rect 25096 15688 25102 15700
rect 25133 15691 25191 15697
rect 25133 15688 25145 15691
rect 25096 15660 25145 15688
rect 25096 15648 25102 15660
rect 25133 15657 25145 15660
rect 25179 15657 25191 15691
rect 25133 15651 25191 15657
rect 26694 15648 26700 15700
rect 26752 15688 26758 15700
rect 26789 15691 26847 15697
rect 26789 15688 26801 15691
rect 26752 15660 26801 15688
rect 26752 15648 26758 15660
rect 26789 15657 26801 15660
rect 26835 15657 26847 15691
rect 27430 15688 27436 15700
rect 27391 15660 27436 15688
rect 26789 15651 26847 15657
rect 27430 15648 27436 15660
rect 27488 15648 27494 15700
rect 27540 15660 46520 15688
rect 2464 15592 2774 15620
rect 2464 15580 2470 15592
rect 18690 15580 18696 15632
rect 18748 15620 18754 15632
rect 27540 15620 27568 15660
rect 29086 15620 29092 15632
rect 18748 15592 27568 15620
rect 27632 15592 29092 15620
rect 18748 15580 18754 15592
rect 7650 15512 7656 15564
rect 7708 15552 7714 15564
rect 18049 15555 18107 15561
rect 18049 15552 18061 15555
rect 7708 15524 18061 15552
rect 7708 15512 7714 15524
rect 18049 15521 18061 15524
rect 18095 15552 18107 15555
rect 18414 15552 18420 15564
rect 18095 15524 18420 15552
rect 18095 15521 18107 15524
rect 18049 15515 18107 15521
rect 18414 15512 18420 15524
rect 18472 15552 18478 15564
rect 27632 15552 27660 15592
rect 29086 15580 29092 15592
rect 29144 15580 29150 15632
rect 32858 15620 32864 15632
rect 32819 15592 32864 15620
rect 32858 15580 32864 15592
rect 32916 15580 32922 15632
rect 18472 15524 27660 15552
rect 18472 15512 18478 15524
rect 28074 15512 28080 15564
rect 28132 15552 28138 15564
rect 28629 15555 28687 15561
rect 28629 15552 28641 15555
rect 28132 15524 28641 15552
rect 28132 15512 28138 15524
rect 28629 15521 28641 15524
rect 28675 15521 28687 15555
rect 46290 15552 46296 15564
rect 46251 15524 46296 15552
rect 28629 15515 28687 15521
rect 46290 15512 46296 15524
rect 46348 15512 46354 15564
rect 46492 15561 46520 15660
rect 46477 15555 46535 15561
rect 46477 15521 46489 15555
rect 46523 15521 46535 15555
rect 48130 15552 48136 15564
rect 48091 15524 48136 15552
rect 46477 15515 46535 15521
rect 48130 15512 48136 15524
rect 48188 15512 48194 15564
rect 17865 15487 17923 15493
rect 17865 15453 17877 15487
rect 17911 15484 17923 15487
rect 18322 15484 18328 15496
rect 17911 15456 18328 15484
rect 17911 15453 17923 15456
rect 17865 15447 17923 15453
rect 18322 15444 18328 15456
rect 18380 15484 18386 15496
rect 19705 15487 19763 15493
rect 19705 15484 19717 15487
rect 18380 15456 19717 15484
rect 18380 15444 18386 15456
rect 19705 15453 19717 15456
rect 19751 15453 19763 15487
rect 20714 15484 20720 15496
rect 20675 15456 20720 15484
rect 19705 15447 19763 15453
rect 20714 15444 20720 15456
rect 20772 15444 20778 15496
rect 20809 15487 20867 15493
rect 20809 15453 20821 15487
rect 20855 15484 20867 15487
rect 20898 15484 20904 15496
rect 20855 15456 20904 15484
rect 20855 15453 20867 15456
rect 20809 15447 20867 15453
rect 20898 15444 20904 15456
rect 20956 15444 20962 15496
rect 21082 15484 21088 15496
rect 21043 15456 21088 15484
rect 21082 15444 21088 15456
rect 21140 15444 21146 15496
rect 24854 15444 24860 15496
rect 24912 15484 24918 15496
rect 25041 15487 25099 15493
rect 25041 15484 25053 15487
rect 24912 15456 25053 15484
rect 24912 15444 24918 15456
rect 25041 15453 25053 15456
rect 25087 15453 25099 15487
rect 26602 15484 26608 15496
rect 26563 15456 26608 15484
rect 25041 15447 25099 15453
rect 26602 15444 26608 15456
rect 26660 15444 26666 15496
rect 26878 15484 26884 15496
rect 26839 15456 26884 15484
rect 26878 15444 26884 15456
rect 26936 15444 26942 15496
rect 27341 15487 27399 15493
rect 27341 15453 27353 15487
rect 27387 15453 27399 15487
rect 27341 15447 27399 15453
rect 27433 15487 27491 15493
rect 27433 15453 27445 15487
rect 27479 15453 27491 15487
rect 28261 15487 28319 15493
rect 28261 15484 28273 15487
rect 27433 15447 27491 15453
rect 27724 15456 28273 15484
rect 22373 15419 22431 15425
rect 22373 15385 22385 15419
rect 22419 15416 22431 15419
rect 24872 15416 24900 15444
rect 22419 15388 24900 15416
rect 26421 15419 26479 15425
rect 22419 15385 22431 15388
rect 22373 15379 22431 15385
rect 26421 15385 26433 15419
rect 26467 15416 26479 15419
rect 27356 15416 27384 15447
rect 26467 15388 27384 15416
rect 26467 15385 26479 15388
rect 26421 15379 26479 15385
rect 19426 15308 19432 15360
rect 19484 15348 19490 15360
rect 19797 15351 19855 15357
rect 19797 15348 19809 15351
rect 19484 15320 19809 15348
rect 19484 15308 19490 15320
rect 19797 15317 19809 15320
rect 19843 15317 19855 15351
rect 20530 15348 20536 15360
rect 20491 15320 20536 15348
rect 19797 15311 19855 15317
rect 20530 15308 20536 15320
rect 20588 15308 20594 15360
rect 22186 15308 22192 15360
rect 22244 15348 22250 15360
rect 22573 15351 22631 15357
rect 22573 15348 22585 15351
rect 22244 15320 22585 15348
rect 22244 15308 22250 15320
rect 22573 15317 22585 15320
rect 22619 15317 22631 15351
rect 22573 15311 22631 15317
rect 22741 15351 22799 15357
rect 22741 15317 22753 15351
rect 22787 15348 22799 15351
rect 23566 15348 23572 15360
rect 22787 15320 23572 15348
rect 22787 15317 22799 15320
rect 22741 15311 22799 15317
rect 23566 15308 23572 15320
rect 23624 15308 23630 15360
rect 23658 15308 23664 15360
rect 23716 15348 23722 15360
rect 24946 15348 24952 15360
rect 23716 15320 24952 15348
rect 23716 15308 23722 15320
rect 24946 15308 24952 15320
rect 25004 15308 25010 15360
rect 25866 15308 25872 15360
rect 25924 15348 25930 15360
rect 26142 15348 26148 15360
rect 25924 15320 26148 15348
rect 25924 15308 25930 15320
rect 26142 15308 26148 15320
rect 26200 15348 26206 15360
rect 27448 15348 27476 15447
rect 27724 15357 27752 15456
rect 28261 15453 28273 15456
rect 28307 15453 28319 15487
rect 28261 15447 28319 15453
rect 28350 15444 28356 15496
rect 28408 15484 28414 15496
rect 28445 15487 28503 15493
rect 28445 15484 28457 15487
rect 28408 15456 28457 15484
rect 28408 15444 28414 15456
rect 28445 15453 28457 15456
rect 28491 15453 28503 15487
rect 28445 15447 28503 15453
rect 28537 15487 28595 15493
rect 28537 15453 28549 15487
rect 28583 15453 28595 15487
rect 28537 15447 28595 15453
rect 28813 15487 28871 15493
rect 28813 15453 28825 15487
rect 28859 15484 28871 15487
rect 29178 15484 29184 15496
rect 28859 15456 29184 15484
rect 28859 15453 28871 15456
rect 28813 15447 28871 15453
rect 26200 15320 27476 15348
rect 27709 15351 27767 15357
rect 26200 15308 26206 15320
rect 27709 15317 27721 15351
rect 27755 15317 27767 15351
rect 28552 15348 28580 15447
rect 29178 15444 29184 15456
rect 29236 15444 29242 15496
rect 29546 15484 29552 15496
rect 29507 15456 29552 15484
rect 29546 15444 29552 15456
rect 29604 15484 29610 15496
rect 31110 15484 31116 15496
rect 29604 15456 31116 15484
rect 29604 15444 29610 15456
rect 31110 15444 31116 15456
rect 31168 15484 31174 15496
rect 31478 15484 31484 15496
rect 31168 15456 31484 15484
rect 31168 15444 31174 15456
rect 31478 15444 31484 15456
rect 31536 15444 31542 15496
rect 31754 15493 31760 15496
rect 31748 15447 31760 15493
rect 31812 15484 31818 15496
rect 31812 15456 31848 15484
rect 31754 15444 31760 15447
rect 31812 15444 31818 15456
rect 28997 15419 29055 15425
rect 28997 15385 29009 15419
rect 29043 15416 29055 15419
rect 29794 15419 29852 15425
rect 29794 15416 29806 15419
rect 29043 15388 29806 15416
rect 29043 15385 29055 15388
rect 28997 15379 29055 15385
rect 29794 15385 29806 15388
rect 29840 15385 29852 15419
rect 29794 15379 29852 15385
rect 28718 15348 28724 15360
rect 28552 15320 28724 15348
rect 27709 15311 27767 15317
rect 28718 15308 28724 15320
rect 28776 15348 28782 15360
rect 30929 15351 30987 15357
rect 30929 15348 30941 15351
rect 28776 15320 30941 15348
rect 28776 15308 28782 15320
rect 30929 15317 30941 15320
rect 30975 15317 30987 15351
rect 30929 15311 30987 15317
rect 1104 15258 48852 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 48852 15258
rect 1104 15184 48852 15206
rect 20257 15147 20315 15153
rect 20257 15113 20269 15147
rect 20303 15144 20315 15147
rect 20530 15144 20536 15156
rect 20303 15116 20536 15144
rect 20303 15113 20315 15116
rect 20257 15107 20315 15113
rect 20530 15104 20536 15116
rect 20588 15104 20594 15156
rect 20714 15104 20720 15156
rect 20772 15144 20778 15156
rect 21177 15147 21235 15153
rect 21177 15144 21189 15147
rect 20772 15116 21189 15144
rect 20772 15104 20778 15116
rect 21177 15113 21189 15116
rect 21223 15113 21235 15147
rect 22186 15144 22192 15156
rect 22147 15116 22192 15144
rect 21177 15107 21235 15113
rect 22186 15104 22192 15116
rect 22244 15104 22250 15156
rect 22554 15104 22560 15156
rect 22612 15144 22618 15156
rect 22741 15147 22799 15153
rect 22741 15144 22753 15147
rect 22612 15116 22753 15144
rect 22612 15104 22618 15116
rect 22741 15113 22753 15116
rect 22787 15113 22799 15147
rect 22741 15107 22799 15113
rect 30929 15147 30987 15153
rect 30929 15113 30941 15147
rect 30975 15144 30987 15147
rect 32214 15144 32220 15156
rect 30975 15116 32220 15144
rect 30975 15113 30987 15116
rect 30929 15107 30987 15113
rect 32214 15104 32220 15116
rect 32272 15104 32278 15156
rect 46658 15104 46664 15156
rect 46716 15144 46722 15156
rect 46845 15147 46903 15153
rect 46845 15144 46857 15147
rect 46716 15116 46857 15144
rect 46716 15104 46722 15116
rect 46845 15113 46857 15116
rect 46891 15113 46903 15147
rect 46845 15107 46903 15113
rect 17678 15076 17684 15088
rect 17639 15048 17684 15076
rect 17678 15036 17684 15048
rect 17736 15036 17742 15088
rect 19150 15076 19156 15088
rect 19111 15048 19156 15076
rect 19150 15036 19156 15048
rect 19208 15036 19214 15088
rect 20165 15079 20223 15085
rect 20165 15045 20177 15079
rect 20211 15076 20223 15079
rect 21634 15076 21640 15088
rect 20211 15048 21640 15076
rect 20211 15045 20223 15048
rect 20165 15039 20223 15045
rect 21634 15036 21640 15048
rect 21692 15036 21698 15088
rect 21821 15079 21879 15085
rect 21821 15045 21833 15079
rect 21867 15076 21879 15079
rect 22094 15076 22100 15088
rect 21867 15048 22100 15076
rect 21867 15045 21879 15048
rect 21821 15039 21879 15045
rect 22094 15036 22100 15048
rect 22152 15076 22158 15088
rect 22152 15048 22692 15076
rect 22152 15036 22158 15048
rect 18322 15008 18328 15020
rect 18283 14980 18328 15008
rect 18322 14968 18328 14980
rect 18380 14968 18386 15020
rect 21085 15011 21143 15017
rect 21085 14977 21097 15011
rect 21131 15008 21143 15011
rect 21174 15008 21180 15020
rect 21131 14980 21180 15008
rect 21131 14977 21143 14980
rect 21085 14971 21143 14977
rect 21174 14968 21180 14980
rect 21232 14968 21238 15020
rect 22664 15017 22692 15048
rect 23382 15036 23388 15088
rect 23440 15076 23446 15088
rect 24029 15079 24087 15085
rect 24029 15076 24041 15079
rect 23440 15048 24041 15076
rect 23440 15036 23446 15048
rect 24029 15045 24041 15048
rect 24075 15045 24087 15079
rect 24029 15039 24087 15045
rect 31018 15036 31024 15088
rect 31076 15076 31082 15088
rect 32309 15079 32367 15085
rect 31076 15048 31340 15076
rect 31076 15036 31082 15048
rect 21269 15011 21327 15017
rect 21269 14977 21281 15011
rect 21315 14977 21327 15011
rect 21269 14971 21327 14977
rect 22005 15011 22063 15017
rect 22005 14977 22017 15011
rect 22051 15008 22063 15011
rect 22649 15011 22707 15017
rect 22051 14980 22416 15008
rect 22051 14977 22063 14980
rect 22005 14971 22063 14977
rect 2866 14900 2872 14952
rect 2924 14940 2930 14952
rect 19150 14940 19156 14952
rect 2924 14912 19156 14940
rect 2924 14900 2930 14912
rect 19150 14900 19156 14912
rect 19208 14900 19214 14952
rect 20441 14943 20499 14949
rect 20441 14909 20453 14943
rect 20487 14909 20499 14943
rect 20441 14903 20499 14909
rect 17862 14872 17868 14884
rect 17823 14844 17868 14872
rect 17862 14832 17868 14844
rect 17920 14832 17926 14884
rect 20456 14872 20484 14903
rect 20714 14900 20720 14952
rect 20772 14940 20778 14952
rect 21284 14940 21312 14971
rect 22186 14940 22192 14952
rect 20772 14912 22192 14940
rect 20772 14900 20778 14912
rect 22186 14900 22192 14912
rect 22244 14900 22250 14952
rect 22388 14940 22416 14980
rect 22649 14977 22661 15011
rect 22695 14977 22707 15011
rect 22649 14971 22707 14977
rect 22833 15011 22891 15017
rect 22833 14977 22845 15011
rect 22879 15008 22891 15011
rect 23566 15008 23572 15020
rect 22879 14980 22913 15008
rect 23527 14980 23572 15008
rect 22879 14977 22891 14980
rect 22833 14971 22891 14977
rect 22848 14940 22876 14971
rect 23566 14968 23572 14980
rect 23624 14968 23630 15020
rect 23661 15011 23719 15017
rect 23661 14977 23673 15011
rect 23707 15008 23719 15011
rect 24578 15008 24584 15020
rect 23707 14980 24584 15008
rect 23707 14977 23719 14980
rect 23661 14971 23719 14977
rect 24578 14968 24584 14980
rect 24636 14968 24642 15020
rect 25130 15008 25136 15020
rect 25091 14980 25136 15008
rect 25130 14968 25136 14980
rect 25188 14968 25194 15020
rect 25958 14968 25964 15020
rect 26016 15008 26022 15020
rect 27341 15011 27399 15017
rect 27341 15008 27353 15011
rect 26016 14980 27353 15008
rect 26016 14968 26022 14980
rect 27341 14977 27353 14980
rect 27387 14977 27399 15011
rect 27341 14971 27399 14977
rect 27617 15011 27675 15017
rect 27617 14977 27629 15011
rect 27663 15008 27675 15011
rect 27982 15008 27988 15020
rect 27663 14980 27988 15008
rect 27663 14977 27675 14980
rect 27617 14971 27675 14977
rect 27982 14968 27988 14980
rect 28040 15008 28046 15020
rect 28442 15008 28448 15020
rect 28040 14980 28448 15008
rect 28040 14968 28046 14980
rect 28442 14968 28448 14980
rect 28500 14968 28506 15020
rect 30834 14968 30840 15020
rect 30892 15008 30898 15020
rect 31312 15017 31340 15048
rect 32309 15045 32321 15079
rect 32355 15076 32367 15079
rect 33502 15076 33508 15088
rect 32355 15048 33508 15076
rect 32355 15045 32367 15048
rect 32309 15039 32367 15045
rect 33502 15036 33508 15048
rect 33560 15036 33566 15088
rect 31205 15011 31263 15017
rect 31205 15008 31217 15011
rect 30892 14980 31217 15008
rect 30892 14968 30898 14980
rect 31205 14977 31217 14980
rect 31251 14977 31263 15011
rect 31205 14971 31263 14977
rect 31297 15011 31355 15017
rect 31297 14977 31309 15011
rect 31343 14977 31355 15011
rect 31297 14971 31355 14977
rect 31389 15011 31447 15017
rect 31389 14977 31401 15011
rect 31435 14977 31447 15011
rect 31570 15008 31576 15020
rect 31531 14980 31576 15008
rect 31389 14971 31447 14977
rect 22922 14940 22928 14952
rect 22388 14912 22928 14940
rect 22922 14900 22928 14912
rect 22980 14900 22986 14952
rect 23937 14943 23995 14949
rect 23937 14909 23949 14943
rect 23983 14940 23995 14943
rect 27522 14940 27528 14952
rect 23983 14912 27528 14940
rect 23983 14909 23995 14912
rect 23937 14903 23995 14909
rect 21450 14872 21456 14884
rect 20456 14844 21456 14872
rect 21450 14832 21456 14844
rect 21508 14832 21514 14884
rect 22278 14832 22284 14884
rect 22336 14872 22342 14884
rect 23952 14872 23980 14903
rect 27522 14900 27528 14912
rect 27580 14900 27586 14952
rect 31404 14940 31432 14971
rect 31570 14968 31576 14980
rect 31628 14968 31634 15020
rect 31662 14968 31668 15020
rect 31720 15008 31726 15020
rect 32125 15011 32183 15017
rect 32125 15008 32137 15011
rect 31720 14980 32137 15008
rect 31720 14968 31726 14980
rect 32125 14977 32137 14980
rect 32171 14977 32183 15011
rect 32125 14971 32183 14977
rect 46842 14968 46848 15020
rect 46900 15008 46906 15020
rect 47029 15011 47087 15017
rect 47029 15008 47041 15011
rect 46900 14980 47041 15008
rect 46900 14968 46906 14980
rect 47029 14977 47041 14980
rect 47075 14977 47087 15011
rect 47578 15008 47584 15020
rect 47539 14980 47584 15008
rect 47029 14971 47087 14977
rect 47578 14968 47584 14980
rect 47636 14968 47642 15020
rect 32493 14943 32551 14949
rect 32493 14940 32505 14943
rect 31404 14912 32505 14940
rect 32493 14909 32505 14912
rect 32539 14909 32551 14943
rect 32493 14903 32551 14909
rect 22336 14844 23980 14872
rect 22336 14832 22342 14844
rect 24946 14832 24952 14884
rect 25004 14872 25010 14884
rect 28258 14872 28264 14884
rect 25004 14844 28264 14872
rect 25004 14832 25010 14844
rect 28258 14832 28264 14844
rect 28316 14832 28322 14884
rect 19426 14764 19432 14816
rect 19484 14804 19490 14816
rect 19797 14807 19855 14813
rect 19797 14804 19809 14807
rect 19484 14776 19809 14804
rect 19484 14764 19490 14776
rect 19797 14773 19809 14776
rect 19843 14773 19855 14807
rect 19797 14767 19855 14773
rect 20622 14764 20628 14816
rect 20680 14804 20686 14816
rect 22296 14804 22324 14832
rect 20680 14776 22324 14804
rect 23385 14807 23443 14813
rect 20680 14764 20686 14776
rect 23385 14773 23397 14807
rect 23431 14804 23443 14807
rect 23474 14804 23480 14816
rect 23431 14776 23480 14804
rect 23431 14773 23443 14776
rect 23385 14767 23443 14773
rect 23474 14764 23480 14776
rect 23532 14764 23538 14816
rect 24854 14764 24860 14816
rect 24912 14804 24918 14816
rect 25317 14807 25375 14813
rect 25317 14804 25329 14807
rect 24912 14776 25329 14804
rect 24912 14764 24918 14776
rect 25317 14773 25329 14776
rect 25363 14773 25375 14807
rect 27154 14804 27160 14816
rect 27115 14776 27160 14804
rect 25317 14767 25375 14773
rect 27154 14764 27160 14776
rect 27212 14764 27218 14816
rect 27525 14807 27583 14813
rect 27525 14773 27537 14807
rect 27571 14804 27583 14807
rect 27614 14804 27620 14816
rect 27571 14776 27620 14804
rect 27571 14773 27583 14776
rect 27525 14767 27583 14773
rect 27614 14764 27620 14776
rect 27672 14764 27678 14816
rect 46474 14764 46480 14816
rect 46532 14804 46538 14816
rect 47673 14807 47731 14813
rect 47673 14804 47685 14807
rect 46532 14776 47685 14804
rect 46532 14764 46538 14776
rect 47673 14773 47685 14776
rect 47719 14773 47731 14807
rect 47673 14767 47731 14773
rect 1104 14714 48852 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 48852 14714
rect 1104 14640 48852 14662
rect 20073 14603 20131 14609
rect 20073 14569 20085 14603
rect 20119 14600 20131 14603
rect 20898 14600 20904 14612
rect 20119 14572 20904 14600
rect 20119 14569 20131 14572
rect 20073 14563 20131 14569
rect 20898 14560 20904 14572
rect 20956 14560 20962 14612
rect 20993 14603 21051 14609
rect 20993 14569 21005 14603
rect 21039 14600 21051 14603
rect 21174 14600 21180 14612
rect 21039 14572 21180 14600
rect 21039 14569 21051 14572
rect 20993 14563 21051 14569
rect 20530 14532 20536 14544
rect 20272 14504 20536 14532
rect 17954 14464 17960 14476
rect 17144 14436 17960 14464
rect 17144 14405 17172 14436
rect 17954 14424 17960 14436
rect 18012 14464 18018 14476
rect 20162 14464 20168 14476
rect 18012 14436 20168 14464
rect 18012 14424 18018 14436
rect 20162 14424 20168 14436
rect 20220 14424 20226 14476
rect 17129 14399 17187 14405
rect 17129 14365 17141 14399
rect 17175 14365 17187 14399
rect 19426 14396 19432 14408
rect 19387 14368 19432 14396
rect 17129 14359 17187 14365
rect 19426 14356 19432 14368
rect 19484 14356 19490 14408
rect 17957 14331 18015 14337
rect 17957 14297 17969 14331
rect 18003 14328 18015 14331
rect 19610 14328 19616 14340
rect 18003 14300 19616 14328
rect 18003 14297 18015 14300
rect 17957 14291 18015 14297
rect 19610 14288 19616 14300
rect 19668 14288 19674 14340
rect 17310 14260 17316 14272
rect 17271 14232 17316 14260
rect 17310 14220 17316 14232
rect 17368 14220 17374 14272
rect 17402 14220 17408 14272
rect 17460 14260 17466 14272
rect 17586 14260 17592 14272
rect 17460 14232 17592 14260
rect 17460 14220 17466 14232
rect 17586 14220 17592 14232
rect 17644 14260 17650 14272
rect 18049 14263 18107 14269
rect 18049 14260 18061 14263
rect 17644 14232 18061 14260
rect 17644 14220 17650 14232
rect 18049 14229 18061 14232
rect 18095 14229 18107 14263
rect 19242 14260 19248 14272
rect 19203 14232 19248 14260
rect 18049 14223 18107 14229
rect 19242 14220 19248 14232
rect 19300 14220 19306 14272
rect 20180 14260 20208 14424
rect 20272 14405 20300 14504
rect 20530 14492 20536 14504
rect 20588 14492 20594 14544
rect 21008 14464 21036 14563
rect 21174 14560 21180 14572
rect 21232 14600 21238 14612
rect 21450 14600 21456 14612
rect 21232 14572 21456 14600
rect 21232 14560 21238 14572
rect 21450 14560 21456 14572
rect 21508 14560 21514 14612
rect 23106 14560 23112 14612
rect 23164 14600 23170 14612
rect 24578 14600 24584 14612
rect 23164 14572 24440 14600
rect 24539 14572 24584 14600
rect 23164 14560 23170 14572
rect 21266 14492 21272 14544
rect 21324 14532 21330 14544
rect 23385 14535 23443 14541
rect 23385 14532 23397 14535
rect 21324 14504 23397 14532
rect 21324 14492 21330 14504
rect 23385 14501 23397 14504
rect 23431 14501 23443 14535
rect 23658 14532 23664 14544
rect 23385 14495 23443 14501
rect 23483 14504 23664 14532
rect 20548 14436 21036 14464
rect 21637 14467 21695 14473
rect 20548 14405 20576 14436
rect 21637 14433 21649 14467
rect 21683 14464 21695 14467
rect 22738 14464 22744 14476
rect 21683 14436 22744 14464
rect 21683 14433 21695 14436
rect 21637 14427 21695 14433
rect 22738 14424 22744 14436
rect 22796 14424 22802 14476
rect 23483 14464 23511 14504
rect 23658 14492 23664 14504
rect 23716 14532 23722 14544
rect 23842 14532 23848 14544
rect 23716 14504 23848 14532
rect 23716 14492 23722 14504
rect 23842 14492 23848 14504
rect 23900 14492 23906 14544
rect 23400 14436 23511 14464
rect 24412 14464 24440 14572
rect 24578 14560 24584 14572
rect 24636 14560 24642 14612
rect 24670 14560 24676 14612
rect 24728 14600 24734 14612
rect 25317 14603 25375 14609
rect 25317 14600 25329 14603
rect 24728 14572 25329 14600
rect 24728 14560 24734 14572
rect 25317 14569 25329 14572
rect 25363 14600 25375 14603
rect 26878 14600 26884 14612
rect 25363 14572 26884 14600
rect 25363 14569 25375 14572
rect 25317 14563 25375 14569
rect 26878 14560 26884 14572
rect 26936 14560 26942 14612
rect 27062 14560 27068 14612
rect 27120 14600 27126 14612
rect 27430 14600 27436 14612
rect 27120 14572 27436 14600
rect 27120 14560 27126 14572
rect 27430 14560 27436 14572
rect 27488 14600 27494 14612
rect 28169 14603 28227 14609
rect 28169 14600 28181 14603
rect 27488 14572 28181 14600
rect 27488 14560 27494 14572
rect 28169 14569 28181 14572
rect 28215 14569 28227 14603
rect 28169 14563 28227 14569
rect 24489 14535 24547 14541
rect 24489 14501 24501 14535
rect 24535 14532 24547 14535
rect 25682 14532 25688 14544
rect 24535 14504 25688 14532
rect 24535 14501 24547 14504
rect 24489 14495 24547 14501
rect 25682 14492 25688 14504
rect 25740 14532 25746 14544
rect 26142 14532 26148 14544
rect 25740 14504 26148 14532
rect 25740 14492 25746 14504
rect 26142 14492 26148 14504
rect 26200 14492 26206 14544
rect 26329 14535 26387 14541
rect 26329 14501 26341 14535
rect 26375 14532 26387 14535
rect 28442 14532 28448 14544
rect 26375 14504 28448 14532
rect 26375 14501 26387 14504
rect 26329 14495 26387 14501
rect 28442 14492 28448 14504
rect 28500 14532 28506 14544
rect 28902 14532 28908 14544
rect 28500 14504 28908 14532
rect 28500 14492 28506 14504
rect 28902 14492 28908 14504
rect 28960 14492 28966 14544
rect 24673 14467 24731 14473
rect 24412 14436 24521 14464
rect 20257 14399 20315 14405
rect 20257 14365 20269 14399
rect 20303 14365 20315 14399
rect 20257 14359 20315 14365
rect 20533 14399 20591 14405
rect 20533 14365 20545 14399
rect 20579 14365 20591 14399
rect 20533 14359 20591 14365
rect 20806 14356 20812 14408
rect 20864 14396 20870 14408
rect 21174 14396 21180 14408
rect 20864 14368 21180 14396
rect 20864 14356 20870 14368
rect 21174 14356 21180 14368
rect 21232 14396 21238 14408
rect 23106 14396 23112 14408
rect 21232 14368 23112 14396
rect 21232 14356 21238 14368
rect 23106 14356 23112 14368
rect 23164 14356 23170 14408
rect 20441 14331 20499 14337
rect 20441 14297 20453 14331
rect 20487 14328 20499 14331
rect 20714 14328 20720 14340
rect 20487 14300 20720 14328
rect 20487 14297 20499 14300
rect 20441 14291 20499 14297
rect 20714 14288 20720 14300
rect 20772 14288 20778 14340
rect 21082 14288 21088 14340
rect 21140 14328 21146 14340
rect 21361 14331 21419 14337
rect 21361 14328 21373 14331
rect 21140 14300 21373 14328
rect 21140 14288 21146 14300
rect 21361 14297 21373 14300
rect 21407 14328 21419 14331
rect 22002 14328 22008 14340
rect 21407 14300 22008 14328
rect 21407 14297 21419 14300
rect 21361 14291 21419 14297
rect 22002 14288 22008 14300
rect 22060 14288 22066 14340
rect 22462 14288 22468 14340
rect 22520 14328 22526 14340
rect 22649 14331 22707 14337
rect 22649 14328 22661 14331
rect 22520 14300 22661 14328
rect 22520 14288 22526 14300
rect 22649 14297 22661 14300
rect 22695 14297 22707 14331
rect 23290 14328 23296 14340
rect 22649 14291 22707 14297
rect 22756 14300 23296 14328
rect 20898 14260 20904 14272
rect 20180 14232 20904 14260
rect 20898 14220 20904 14232
rect 20956 14220 20962 14272
rect 21453 14263 21511 14269
rect 21453 14229 21465 14263
rect 21499 14260 21511 14263
rect 21634 14260 21640 14272
rect 21499 14232 21640 14260
rect 21499 14229 21511 14232
rect 21453 14223 21511 14229
rect 21634 14220 21640 14232
rect 21692 14220 21698 14272
rect 22186 14260 22192 14272
rect 22147 14232 22192 14260
rect 22186 14220 22192 14232
rect 22244 14220 22250 14272
rect 22557 14263 22615 14269
rect 22557 14229 22569 14263
rect 22603 14260 22615 14263
rect 22756 14260 22784 14300
rect 23290 14288 23296 14300
rect 23348 14288 23354 14340
rect 23400 14337 23428 14436
rect 23670 14399 23728 14405
rect 23670 14365 23682 14399
rect 23716 14396 23728 14399
rect 23716 14368 23796 14396
rect 23716 14365 23728 14368
rect 23670 14359 23728 14365
rect 23385 14331 23443 14337
rect 23385 14297 23397 14331
rect 23431 14297 23443 14331
rect 23768 14328 23796 14368
rect 24026 14356 24032 14408
rect 24084 14396 24090 14408
rect 24397 14399 24455 14405
rect 24397 14396 24409 14399
rect 24084 14368 24409 14396
rect 24084 14356 24090 14368
rect 24397 14365 24409 14368
rect 24443 14365 24455 14399
rect 24493 14396 24521 14436
rect 24673 14433 24685 14467
rect 24719 14464 24731 14467
rect 24946 14464 24952 14476
rect 24719 14436 24952 14464
rect 24719 14433 24731 14436
rect 24673 14427 24731 14433
rect 24946 14424 24952 14436
rect 25004 14424 25010 14476
rect 26694 14424 26700 14476
rect 26752 14464 26758 14476
rect 46474 14464 46480 14476
rect 26752 14436 28212 14464
rect 46435 14436 46480 14464
rect 26752 14424 26758 14436
rect 26145 14399 26203 14405
rect 26145 14396 26157 14399
rect 24493 14368 26157 14396
rect 24397 14359 24455 14365
rect 26145 14365 26157 14368
rect 26191 14365 26203 14399
rect 27154 14396 27160 14408
rect 27115 14368 27160 14396
rect 26145 14359 26203 14365
rect 27154 14356 27160 14368
rect 27212 14356 27218 14408
rect 27522 14396 27528 14408
rect 27483 14368 27528 14396
rect 27522 14356 27528 14368
rect 27580 14356 27586 14408
rect 28184 14405 28212 14436
rect 46474 14424 46480 14436
rect 46532 14424 46538 14476
rect 28169 14399 28227 14405
rect 28169 14365 28181 14399
rect 28215 14365 28227 14399
rect 28350 14396 28356 14408
rect 28311 14368 28356 14396
rect 28169 14359 28227 14365
rect 28350 14356 28356 14368
rect 28408 14356 28414 14408
rect 31478 14396 31484 14408
rect 31439 14368 31484 14396
rect 31478 14356 31484 14368
rect 31536 14356 31542 14408
rect 46293 14399 46351 14405
rect 46293 14365 46305 14399
rect 46339 14365 46351 14399
rect 46293 14359 46351 14365
rect 23385 14291 23443 14297
rect 23483 14300 23796 14328
rect 22603 14232 22784 14260
rect 22603 14229 22615 14232
rect 22557 14223 22615 14229
rect 22830 14220 22836 14272
rect 22888 14260 22894 14272
rect 23483 14260 23511 14300
rect 25038 14288 25044 14340
rect 25096 14328 25102 14340
rect 25225 14331 25283 14337
rect 25225 14328 25237 14331
rect 25096 14300 25237 14328
rect 25096 14288 25102 14300
rect 25225 14297 25237 14300
rect 25271 14297 25283 14331
rect 25225 14291 25283 14297
rect 27341 14331 27399 14337
rect 27341 14297 27353 14331
rect 27387 14297 27399 14331
rect 27341 14291 27399 14297
rect 27433 14331 27491 14337
rect 27433 14297 27445 14331
rect 27479 14297 27491 14331
rect 46308 14328 46336 14359
rect 47670 14328 47676 14340
rect 46308 14300 47676 14328
rect 27433 14291 27491 14297
rect 22888 14232 23511 14260
rect 23569 14263 23627 14269
rect 22888 14220 22894 14232
rect 23569 14229 23581 14263
rect 23615 14260 23627 14263
rect 24394 14260 24400 14272
rect 23615 14232 24400 14260
rect 23615 14229 23627 14232
rect 23569 14223 23627 14229
rect 24394 14220 24400 14232
rect 24452 14260 24458 14272
rect 24670 14260 24676 14272
rect 24452 14232 24676 14260
rect 24452 14220 24458 14232
rect 24670 14220 24676 14232
rect 24728 14220 24734 14272
rect 27154 14220 27160 14272
rect 27212 14260 27218 14272
rect 27356 14260 27384 14291
rect 27212 14232 27384 14260
rect 27448 14260 27476 14291
rect 47670 14288 47676 14300
rect 47728 14288 47734 14340
rect 48130 14328 48136 14340
rect 48091 14300 48136 14328
rect 48130 14288 48136 14300
rect 48188 14288 48194 14340
rect 27614 14260 27620 14272
rect 27448 14232 27620 14260
rect 27212 14220 27218 14232
rect 27614 14220 27620 14232
rect 27672 14220 27678 14272
rect 27709 14263 27767 14269
rect 27709 14229 27721 14263
rect 27755 14260 27767 14263
rect 28074 14260 28080 14272
rect 27755 14232 28080 14260
rect 27755 14229 27767 14232
rect 27709 14223 27767 14229
rect 28074 14220 28080 14232
rect 28132 14220 28138 14272
rect 31573 14263 31631 14269
rect 31573 14229 31585 14263
rect 31619 14260 31631 14263
rect 32398 14260 32404 14272
rect 31619 14232 32404 14260
rect 31619 14229 31631 14232
rect 31573 14223 31631 14229
rect 32398 14220 32404 14232
rect 32456 14220 32462 14272
rect 1104 14170 48852 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 48852 14170
rect 1104 14096 48852 14118
rect 21266 14056 21272 14068
rect 20364 14028 21272 14056
rect 18500 13991 18558 13997
rect 18500 13957 18512 13991
rect 18546 13988 18558 13991
rect 19242 13988 19248 14000
rect 18546 13960 19248 13988
rect 18546 13957 18558 13960
rect 18500 13951 18558 13957
rect 19242 13948 19248 13960
rect 19300 13948 19306 14000
rect 2038 13920 2044 13932
rect 1999 13892 2044 13920
rect 2038 13880 2044 13892
rect 2096 13880 2102 13932
rect 17402 13920 17408 13932
rect 17363 13892 17408 13920
rect 17402 13880 17408 13892
rect 17460 13880 17466 13932
rect 17494 13880 17500 13932
rect 17552 13920 17558 13932
rect 17681 13923 17739 13929
rect 17552 13892 17597 13920
rect 17552 13880 17558 13892
rect 17681 13889 17693 13923
rect 17727 13889 17739 13923
rect 17681 13883 17739 13889
rect 17773 13923 17831 13929
rect 17773 13889 17785 13923
rect 17819 13920 17831 13923
rect 17954 13920 17960 13932
rect 17819 13892 17960 13920
rect 17819 13889 17831 13892
rect 17773 13883 17831 13889
rect 17696 13852 17724 13883
rect 17954 13880 17960 13892
rect 18012 13880 18018 13932
rect 20364 13929 20392 14028
rect 21266 14016 21272 14028
rect 21324 14016 21330 14068
rect 22462 14016 22468 14068
rect 22520 14056 22526 14068
rect 23382 14056 23388 14068
rect 22520 14028 23388 14056
rect 22520 14016 22526 14028
rect 23382 14016 23388 14028
rect 23440 14056 23446 14068
rect 24581 14059 24639 14065
rect 24581 14056 24593 14059
rect 23440 14028 24593 14056
rect 23440 14016 23446 14028
rect 24581 14025 24593 14028
rect 24627 14025 24639 14059
rect 24581 14019 24639 14025
rect 26973 14059 27031 14065
rect 26973 14025 26985 14059
rect 27019 14056 27031 14059
rect 27154 14056 27160 14068
rect 27019 14028 27160 14056
rect 27019 14025 27031 14028
rect 26973 14019 27031 14025
rect 27154 14016 27160 14028
rect 27212 14016 27218 14068
rect 27264 14028 27568 14056
rect 20622 13988 20628 14000
rect 20583 13960 20628 13988
rect 20622 13948 20628 13960
rect 20680 13948 20686 14000
rect 20717 13991 20775 13997
rect 20717 13957 20729 13991
rect 20763 13988 20775 13991
rect 20763 13960 21036 13988
rect 20763 13957 20775 13960
rect 20717 13951 20775 13957
rect 20530 13929 20536 13932
rect 20349 13923 20407 13929
rect 20349 13889 20361 13923
rect 20395 13889 20407 13923
rect 20349 13883 20407 13889
rect 20497 13923 20536 13929
rect 20497 13889 20509 13923
rect 20497 13883 20536 13889
rect 20530 13880 20536 13883
rect 20588 13880 20594 13932
rect 18138 13852 18144 13864
rect 17696 13824 18144 13852
rect 18138 13812 18144 13824
rect 18196 13812 18202 13864
rect 18233 13855 18291 13861
rect 18233 13821 18245 13855
rect 18279 13821 18291 13855
rect 18233 13815 18291 13821
rect 19628 13824 20576 13852
rect 1578 13676 1584 13728
rect 1636 13716 1642 13728
rect 2133 13719 2191 13725
rect 2133 13716 2145 13719
rect 1636 13688 2145 13716
rect 1636 13676 1642 13688
rect 2133 13685 2145 13688
rect 2179 13685 2191 13719
rect 2866 13716 2872 13728
rect 2827 13688 2872 13716
rect 2133 13679 2191 13685
rect 2866 13676 2872 13688
rect 2924 13676 2930 13728
rect 17218 13716 17224 13728
rect 17179 13688 17224 13716
rect 17218 13676 17224 13688
rect 17276 13676 17282 13728
rect 18248 13716 18276 13815
rect 19628 13793 19656 13824
rect 19613 13787 19671 13793
rect 19613 13753 19625 13787
rect 19659 13753 19671 13787
rect 19613 13747 19671 13753
rect 19242 13716 19248 13728
rect 18248 13688 19248 13716
rect 19242 13676 19248 13688
rect 19300 13676 19306 13728
rect 20548 13716 20576 13824
rect 20622 13812 20628 13864
rect 20680 13852 20686 13864
rect 20732 13852 20760 13951
rect 20898 13929 20904 13932
rect 20855 13923 20904 13929
rect 20855 13889 20867 13923
rect 20901 13889 20904 13923
rect 20855 13883 20904 13889
rect 20898 13880 20904 13883
rect 20956 13880 20962 13932
rect 21008 13920 21036 13960
rect 22002 13948 22008 14000
rect 22060 13988 22066 14000
rect 22060 13960 23244 13988
rect 22060 13948 22066 13960
rect 23216 13929 23244 13960
rect 23290 13948 23296 14000
rect 23348 13988 23354 14000
rect 23658 13988 23664 14000
rect 23348 13960 23664 13988
rect 23348 13948 23354 13960
rect 23658 13948 23664 13960
rect 23716 13988 23722 14000
rect 24026 13988 24032 14000
rect 23716 13960 24032 13988
rect 23716 13948 23722 13960
rect 24026 13948 24032 13960
rect 24084 13948 24090 14000
rect 23474 13929 23480 13932
rect 22189 13923 22247 13929
rect 22189 13920 22201 13923
rect 21008 13892 22201 13920
rect 22189 13889 22201 13892
rect 22235 13889 22247 13923
rect 22189 13883 22247 13889
rect 23201 13923 23259 13929
rect 23201 13889 23213 13923
rect 23247 13889 23259 13923
rect 23468 13920 23480 13929
rect 23435 13892 23480 13920
rect 23201 13883 23259 13889
rect 23468 13883 23480 13892
rect 23474 13880 23480 13883
rect 23532 13880 23538 13932
rect 27154 13920 27160 13932
rect 27115 13892 27160 13920
rect 27154 13880 27160 13892
rect 27212 13880 27218 13932
rect 27264 13929 27292 14028
rect 27540 13988 27568 14028
rect 27614 14016 27620 14068
rect 27672 14056 27678 14068
rect 29365 14059 29423 14065
rect 29365 14056 29377 14059
rect 27672 14028 29377 14056
rect 27672 14016 27678 14028
rect 29365 14025 29377 14028
rect 29411 14025 29423 14059
rect 29365 14019 29423 14025
rect 31018 14016 31024 14068
rect 31076 14016 31082 14068
rect 31846 14016 31852 14068
rect 31904 14056 31910 14068
rect 31904 14028 33640 14056
rect 31904 14016 31910 14028
rect 29546 13988 29552 14000
rect 27540 13960 27936 13988
rect 27249 13923 27307 13929
rect 27249 13889 27261 13923
rect 27295 13889 27307 13923
rect 27430 13920 27436 13932
rect 27391 13892 27436 13920
rect 27249 13883 27307 13889
rect 27430 13880 27436 13892
rect 27488 13880 27494 13932
rect 27525 13923 27583 13929
rect 27525 13889 27537 13923
rect 27571 13920 27583 13923
rect 27571 13892 27660 13920
rect 27571 13889 27583 13892
rect 27525 13883 27583 13889
rect 22278 13852 22284 13864
rect 20680 13824 20760 13852
rect 22239 13824 22284 13852
rect 20680 13812 20686 13824
rect 22278 13812 22284 13824
rect 22336 13812 22342 13864
rect 22465 13855 22523 13861
rect 22465 13821 22477 13855
rect 22511 13821 22523 13855
rect 22465 13815 22523 13821
rect 21634 13784 21640 13796
rect 20824 13756 21640 13784
rect 20824 13716 20852 13756
rect 21634 13744 21640 13756
rect 21692 13744 21698 13796
rect 20990 13716 20996 13728
rect 20548 13688 20852 13716
rect 20951 13688 20996 13716
rect 20990 13676 20996 13688
rect 21048 13676 21054 13728
rect 21542 13676 21548 13728
rect 21600 13716 21606 13728
rect 21821 13719 21879 13725
rect 21821 13716 21833 13719
rect 21600 13688 21833 13716
rect 21600 13676 21606 13688
rect 21821 13685 21833 13688
rect 21867 13685 21879 13719
rect 22480 13716 22508 13815
rect 25590 13812 25596 13864
rect 25648 13852 25654 13864
rect 25648 13824 27200 13852
rect 25648 13812 25654 13824
rect 27172 13784 27200 13824
rect 27632 13784 27660 13892
rect 27172 13756 27660 13784
rect 27908 13784 27936 13960
rect 28000 13960 29552 13988
rect 28000 13929 28028 13960
rect 29546 13948 29552 13960
rect 29604 13948 29610 14000
rect 31036 13988 31064 14016
rect 32398 13988 32404 14000
rect 31036 13960 31156 13988
rect 32359 13960 32404 13988
rect 27985 13923 28043 13929
rect 27985 13889 27997 13923
rect 28031 13889 28043 13923
rect 27985 13883 28043 13889
rect 28074 13880 28080 13932
rect 28132 13920 28138 13932
rect 28241 13923 28299 13929
rect 28241 13920 28253 13923
rect 28132 13892 28253 13920
rect 28132 13880 28138 13892
rect 28241 13889 28253 13892
rect 28287 13889 28299 13923
rect 28241 13883 28299 13889
rect 28626 13880 28632 13932
rect 28684 13920 28690 13932
rect 31128 13929 31156 13960
rect 32398 13948 32404 13960
rect 32456 13948 32462 14000
rect 31021 13923 31079 13929
rect 31021 13920 31033 13923
rect 28684 13892 31033 13920
rect 28684 13880 28690 13892
rect 31021 13889 31033 13892
rect 31067 13889 31079 13923
rect 31021 13883 31079 13889
rect 31113 13923 31171 13929
rect 31113 13889 31125 13923
rect 31159 13889 31171 13923
rect 31113 13883 31171 13889
rect 31205 13923 31263 13929
rect 31205 13889 31217 13923
rect 31251 13889 31263 13923
rect 31205 13883 31263 13889
rect 31389 13923 31447 13929
rect 31389 13889 31401 13923
rect 31435 13920 31447 13923
rect 31570 13920 31576 13932
rect 31435 13892 31576 13920
rect 31435 13889 31447 13892
rect 31389 13883 31447 13889
rect 31220 13852 31248 13883
rect 31570 13880 31576 13892
rect 31628 13880 31634 13932
rect 32030 13852 32036 13864
rect 31220 13824 32036 13852
rect 32030 13812 32036 13824
rect 32088 13812 32094 13864
rect 32214 13852 32220 13864
rect 32175 13824 32220 13852
rect 32214 13812 32220 13824
rect 32272 13812 32278 13864
rect 33612 13852 33640 14028
rect 34057 13923 34115 13929
rect 34057 13889 34069 13923
rect 34103 13920 34115 13923
rect 46198 13920 46204 13932
rect 34103 13892 46204 13920
rect 34103 13889 34115 13892
rect 34057 13883 34115 13889
rect 46198 13880 46204 13892
rect 46256 13880 46262 13932
rect 47854 13920 47860 13932
rect 47815 13892 47860 13920
rect 47854 13880 47860 13892
rect 47912 13880 47918 13932
rect 33612 13824 48084 13852
rect 48056 13793 48084 13824
rect 48041 13787 48099 13793
rect 27908 13756 28028 13784
rect 25314 13716 25320 13728
rect 22480 13688 25320 13716
rect 21821 13679 21879 13685
rect 25314 13676 25320 13688
rect 25372 13716 25378 13728
rect 27890 13716 27896 13728
rect 25372 13688 27896 13716
rect 25372 13676 25378 13688
rect 27890 13676 27896 13688
rect 27948 13676 27954 13728
rect 28000 13716 28028 13756
rect 48041 13753 48053 13787
rect 48087 13753 48099 13787
rect 48041 13747 48099 13753
rect 28902 13716 28908 13728
rect 28000 13688 28908 13716
rect 28902 13676 28908 13688
rect 28960 13676 28966 13728
rect 30742 13716 30748 13728
rect 30703 13688 30748 13716
rect 30742 13676 30748 13688
rect 30800 13676 30806 13728
rect 1104 13626 48852 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 48852 13626
rect 1104 13552 48852 13574
rect 20530 13472 20536 13524
rect 20588 13512 20594 13524
rect 20625 13515 20683 13521
rect 20625 13512 20637 13515
rect 20588 13484 20637 13512
rect 20588 13472 20594 13484
rect 20625 13481 20637 13484
rect 20671 13512 20683 13515
rect 22278 13512 22284 13524
rect 20671 13484 22284 13512
rect 20671 13481 20683 13484
rect 20625 13475 20683 13481
rect 22278 13472 22284 13484
rect 22336 13472 22342 13524
rect 23477 13515 23535 13521
rect 23477 13481 23489 13515
rect 23523 13512 23535 13515
rect 23566 13512 23572 13524
rect 23523 13484 23572 13512
rect 23523 13481 23535 13484
rect 23477 13475 23535 13481
rect 23566 13472 23572 13484
rect 23624 13472 23630 13524
rect 25130 13472 25136 13524
rect 25188 13512 25194 13524
rect 26329 13515 26387 13521
rect 26329 13512 26341 13515
rect 25188 13484 26341 13512
rect 25188 13472 25194 13484
rect 26329 13481 26341 13484
rect 26375 13481 26387 13515
rect 26329 13475 26387 13481
rect 26694 13472 26700 13524
rect 26752 13512 26758 13524
rect 26789 13515 26847 13521
rect 26789 13512 26801 13515
rect 26752 13484 26801 13512
rect 26752 13472 26758 13484
rect 26789 13481 26801 13484
rect 26835 13481 26847 13515
rect 26789 13475 26847 13481
rect 32214 13472 32220 13524
rect 32272 13512 32278 13524
rect 32493 13515 32551 13521
rect 32493 13512 32505 13515
rect 32272 13484 32505 13512
rect 32272 13472 32278 13484
rect 32493 13481 32505 13484
rect 32539 13481 32551 13515
rect 47670 13512 47676 13524
rect 47631 13484 47676 13512
rect 32493 13475 32551 13481
rect 47670 13472 47676 13484
rect 47728 13472 47734 13524
rect 2866 13444 2872 13456
rect 1412 13416 2872 13444
rect 1412 13385 1440 13416
rect 2866 13404 2872 13416
rect 2924 13404 2930 13456
rect 4062 13404 4068 13456
rect 4120 13444 4126 13456
rect 6914 13444 6920 13456
rect 4120 13416 6920 13444
rect 4120 13404 4126 13416
rect 6914 13404 6920 13416
rect 6972 13404 6978 13456
rect 21453 13447 21511 13453
rect 21453 13413 21465 13447
rect 21499 13444 21511 13447
rect 22830 13444 22836 13456
rect 21499 13416 22836 13444
rect 21499 13413 21511 13416
rect 21453 13407 21511 13413
rect 22830 13404 22836 13416
rect 22888 13404 22894 13456
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13345 1455 13379
rect 1578 13376 1584 13388
rect 1539 13348 1584 13376
rect 1397 13339 1455 13345
rect 1578 13336 1584 13348
rect 1636 13336 1642 13388
rect 2774 13336 2780 13388
rect 2832 13376 2838 13388
rect 2832 13348 2877 13376
rect 2832 13336 2838 13348
rect 12526 13336 12532 13388
rect 12584 13376 12590 13388
rect 14553 13379 14611 13385
rect 14553 13376 14565 13379
rect 12584 13348 14565 13376
rect 12584 13336 12590 13348
rect 14553 13345 14565 13348
rect 14599 13345 14611 13379
rect 14553 13339 14611 13345
rect 20714 13336 20720 13388
rect 20772 13376 20778 13388
rect 21542 13376 21548 13388
rect 20772 13348 21312 13376
rect 21503 13348 21548 13376
rect 20772 13336 20778 13348
rect 14093 13311 14151 13317
rect 14093 13308 14105 13311
rect 13924 13280 14105 13308
rect 13924 13172 13952 13280
rect 14093 13277 14105 13280
rect 14139 13277 14151 13311
rect 14093 13271 14151 13277
rect 16853 13311 16911 13317
rect 16853 13277 16865 13311
rect 16899 13308 16911 13311
rect 19242 13308 19248 13320
rect 16899 13280 19248 13308
rect 16899 13277 16911 13280
rect 16853 13271 16911 13277
rect 19242 13268 19248 13280
rect 19300 13268 19306 13320
rect 19512 13311 19570 13317
rect 19512 13277 19524 13311
rect 19558 13308 19570 13311
rect 20990 13308 20996 13320
rect 19558 13280 20996 13308
rect 19558 13277 19570 13280
rect 19512 13271 19570 13277
rect 20990 13268 20996 13280
rect 21048 13268 21054 13320
rect 21284 13317 21312 13348
rect 21542 13336 21548 13348
rect 21600 13336 21606 13388
rect 21634 13336 21640 13388
rect 21692 13376 21698 13388
rect 22281 13379 22339 13385
rect 22281 13376 22293 13379
rect 21692 13348 22293 13376
rect 21692 13336 21698 13348
rect 22281 13345 22293 13348
rect 22327 13345 22339 13379
rect 22281 13339 22339 13345
rect 26513 13379 26571 13385
rect 26513 13345 26525 13379
rect 26559 13376 26571 13379
rect 27338 13376 27344 13388
rect 26559 13348 27344 13376
rect 26559 13345 26571 13348
rect 26513 13339 26571 13345
rect 27338 13336 27344 13348
rect 27396 13336 27402 13388
rect 27890 13336 27896 13388
rect 27948 13376 27954 13388
rect 28169 13379 28227 13385
rect 28169 13376 28181 13379
rect 27948 13348 28181 13376
rect 27948 13336 27954 13348
rect 28169 13345 28181 13348
rect 28215 13376 28227 13379
rect 28534 13376 28540 13388
rect 28215 13348 28540 13376
rect 28215 13345 28227 13348
rect 28169 13339 28227 13345
rect 28534 13336 28540 13348
rect 28592 13336 28598 13388
rect 31110 13376 31116 13388
rect 31071 13348 31116 13376
rect 31110 13336 31116 13348
rect 31168 13336 31174 13388
rect 21269 13311 21327 13317
rect 21269 13277 21281 13311
rect 21315 13277 21327 13311
rect 21269 13271 21327 13277
rect 21361 13311 21419 13317
rect 21361 13277 21373 13311
rect 21407 13308 21419 13311
rect 21450 13308 21456 13320
rect 21407 13280 21456 13308
rect 21407 13277 21419 13280
rect 21361 13271 21419 13277
rect 21450 13268 21456 13280
rect 21508 13268 21514 13320
rect 22462 13308 22468 13320
rect 22423 13280 22468 13308
rect 22462 13268 22468 13280
rect 22520 13268 22526 13320
rect 23658 13268 23664 13320
rect 23716 13308 23722 13320
rect 24210 13308 24216 13320
rect 23716 13280 24216 13308
rect 23716 13268 23722 13280
rect 24210 13268 24216 13280
rect 24268 13268 24274 13320
rect 25314 13268 25320 13320
rect 25372 13308 25378 13320
rect 26605 13311 26663 13317
rect 26605 13308 26617 13311
rect 25372 13280 26617 13308
rect 25372 13268 25378 13280
rect 26605 13277 26617 13280
rect 26651 13277 26663 13311
rect 26605 13271 26663 13277
rect 27614 13268 27620 13320
rect 27672 13308 27678 13320
rect 28077 13311 28135 13317
rect 28077 13308 28089 13311
rect 27672 13280 28089 13308
rect 27672 13268 27678 13280
rect 28077 13277 28089 13280
rect 28123 13277 28135 13311
rect 28077 13271 28135 13277
rect 30466 13268 30472 13320
rect 30524 13308 30530 13320
rect 30653 13311 30711 13317
rect 30653 13308 30665 13311
rect 30524 13280 30665 13308
rect 30524 13268 30530 13280
rect 30653 13277 30665 13280
rect 30699 13277 30711 13311
rect 30653 13271 30711 13277
rect 30742 13268 30748 13320
rect 30800 13308 30806 13320
rect 31369 13311 31427 13317
rect 31369 13308 31381 13311
rect 30800 13280 31381 13308
rect 30800 13268 30806 13280
rect 31369 13277 31381 13280
rect 31415 13277 31427 13311
rect 31369 13271 31427 13277
rect 13998 13200 14004 13252
rect 14056 13240 14062 13252
rect 14277 13243 14335 13249
rect 14277 13240 14289 13243
rect 14056 13212 14289 13240
rect 14056 13200 14062 13212
rect 14277 13209 14289 13212
rect 14323 13209 14335 13243
rect 14277 13203 14335 13209
rect 17120 13243 17178 13249
rect 17120 13209 17132 13243
rect 17166 13240 17178 13243
rect 17218 13240 17224 13252
rect 17166 13212 17224 13240
rect 17166 13209 17178 13212
rect 17120 13203 17178 13209
rect 17218 13200 17224 13212
rect 17276 13200 17282 13252
rect 21818 13200 21824 13252
rect 21876 13240 21882 13252
rect 22005 13243 22063 13249
rect 22005 13240 22017 13243
rect 21876 13212 22017 13240
rect 21876 13200 21882 13212
rect 22005 13209 22017 13212
rect 22051 13209 22063 13243
rect 22005 13203 22063 13209
rect 23109 13243 23167 13249
rect 23109 13209 23121 13243
rect 23155 13209 23167 13243
rect 23290 13240 23296 13252
rect 23251 13212 23296 13240
rect 23109 13203 23167 13209
rect 17310 13172 17316 13184
rect 13924 13144 17316 13172
rect 17310 13132 17316 13144
rect 17368 13132 17374 13184
rect 18046 13132 18052 13184
rect 18104 13172 18110 13184
rect 18233 13175 18291 13181
rect 18233 13172 18245 13175
rect 18104 13144 18245 13172
rect 18104 13132 18110 13144
rect 18233 13141 18245 13144
rect 18279 13172 18291 13175
rect 18690 13172 18696 13184
rect 18279 13144 18696 13172
rect 18279 13141 18291 13144
rect 18233 13135 18291 13141
rect 18690 13132 18696 13144
rect 18748 13172 18754 13184
rect 20622 13172 20628 13184
rect 18748 13144 20628 13172
rect 18748 13132 18754 13144
rect 20622 13132 20628 13144
rect 20680 13132 20686 13184
rect 22649 13175 22707 13181
rect 22649 13141 22661 13175
rect 22695 13172 22707 13175
rect 23124 13172 23152 13203
rect 23290 13200 23296 13212
rect 23348 13200 23354 13252
rect 26329 13243 26387 13249
rect 26329 13209 26341 13243
rect 26375 13240 26387 13243
rect 27154 13240 27160 13252
rect 26375 13212 27160 13240
rect 26375 13209 26387 13212
rect 26329 13203 26387 13209
rect 27154 13200 27160 13212
rect 27212 13240 27218 13252
rect 27982 13240 27988 13252
rect 27212 13212 27660 13240
rect 27943 13212 27988 13240
rect 27212 13200 27218 13212
rect 22695 13144 23152 13172
rect 22695 13141 22707 13144
rect 22649 13135 22707 13141
rect 23842 13132 23848 13184
rect 23900 13172 23906 13184
rect 26970 13172 26976 13184
rect 23900 13144 26976 13172
rect 23900 13132 23906 13144
rect 26970 13132 26976 13144
rect 27028 13132 27034 13184
rect 27632 13181 27660 13212
rect 27982 13200 27988 13212
rect 28040 13200 28046 13252
rect 27617 13175 27675 13181
rect 27617 13141 27629 13175
rect 27663 13141 27675 13175
rect 27617 13135 27675 13141
rect 27706 13132 27712 13184
rect 27764 13172 27770 13184
rect 28534 13172 28540 13184
rect 27764 13144 28540 13172
rect 27764 13132 27770 13144
rect 28534 13132 28540 13144
rect 28592 13132 28598 13184
rect 30469 13175 30527 13181
rect 30469 13141 30481 13175
rect 30515 13172 30527 13175
rect 30558 13172 30564 13184
rect 30515 13144 30564 13172
rect 30515 13141 30527 13144
rect 30469 13135 30527 13141
rect 30558 13132 30564 13144
rect 30616 13172 30622 13184
rect 31662 13172 31668 13184
rect 30616 13144 31668 13172
rect 30616 13132 30622 13144
rect 31662 13132 31668 13144
rect 31720 13132 31726 13184
rect 1104 13082 48852 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 48852 13082
rect 1104 13008 48852 13030
rect 13998 12968 14004 12980
rect 13959 12940 14004 12968
rect 13998 12928 14004 12940
rect 14056 12928 14062 12980
rect 18138 12968 18144 12980
rect 18099 12940 18144 12968
rect 18138 12928 18144 12940
rect 18196 12928 18202 12980
rect 21174 12968 21180 12980
rect 21135 12940 21180 12968
rect 21174 12928 21180 12940
rect 21232 12928 21238 12980
rect 22465 12971 22523 12977
rect 22465 12937 22477 12971
rect 22511 12968 22523 12971
rect 22511 12940 23244 12968
rect 22511 12937 22523 12940
rect 22465 12931 22523 12937
rect 18046 12900 18052 12912
rect 17880 12872 18052 12900
rect 1673 12835 1731 12841
rect 1673 12801 1685 12835
rect 1719 12832 1731 12835
rect 8478 12832 8484 12844
rect 1719 12804 8484 12832
rect 1719 12801 1731 12804
rect 1673 12795 1731 12801
rect 8478 12792 8484 12804
rect 8536 12792 8542 12844
rect 9766 12832 9772 12844
rect 9679 12804 9772 12832
rect 9766 12792 9772 12804
rect 9824 12832 9830 12844
rect 11606 12832 11612 12844
rect 9824 12804 11612 12832
rect 9824 12792 9830 12804
rect 11606 12792 11612 12804
rect 11664 12832 11670 12844
rect 13909 12835 13967 12841
rect 13909 12832 13921 12835
rect 11664 12804 13921 12832
rect 11664 12792 11670 12804
rect 13909 12801 13921 12804
rect 13955 12832 13967 12835
rect 15470 12832 15476 12844
rect 13955 12804 15476 12832
rect 13955 12801 13967 12804
rect 13909 12795 13967 12801
rect 15470 12792 15476 12804
rect 15528 12792 15534 12844
rect 17880 12841 17908 12872
rect 18046 12860 18052 12872
rect 18104 12860 18110 12912
rect 19610 12860 19616 12912
rect 19668 12900 19674 12912
rect 20070 12900 20076 12912
rect 19668 12872 20076 12900
rect 19668 12860 19674 12872
rect 20070 12860 20076 12872
rect 20128 12860 20134 12912
rect 21085 12903 21143 12909
rect 21085 12869 21097 12903
rect 21131 12900 21143 12903
rect 22646 12900 22652 12912
rect 21131 12872 22652 12900
rect 21131 12869 21143 12872
rect 21085 12863 21143 12869
rect 22646 12860 22652 12872
rect 22704 12860 22710 12912
rect 17865 12835 17923 12841
rect 17865 12801 17877 12835
rect 17911 12801 17923 12835
rect 17865 12795 17923 12801
rect 17957 12835 18015 12841
rect 17957 12801 17969 12835
rect 18003 12801 18015 12835
rect 17957 12795 18015 12801
rect 1394 12764 1400 12776
rect 1355 12736 1400 12764
rect 1394 12724 1400 12736
rect 1452 12724 1458 12776
rect 7926 12724 7932 12776
rect 7984 12764 7990 12776
rect 10045 12767 10103 12773
rect 10045 12764 10057 12767
rect 7984 12736 10057 12764
rect 7984 12724 7990 12736
rect 10045 12733 10057 12736
rect 10091 12764 10103 12767
rect 10502 12764 10508 12776
rect 10091 12736 10508 12764
rect 10091 12733 10103 12736
rect 10045 12727 10103 12733
rect 10502 12724 10508 12736
rect 10560 12724 10566 12776
rect 17972 12696 18000 12795
rect 21542 12792 21548 12844
rect 21600 12832 21606 12844
rect 22005 12835 22063 12841
rect 22005 12832 22017 12835
rect 21600 12804 22017 12832
rect 21600 12792 21606 12804
rect 22005 12801 22017 12804
rect 22051 12801 22063 12835
rect 22005 12795 22063 12801
rect 22281 12835 22339 12841
rect 22281 12801 22293 12835
rect 22327 12832 22339 12835
rect 22462 12832 22468 12844
rect 22327 12804 22468 12832
rect 22327 12801 22339 12804
rect 22281 12795 22339 12801
rect 22462 12792 22468 12804
rect 22520 12832 22526 12844
rect 22922 12832 22928 12844
rect 22520 12804 22928 12832
rect 22520 12792 22526 12804
rect 22922 12792 22928 12804
rect 22980 12792 22986 12844
rect 23216 12832 23244 12940
rect 23290 12928 23296 12980
rect 23348 12968 23354 12980
rect 26421 12971 26479 12977
rect 26421 12968 26433 12971
rect 23348 12940 26433 12968
rect 23348 12928 23354 12940
rect 26421 12937 26433 12940
rect 26467 12937 26479 12971
rect 27338 12968 27344 12980
rect 27299 12940 27344 12968
rect 26421 12931 26479 12937
rect 27338 12928 27344 12940
rect 27396 12968 27402 12980
rect 28902 12968 28908 12980
rect 27396 12940 28580 12968
rect 28863 12940 28908 12968
rect 27396 12928 27402 12940
rect 23842 12860 23848 12912
rect 23900 12900 23906 12912
rect 24213 12903 24271 12909
rect 24213 12900 24225 12903
rect 23900 12872 24225 12900
rect 23900 12860 23906 12872
rect 24213 12869 24225 12872
rect 24259 12869 24271 12903
rect 24394 12900 24400 12912
rect 24355 12872 24400 12900
rect 24213 12863 24271 12869
rect 24394 12860 24400 12872
rect 24452 12860 24458 12912
rect 25314 12900 25320 12912
rect 24504 12872 25320 12900
rect 24504 12841 24532 12872
rect 25314 12860 25320 12872
rect 25372 12860 25378 12912
rect 25961 12903 26019 12909
rect 25961 12869 25973 12903
rect 26007 12900 26019 12903
rect 27798 12900 27804 12912
rect 26007 12872 27804 12900
rect 26007 12869 26019 12872
rect 25961 12863 26019 12869
rect 27798 12860 27804 12872
rect 27856 12860 27862 12912
rect 28552 12909 28580 12940
rect 28902 12928 28908 12940
rect 28960 12928 28966 12980
rect 32030 12928 32036 12980
rect 32088 12968 32094 12980
rect 32493 12971 32551 12977
rect 32493 12968 32505 12971
rect 32088 12940 32505 12968
rect 32088 12928 32094 12940
rect 32493 12937 32505 12940
rect 32539 12937 32551 12971
rect 32493 12931 32551 12937
rect 28537 12903 28595 12909
rect 28537 12869 28549 12903
rect 28583 12869 28595 12903
rect 28537 12863 28595 12869
rect 31662 12860 31668 12912
rect 31720 12900 31726 12912
rect 32125 12903 32183 12909
rect 32125 12900 32137 12903
rect 31720 12872 32137 12900
rect 31720 12860 31726 12872
rect 32125 12869 32137 12872
rect 32171 12869 32183 12903
rect 32125 12863 32183 12869
rect 32214 12860 32220 12912
rect 32272 12900 32278 12912
rect 32309 12903 32367 12909
rect 32309 12900 32321 12903
rect 32272 12872 32321 12900
rect 32272 12860 32278 12872
rect 32309 12869 32321 12872
rect 32355 12869 32367 12903
rect 32309 12863 32367 12869
rect 24489 12835 24547 12841
rect 23216 12804 24440 12832
rect 21450 12724 21456 12776
rect 21508 12764 21514 12776
rect 22097 12767 22155 12773
rect 22097 12764 22109 12767
rect 21508 12736 22109 12764
rect 21508 12724 21514 12736
rect 22097 12733 22109 12736
rect 22143 12733 22155 12767
rect 23658 12764 23664 12776
rect 22097 12727 22155 12733
rect 22480 12736 23664 12764
rect 22480 12696 22508 12736
rect 23658 12724 23664 12736
rect 23716 12724 23722 12776
rect 24412 12764 24440 12804
rect 24489 12801 24501 12835
rect 24535 12801 24547 12835
rect 25130 12832 25136 12844
rect 25091 12804 25136 12832
rect 24489 12795 24547 12801
rect 25130 12792 25136 12804
rect 25188 12792 25194 12844
rect 26237 12835 26295 12841
rect 26237 12801 26249 12835
rect 26283 12832 26295 12835
rect 26694 12832 26700 12844
rect 26283 12804 26700 12832
rect 26283 12801 26295 12804
rect 26237 12795 26295 12801
rect 26694 12792 26700 12804
rect 26752 12792 26758 12844
rect 27706 12832 27712 12844
rect 27667 12804 27712 12832
rect 27706 12792 27712 12804
rect 27764 12832 27770 12844
rect 28626 12832 28632 12844
rect 27764 12804 28632 12832
rect 27764 12792 27770 12804
rect 28626 12792 28632 12804
rect 28684 12792 28690 12844
rect 28721 12835 28779 12841
rect 28721 12801 28733 12835
rect 28767 12801 28779 12835
rect 28721 12795 28779 12801
rect 30561 12835 30619 12841
rect 30561 12801 30573 12835
rect 30607 12832 30619 12835
rect 30834 12832 30840 12844
rect 30607 12804 30840 12832
rect 30607 12801 30619 12804
rect 30561 12795 30619 12801
rect 25038 12764 25044 12776
rect 24412 12736 25044 12764
rect 25038 12724 25044 12736
rect 25096 12764 25102 12776
rect 25225 12767 25283 12773
rect 25225 12764 25237 12767
rect 25096 12736 25237 12764
rect 25096 12724 25102 12736
rect 25225 12733 25237 12736
rect 25271 12733 25283 12767
rect 25225 12727 25283 12733
rect 26145 12767 26203 12773
rect 26145 12733 26157 12767
rect 26191 12764 26203 12767
rect 27614 12764 27620 12776
rect 26191 12736 27620 12764
rect 26191 12733 26203 12736
rect 26145 12727 26203 12733
rect 27614 12724 27620 12736
rect 27672 12724 27678 12776
rect 27890 12764 27896 12776
rect 27851 12736 27896 12764
rect 27890 12724 27896 12736
rect 27948 12724 27954 12776
rect 17972 12668 22508 12696
rect 22554 12656 22560 12708
rect 22612 12696 22618 12708
rect 22612 12668 26087 12696
rect 22612 12656 22618 12668
rect 18598 12588 18604 12640
rect 18656 12628 18662 12640
rect 19426 12628 19432 12640
rect 18656 12600 19432 12628
rect 18656 12588 18662 12600
rect 19426 12588 19432 12600
rect 19484 12588 19490 12640
rect 22186 12628 22192 12640
rect 22147 12600 22192 12628
rect 22186 12588 22192 12600
rect 22244 12588 22250 12640
rect 23842 12588 23848 12640
rect 23900 12628 23906 12640
rect 24213 12631 24271 12637
rect 24213 12628 24225 12631
rect 23900 12600 24225 12628
rect 23900 12588 23906 12600
rect 24213 12597 24225 12600
rect 24259 12597 24271 12631
rect 25314 12628 25320 12640
rect 25275 12600 25320 12628
rect 24213 12591 24271 12597
rect 25314 12588 25320 12600
rect 25372 12588 25378 12640
rect 25501 12631 25559 12637
rect 25501 12597 25513 12631
rect 25547 12628 25559 12631
rect 25682 12628 25688 12640
rect 25547 12600 25688 12628
rect 25547 12597 25559 12600
rect 25501 12591 25559 12597
rect 25682 12588 25688 12600
rect 25740 12588 25746 12640
rect 25958 12628 25964 12640
rect 25919 12600 25964 12628
rect 25958 12588 25964 12600
rect 26016 12588 26022 12640
rect 26059 12628 26087 12668
rect 26326 12656 26332 12708
rect 26384 12696 26390 12708
rect 27522 12696 27528 12708
rect 26384 12668 27528 12696
rect 26384 12656 26390 12668
rect 27522 12656 27528 12668
rect 27580 12696 27586 12708
rect 28736 12696 28764 12795
rect 30834 12792 30840 12804
rect 30892 12832 30898 12844
rect 31018 12832 31024 12844
rect 30892 12804 31024 12832
rect 30892 12792 30898 12804
rect 31018 12792 31024 12804
rect 31076 12792 31082 12844
rect 30285 12767 30343 12773
rect 30285 12733 30297 12767
rect 30331 12733 30343 12767
rect 30285 12727 30343 12733
rect 27580 12668 28764 12696
rect 27580 12656 27586 12668
rect 30300 12628 30328 12727
rect 42794 12656 42800 12708
rect 42852 12696 42858 12708
rect 46842 12696 46848 12708
rect 42852 12668 46848 12696
rect 42852 12656 42858 12668
rect 46842 12656 46848 12668
rect 46900 12656 46906 12708
rect 26059 12600 30328 12628
rect 1104 12538 48852 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 48852 12538
rect 1104 12464 48852 12486
rect 23382 12384 23388 12436
rect 23440 12424 23446 12436
rect 23753 12427 23811 12433
rect 23753 12424 23765 12427
rect 23440 12396 23765 12424
rect 23440 12384 23446 12396
rect 23753 12393 23765 12396
rect 23799 12393 23811 12427
rect 23753 12387 23811 12393
rect 25133 12427 25191 12433
rect 25133 12393 25145 12427
rect 25179 12424 25191 12427
rect 25314 12424 25320 12436
rect 25179 12396 25320 12424
rect 25179 12393 25191 12396
rect 25133 12387 25191 12393
rect 18601 12359 18659 12365
rect 18601 12325 18613 12359
rect 18647 12356 18659 12359
rect 19242 12356 19248 12368
rect 18647 12328 19248 12356
rect 18647 12325 18659 12328
rect 18601 12319 18659 12325
rect 19242 12316 19248 12328
rect 19300 12316 19306 12368
rect 20070 12356 20076 12368
rect 19720 12328 20076 12356
rect 11606 12220 11612 12232
rect 11567 12192 11612 12220
rect 11606 12180 11612 12192
rect 11664 12180 11670 12232
rect 17862 12180 17868 12232
rect 17920 12220 17926 12232
rect 19720 12229 19748 12328
rect 20070 12316 20076 12328
rect 20128 12356 20134 12368
rect 22554 12356 22560 12368
rect 20128 12328 22560 12356
rect 20128 12316 20134 12328
rect 22554 12316 22560 12328
rect 22612 12316 22618 12368
rect 24118 12356 24124 12368
rect 23676 12328 24124 12356
rect 21082 12248 21088 12300
rect 21140 12288 21146 12300
rect 21140 12260 21772 12288
rect 21140 12248 21146 12260
rect 18417 12223 18475 12229
rect 18417 12220 18429 12223
rect 17920 12192 18429 12220
rect 17920 12180 17926 12192
rect 18417 12189 18429 12192
rect 18463 12189 18475 12223
rect 18417 12183 18475 12189
rect 19705 12223 19763 12229
rect 19705 12189 19717 12223
rect 19751 12189 19763 12223
rect 21542 12220 21548 12232
rect 21503 12192 21548 12220
rect 19705 12183 19763 12189
rect 21542 12180 21548 12192
rect 21600 12180 21606 12232
rect 21744 12229 21772 12260
rect 21818 12248 21824 12300
rect 21876 12288 21882 12300
rect 23014 12288 23020 12300
rect 21876 12260 21921 12288
rect 22020 12260 23020 12288
rect 21876 12248 21882 12260
rect 21729 12223 21787 12229
rect 21729 12189 21741 12223
rect 21775 12189 21787 12223
rect 21729 12183 21787 12189
rect 21913 12223 21971 12229
rect 21913 12189 21925 12223
rect 21959 12220 21971 12223
rect 22020 12220 22048 12260
rect 23014 12248 23020 12260
rect 23072 12248 23078 12300
rect 23676 12297 23704 12328
rect 24118 12316 24124 12328
rect 24176 12356 24182 12368
rect 25148 12356 25176 12387
rect 25314 12384 25320 12396
rect 25372 12384 25378 12436
rect 25590 12384 25596 12436
rect 25648 12424 25654 12436
rect 25777 12427 25835 12433
rect 25777 12424 25789 12427
rect 25648 12396 25789 12424
rect 25648 12384 25654 12396
rect 25777 12393 25789 12396
rect 25823 12424 25835 12427
rect 25866 12424 25872 12436
rect 25823 12396 25872 12424
rect 25823 12393 25835 12396
rect 25777 12387 25835 12393
rect 25866 12384 25872 12396
rect 25924 12384 25930 12436
rect 26602 12384 26608 12436
rect 26660 12424 26666 12436
rect 30466 12424 30472 12436
rect 26660 12396 30472 12424
rect 26660 12384 26666 12396
rect 30466 12384 30472 12396
rect 30524 12384 30530 12436
rect 38470 12384 38476 12436
rect 38528 12424 38534 12436
rect 46842 12424 46848 12436
rect 38528 12396 46848 12424
rect 38528 12384 38534 12396
rect 46842 12384 46848 12396
rect 46900 12384 46906 12436
rect 24176 12328 25176 12356
rect 24176 12316 24182 12328
rect 27062 12316 27068 12368
rect 27120 12356 27126 12368
rect 28534 12356 28540 12368
rect 27120 12328 28540 12356
rect 27120 12316 27126 12328
rect 28534 12316 28540 12328
rect 28592 12316 28598 12368
rect 30374 12316 30380 12368
rect 30432 12356 30438 12368
rect 30834 12356 30840 12368
rect 30432 12328 30840 12356
rect 30432 12316 30438 12328
rect 30834 12316 30840 12328
rect 30892 12356 30898 12368
rect 30892 12328 31754 12356
rect 30892 12316 30898 12328
rect 23842 12297 23848 12300
rect 23661 12291 23719 12297
rect 23661 12257 23673 12291
rect 23707 12257 23719 12291
rect 23841 12288 23848 12297
rect 23803 12260 23848 12288
rect 23661 12251 23719 12257
rect 23841 12251 23848 12260
rect 23842 12248 23848 12251
rect 23900 12248 23906 12300
rect 24765 12291 24823 12297
rect 24765 12257 24777 12291
rect 24811 12288 24823 12291
rect 25961 12291 26019 12297
rect 25961 12288 25973 12291
rect 24811 12260 25973 12288
rect 24811 12257 24823 12260
rect 24765 12251 24823 12257
rect 25961 12257 25973 12260
rect 26007 12257 26019 12291
rect 25961 12251 26019 12257
rect 26142 12248 26148 12300
rect 26200 12288 26206 12300
rect 27525 12291 27583 12297
rect 27525 12288 27537 12291
rect 26200 12260 27537 12288
rect 26200 12248 26206 12260
rect 27525 12257 27537 12260
rect 27571 12257 27583 12291
rect 27890 12288 27896 12300
rect 27525 12251 27583 12257
rect 27632 12260 27896 12288
rect 21959 12192 22048 12220
rect 22097 12223 22155 12229
rect 21959 12189 21971 12192
rect 21913 12183 21971 12189
rect 22097 12189 22109 12223
rect 22143 12220 22155 12223
rect 22186 12220 22192 12232
rect 22143 12192 22192 12220
rect 22143 12189 22155 12192
rect 22097 12183 22155 12189
rect 19610 12112 19616 12164
rect 19668 12152 19674 12164
rect 20070 12152 20076 12164
rect 19668 12124 20076 12152
rect 19668 12112 19674 12124
rect 20070 12112 20076 12124
rect 20128 12112 20134 12164
rect 21744 12152 21772 12183
rect 22186 12180 22192 12192
rect 22244 12220 22250 12232
rect 23198 12220 23204 12232
rect 22244 12192 23204 12220
rect 22244 12180 22250 12192
rect 23198 12180 23204 12192
rect 23256 12180 23262 12232
rect 23569 12223 23627 12229
rect 23569 12189 23581 12223
rect 23615 12189 23627 12223
rect 24946 12220 24952 12232
rect 24907 12192 24952 12220
rect 23569 12183 23627 12189
rect 23474 12152 23480 12164
rect 21744 12124 23480 12152
rect 23474 12112 23480 12124
rect 23532 12112 23538 12164
rect 23584 12152 23612 12183
rect 24946 12180 24952 12192
rect 25004 12220 25010 12232
rect 25130 12220 25136 12232
rect 25004 12192 25136 12220
rect 25004 12180 25010 12192
rect 25130 12180 25136 12192
rect 25188 12180 25194 12232
rect 25225 12223 25283 12229
rect 25225 12189 25237 12223
rect 25271 12189 25283 12223
rect 25682 12220 25688 12232
rect 25643 12192 25688 12220
rect 25225 12183 25283 12189
rect 24394 12152 24400 12164
rect 23584 12124 24400 12152
rect 24394 12112 24400 12124
rect 24452 12152 24458 12164
rect 25240 12152 25268 12183
rect 25682 12180 25688 12192
rect 25740 12220 25746 12232
rect 26326 12220 26332 12232
rect 25740 12192 26332 12220
rect 25740 12180 25746 12192
rect 26326 12180 26332 12192
rect 26384 12180 26390 12232
rect 27154 12220 27160 12232
rect 27115 12192 27160 12220
rect 27154 12180 27160 12192
rect 27212 12180 27218 12232
rect 27341 12223 27399 12229
rect 27341 12189 27353 12223
rect 27387 12189 27399 12223
rect 27341 12183 27399 12189
rect 27433 12223 27491 12229
rect 27433 12189 27445 12223
rect 27479 12220 27491 12223
rect 27632 12220 27660 12260
rect 27890 12248 27896 12260
rect 27948 12248 27954 12300
rect 27982 12248 27988 12300
rect 28040 12288 28046 12300
rect 31726 12288 31754 12328
rect 28040 12260 30512 12288
rect 31726 12260 31800 12288
rect 28040 12248 28046 12260
rect 27479 12192 27660 12220
rect 27479 12189 27491 12192
rect 27433 12183 27491 12189
rect 24452 12124 25268 12152
rect 26068 12124 26372 12152
rect 24452 12112 24458 12124
rect 11698 12084 11704 12096
rect 11659 12056 11704 12084
rect 11698 12044 11704 12056
rect 11756 12044 11762 12096
rect 19334 12044 19340 12096
rect 19392 12084 19398 12096
rect 19797 12087 19855 12093
rect 19797 12084 19809 12087
rect 19392 12056 19809 12084
rect 19392 12044 19398 12056
rect 19797 12053 19809 12056
rect 19843 12053 19855 12087
rect 22278 12084 22284 12096
rect 22239 12056 22284 12084
rect 19797 12047 19855 12053
rect 22278 12044 22284 12056
rect 22336 12044 22342 12096
rect 22646 12044 22652 12096
rect 22704 12084 22710 12096
rect 26068 12084 26096 12124
rect 26234 12084 26240 12096
rect 22704 12056 26096 12084
rect 26195 12056 26240 12084
rect 22704 12044 22710 12056
rect 26234 12044 26240 12056
rect 26292 12044 26298 12096
rect 26344 12084 26372 12124
rect 26418 12112 26424 12164
rect 26476 12152 26482 12164
rect 27356 12152 27384 12183
rect 27706 12180 27712 12232
rect 27764 12220 27770 12232
rect 28258 12220 28264 12232
rect 27764 12192 28264 12220
rect 27764 12180 27770 12192
rect 28258 12180 28264 12192
rect 28316 12180 28322 12232
rect 28442 12220 28448 12232
rect 28403 12192 28448 12220
rect 28442 12180 28448 12192
rect 28500 12180 28506 12232
rect 28534 12180 28540 12232
rect 28592 12220 28598 12232
rect 30101 12223 30159 12229
rect 30101 12220 30113 12223
rect 28592 12192 30113 12220
rect 28592 12180 28598 12192
rect 30101 12189 30113 12192
rect 30147 12189 30159 12223
rect 30101 12183 30159 12189
rect 30377 12223 30435 12229
rect 30377 12189 30389 12223
rect 30423 12189 30435 12223
rect 30484 12220 30512 12260
rect 31772 12229 31800 12260
rect 31665 12223 31723 12229
rect 31665 12220 31677 12223
rect 30484 12192 31677 12220
rect 30377 12183 30435 12189
rect 31665 12189 31677 12192
rect 31711 12189 31723 12223
rect 31665 12183 31723 12189
rect 31757 12223 31815 12229
rect 31757 12189 31769 12223
rect 31803 12189 31815 12223
rect 31757 12183 31815 12189
rect 28629 12155 28687 12161
rect 28629 12152 28641 12155
rect 26476 12124 27384 12152
rect 27540 12124 28641 12152
rect 26476 12112 26482 12124
rect 27540 12096 27568 12124
rect 28629 12121 28641 12124
rect 28675 12121 28687 12155
rect 30392 12152 30420 12183
rect 31846 12180 31852 12232
rect 31904 12220 31910 12232
rect 32033 12223 32091 12229
rect 31904 12192 31949 12220
rect 31904 12180 31910 12192
rect 32033 12189 32045 12223
rect 32079 12189 32091 12223
rect 32033 12183 32091 12189
rect 30650 12152 30656 12164
rect 30392 12124 30656 12152
rect 28629 12115 28687 12121
rect 30650 12112 30656 12124
rect 30708 12152 30714 12164
rect 31570 12152 31576 12164
rect 30708 12124 31576 12152
rect 30708 12112 30714 12124
rect 31570 12112 31576 12124
rect 31628 12152 31634 12164
rect 32048 12152 32076 12183
rect 31628 12124 32076 12152
rect 31628 12112 31634 12124
rect 27062 12084 27068 12096
rect 26344 12056 27068 12084
rect 27062 12044 27068 12056
rect 27120 12044 27126 12096
rect 27522 12044 27528 12096
rect 27580 12044 27586 12096
rect 27893 12087 27951 12093
rect 27893 12053 27905 12087
rect 27939 12084 27951 12087
rect 28074 12084 28080 12096
rect 27939 12056 28080 12084
rect 27939 12053 27951 12056
rect 27893 12047 27951 12053
rect 28074 12044 28080 12056
rect 28132 12044 28138 12096
rect 30742 12044 30748 12096
rect 30800 12084 30806 12096
rect 31389 12087 31447 12093
rect 31389 12084 31401 12087
rect 30800 12056 31401 12084
rect 30800 12044 30806 12056
rect 31389 12053 31401 12056
rect 31435 12053 31447 12087
rect 31389 12047 31447 12053
rect 1104 11994 48852 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 48852 11994
rect 1104 11920 48852 11942
rect 12710 11840 12716 11892
rect 12768 11880 12774 11892
rect 18417 11883 18475 11889
rect 18417 11880 18429 11883
rect 12768 11852 18429 11880
rect 12768 11840 12774 11852
rect 18417 11849 18429 11852
rect 18463 11849 18475 11883
rect 18417 11843 18475 11849
rect 18432 11744 18460 11843
rect 21542 11840 21548 11892
rect 21600 11880 21606 11892
rect 23477 11883 23535 11889
rect 23477 11880 23489 11883
rect 21600 11852 23489 11880
rect 21600 11840 21606 11852
rect 23477 11849 23489 11852
rect 23523 11849 23535 11883
rect 23477 11843 23535 11849
rect 24029 11883 24087 11889
rect 24029 11849 24041 11883
rect 24075 11880 24087 11883
rect 24118 11880 24124 11892
rect 24075 11852 24124 11880
rect 24075 11849 24087 11852
rect 24029 11843 24087 11849
rect 24118 11840 24124 11852
rect 24176 11840 24182 11892
rect 24946 11840 24952 11892
rect 25004 11880 25010 11892
rect 25501 11883 25559 11889
rect 25501 11880 25513 11883
rect 25004 11852 25513 11880
rect 25004 11840 25010 11852
rect 25501 11849 25513 11852
rect 25547 11849 25559 11883
rect 25501 11843 25559 11849
rect 27157 11883 27215 11889
rect 27157 11849 27169 11883
rect 27203 11880 27215 11883
rect 27430 11880 27436 11892
rect 27203 11852 27436 11880
rect 27203 11849 27215 11852
rect 27157 11843 27215 11849
rect 27430 11840 27436 11852
rect 27488 11840 27494 11892
rect 31481 11883 31539 11889
rect 29196 11852 30604 11880
rect 21818 11772 21824 11824
rect 21876 11812 21882 11824
rect 22281 11815 22339 11821
rect 22281 11812 22293 11815
rect 21876 11784 22293 11812
rect 21876 11772 21882 11784
rect 22281 11781 22293 11784
rect 22327 11781 22339 11815
rect 22281 11775 22339 11781
rect 25869 11815 25927 11821
rect 25869 11781 25881 11815
rect 25915 11812 25927 11815
rect 26786 11812 26792 11824
rect 25915 11784 26792 11812
rect 25915 11781 25927 11784
rect 25869 11775 25927 11781
rect 26786 11772 26792 11784
rect 26844 11772 26850 11824
rect 26970 11812 26976 11824
rect 26931 11784 26976 11812
rect 26970 11772 26976 11784
rect 27028 11772 27034 11824
rect 27890 11772 27896 11824
rect 27948 11812 27954 11824
rect 27948 11784 28028 11812
rect 27948 11772 27954 11784
rect 18785 11747 18843 11753
rect 18785 11744 18797 11747
rect 18432 11716 18797 11744
rect 18785 11713 18797 11716
rect 18831 11744 18843 11747
rect 19886 11744 19892 11756
rect 18831 11716 19892 11744
rect 18831 11713 18843 11716
rect 18785 11707 18843 11713
rect 19886 11704 19892 11716
rect 19944 11704 19950 11756
rect 20165 11747 20223 11753
rect 20165 11713 20177 11747
rect 20211 11713 20223 11747
rect 20165 11707 20223 11713
rect 20349 11747 20407 11753
rect 20349 11713 20361 11747
rect 20395 11744 20407 11747
rect 20530 11744 20536 11756
rect 20395 11716 20536 11744
rect 20395 11713 20407 11716
rect 20349 11707 20407 11713
rect 19058 11676 19064 11688
rect 19019 11648 19064 11676
rect 19058 11636 19064 11648
rect 19116 11676 19122 11688
rect 20180 11676 20208 11707
rect 20530 11704 20536 11716
rect 20588 11704 20594 11756
rect 22186 11744 22192 11756
rect 22147 11716 22192 11744
rect 22186 11704 22192 11716
rect 22244 11704 22250 11756
rect 23017 11747 23075 11753
rect 23017 11713 23029 11747
rect 23063 11713 23075 11747
rect 24394 11744 24400 11756
rect 24355 11716 24400 11744
rect 23017 11707 23075 11713
rect 19116 11648 20208 11676
rect 22373 11679 22431 11685
rect 19116 11636 19122 11648
rect 22373 11645 22385 11679
rect 22419 11676 22431 11679
rect 22738 11676 22744 11688
rect 22419 11648 22744 11676
rect 22419 11645 22431 11648
rect 22373 11639 22431 11645
rect 22738 11636 22744 11648
rect 22796 11636 22802 11688
rect 21821 11611 21879 11617
rect 18984 11580 20668 11608
rect 18984 11552 19012 11580
rect 17034 11500 17040 11552
rect 17092 11540 17098 11552
rect 18966 11540 18972 11552
rect 17092 11512 18972 11540
rect 17092 11500 17098 11512
rect 18966 11500 18972 11512
rect 19024 11500 19030 11552
rect 20530 11540 20536 11552
rect 20491 11512 20536 11540
rect 20530 11500 20536 11512
rect 20588 11500 20594 11552
rect 20640 11540 20668 11580
rect 21821 11577 21833 11611
rect 21867 11608 21879 11611
rect 22462 11608 22468 11620
rect 21867 11580 22468 11608
rect 21867 11577 21879 11580
rect 21821 11571 21879 11577
rect 22462 11568 22468 11580
rect 22520 11608 22526 11620
rect 23032 11608 23060 11707
rect 24394 11704 24400 11716
rect 24452 11704 24458 11756
rect 24489 11747 24547 11753
rect 24489 11713 24501 11747
rect 24535 11744 24547 11747
rect 25774 11744 25780 11756
rect 24535 11716 25780 11744
rect 24535 11713 24547 11716
rect 24489 11707 24547 11713
rect 24210 11636 24216 11688
rect 24268 11676 24274 11688
rect 24504 11676 24532 11707
rect 25774 11704 25780 11716
rect 25832 11704 25838 11756
rect 25961 11747 26019 11753
rect 25961 11713 25973 11747
rect 26007 11744 26019 11747
rect 26326 11744 26332 11756
rect 26007 11716 26332 11744
rect 26007 11713 26019 11716
rect 25961 11707 26019 11713
rect 26326 11704 26332 11716
rect 26384 11744 26390 11756
rect 26694 11744 26700 11756
rect 26384 11716 26700 11744
rect 26384 11704 26390 11716
rect 26694 11704 26700 11716
rect 26752 11704 26758 11756
rect 27249 11747 27307 11753
rect 27249 11713 27261 11747
rect 27295 11744 27307 11747
rect 27338 11744 27344 11756
rect 27295 11716 27344 11744
rect 27295 11713 27307 11716
rect 27249 11707 27307 11713
rect 27338 11704 27344 11716
rect 27396 11704 27402 11756
rect 28000 11753 28028 11784
rect 28074 11772 28080 11824
rect 28132 11812 28138 11824
rect 29196 11812 29224 11852
rect 28132 11784 29224 11812
rect 30576 11812 30604 11852
rect 31481 11849 31493 11883
rect 31527 11880 31539 11883
rect 31846 11880 31852 11892
rect 31527 11852 31852 11880
rect 31527 11849 31539 11852
rect 31481 11843 31539 11849
rect 31846 11840 31852 11852
rect 31904 11840 31910 11892
rect 39117 11815 39175 11821
rect 28132 11772 28138 11784
rect 27976 11747 28034 11753
rect 27976 11713 27988 11747
rect 28022 11713 28034 11747
rect 27976 11707 28034 11713
rect 28350 11704 28356 11756
rect 28408 11744 28414 11756
rect 30285 11747 30343 11753
rect 30285 11744 30297 11747
rect 28408 11716 30297 11744
rect 28408 11704 28414 11716
rect 30285 11713 30297 11716
rect 30331 11713 30343 11747
rect 30374 11738 30380 11790
rect 30432 11738 30438 11790
rect 30576 11784 31754 11812
rect 30285 11707 30343 11713
rect 30377 11713 30389 11738
rect 30423 11713 30435 11738
rect 30377 11707 30435 11713
rect 30466 11704 30472 11756
rect 30524 11744 30530 11756
rect 30524 11716 30569 11744
rect 30524 11704 30530 11716
rect 30650 11704 30656 11756
rect 30708 11744 30714 11756
rect 31113 11747 31171 11753
rect 30708 11716 30753 11744
rect 30708 11704 30714 11716
rect 31113 11713 31125 11747
rect 31159 11713 31171 11747
rect 31113 11707 31171 11713
rect 31297 11747 31355 11753
rect 31297 11713 31309 11747
rect 31343 11713 31355 11747
rect 31726 11744 31754 11784
rect 39117 11781 39129 11815
rect 39163 11812 39175 11815
rect 42794 11812 42800 11824
rect 39163 11784 42800 11812
rect 39163 11781 39175 11784
rect 39117 11775 39175 11781
rect 42794 11772 42800 11784
rect 42852 11772 42858 11824
rect 37277 11747 37335 11753
rect 37277 11744 37289 11747
rect 31726 11716 37289 11744
rect 31297 11707 31355 11713
rect 37277 11713 37289 11716
rect 37323 11713 37335 11747
rect 37277 11707 37335 11713
rect 24268 11648 24532 11676
rect 24581 11679 24639 11685
rect 24268 11636 24274 11648
rect 24581 11645 24593 11679
rect 24627 11676 24639 11679
rect 25038 11676 25044 11688
rect 24627 11648 25044 11676
rect 24627 11645 24639 11648
rect 24581 11639 24639 11645
rect 24596 11608 24624 11639
rect 25038 11636 25044 11648
rect 25096 11676 25102 11688
rect 26053 11679 26111 11685
rect 26053 11676 26065 11679
rect 25096 11648 26065 11676
rect 25096 11636 25102 11648
rect 26053 11645 26065 11648
rect 26099 11645 26111 11679
rect 26053 11639 26111 11645
rect 27709 11679 27767 11685
rect 27709 11645 27721 11679
rect 27755 11645 27767 11679
rect 27709 11639 27767 11645
rect 22520 11580 23060 11608
rect 23124 11580 24624 11608
rect 22520 11568 22526 11580
rect 22646 11540 22652 11552
rect 20640 11512 22652 11540
rect 22646 11500 22652 11512
rect 22704 11500 22710 11552
rect 22738 11500 22744 11552
rect 22796 11540 22802 11552
rect 23124 11540 23152 11580
rect 22796 11512 23152 11540
rect 23293 11543 23351 11549
rect 22796 11500 22802 11512
rect 23293 11509 23305 11543
rect 23339 11540 23351 11543
rect 25590 11540 25596 11552
rect 23339 11512 25596 11540
rect 23339 11509 23351 11512
rect 23293 11503 23351 11509
rect 25590 11500 25596 11512
rect 25648 11500 25654 11552
rect 26970 11540 26976 11552
rect 26931 11512 26976 11540
rect 26970 11500 26976 11512
rect 27028 11500 27034 11552
rect 27724 11540 27752 11639
rect 29638 11636 29644 11688
rect 29696 11676 29702 11688
rect 30558 11676 30564 11688
rect 29696 11648 30564 11676
rect 29696 11636 29702 11648
rect 30558 11636 30564 11648
rect 30616 11676 30622 11688
rect 31128 11676 31156 11707
rect 30616 11648 31156 11676
rect 30616 11636 30622 11648
rect 31312 11620 31340 11707
rect 37458 11676 37464 11688
rect 37419 11648 37464 11676
rect 37458 11636 37464 11648
rect 37516 11636 37522 11688
rect 29730 11568 29736 11620
rect 29788 11608 29794 11620
rect 31294 11608 31300 11620
rect 29788 11580 31300 11608
rect 29788 11568 29794 11580
rect 31294 11568 31300 11580
rect 31352 11568 31358 11620
rect 37274 11608 37280 11620
rect 31726 11580 37280 11608
rect 27890 11540 27896 11552
rect 27724 11512 27896 11540
rect 27890 11500 27896 11512
rect 27948 11500 27954 11552
rect 27982 11500 27988 11552
rect 28040 11540 28046 11552
rect 29089 11543 29147 11549
rect 29089 11540 29101 11543
rect 28040 11512 29101 11540
rect 28040 11500 28046 11512
rect 29089 11509 29101 11512
rect 29135 11509 29147 11543
rect 30006 11540 30012 11552
rect 29967 11512 30012 11540
rect 29089 11503 29147 11509
rect 30006 11500 30012 11512
rect 30064 11500 30070 11552
rect 30098 11500 30104 11552
rect 30156 11540 30162 11552
rect 31726 11540 31754 11580
rect 37274 11568 37280 11580
rect 37332 11568 37338 11620
rect 30156 11512 31754 11540
rect 30156 11500 30162 11512
rect 1104 11450 48852 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 48852 11450
rect 1104 11376 48852 11398
rect 18046 11336 18052 11348
rect 11532 11308 18052 11336
rect 11532 11209 11560 11308
rect 18046 11296 18052 11308
rect 18104 11336 18110 11348
rect 18693 11339 18751 11345
rect 18693 11336 18705 11339
rect 18104 11308 18705 11336
rect 18104 11296 18110 11308
rect 18693 11305 18705 11308
rect 18739 11305 18751 11339
rect 18693 11299 18751 11305
rect 21818 11296 21824 11348
rect 21876 11336 21882 11348
rect 22557 11339 22615 11345
rect 22557 11336 22569 11339
rect 21876 11308 22569 11336
rect 21876 11296 21882 11308
rect 22557 11305 22569 11308
rect 22603 11305 22615 11339
rect 22557 11299 22615 11305
rect 23474 11296 23480 11348
rect 23532 11336 23538 11348
rect 25777 11339 25835 11345
rect 23532 11308 25452 11336
rect 23532 11296 23538 11308
rect 2041 11203 2099 11209
rect 2041 11169 2053 11203
rect 2087 11200 2099 11203
rect 11517 11203 11575 11209
rect 2087 11172 2774 11200
rect 2087 11169 2099 11172
rect 2041 11163 2099 11169
rect 2498 11132 2504 11144
rect 2459 11104 2504 11132
rect 2498 11092 2504 11104
rect 2556 11092 2562 11144
rect 1854 11064 1860 11076
rect 1815 11036 1860 11064
rect 1854 11024 1860 11036
rect 1912 11024 1918 11076
rect 2746 11064 2774 11172
rect 11517 11169 11529 11203
rect 11563 11169 11575 11203
rect 11698 11200 11704 11212
rect 11659 11172 11704 11200
rect 11517 11163 11575 11169
rect 11698 11160 11704 11172
rect 11756 11160 11762 11212
rect 13078 11200 13084 11212
rect 13039 11172 13084 11200
rect 13078 11160 13084 11172
rect 13136 11160 13142 11212
rect 18966 11160 18972 11212
rect 19024 11200 19030 11212
rect 19245 11203 19303 11209
rect 19245 11200 19257 11203
rect 19024 11172 19257 11200
rect 19024 11160 19030 11172
rect 19245 11169 19257 11172
rect 19291 11169 19303 11203
rect 19245 11163 19303 11169
rect 20254 11160 20260 11212
rect 20312 11200 20318 11212
rect 20714 11200 20720 11212
rect 20312 11172 20720 11200
rect 20312 11160 20318 11172
rect 20714 11160 20720 11172
rect 20772 11160 20778 11212
rect 14182 11132 14188 11144
rect 13280 11104 14188 11132
rect 13280 11064 13308 11104
rect 14182 11092 14188 11104
rect 14240 11092 14246 11144
rect 17313 11135 17371 11141
rect 17313 11101 17325 11135
rect 17359 11132 17371 11135
rect 17954 11132 17960 11144
rect 17359 11104 17960 11132
rect 17359 11101 17371 11104
rect 17313 11095 17371 11101
rect 17954 11092 17960 11104
rect 18012 11132 18018 11144
rect 18012 11104 19288 11132
rect 18012 11092 18018 11104
rect 19260 11076 19288 11104
rect 19426 11092 19432 11144
rect 19484 11132 19490 11144
rect 19521 11135 19579 11141
rect 19521 11132 19533 11135
rect 19484 11104 19533 11132
rect 19484 11092 19490 11104
rect 19521 11101 19533 11104
rect 19567 11101 19579 11135
rect 19521 11095 19579 11101
rect 21177 11135 21235 11141
rect 21177 11101 21189 11135
rect 21223 11132 21235 11135
rect 22002 11132 22008 11144
rect 21223 11104 22008 11132
rect 21223 11101 21235 11104
rect 21177 11095 21235 11101
rect 22002 11092 22008 11104
rect 22060 11132 22066 11144
rect 24397 11135 24455 11141
rect 24397 11132 24409 11135
rect 22060 11104 24409 11132
rect 22060 11092 22066 11104
rect 24397 11101 24409 11104
rect 24443 11132 24455 11135
rect 24443 11104 24808 11132
rect 24443 11101 24455 11104
rect 24397 11095 24455 11101
rect 2746 11036 13308 11064
rect 17580 11067 17638 11073
rect 17580 11033 17592 11067
rect 17626 11064 17638 11067
rect 18782 11064 18788 11076
rect 17626 11036 18788 11064
rect 17626 11033 17638 11036
rect 17580 11027 17638 11033
rect 18782 11024 18788 11036
rect 18840 11024 18846 11076
rect 19242 11024 19248 11076
rect 19300 11024 19306 11076
rect 21444 11067 21502 11073
rect 21444 11033 21456 11067
rect 21490 11064 21502 11067
rect 22278 11064 22284 11076
rect 21490 11036 22284 11064
rect 21490 11033 21502 11036
rect 21444 11027 21502 11033
rect 22278 11024 22284 11036
rect 22336 11024 22342 11076
rect 24670 11073 24676 11076
rect 24664 11064 24676 11073
rect 24631 11036 24676 11064
rect 24664 11027 24676 11036
rect 24670 11024 24676 11027
rect 24728 11024 24734 11076
rect 24780 11064 24808 11104
rect 25424 11064 25452 11308
rect 25777 11305 25789 11339
rect 25823 11336 25835 11339
rect 25958 11336 25964 11348
rect 25823 11308 25964 11336
rect 25823 11305 25835 11308
rect 25777 11299 25835 11305
rect 25958 11296 25964 11308
rect 26016 11296 26022 11348
rect 27154 11296 27160 11348
rect 27212 11336 27218 11348
rect 28813 11339 28871 11345
rect 28813 11336 28825 11339
rect 27212 11308 28825 11336
rect 27212 11296 27218 11308
rect 28813 11305 28825 11308
rect 28859 11305 28871 11339
rect 28813 11299 28871 11305
rect 30009 11339 30067 11345
rect 30009 11305 30021 11339
rect 30055 11336 30067 11339
rect 30466 11336 30472 11348
rect 30055 11308 30472 11336
rect 30055 11305 30067 11308
rect 30009 11299 30067 11305
rect 30466 11296 30472 11308
rect 30524 11296 30530 11348
rect 37369 11339 37427 11345
rect 37369 11305 37381 11339
rect 37415 11336 37427 11339
rect 37458 11336 37464 11348
rect 37415 11308 37464 11336
rect 37415 11305 37427 11308
rect 37369 11299 37427 11305
rect 37458 11296 37464 11308
rect 37516 11296 37522 11348
rect 26142 11228 26148 11280
rect 26200 11268 26206 11280
rect 30098 11268 30104 11280
rect 26200 11240 30104 11268
rect 26200 11228 26206 11240
rect 30098 11228 30104 11240
rect 30156 11228 30162 11280
rect 26326 11160 26332 11212
rect 26384 11200 26390 11212
rect 26513 11203 26571 11209
rect 26513 11200 26525 11203
rect 26384 11172 26525 11200
rect 26384 11160 26390 11172
rect 26513 11169 26525 11172
rect 26559 11200 26571 11203
rect 27154 11200 27160 11212
rect 26559 11172 27160 11200
rect 26559 11169 26571 11172
rect 26513 11163 26571 11169
rect 27154 11160 27160 11172
rect 27212 11160 27218 11212
rect 27890 11160 27896 11212
rect 27948 11200 27954 11212
rect 28261 11203 28319 11209
rect 28261 11200 28273 11203
rect 27948 11172 28273 11200
rect 27948 11160 27954 11172
rect 28261 11169 28273 11172
rect 28307 11200 28319 11203
rect 29546 11200 29552 11212
rect 28307 11172 29552 11200
rect 28307 11169 28319 11172
rect 28261 11163 28319 11169
rect 29546 11160 29552 11172
rect 29604 11160 29610 11212
rect 26234 11132 26240 11144
rect 26195 11104 26240 11132
rect 26234 11092 26240 11104
rect 26292 11092 26298 11144
rect 26418 11092 26424 11144
rect 26476 11132 26482 11144
rect 26476 11104 26569 11132
rect 26476 11092 26482 11104
rect 26602 11092 26608 11144
rect 26660 11132 26666 11144
rect 26660 11104 26705 11132
rect 26660 11092 26666 11104
rect 26786 11092 26792 11144
rect 26844 11132 26850 11144
rect 26844 11104 26937 11132
rect 26844 11092 26850 11104
rect 26970 11092 26976 11144
rect 27028 11132 27034 11144
rect 28721 11135 28779 11141
rect 28721 11132 28733 11135
rect 27028 11104 28733 11132
rect 27028 11092 27034 11104
rect 28721 11101 28733 11104
rect 28767 11101 28779 11135
rect 28902 11132 28908 11144
rect 28863 11104 28908 11132
rect 28721 11095 28779 11101
rect 28902 11092 28908 11104
rect 28960 11092 28966 11144
rect 29564 11132 29592 11160
rect 30742 11141 30748 11144
rect 30469 11135 30527 11141
rect 30469 11132 30481 11135
rect 29564 11104 30481 11132
rect 30469 11101 30481 11104
rect 30515 11101 30527 11135
rect 30736 11132 30748 11141
rect 30703 11104 30748 11132
rect 30469 11095 30527 11101
rect 30736 11095 30748 11104
rect 30742 11092 30748 11095
rect 30800 11092 30806 11144
rect 37274 11132 37280 11144
rect 37235 11104 37280 11132
rect 37274 11092 37280 11104
rect 37332 11092 37338 11144
rect 47118 11132 47124 11144
rect 47079 11104 47124 11132
rect 47118 11092 47124 11104
rect 47176 11092 47182 11144
rect 47946 11132 47952 11144
rect 47907 11104 47952 11132
rect 47946 11092 47952 11104
rect 48004 11092 48010 11144
rect 26436 11064 26464 11092
rect 24780 11036 24900 11064
rect 25424 11036 26464 11064
rect 26804 11064 26832 11092
rect 26804 11036 27108 11064
rect 2590 10996 2596 11008
rect 2551 10968 2596 10996
rect 2590 10956 2596 10968
rect 2648 10956 2654 11008
rect 18322 10956 18328 11008
rect 18380 10996 18386 11008
rect 19150 10996 19156 11008
rect 18380 10968 19156 10996
rect 18380 10956 18386 10968
rect 19150 10956 19156 10968
rect 19208 10956 19214 11008
rect 24872 10996 24900 11036
rect 25314 10996 25320 11008
rect 24872 10968 25320 10996
rect 25314 10956 25320 10968
rect 25372 10956 25378 11008
rect 26970 10996 26976 11008
rect 26931 10968 26976 10996
rect 26970 10956 26976 10968
rect 27028 10956 27034 11008
rect 27080 10996 27108 11036
rect 27522 11024 27528 11076
rect 27580 11064 27586 11076
rect 28077 11067 28135 11073
rect 28077 11064 28089 11067
rect 27580 11036 28089 11064
rect 27580 11024 27586 11036
rect 28077 11033 28089 11036
rect 28123 11033 28135 11067
rect 29638 11064 29644 11076
rect 29599 11036 29644 11064
rect 28077 11027 28135 11033
rect 29638 11024 29644 11036
rect 29696 11024 29702 11076
rect 29825 11067 29883 11073
rect 29825 11033 29837 11067
rect 29871 11064 29883 11067
rect 30374 11064 30380 11076
rect 29871 11036 30380 11064
rect 29871 11033 29883 11036
rect 29825 11027 29883 11033
rect 30374 11024 30380 11036
rect 30432 11024 30438 11076
rect 31294 11024 31300 11076
rect 31352 11064 31358 11076
rect 31352 11036 31892 11064
rect 31352 11024 31358 11036
rect 28350 10996 28356 11008
rect 27080 10968 28356 10996
rect 28350 10956 28356 10968
rect 28408 10956 28414 11008
rect 31864 11005 31892 11036
rect 31849 10999 31907 11005
rect 31849 10965 31861 10999
rect 31895 10965 31907 10999
rect 47210 10996 47216 11008
rect 47171 10968 47216 10996
rect 31849 10959 31907 10965
rect 47210 10956 47216 10968
rect 47268 10956 47274 11008
rect 1104 10906 48852 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 48852 10906
rect 1104 10832 48852 10854
rect 18782 10792 18788 10804
rect 18743 10764 18788 10792
rect 18782 10752 18788 10764
rect 18840 10752 18846 10804
rect 19242 10752 19248 10804
rect 19300 10792 19306 10804
rect 21266 10792 21272 10804
rect 19300 10764 19840 10792
rect 21227 10764 21272 10792
rect 19300 10752 19306 10764
rect 1949 10727 2007 10733
rect 1949 10693 1961 10727
rect 1995 10724 2007 10727
rect 2590 10724 2596 10736
rect 1995 10696 2596 10724
rect 1995 10693 2007 10696
rect 1949 10687 2007 10693
rect 2590 10684 2596 10696
rect 2648 10684 2654 10736
rect 18046 10684 18052 10736
rect 18104 10724 18110 10736
rect 18141 10727 18199 10733
rect 18141 10724 18153 10727
rect 18104 10696 18153 10724
rect 18104 10684 18110 10696
rect 18141 10693 18153 10696
rect 18187 10693 18199 10727
rect 18141 10687 18199 10693
rect 18325 10727 18383 10733
rect 18325 10693 18337 10727
rect 18371 10724 18383 10727
rect 19812 10724 19840 10764
rect 21266 10752 21272 10764
rect 21324 10752 21330 10804
rect 24670 10792 24676 10804
rect 24631 10764 24676 10792
rect 24670 10752 24676 10764
rect 24728 10752 24734 10804
rect 25314 10792 25320 10804
rect 25275 10764 25320 10792
rect 25314 10752 25320 10764
rect 25372 10752 25378 10804
rect 18371 10696 19288 10724
rect 19812 10696 19932 10724
rect 18371 10693 18383 10696
rect 18325 10687 18383 10693
rect 17957 10659 18015 10665
rect 17957 10625 17969 10659
rect 18003 10656 18015 10659
rect 18966 10656 18972 10668
rect 18003 10628 18972 10656
rect 18003 10625 18015 10628
rect 17957 10619 18015 10625
rect 18966 10616 18972 10628
rect 19024 10616 19030 10668
rect 19260 10665 19288 10696
rect 19061 10659 19119 10665
rect 19061 10625 19073 10659
rect 19107 10625 19119 10659
rect 19061 10619 19119 10625
rect 19153 10659 19211 10665
rect 19153 10625 19165 10659
rect 19199 10625 19211 10659
rect 19153 10619 19211 10625
rect 19245 10659 19303 10665
rect 19245 10625 19257 10659
rect 19291 10625 19303 10659
rect 19426 10656 19432 10668
rect 19387 10628 19432 10656
rect 19245 10619 19303 10625
rect 1578 10548 1584 10600
rect 1636 10588 1642 10600
rect 1765 10591 1823 10597
rect 1765 10588 1777 10591
rect 1636 10560 1777 10588
rect 1636 10548 1642 10560
rect 1765 10557 1777 10560
rect 1811 10557 1823 10591
rect 2958 10588 2964 10600
rect 2919 10560 2964 10588
rect 1765 10551 1823 10557
rect 2958 10548 2964 10560
rect 3016 10548 3022 10600
rect 19076 10452 19104 10619
rect 19168 10588 19196 10619
rect 19426 10616 19432 10628
rect 19484 10656 19490 10668
rect 19794 10656 19800 10668
rect 19484 10628 19800 10656
rect 19484 10616 19490 10628
rect 19794 10616 19800 10628
rect 19852 10616 19858 10668
rect 19904 10665 19932 10696
rect 20070 10684 20076 10736
rect 20128 10724 20134 10736
rect 20898 10724 20904 10736
rect 20128 10696 20904 10724
rect 20128 10684 20134 10696
rect 20898 10684 20904 10696
rect 20956 10684 20962 10736
rect 21726 10684 21732 10736
rect 21784 10724 21790 10736
rect 25225 10727 25283 10733
rect 21784 10696 25176 10724
rect 21784 10684 21790 10696
rect 20162 10665 20168 10668
rect 19889 10659 19947 10665
rect 19889 10625 19901 10659
rect 19935 10625 19947 10659
rect 19889 10619 19947 10625
rect 20156 10619 20168 10665
rect 20220 10656 20226 10668
rect 20220 10628 20256 10656
rect 20162 10616 20168 10619
rect 20220 10616 20226 10628
rect 23382 10616 23388 10668
rect 23440 10656 23446 10668
rect 23937 10659 23995 10665
rect 23937 10656 23949 10659
rect 23440 10628 23949 10656
rect 23440 10616 23446 10628
rect 23937 10625 23949 10628
rect 23983 10625 23995 10659
rect 23937 10619 23995 10625
rect 24121 10659 24179 10665
rect 24121 10625 24133 10659
rect 24167 10625 24179 10659
rect 24121 10619 24179 10625
rect 19334 10588 19340 10600
rect 19168 10560 19340 10588
rect 19334 10548 19340 10560
rect 19392 10548 19398 10600
rect 23474 10548 23480 10600
rect 23532 10588 23538 10600
rect 24136 10588 24164 10619
rect 24210 10616 24216 10668
rect 24268 10656 24274 10668
rect 24268 10628 24313 10656
rect 24268 10616 24274 10628
rect 24394 10616 24400 10668
rect 24452 10656 24458 10668
rect 24489 10659 24547 10665
rect 24489 10656 24501 10659
rect 24452 10628 24501 10656
rect 24452 10616 24458 10628
rect 24489 10625 24501 10628
rect 24535 10625 24547 10659
rect 25148 10656 25176 10696
rect 25225 10693 25237 10727
rect 25271 10724 25283 10727
rect 27522 10724 27528 10736
rect 25271 10696 27528 10724
rect 25271 10693 25283 10696
rect 25225 10687 25283 10693
rect 27522 10684 27528 10696
rect 27580 10684 27586 10736
rect 30006 10733 30012 10736
rect 30000 10724 30012 10733
rect 29967 10696 30012 10724
rect 30000 10687 30012 10696
rect 30006 10684 30012 10687
rect 30064 10684 30070 10736
rect 47762 10656 47768 10668
rect 25148 10628 31754 10656
rect 47723 10628 47768 10656
rect 24489 10619 24547 10625
rect 23532 10560 24164 10588
rect 24305 10591 24363 10597
rect 23532 10548 23538 10560
rect 24305 10557 24317 10591
rect 24351 10588 24363 10591
rect 26602 10588 26608 10600
rect 24351 10560 26608 10588
rect 24351 10557 24363 10560
rect 24305 10551 24363 10557
rect 22186 10520 22192 10532
rect 21192 10492 22192 10520
rect 21192 10452 21220 10492
rect 22186 10480 22192 10492
rect 22244 10480 22250 10532
rect 24210 10480 24216 10532
rect 24268 10520 24274 10532
rect 24394 10520 24400 10532
rect 24268 10492 24400 10520
rect 24268 10480 24274 10492
rect 24394 10480 24400 10492
rect 24452 10480 24458 10532
rect 19076 10424 21220 10452
rect 23014 10412 23020 10464
rect 23072 10452 23078 10464
rect 24493 10452 24521 10560
rect 26602 10548 26608 10560
rect 26660 10548 26666 10600
rect 29546 10548 29552 10600
rect 29604 10588 29610 10600
rect 29733 10591 29791 10597
rect 29733 10588 29745 10591
rect 29604 10560 29745 10588
rect 29604 10548 29610 10560
rect 29733 10557 29745 10560
rect 29779 10557 29791 10591
rect 29733 10551 29791 10557
rect 23072 10424 24521 10452
rect 23072 10412 23078 10424
rect 30374 10412 30380 10464
rect 30432 10452 30438 10464
rect 31113 10455 31171 10461
rect 31113 10452 31125 10455
rect 30432 10424 31125 10452
rect 30432 10412 30438 10424
rect 31113 10421 31125 10424
rect 31159 10421 31171 10455
rect 31726 10452 31754 10628
rect 47762 10616 47768 10628
rect 47820 10616 47826 10668
rect 47857 10455 47915 10461
rect 47857 10452 47869 10455
rect 31726 10424 47869 10452
rect 31113 10415 31171 10421
rect 47857 10421 47869 10424
rect 47903 10421 47915 10455
rect 47857 10415 47915 10421
rect 1104 10362 48852 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 48852 10362
rect 1104 10288 48852 10310
rect 1578 10248 1584 10260
rect 1539 10220 1584 10248
rect 1578 10208 1584 10220
rect 1636 10208 1642 10260
rect 20073 10251 20131 10257
rect 20073 10217 20085 10251
rect 20119 10248 20131 10251
rect 20162 10248 20168 10260
rect 20119 10220 20168 10248
rect 20119 10217 20131 10220
rect 20073 10211 20131 10217
rect 20162 10208 20168 10220
rect 20220 10208 20226 10260
rect 27154 10248 27160 10260
rect 27115 10220 27160 10248
rect 27154 10208 27160 10220
rect 27212 10208 27218 10260
rect 19334 10140 19340 10192
rect 19392 10180 19398 10192
rect 20438 10180 20444 10192
rect 19392 10152 20444 10180
rect 19392 10140 19398 10152
rect 20272 10112 20300 10152
rect 20438 10140 20444 10152
rect 20496 10140 20502 10192
rect 20530 10140 20536 10192
rect 20588 10180 20594 10192
rect 47946 10180 47952 10192
rect 20588 10152 20668 10180
rect 20588 10140 20594 10152
rect 20272 10084 20484 10112
rect 1946 10004 1952 10056
rect 2004 10044 2010 10056
rect 2225 10047 2283 10053
rect 2225 10044 2237 10047
rect 2004 10016 2237 10044
rect 2004 10004 2010 10016
rect 2225 10013 2237 10016
rect 2271 10013 2283 10047
rect 2225 10007 2283 10013
rect 2685 10047 2743 10053
rect 2685 10013 2697 10047
rect 2731 10044 2743 10047
rect 3050 10044 3056 10056
rect 2731 10016 3056 10044
rect 2731 10013 2743 10016
rect 2685 10007 2743 10013
rect 3050 10004 3056 10016
rect 3108 10004 3114 10056
rect 20456 10053 20484 10084
rect 20329 10047 20387 10053
rect 20329 10013 20341 10047
rect 20375 10044 20387 10047
rect 20422 10047 20484 10053
rect 20375 10013 20392 10044
rect 20329 10007 20392 10013
rect 20422 10013 20434 10047
rect 20468 10016 20484 10047
rect 20538 10044 20596 10050
rect 20468 10013 20480 10016
rect 20422 10007 20480 10013
rect 20538 10010 20550 10044
rect 20584 10010 20596 10044
rect 19150 9936 19156 9988
rect 19208 9976 19214 9988
rect 19245 9979 19303 9985
rect 19245 9976 19257 9979
rect 19208 9948 19257 9976
rect 19208 9936 19214 9948
rect 19245 9945 19257 9948
rect 19291 9945 19303 9979
rect 19426 9976 19432 9988
rect 19387 9948 19432 9976
rect 19245 9939 19303 9945
rect 19426 9936 19432 9948
rect 19484 9936 19490 9988
rect 2774 9868 2780 9920
rect 2832 9908 2838 9920
rect 2832 9880 2877 9908
rect 2832 9868 2838 9880
rect 19334 9868 19340 9920
rect 19392 9908 19398 9920
rect 19613 9911 19671 9917
rect 19613 9908 19625 9911
rect 19392 9880 19625 9908
rect 19392 9868 19398 9880
rect 19613 9877 19625 9880
rect 19659 9877 19671 9911
rect 20364 9908 20392 10007
rect 20538 10004 20596 10010
rect 20548 9976 20576 10004
rect 20640 9976 20668 10152
rect 46308 10152 47952 10180
rect 25314 10072 25320 10124
rect 25372 10112 25378 10124
rect 46308 10121 46336 10152
rect 47946 10140 47952 10152
rect 48004 10140 48010 10192
rect 25777 10115 25835 10121
rect 25777 10112 25789 10115
rect 25372 10084 25789 10112
rect 25372 10072 25378 10084
rect 25777 10081 25789 10084
rect 25823 10081 25835 10115
rect 25777 10075 25835 10081
rect 46293 10115 46351 10121
rect 46293 10081 46305 10115
rect 46339 10081 46351 10115
rect 46293 10075 46351 10081
rect 46477 10115 46535 10121
rect 46477 10081 46489 10115
rect 46523 10112 46535 10115
rect 47210 10112 47216 10124
rect 46523 10084 47216 10112
rect 46523 10081 46535 10084
rect 46477 10075 46535 10081
rect 47210 10072 47216 10084
rect 47268 10072 47274 10124
rect 48130 10112 48136 10124
rect 48091 10084 48136 10112
rect 48130 10072 48136 10084
rect 48188 10072 48194 10124
rect 20717 10047 20775 10053
rect 20717 10013 20729 10047
rect 20763 10044 20775 10047
rect 20990 10044 20996 10056
rect 20763 10016 20996 10044
rect 20763 10013 20775 10016
rect 20717 10007 20775 10013
rect 20990 10004 20996 10016
rect 21048 10004 21054 10056
rect 26044 10047 26102 10053
rect 26044 10013 26056 10047
rect 26090 10044 26102 10047
rect 26970 10044 26976 10056
rect 26090 10016 26976 10044
rect 26090 10013 26102 10016
rect 26044 10007 26102 10013
rect 26970 10004 26976 10016
rect 27028 10004 27034 10056
rect 20548 9948 20668 9976
rect 22094 9908 22100 9920
rect 20364 9880 22100 9908
rect 19613 9871 19671 9877
rect 22094 9868 22100 9880
rect 22152 9908 22158 9920
rect 26602 9908 26608 9920
rect 22152 9880 26608 9908
rect 22152 9868 22158 9880
rect 26602 9868 26608 9880
rect 26660 9868 26666 9920
rect 1104 9818 48852 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 48852 9818
rect 1104 9744 48852 9766
rect 18598 9664 18604 9716
rect 18656 9704 18662 9716
rect 18656 9676 19748 9704
rect 18656 9664 18662 9676
rect 2133 9639 2191 9645
rect 2133 9605 2145 9639
rect 2179 9636 2191 9639
rect 2774 9636 2780 9648
rect 2179 9608 2780 9636
rect 2179 9605 2191 9608
rect 2133 9599 2191 9605
rect 2774 9596 2780 9608
rect 2832 9596 2838 9648
rect 4062 9596 4068 9648
rect 4120 9636 4126 9648
rect 12526 9636 12532 9648
rect 4120 9608 12532 9636
rect 4120 9596 4126 9608
rect 12526 9596 12532 9608
rect 12584 9596 12590 9648
rect 17954 9636 17960 9648
rect 17328 9608 17960 9636
rect 1946 9568 1952 9580
rect 1907 9540 1952 9568
rect 1946 9528 1952 9540
rect 2004 9528 2010 9580
rect 17328 9577 17356 9608
rect 17954 9596 17960 9608
rect 18012 9596 18018 9648
rect 19720 9636 19748 9676
rect 19978 9664 19984 9716
rect 20036 9704 20042 9716
rect 20990 9704 20996 9716
rect 20036 9676 20996 9704
rect 20036 9664 20042 9676
rect 20990 9664 20996 9676
rect 21048 9664 21054 9716
rect 27816 9676 28304 9704
rect 19720 9608 23612 9636
rect 17313 9571 17371 9577
rect 17313 9537 17325 9571
rect 17359 9537 17371 9571
rect 17313 9531 17371 9537
rect 17580 9571 17638 9577
rect 17580 9537 17592 9571
rect 17626 9568 17638 9571
rect 17626 9540 18552 9568
rect 17626 9537 17638 9540
rect 17580 9531 17638 9537
rect 2866 9500 2872 9512
rect 2827 9472 2872 9500
rect 2866 9460 2872 9472
rect 2924 9460 2930 9512
rect 18524 9432 18552 9540
rect 18690 9528 18696 9580
rect 18748 9568 18754 9580
rect 19429 9574 19487 9577
rect 19260 9571 19487 9574
rect 19260 9568 19441 9571
rect 18748 9546 19441 9568
rect 18748 9540 19288 9546
rect 18748 9528 18754 9540
rect 19429 9537 19441 9546
rect 19475 9537 19487 9571
rect 19429 9531 19487 9537
rect 19521 9571 19579 9577
rect 19521 9537 19533 9571
rect 19567 9537 19579 9571
rect 19521 9531 19579 9537
rect 19536 9500 19564 9531
rect 19610 9528 19616 9580
rect 19668 9568 19674 9580
rect 19797 9571 19855 9577
rect 19668 9540 19713 9568
rect 19668 9528 19674 9540
rect 19797 9537 19809 9571
rect 19843 9568 19855 9571
rect 19978 9568 19984 9580
rect 19843 9540 19984 9568
rect 19843 9537 19855 9540
rect 19797 9531 19855 9537
rect 19978 9528 19984 9540
rect 20036 9528 20042 9580
rect 20254 9528 20260 9580
rect 20312 9568 20318 9580
rect 23017 9571 23075 9577
rect 23017 9568 23029 9571
rect 20312 9540 23029 9568
rect 20312 9528 20318 9540
rect 23017 9537 23029 9540
rect 23063 9537 23075 9571
rect 23584 9568 23612 9608
rect 23658 9596 23664 9648
rect 23716 9636 23722 9648
rect 24397 9639 24455 9645
rect 24397 9636 24409 9639
rect 23716 9608 24409 9636
rect 23716 9596 23722 9608
rect 24397 9605 24409 9608
rect 24443 9605 24455 9639
rect 27816 9636 27844 9676
rect 24397 9599 24455 9605
rect 26344 9608 27844 9636
rect 26344 9568 26372 9608
rect 23584 9540 26372 9568
rect 23017 9531 23075 9537
rect 26418 9528 26424 9580
rect 26476 9568 26482 9580
rect 27065 9571 27123 9577
rect 27065 9568 27077 9571
rect 26476 9540 27077 9568
rect 26476 9528 26482 9540
rect 27065 9537 27077 9540
rect 27111 9537 27123 9571
rect 27065 9531 27123 9537
rect 27249 9571 27307 9577
rect 27249 9537 27261 9571
rect 27295 9568 27307 9571
rect 27798 9568 27804 9580
rect 27295 9540 27804 9568
rect 27295 9537 27307 9540
rect 27249 9531 27307 9537
rect 27798 9528 27804 9540
rect 27856 9528 27862 9580
rect 27982 9528 27988 9580
rect 28040 9568 28046 9580
rect 28149 9571 28207 9577
rect 28149 9568 28161 9571
rect 28040 9540 28161 9568
rect 28040 9528 28046 9540
rect 28149 9537 28161 9540
rect 28195 9537 28207 9571
rect 28276 9568 28304 9676
rect 38562 9596 38568 9648
rect 38620 9636 38626 9648
rect 46842 9636 46848 9648
rect 38620 9608 46848 9636
rect 38620 9596 38626 9608
rect 46842 9596 46848 9608
rect 46900 9596 46906 9648
rect 29917 9571 29975 9577
rect 29917 9568 29929 9571
rect 28276 9540 29929 9568
rect 28149 9531 28207 9537
rect 29917 9537 29929 9540
rect 29963 9568 29975 9571
rect 30561 9571 30619 9577
rect 30561 9568 30573 9571
rect 29963 9540 30573 9568
rect 29963 9537 29975 9540
rect 29917 9531 29975 9537
rect 30561 9537 30573 9540
rect 30607 9568 30619 9571
rect 31478 9568 31484 9580
rect 30607 9540 31484 9568
rect 30607 9537 30619 9540
rect 30561 9531 30619 9537
rect 31478 9528 31484 9540
rect 31536 9528 31542 9580
rect 20438 9500 20444 9512
rect 19536 9472 20444 9500
rect 20438 9460 20444 9472
rect 20496 9460 20502 9512
rect 23293 9503 23351 9509
rect 23293 9469 23305 9503
rect 23339 9500 23351 9503
rect 23382 9500 23388 9512
rect 23339 9472 23388 9500
rect 23339 9469 23351 9472
rect 23293 9463 23351 9469
rect 23382 9460 23388 9472
rect 23440 9460 23446 9512
rect 26970 9460 26976 9512
rect 27028 9500 27034 9512
rect 27890 9500 27896 9512
rect 27028 9472 27896 9500
rect 27028 9460 27034 9472
rect 27890 9460 27896 9472
rect 27948 9460 27954 9512
rect 19153 9435 19211 9441
rect 19153 9432 19165 9435
rect 18524 9404 19165 9432
rect 19153 9401 19165 9404
rect 19199 9401 19211 9435
rect 19153 9395 19211 9401
rect 17954 9324 17960 9376
rect 18012 9364 18018 9376
rect 18693 9367 18751 9373
rect 18693 9364 18705 9367
rect 18012 9336 18705 9364
rect 18012 9324 18018 9336
rect 18693 9333 18705 9336
rect 18739 9364 18751 9367
rect 19426 9364 19432 9376
rect 18739 9336 19432 9364
rect 18739 9333 18751 9336
rect 18693 9327 18751 9333
rect 19426 9324 19432 9336
rect 19484 9324 19490 9376
rect 23842 9324 23848 9376
rect 23900 9364 23906 9376
rect 24489 9367 24547 9373
rect 24489 9364 24501 9367
rect 23900 9336 24501 9364
rect 23900 9324 23906 9336
rect 24489 9333 24501 9336
rect 24535 9364 24547 9367
rect 24946 9364 24952 9376
rect 24535 9336 24952 9364
rect 24535 9333 24547 9336
rect 24489 9327 24547 9333
rect 24946 9324 24952 9336
rect 25004 9324 25010 9376
rect 27433 9367 27491 9373
rect 27433 9333 27445 9367
rect 27479 9364 27491 9367
rect 27706 9364 27712 9376
rect 27479 9336 27712 9364
rect 27479 9333 27491 9336
rect 27433 9327 27491 9333
rect 27706 9324 27712 9336
rect 27764 9324 27770 9376
rect 27798 9324 27804 9376
rect 27856 9364 27862 9376
rect 28258 9364 28264 9376
rect 27856 9336 28264 9364
rect 27856 9324 27862 9336
rect 28258 9324 28264 9336
rect 28316 9364 28322 9376
rect 29273 9367 29331 9373
rect 29273 9364 29285 9367
rect 28316 9336 29285 9364
rect 28316 9324 28322 9336
rect 29273 9333 29285 9336
rect 29319 9333 29331 9367
rect 30006 9364 30012 9376
rect 29967 9336 30012 9364
rect 29273 9327 29331 9333
rect 30006 9324 30012 9336
rect 30064 9324 30070 9376
rect 30650 9364 30656 9376
rect 30611 9336 30656 9364
rect 30650 9324 30656 9336
rect 30708 9324 30714 9376
rect 1104 9274 48852 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 48852 9274
rect 1104 9200 48852 9222
rect 17770 9120 17776 9172
rect 17828 9160 17834 9172
rect 22370 9160 22376 9172
rect 17828 9132 22376 9160
rect 17828 9120 17834 9132
rect 22370 9120 22376 9132
rect 22428 9120 22434 9172
rect 27249 9163 27307 9169
rect 27249 9129 27261 9163
rect 27295 9160 27307 9163
rect 27982 9160 27988 9172
rect 27295 9132 27988 9160
rect 27295 9129 27307 9132
rect 27249 9123 27307 9129
rect 27982 9120 27988 9132
rect 28040 9120 28046 9172
rect 24946 9052 24952 9104
rect 25004 9052 25010 9104
rect 48038 9092 48044 9104
rect 27356 9064 48044 9092
rect 19242 9024 19248 9036
rect 19203 8996 19248 9024
rect 19242 8984 19248 8996
rect 19300 8984 19306 9036
rect 22833 9027 22891 9033
rect 22833 8993 22845 9027
rect 22879 9024 22891 9027
rect 24486 9024 24492 9036
rect 22879 8996 24492 9024
rect 22879 8993 22891 8996
rect 22833 8987 22891 8993
rect 24486 8984 24492 8996
rect 24544 8984 24550 9036
rect 24964 9024 24992 9052
rect 24872 8996 24992 9024
rect 19150 8916 19156 8968
rect 19208 8956 19214 8968
rect 21269 8959 21327 8965
rect 19208 8928 21128 8956
rect 19208 8916 19214 8928
rect 19512 8891 19570 8897
rect 19512 8857 19524 8891
rect 19558 8857 19570 8891
rect 19512 8851 19570 8857
rect 19426 8780 19432 8832
rect 19484 8820 19490 8832
rect 19536 8820 19564 8851
rect 19978 8848 19984 8900
rect 20036 8888 20042 8900
rect 20990 8888 20996 8900
rect 20036 8860 20996 8888
rect 20036 8848 20042 8860
rect 20990 8848 20996 8860
rect 21048 8848 21054 8900
rect 21100 8897 21128 8928
rect 21269 8925 21281 8959
rect 21315 8956 21327 8959
rect 22922 8956 22928 8968
rect 21315 8928 22928 8956
rect 21315 8925 21327 8928
rect 21269 8919 21327 8925
rect 22922 8916 22928 8928
rect 22980 8916 22986 8968
rect 23109 8959 23167 8965
rect 23109 8925 23121 8959
rect 23155 8956 23167 8959
rect 23290 8956 23296 8968
rect 23155 8928 23296 8956
rect 23155 8925 23167 8928
rect 23109 8919 23167 8925
rect 23290 8916 23296 8928
rect 23348 8916 23354 8968
rect 23658 8916 23664 8968
rect 23716 8956 23722 8968
rect 24872 8965 24900 8996
rect 24719 8959 24777 8965
rect 24719 8956 24731 8959
rect 23716 8928 24731 8956
rect 23716 8916 23722 8928
rect 24719 8925 24731 8928
rect 24765 8925 24777 8959
rect 24719 8919 24777 8925
rect 24854 8959 24912 8965
rect 24854 8925 24866 8959
rect 24900 8925 24912 8959
rect 24854 8919 24912 8925
rect 24949 8959 25007 8965
rect 24949 8925 24961 8959
rect 24995 8956 25007 8959
rect 25038 8956 25044 8968
rect 24995 8928 25044 8956
rect 24995 8925 25007 8928
rect 24949 8919 25007 8925
rect 25038 8916 25044 8928
rect 25096 8916 25102 8968
rect 25130 8916 25136 8968
rect 25188 8956 25194 8968
rect 26418 8956 26424 8968
rect 25188 8928 25233 8956
rect 26379 8928 26424 8956
rect 25188 8916 25194 8928
rect 26418 8916 26424 8928
rect 26476 8916 26482 8968
rect 27356 8956 27384 9064
rect 48038 9052 48044 9064
rect 48096 9052 48102 9104
rect 27798 9024 27804 9036
rect 27632 8996 27804 9024
rect 27632 8965 27660 8996
rect 27798 8984 27804 8996
rect 27856 8984 27862 9036
rect 30006 9024 30012 9036
rect 29967 8996 30012 9024
rect 30006 8984 30012 8996
rect 30064 8984 30070 9036
rect 30282 9024 30288 9036
rect 30243 8996 30288 9024
rect 30282 8984 30288 8996
rect 30340 8984 30346 9036
rect 27479 8959 27537 8965
rect 27479 8956 27491 8959
rect 27356 8928 27491 8956
rect 27479 8925 27491 8928
rect 27525 8925 27537 8959
rect 27479 8919 27537 8925
rect 27614 8959 27672 8965
rect 27614 8925 27626 8959
rect 27660 8925 27672 8959
rect 27614 8919 27672 8925
rect 27706 8916 27712 8968
rect 27764 8956 27770 8968
rect 27764 8928 27809 8956
rect 27764 8916 27770 8928
rect 27890 8916 27896 8968
rect 27948 8956 27954 8968
rect 29825 8959 29883 8965
rect 27948 8928 27993 8956
rect 27948 8916 27954 8928
rect 29825 8925 29837 8959
rect 29871 8925 29883 8959
rect 29825 8919 29883 8925
rect 21085 8891 21143 8897
rect 21085 8857 21097 8891
rect 21131 8888 21143 8891
rect 21174 8888 21180 8900
rect 21131 8860 21180 8888
rect 21131 8857 21143 8860
rect 21085 8851 21143 8857
rect 21174 8848 21180 8860
rect 21232 8848 21238 8900
rect 22005 8891 22063 8897
rect 22005 8857 22017 8891
rect 22051 8857 22063 8891
rect 22186 8888 22192 8900
rect 22147 8860 22192 8888
rect 22005 8851 22063 8857
rect 20622 8820 20628 8832
rect 19484 8792 19564 8820
rect 20583 8792 20628 8820
rect 19484 8780 19490 8792
rect 20622 8780 20628 8792
rect 20680 8780 20686 8832
rect 20806 8780 20812 8832
rect 20864 8820 20870 8832
rect 21453 8823 21511 8829
rect 21453 8820 21465 8823
rect 20864 8792 21465 8820
rect 20864 8780 20870 8792
rect 21453 8789 21465 8792
rect 21499 8789 21511 8823
rect 22020 8820 22048 8851
rect 22186 8848 22192 8860
rect 22244 8848 22250 8900
rect 23382 8888 23388 8900
rect 22296 8860 23388 8888
rect 22296 8820 22324 8860
rect 23382 8848 23388 8860
rect 23440 8848 23446 8900
rect 26602 8888 26608 8900
rect 26563 8860 26608 8888
rect 26602 8848 26608 8860
rect 26660 8848 26666 8900
rect 29840 8888 29868 8919
rect 30374 8888 30380 8900
rect 29840 8860 30380 8888
rect 30374 8848 30380 8860
rect 30432 8848 30438 8900
rect 47946 8888 47952 8900
rect 47907 8860 47952 8888
rect 47946 8848 47952 8860
rect 48004 8848 48010 8900
rect 22020 8792 22324 8820
rect 22373 8823 22431 8829
rect 21453 8783 21511 8789
rect 22373 8789 22385 8823
rect 22419 8820 22431 8823
rect 23198 8820 23204 8832
rect 22419 8792 23204 8820
rect 22419 8789 22431 8792
rect 22373 8783 22431 8789
rect 23198 8780 23204 8792
rect 23256 8780 23262 8832
rect 24489 8823 24547 8829
rect 24489 8789 24501 8823
rect 24535 8820 24547 8823
rect 24946 8820 24952 8832
rect 24535 8792 24952 8820
rect 24535 8789 24547 8792
rect 24489 8783 24547 8789
rect 24946 8780 24952 8792
rect 25004 8780 25010 8832
rect 26789 8823 26847 8829
rect 26789 8789 26801 8823
rect 26835 8820 26847 8823
rect 27062 8820 27068 8832
rect 26835 8792 27068 8820
rect 26835 8789 26847 8792
rect 26789 8783 26847 8789
rect 27062 8780 27068 8792
rect 27120 8780 27126 8832
rect 38286 8780 38292 8832
rect 38344 8820 38350 8832
rect 48041 8823 48099 8829
rect 48041 8820 48053 8823
rect 38344 8792 48053 8820
rect 38344 8780 38350 8792
rect 48041 8789 48053 8792
rect 48087 8789 48099 8823
rect 48041 8783 48099 8789
rect 1104 8730 48852 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 48852 8730
rect 1104 8656 48852 8678
rect 3602 8576 3608 8628
rect 3660 8616 3666 8628
rect 30282 8616 30288 8628
rect 3660 8588 30288 8616
rect 3660 8576 3666 8588
rect 30282 8576 30288 8588
rect 30340 8576 30346 8628
rect 47857 8619 47915 8625
rect 47857 8616 47869 8619
rect 31726 8588 47869 8616
rect 20438 8508 20444 8560
rect 20496 8548 20502 8560
rect 20496 8520 20757 8548
rect 20496 8508 20502 8520
rect 1854 8480 1860 8492
rect 1815 8452 1860 8480
rect 1854 8440 1860 8452
rect 1912 8440 1918 8492
rect 17954 8480 17960 8492
rect 17915 8452 17960 8480
rect 17954 8440 17960 8452
rect 18012 8440 18018 8492
rect 20729 8489 20757 8520
rect 21542 8508 21548 8560
rect 21600 8548 21606 8560
rect 22005 8551 22063 8557
rect 22005 8548 22017 8551
rect 21600 8520 22017 8548
rect 21600 8508 21606 8520
rect 22005 8517 22017 8520
rect 22051 8517 22063 8551
rect 22005 8511 22063 8517
rect 22094 8508 22100 8560
rect 22152 8548 22158 8560
rect 23106 8557 23112 8560
rect 22152 8520 23060 8548
rect 22152 8508 22158 8520
rect 20579 8483 20637 8489
rect 20579 8480 20591 8483
rect 20364 8452 20591 8480
rect 18138 8412 18144 8424
rect 18099 8384 18144 8412
rect 18138 8372 18144 8384
rect 18196 8372 18202 8424
rect 19334 8412 19340 8424
rect 19295 8384 19340 8412
rect 19334 8372 19340 8384
rect 19392 8372 19398 8424
rect 2133 8347 2191 8353
rect 2133 8313 2145 8347
rect 2179 8344 2191 8347
rect 20254 8344 20260 8356
rect 2179 8316 20260 8344
rect 2179 8313 2191 8316
rect 2133 8307 2191 8313
rect 20254 8304 20260 8316
rect 20312 8304 20318 8356
rect 20364 8344 20392 8452
rect 20579 8449 20591 8452
rect 20625 8449 20637 8483
rect 20579 8443 20637 8449
rect 20698 8483 20757 8489
rect 20698 8449 20710 8483
rect 20744 8452 20757 8483
rect 20744 8449 20756 8452
rect 20698 8443 20756 8449
rect 20806 8440 20812 8492
rect 20864 8480 20870 8492
rect 20864 8452 20909 8480
rect 20864 8440 20870 8452
rect 20990 8440 20996 8492
rect 21048 8480 21054 8492
rect 21048 8452 21093 8480
rect 21048 8440 21054 8452
rect 21174 8440 21180 8492
rect 21232 8480 21238 8492
rect 22848 8489 22876 8520
rect 21821 8483 21879 8489
rect 21821 8480 21833 8483
rect 21232 8452 21833 8480
rect 21232 8440 21238 8452
rect 21821 8449 21833 8452
rect 21867 8449 21879 8483
rect 21821 8443 21879 8449
rect 22833 8483 22891 8489
rect 22833 8449 22845 8483
rect 22879 8449 22891 8483
rect 23032 8480 23060 8520
rect 23100 8511 23112 8557
rect 23164 8548 23170 8560
rect 23164 8520 23200 8548
rect 23106 8508 23112 8511
rect 23164 8508 23170 8520
rect 25682 8508 25688 8560
rect 25740 8548 25746 8560
rect 29917 8551 29975 8557
rect 25740 8520 28028 8548
rect 25740 8508 25746 8520
rect 24857 8483 24915 8489
rect 24857 8480 24869 8483
rect 23032 8452 24869 8480
rect 22833 8443 22891 8449
rect 24857 8449 24869 8452
rect 24903 8449 24915 8483
rect 24857 8443 24915 8449
rect 24946 8440 24952 8492
rect 25004 8480 25010 8492
rect 25113 8483 25171 8489
rect 25113 8480 25125 8483
rect 25004 8452 25125 8480
rect 25004 8440 25010 8452
rect 25113 8449 25125 8452
rect 25159 8449 25171 8483
rect 26970 8480 26976 8492
rect 26931 8452 26976 8480
rect 25113 8443 25171 8449
rect 26970 8440 26976 8452
rect 27028 8440 27034 8492
rect 27246 8489 27252 8492
rect 27240 8443 27252 8489
rect 27304 8480 27310 8492
rect 27304 8452 27340 8480
rect 27246 8440 27252 8443
rect 27304 8440 27310 8452
rect 28000 8412 28028 8520
rect 29917 8517 29929 8551
rect 29963 8548 29975 8551
rect 30650 8548 30656 8560
rect 29963 8520 30656 8548
rect 29963 8517 29975 8520
rect 29917 8511 29975 8517
rect 30650 8508 30656 8520
rect 30708 8508 30714 8560
rect 31726 8548 31754 8588
rect 47857 8585 47869 8588
rect 47903 8585 47915 8619
rect 47857 8579 47915 8585
rect 31128 8520 31754 8548
rect 29730 8480 29736 8492
rect 29691 8452 29736 8480
rect 29730 8440 29736 8452
rect 29788 8440 29794 8492
rect 31128 8412 31156 8520
rect 47762 8480 47768 8492
rect 47723 8452 47768 8480
rect 47762 8440 47768 8452
rect 47820 8440 47826 8492
rect 28000 8384 31156 8412
rect 31205 8415 31263 8421
rect 31205 8381 31217 8415
rect 31251 8381 31263 8415
rect 31205 8375 31263 8381
rect 21818 8344 21824 8356
rect 20364 8316 21824 8344
rect 21818 8304 21824 8316
rect 21876 8304 21882 8356
rect 21910 8304 21916 8356
rect 21968 8344 21974 8356
rect 22189 8347 22247 8353
rect 22189 8344 22201 8347
rect 21968 8316 22201 8344
rect 21968 8304 21974 8316
rect 22189 8313 22201 8316
rect 22235 8313 22247 8347
rect 24210 8344 24216 8356
rect 24123 8316 24216 8344
rect 22189 8307 22247 8313
rect 24210 8304 24216 8316
rect 24268 8304 24274 8356
rect 26234 8344 26240 8356
rect 26147 8316 26240 8344
rect 26234 8304 26240 8316
rect 26292 8344 26298 8356
rect 26786 8344 26792 8356
rect 26292 8316 26792 8344
rect 26292 8304 26298 8316
rect 26786 8304 26792 8316
rect 26844 8304 26850 8356
rect 29822 8304 29828 8356
rect 29880 8344 29886 8356
rect 31220 8344 31248 8375
rect 29880 8316 31248 8344
rect 29880 8304 29886 8316
rect 20346 8276 20352 8288
rect 20307 8248 20352 8276
rect 20346 8236 20352 8248
rect 20404 8236 20410 8288
rect 20622 8236 20628 8288
rect 20680 8276 20686 8288
rect 21542 8276 21548 8288
rect 20680 8248 21548 8276
rect 20680 8236 20686 8248
rect 21542 8236 21548 8248
rect 21600 8236 21606 8288
rect 22278 8236 22284 8288
rect 22336 8276 22342 8288
rect 24228 8276 24256 8304
rect 22336 8248 24256 8276
rect 22336 8236 22342 8248
rect 26602 8236 26608 8288
rect 26660 8276 26666 8288
rect 28353 8279 28411 8285
rect 28353 8276 28365 8279
rect 26660 8248 28365 8276
rect 26660 8236 26666 8248
rect 28353 8245 28365 8248
rect 28399 8245 28411 8279
rect 28353 8239 28411 8245
rect 1104 8186 48852 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 48852 8186
rect 1104 8112 48852 8134
rect 18138 8032 18144 8084
rect 18196 8072 18202 8084
rect 18509 8075 18567 8081
rect 18509 8072 18521 8075
rect 18196 8044 18521 8072
rect 18196 8032 18202 8044
rect 18509 8041 18521 8044
rect 18555 8041 18567 8075
rect 18509 8035 18567 8041
rect 20346 8032 20352 8084
rect 20404 8072 20410 8084
rect 22922 8072 22928 8084
rect 20404 8044 21588 8072
rect 22835 8044 22928 8072
rect 20404 8032 20410 8044
rect 2130 7964 2136 8016
rect 2188 8004 2194 8016
rect 7742 8004 7748 8016
rect 2188 7976 7748 8004
rect 2188 7964 2194 7976
rect 7742 7964 7748 7976
rect 7800 7964 7806 8016
rect 18690 7964 18696 8016
rect 18748 8004 18754 8016
rect 18748 7976 20760 8004
rect 18748 7964 18754 7976
rect 19245 7939 19303 7945
rect 19245 7905 19257 7939
rect 19291 7936 19303 7939
rect 20622 7936 20628 7948
rect 19291 7908 20628 7936
rect 19291 7905 19303 7908
rect 19245 7899 19303 7905
rect 20622 7896 20628 7908
rect 20680 7896 20686 7948
rect 20732 7945 20760 7976
rect 20717 7939 20775 7945
rect 20717 7905 20729 7939
rect 20763 7905 20775 7939
rect 21560 7936 21588 8044
rect 22922 8032 22928 8044
rect 22980 8072 22986 8084
rect 22980 8044 24992 8072
rect 22980 8032 22986 8044
rect 24964 8004 24992 8044
rect 25038 8032 25044 8084
rect 25096 8072 25102 8084
rect 25869 8075 25927 8081
rect 25869 8072 25881 8075
rect 25096 8044 25881 8072
rect 25096 8032 25102 8044
rect 25869 8041 25881 8044
rect 25915 8041 25927 8075
rect 25869 8035 25927 8041
rect 26605 8075 26663 8081
rect 26605 8041 26617 8075
rect 26651 8072 26663 8075
rect 27246 8072 27252 8084
rect 26651 8044 27252 8072
rect 26651 8041 26663 8044
rect 26605 8035 26663 8041
rect 27246 8032 27252 8044
rect 27304 8032 27310 8084
rect 24964 7976 31754 8004
rect 21560 7908 21680 7936
rect 20717 7899 20775 7905
rect 1394 7868 1400 7880
rect 1355 7840 1400 7868
rect 1394 7828 1400 7840
rect 1452 7828 1458 7880
rect 18417 7871 18475 7877
rect 18417 7837 18429 7871
rect 18463 7868 18475 7871
rect 18598 7868 18604 7880
rect 18463 7840 18604 7868
rect 18463 7837 18475 7840
rect 18417 7831 18475 7837
rect 18598 7828 18604 7840
rect 18656 7828 18662 7880
rect 21545 7871 21603 7877
rect 21545 7837 21557 7871
rect 21591 7837 21603 7871
rect 21652 7868 21680 7908
rect 23842 7896 23848 7948
rect 23900 7936 23906 7948
rect 27798 7936 27804 7948
rect 23900 7908 27804 7936
rect 23900 7896 23906 7908
rect 21801 7871 21859 7877
rect 21801 7868 21813 7871
rect 21652 7840 21813 7868
rect 21545 7831 21603 7837
rect 21801 7837 21813 7840
rect 21847 7837 21859 7871
rect 21801 7831 21859 7837
rect 18874 7760 18880 7812
rect 18932 7800 18938 7812
rect 19429 7803 19487 7809
rect 19429 7800 19441 7803
rect 18932 7772 19441 7800
rect 18932 7760 18938 7772
rect 19429 7769 19441 7772
rect 19475 7769 19487 7803
rect 19429 7763 19487 7769
rect 1581 7735 1639 7741
rect 1581 7701 1593 7735
rect 1627 7732 1639 7735
rect 16666 7732 16672 7744
rect 1627 7704 16672 7732
rect 1627 7701 1639 7704
rect 1581 7695 1639 7701
rect 16666 7692 16672 7704
rect 16724 7692 16730 7744
rect 21560 7732 21588 7831
rect 23014 7828 23020 7880
rect 23072 7868 23078 7880
rect 24761 7877 24789 7908
rect 24627 7871 24685 7877
rect 24627 7868 24639 7871
rect 23072 7840 24639 7868
rect 23072 7828 23078 7840
rect 24627 7837 24639 7840
rect 24673 7837 24685 7871
rect 24627 7831 24685 7837
rect 24746 7871 24804 7877
rect 24746 7837 24758 7871
rect 24792 7837 24804 7871
rect 24746 7831 24804 7837
rect 24862 7871 24920 7877
rect 24862 7837 24874 7871
rect 24908 7837 24920 7871
rect 25038 7868 25044 7880
rect 24999 7840 25044 7868
rect 24862 7831 24920 7837
rect 23382 7800 23388 7812
rect 23343 7772 23388 7800
rect 23382 7760 23388 7772
rect 23440 7760 23446 7812
rect 23566 7800 23572 7812
rect 23527 7772 23572 7800
rect 23566 7760 23572 7772
rect 23624 7760 23630 7812
rect 23753 7803 23811 7809
rect 23753 7769 23765 7803
rect 23799 7800 23811 7803
rect 24872 7800 24900 7831
rect 25038 7828 25044 7840
rect 25096 7828 25102 7880
rect 25314 7828 25320 7880
rect 25372 7868 25378 7880
rect 25501 7871 25559 7877
rect 25501 7868 25513 7871
rect 25372 7840 25513 7868
rect 25372 7828 25378 7840
rect 25501 7837 25513 7840
rect 25547 7868 25559 7871
rect 26418 7868 26424 7880
rect 25547 7840 26424 7868
rect 25547 7837 25559 7840
rect 25501 7831 25559 7837
rect 26418 7828 26424 7840
rect 26476 7828 26482 7880
rect 26878 7868 26884 7880
rect 26839 7840 26884 7868
rect 26878 7828 26884 7840
rect 26936 7828 26942 7880
rect 26988 7877 27016 7908
rect 27798 7896 27804 7908
rect 27856 7896 27862 7948
rect 26973 7871 27031 7877
rect 26973 7837 26985 7871
rect 27019 7837 27031 7871
rect 26973 7831 27031 7837
rect 27062 7828 27068 7880
rect 27120 7877 27126 7880
rect 27120 7868 27128 7877
rect 27120 7840 27165 7868
rect 27120 7831 27128 7840
rect 27120 7828 27126 7831
rect 27246 7828 27252 7880
rect 27304 7868 27310 7880
rect 27890 7868 27896 7880
rect 27304 7840 27896 7868
rect 27304 7828 27310 7840
rect 27890 7828 27896 7840
rect 27948 7828 27954 7880
rect 31726 7868 31754 7976
rect 37274 7868 37280 7880
rect 31726 7840 37280 7868
rect 37274 7828 37280 7840
rect 37332 7828 37338 7880
rect 46290 7868 46296 7880
rect 46251 7840 46296 7868
rect 46290 7828 46296 7840
rect 46348 7828 46354 7880
rect 23799 7772 24900 7800
rect 25685 7803 25743 7809
rect 23799 7769 23811 7772
rect 23753 7763 23811 7769
rect 25685 7769 25697 7803
rect 25731 7800 25743 7803
rect 26234 7800 26240 7812
rect 25731 7772 26240 7800
rect 25731 7769 25743 7772
rect 25685 7763 25743 7769
rect 26234 7760 26240 7772
rect 26292 7760 26298 7812
rect 27154 7760 27160 7812
rect 27212 7800 27218 7812
rect 35894 7800 35900 7812
rect 27212 7772 35900 7800
rect 27212 7760 27218 7772
rect 35894 7760 35900 7772
rect 35952 7760 35958 7812
rect 46477 7803 46535 7809
rect 46477 7769 46489 7803
rect 46523 7800 46535 7803
rect 46750 7800 46756 7812
rect 46523 7772 46756 7800
rect 46523 7769 46535 7772
rect 46477 7763 46535 7769
rect 46750 7760 46756 7772
rect 46808 7760 46814 7812
rect 48130 7800 48136 7812
rect 48091 7772 48136 7800
rect 48130 7760 48136 7772
rect 48188 7760 48194 7812
rect 22002 7732 22008 7744
rect 21560 7704 22008 7732
rect 22002 7692 22008 7704
rect 22060 7692 22066 7744
rect 24394 7732 24400 7744
rect 24355 7704 24400 7732
rect 24394 7692 24400 7704
rect 24452 7692 24458 7744
rect 1104 7642 48852 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 48852 7642
rect 1104 7568 48852 7590
rect 18874 7528 18880 7540
rect 18835 7500 18880 7528
rect 18874 7488 18880 7500
rect 18932 7488 18938 7540
rect 19426 7528 19432 7540
rect 19387 7500 19432 7528
rect 19426 7488 19432 7500
rect 19484 7488 19490 7540
rect 20438 7528 20444 7540
rect 19812 7500 20444 7528
rect 18598 7352 18604 7404
rect 18656 7392 18662 7404
rect 19812 7401 19840 7500
rect 20438 7488 20444 7500
rect 20496 7488 20502 7540
rect 21818 7488 21824 7540
rect 21876 7528 21882 7540
rect 23566 7528 23572 7540
rect 21876 7500 23572 7528
rect 21876 7488 21882 7500
rect 23566 7488 23572 7500
rect 23624 7528 23630 7540
rect 24121 7531 24179 7537
rect 24121 7528 24133 7531
rect 23624 7500 24133 7528
rect 23624 7488 23630 7500
rect 24121 7497 24133 7500
rect 24167 7497 24179 7531
rect 24121 7491 24179 7497
rect 31202 7488 31208 7540
rect 31260 7528 31266 7540
rect 46750 7528 46756 7540
rect 31260 7500 45554 7528
rect 46711 7500 46756 7528
rect 31260 7488 31266 7500
rect 21910 7460 21916 7472
rect 19904 7432 21916 7460
rect 19904 7401 19932 7432
rect 21910 7420 21916 7432
rect 21968 7420 21974 7472
rect 23008 7463 23066 7469
rect 23008 7429 23020 7463
rect 23054 7460 23066 7463
rect 24394 7460 24400 7472
rect 23054 7432 24400 7460
rect 23054 7429 23066 7432
rect 23008 7423 23066 7429
rect 24394 7420 24400 7432
rect 24452 7420 24458 7472
rect 36633 7463 36691 7469
rect 36633 7429 36645 7463
rect 36679 7460 36691 7463
rect 37461 7463 37519 7469
rect 37461 7460 37473 7463
rect 36679 7432 37473 7460
rect 36679 7429 36691 7432
rect 36633 7423 36691 7429
rect 37461 7429 37473 7432
rect 37507 7429 37519 7463
rect 37461 7423 37519 7429
rect 18785 7395 18843 7401
rect 18785 7392 18797 7395
rect 18656 7364 18797 7392
rect 18656 7352 18662 7364
rect 18785 7361 18797 7364
rect 18831 7361 18843 7395
rect 18785 7355 18843 7361
rect 19705 7395 19763 7401
rect 19705 7361 19717 7395
rect 19751 7361 19763 7395
rect 19705 7355 19763 7361
rect 19797 7395 19855 7401
rect 19797 7361 19809 7395
rect 19843 7361 19855 7395
rect 19797 7355 19855 7361
rect 19889 7395 19947 7401
rect 19889 7361 19901 7395
rect 19935 7361 19947 7395
rect 19889 7355 19947 7361
rect 19720 7324 19748 7355
rect 19978 7352 19984 7404
rect 20036 7392 20042 7404
rect 20073 7395 20131 7401
rect 20073 7392 20085 7395
rect 20036 7364 20085 7392
rect 20036 7352 20042 7364
rect 20073 7361 20085 7364
rect 20119 7361 20131 7395
rect 20073 7355 20131 7361
rect 22002 7352 22008 7404
rect 22060 7392 22066 7404
rect 22741 7395 22799 7401
rect 22741 7392 22753 7395
rect 22060 7364 22753 7392
rect 22060 7352 22066 7364
rect 22741 7361 22753 7364
rect 22787 7361 22799 7395
rect 22741 7355 22799 7361
rect 36541 7395 36599 7401
rect 36541 7361 36553 7395
rect 36587 7361 36599 7395
rect 37274 7392 37280 7404
rect 37235 7364 37280 7392
rect 36541 7355 36599 7361
rect 22186 7324 22192 7336
rect 19720 7296 22192 7324
rect 22186 7284 22192 7296
rect 22244 7284 22250 7336
rect 36556 7324 36584 7355
rect 37274 7352 37280 7364
rect 37332 7352 37338 7404
rect 45526 7392 45554 7500
rect 46750 7488 46756 7500
rect 46808 7488 46814 7540
rect 46290 7420 46296 7472
rect 46348 7460 46354 7472
rect 46348 7432 47808 7460
rect 46348 7420 46354 7432
rect 45646 7392 45652 7404
rect 45526 7364 45652 7392
rect 45646 7352 45652 7364
rect 45704 7392 45710 7404
rect 47780 7401 47808 7432
rect 46661 7395 46719 7401
rect 46661 7392 46673 7395
rect 45704 7364 46673 7392
rect 45704 7352 45710 7364
rect 46661 7361 46673 7364
rect 46707 7361 46719 7395
rect 46661 7355 46719 7361
rect 47765 7395 47823 7401
rect 47765 7361 47777 7395
rect 47811 7361 47823 7395
rect 47765 7355 47823 7361
rect 38010 7324 38016 7336
rect 36556 7296 37412 7324
rect 37971 7296 38016 7324
rect 37384 7268 37412 7296
rect 38010 7284 38016 7296
rect 38068 7284 38074 7336
rect 37366 7216 37372 7268
rect 37424 7216 37430 7268
rect 2038 7188 2044 7200
rect 1999 7160 2044 7188
rect 2038 7148 2044 7160
rect 2096 7148 2102 7200
rect 1104 7098 48852 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 48852 7098
rect 1104 7024 48852 7046
rect 19306 6956 28994 6984
rect 1397 6851 1455 6857
rect 1397 6817 1409 6851
rect 1443 6848 1455 6851
rect 2038 6848 2044 6860
rect 1443 6820 2044 6848
rect 1443 6817 1455 6820
rect 1397 6811 1455 6817
rect 2038 6808 2044 6820
rect 2096 6808 2102 6860
rect 2774 6808 2780 6860
rect 2832 6848 2838 6860
rect 2832 6820 2877 6848
rect 2832 6808 2838 6820
rect 1581 6715 1639 6721
rect 1581 6681 1593 6715
rect 1627 6712 1639 6715
rect 2222 6712 2228 6724
rect 1627 6684 2228 6712
rect 1627 6681 1639 6684
rect 1581 6675 1639 6681
rect 2222 6672 2228 6684
rect 2280 6672 2286 6724
rect 18966 6672 18972 6724
rect 19024 6712 19030 6724
rect 19306 6712 19334 6956
rect 23198 6916 23204 6928
rect 23115 6888 23204 6916
rect 22738 6740 22744 6792
rect 22796 6780 22802 6792
rect 23115 6789 23143 6888
rect 23198 6876 23204 6888
rect 23256 6876 23262 6928
rect 28966 6848 28994 6956
rect 45833 6851 45891 6857
rect 45833 6848 45845 6851
rect 28966 6820 45845 6848
rect 45833 6817 45845 6820
rect 45879 6817 45891 6851
rect 45833 6811 45891 6817
rect 22879 6783 22937 6789
rect 22879 6780 22891 6783
rect 22796 6752 22891 6780
rect 22796 6740 22802 6752
rect 22879 6749 22891 6752
rect 22925 6749 22937 6783
rect 22879 6743 22937 6749
rect 22998 6783 23056 6789
rect 22998 6749 23010 6783
rect 23044 6749 23056 6783
rect 22998 6743 23056 6749
rect 23098 6783 23156 6789
rect 23098 6749 23110 6783
rect 23144 6749 23156 6783
rect 23098 6743 23156 6749
rect 19024 6684 19334 6712
rect 23013 6712 23041 6743
rect 23290 6740 23296 6792
rect 23348 6780 23354 6792
rect 23348 6752 23393 6780
rect 23348 6740 23354 6752
rect 23842 6712 23848 6724
rect 23013 6684 23848 6712
rect 19024 6672 19030 6684
rect 23842 6672 23848 6684
rect 23900 6672 23906 6724
rect 46014 6712 46020 6724
rect 45975 6684 46020 6712
rect 46014 6672 46020 6684
rect 46072 6672 46078 6724
rect 47670 6712 47676 6724
rect 47631 6684 47676 6712
rect 47670 6672 47676 6684
rect 47728 6672 47734 6724
rect 22649 6647 22707 6653
rect 22649 6613 22661 6647
rect 22695 6644 22707 6647
rect 23106 6644 23112 6656
rect 22695 6616 23112 6644
rect 22695 6613 22707 6616
rect 22649 6607 22707 6613
rect 23106 6604 23112 6616
rect 23164 6604 23170 6656
rect 1104 6554 48852 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 48852 6554
rect 1104 6480 48852 6502
rect 2222 6440 2228 6452
rect 2183 6412 2228 6440
rect 2222 6400 2228 6412
rect 2280 6400 2286 6452
rect 45925 6443 45983 6449
rect 45925 6409 45937 6443
rect 45971 6440 45983 6443
rect 46014 6440 46020 6452
rect 45971 6412 46020 6440
rect 45971 6409 45983 6412
rect 45925 6403 45983 6409
rect 46014 6400 46020 6412
rect 46072 6400 46078 6452
rect 1486 6264 1492 6316
rect 1544 6304 1550 6316
rect 2133 6307 2191 6313
rect 2133 6304 2145 6307
rect 1544 6276 2145 6304
rect 1544 6264 1550 6276
rect 2133 6273 2145 6276
rect 2179 6273 2191 6307
rect 45830 6304 45836 6316
rect 45791 6276 45836 6304
rect 2133 6267 2191 6273
rect 45830 6264 45836 6276
rect 45888 6264 45894 6316
rect 9122 6128 9128 6180
rect 9180 6168 9186 6180
rect 26050 6168 26056 6180
rect 9180 6140 26056 6168
rect 9180 6128 9186 6140
rect 26050 6128 26056 6140
rect 26108 6128 26114 6180
rect 46290 6060 46296 6112
rect 46348 6100 46354 6112
rect 47765 6103 47823 6109
rect 47765 6100 47777 6103
rect 46348 6072 47777 6100
rect 46348 6060 46354 6072
rect 47765 6069 47777 6072
rect 47811 6069 47823 6103
rect 47765 6063 47823 6069
rect 1104 6010 48852 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 48852 6010
rect 1104 5936 48852 5958
rect 24670 5896 24676 5908
rect 24631 5868 24676 5896
rect 24670 5856 24676 5868
rect 24728 5896 24734 5908
rect 25041 5899 25099 5905
rect 25041 5896 25053 5899
rect 24728 5868 25053 5896
rect 24728 5856 24734 5868
rect 25041 5865 25053 5868
rect 25087 5865 25099 5899
rect 25498 5896 25504 5908
rect 25459 5868 25504 5896
rect 25041 5859 25099 5865
rect 25498 5856 25504 5868
rect 25556 5856 25562 5908
rect 46290 5760 46296 5772
rect 46251 5732 46296 5760
rect 46290 5720 46296 5732
rect 46348 5720 46354 5772
rect 1762 5692 1768 5704
rect 1723 5664 1768 5692
rect 1762 5652 1768 5664
rect 1820 5652 1826 5704
rect 2225 5695 2283 5701
rect 2225 5661 2237 5695
rect 2271 5692 2283 5695
rect 2314 5692 2320 5704
rect 2271 5664 2320 5692
rect 2271 5661 2283 5664
rect 2225 5655 2283 5661
rect 2314 5652 2320 5664
rect 2372 5652 2378 5704
rect 2961 5695 3019 5701
rect 2961 5661 2973 5695
rect 3007 5692 3019 5695
rect 20162 5692 20168 5704
rect 3007 5664 20168 5692
rect 3007 5661 3019 5664
rect 2961 5655 3019 5661
rect 20162 5652 20168 5664
rect 20220 5652 20226 5704
rect 25222 5692 25228 5704
rect 25183 5664 25228 5692
rect 25222 5652 25228 5664
rect 25280 5652 25286 5704
rect 25317 5695 25375 5701
rect 25317 5661 25329 5695
rect 25363 5692 25375 5695
rect 25866 5692 25872 5704
rect 25363 5664 25872 5692
rect 25363 5661 25375 5664
rect 25317 5655 25375 5661
rect 25866 5652 25872 5664
rect 25924 5652 25930 5704
rect 25041 5627 25099 5633
rect 25041 5593 25053 5627
rect 25087 5624 25099 5627
rect 34514 5624 34520 5636
rect 25087 5596 34520 5624
rect 25087 5593 25099 5596
rect 25041 5587 25099 5593
rect 34514 5584 34520 5596
rect 34572 5584 34578 5636
rect 46477 5627 46535 5633
rect 46477 5593 46489 5627
rect 46523 5624 46535 5627
rect 46934 5624 46940 5636
rect 46523 5596 46940 5624
rect 46523 5593 46535 5596
rect 46477 5587 46535 5593
rect 46934 5584 46940 5596
rect 46992 5584 46998 5636
rect 48130 5624 48136 5636
rect 48091 5596 48136 5624
rect 48130 5584 48136 5596
rect 48188 5584 48194 5636
rect 1578 5516 1584 5568
rect 1636 5556 1642 5568
rect 2317 5559 2375 5565
rect 2317 5556 2329 5559
rect 1636 5528 2329 5556
rect 1636 5516 1642 5528
rect 2317 5525 2329 5528
rect 2363 5525 2375 5559
rect 3050 5556 3056 5568
rect 3011 5528 3056 5556
rect 2317 5519 2375 5525
rect 3050 5516 3056 5528
rect 3108 5516 3114 5568
rect 39114 5516 39120 5568
rect 39172 5556 39178 5568
rect 47026 5556 47032 5568
rect 39172 5528 47032 5556
rect 39172 5516 39178 5528
rect 47026 5516 47032 5528
rect 47084 5516 47090 5568
rect 1104 5466 48852 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 48852 5466
rect 1104 5392 48852 5414
rect 46934 5352 46940 5364
rect 46895 5324 46940 5352
rect 46934 5312 46940 5324
rect 46992 5312 46998 5364
rect 2317 5287 2375 5293
rect 2317 5253 2329 5287
rect 2363 5284 2375 5287
rect 3050 5284 3056 5296
rect 2363 5256 3056 5284
rect 2363 5253 2375 5256
rect 2317 5247 2375 5253
rect 3050 5244 3056 5256
rect 3108 5244 3114 5296
rect 31481 5287 31539 5293
rect 31481 5253 31493 5287
rect 31527 5284 31539 5287
rect 32401 5287 32459 5293
rect 32401 5284 32413 5287
rect 31527 5256 32413 5284
rect 31527 5253 31539 5256
rect 31481 5247 31539 5253
rect 32401 5253 32413 5256
rect 32447 5253 32459 5287
rect 47946 5284 47952 5296
rect 47907 5256 47952 5284
rect 32401 5247 32459 5253
rect 47946 5244 47952 5256
rect 48004 5244 48010 5296
rect 1762 5176 1768 5228
rect 1820 5216 1826 5228
rect 2133 5219 2191 5225
rect 2133 5216 2145 5219
rect 1820 5188 2145 5216
rect 1820 5176 1826 5188
rect 2133 5185 2145 5188
rect 2179 5185 2191 5219
rect 2133 5179 2191 5185
rect 17862 5176 17868 5228
rect 17920 5216 17926 5228
rect 30742 5216 30748 5228
rect 17920 5188 30748 5216
rect 17920 5176 17926 5188
rect 30742 5176 30748 5188
rect 30800 5216 30806 5228
rect 31389 5219 31447 5225
rect 31389 5216 31401 5219
rect 30800 5188 31401 5216
rect 30800 5176 30806 5188
rect 31389 5185 31401 5188
rect 31435 5185 31447 5219
rect 31389 5179 31447 5185
rect 46658 5176 46664 5228
rect 46716 5216 46722 5228
rect 46845 5219 46903 5225
rect 46845 5216 46857 5219
rect 46716 5188 46857 5216
rect 46716 5176 46722 5188
rect 46845 5185 46857 5188
rect 46891 5216 46903 5219
rect 47210 5216 47216 5228
rect 46891 5188 47216 5216
rect 46891 5185 46903 5188
rect 46845 5179 46903 5185
rect 47210 5176 47216 5188
rect 47268 5176 47274 5228
rect 2774 5108 2780 5160
rect 2832 5148 2838 5160
rect 32217 5151 32275 5157
rect 2832 5120 2877 5148
rect 2832 5108 2838 5120
rect 32217 5117 32229 5151
rect 32263 5148 32275 5151
rect 32582 5148 32588 5160
rect 32263 5120 32588 5148
rect 32263 5117 32275 5120
rect 32217 5111 32275 5117
rect 32582 5108 32588 5120
rect 32640 5108 32646 5160
rect 34057 5151 34115 5157
rect 34057 5117 34069 5151
rect 34103 5148 34115 5151
rect 46750 5148 46756 5160
rect 34103 5120 46756 5148
rect 34103 5117 34115 5120
rect 34057 5111 34115 5117
rect 46750 5108 46756 5120
rect 46808 5108 46814 5160
rect 25222 5040 25228 5092
rect 25280 5080 25286 5092
rect 48133 5083 48191 5089
rect 48133 5080 48145 5083
rect 25280 5052 48145 5080
rect 25280 5040 25286 5052
rect 48133 5049 48145 5052
rect 48179 5049 48191 5083
rect 48133 5043 48191 5049
rect 1394 4972 1400 5024
rect 1452 5012 1458 5024
rect 1673 5015 1731 5021
rect 1673 5012 1685 5015
rect 1452 4984 1685 5012
rect 1452 4972 1458 4984
rect 1673 4981 1685 4984
rect 1719 4981 1731 5015
rect 1673 4975 1731 4981
rect 1104 4922 48852 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 48852 4922
rect 1104 4848 48852 4870
rect 2682 4768 2688 4820
rect 2740 4808 2746 4820
rect 17126 4808 17132 4820
rect 2740 4780 17132 4808
rect 2740 4768 2746 4780
rect 17126 4768 17132 4780
rect 17184 4768 17190 4820
rect 18506 4768 18512 4820
rect 18564 4808 18570 4820
rect 32214 4808 32220 4820
rect 18564 4780 32220 4808
rect 18564 4768 18570 4780
rect 32214 4768 32220 4780
rect 32272 4768 32278 4820
rect 32950 4768 32956 4820
rect 33008 4808 33014 4820
rect 46842 4808 46848 4820
rect 33008 4780 46848 4808
rect 33008 4768 33014 4780
rect 46842 4768 46848 4780
rect 46900 4768 46906 4820
rect 1394 4672 1400 4684
rect 1355 4644 1400 4672
rect 1394 4632 1400 4644
rect 1452 4632 1458 4684
rect 1578 4672 1584 4684
rect 1539 4644 1584 4672
rect 1578 4632 1584 4644
rect 1636 4632 1642 4684
rect 2774 4632 2780 4684
rect 2832 4672 2838 4684
rect 2832 4644 2877 4672
rect 2832 4632 2838 4644
rect 45002 4564 45008 4616
rect 45060 4604 45066 4616
rect 45189 4607 45247 4613
rect 45189 4604 45201 4607
rect 45060 4576 45201 4604
rect 45060 4564 45066 4576
rect 45189 4573 45201 4576
rect 45235 4573 45247 4607
rect 45189 4567 45247 4573
rect 45833 4607 45891 4613
rect 45833 4573 45845 4607
rect 45879 4604 45891 4607
rect 46293 4607 46351 4613
rect 46293 4604 46305 4607
rect 45879 4576 46305 4604
rect 45879 4573 45891 4576
rect 45833 4567 45891 4573
rect 46293 4573 46305 4576
rect 46339 4573 46351 4607
rect 46293 4567 46351 4573
rect 46477 4539 46535 4545
rect 46477 4505 46489 4539
rect 46523 4536 46535 4539
rect 46934 4536 46940 4548
rect 46523 4508 46940 4536
rect 46523 4505 46535 4508
rect 46477 4499 46535 4505
rect 46934 4496 46940 4508
rect 46992 4496 46998 4548
rect 48133 4539 48191 4545
rect 48133 4505 48145 4539
rect 48179 4536 48191 4539
rect 48314 4536 48320 4548
rect 48179 4508 48320 4536
rect 48179 4505 48191 4508
rect 48133 4499 48191 4505
rect 48314 4496 48320 4508
rect 48372 4496 48378 4548
rect 3694 4428 3700 4480
rect 3752 4468 3758 4480
rect 8018 4468 8024 4480
rect 3752 4440 8024 4468
rect 3752 4428 3758 4440
rect 8018 4428 8024 4440
rect 8076 4428 8082 4480
rect 1104 4378 48852 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 48852 4378
rect 1104 4304 48852 4326
rect 6656 4168 7696 4196
rect 2038 4128 2044 4140
rect 1999 4100 2044 4128
rect 2038 4088 2044 4100
rect 2096 4088 2102 4140
rect 2685 4131 2743 4137
rect 2685 4097 2697 4131
rect 2731 4097 2743 4131
rect 2685 4091 2743 4097
rect 2700 3992 2728 4091
rect 3786 4088 3792 4140
rect 3844 4128 3850 4140
rect 4893 4131 4951 4137
rect 4893 4128 4905 4131
rect 3844 4100 4905 4128
rect 3844 4088 3850 4100
rect 4893 4097 4905 4100
rect 4939 4128 4951 4131
rect 6656 4128 6684 4168
rect 4939 4100 6684 4128
rect 4939 4097 4951 4100
rect 4893 4091 4951 4097
rect 6730 4088 6736 4140
rect 6788 4128 6794 4140
rect 6788 4100 6833 4128
rect 6788 4088 6794 4100
rect 7374 4088 7380 4140
rect 7432 4128 7438 4140
rect 7469 4131 7527 4137
rect 7469 4128 7481 4131
rect 7432 4100 7481 4128
rect 7432 4088 7438 4100
rect 7469 4097 7481 4100
rect 7515 4097 7527 4131
rect 7668 4128 7696 4168
rect 20070 4156 20076 4208
rect 20128 4196 20134 4208
rect 23566 4196 23572 4208
rect 20128 4168 23572 4196
rect 20128 4156 20134 4168
rect 23566 4156 23572 4168
rect 23624 4156 23630 4208
rect 9950 4128 9956 4140
rect 7668 4100 9956 4128
rect 7469 4091 7527 4097
rect 9950 4088 9956 4100
rect 10008 4088 10014 4140
rect 10318 4088 10324 4140
rect 10376 4128 10382 4140
rect 11330 4128 11336 4140
rect 10376 4100 11336 4128
rect 10376 4088 10382 4100
rect 11330 4088 11336 4100
rect 11388 4088 11394 4140
rect 11885 4131 11943 4137
rect 11885 4128 11897 4131
rect 11440 4100 11897 4128
rect 7742 4020 7748 4072
rect 7800 4060 7806 4072
rect 11440 4060 11468 4100
rect 11885 4097 11897 4100
rect 11931 4097 11943 4131
rect 11885 4091 11943 4097
rect 12621 4131 12679 4137
rect 12621 4097 12633 4131
rect 12667 4128 12679 4131
rect 18414 4128 18420 4140
rect 12667 4100 18420 4128
rect 12667 4097 12679 4100
rect 12621 4091 12679 4097
rect 18414 4088 18420 4100
rect 18472 4088 18478 4140
rect 20622 4128 20628 4140
rect 20456 4100 20628 4128
rect 20456 4060 20484 4100
rect 20622 4088 20628 4100
rect 20680 4088 20686 4140
rect 30742 4128 30748 4140
rect 30703 4100 30748 4128
rect 30742 4088 30748 4100
rect 30800 4088 30806 4140
rect 32125 4131 32183 4137
rect 32125 4128 32137 4131
rect 31726 4100 32137 4128
rect 7800 4032 11468 4060
rect 12406 4032 20484 4060
rect 7800 4020 7806 4032
rect 12406 3992 12434 4032
rect 20530 4020 20536 4072
rect 20588 4060 20594 4072
rect 28810 4060 28816 4072
rect 20588 4032 28816 4060
rect 20588 4020 20594 4032
rect 28810 4020 28816 4032
rect 28868 4020 28874 4072
rect 28902 4020 28908 4072
rect 28960 4060 28966 4072
rect 31726 4060 31754 4100
rect 32125 4097 32137 4100
rect 32171 4097 32183 4131
rect 32125 4091 32183 4097
rect 36173 4131 36231 4137
rect 36173 4097 36185 4131
rect 36219 4128 36231 4131
rect 37918 4128 37924 4140
rect 36219 4100 37924 4128
rect 36219 4097 36231 4100
rect 36173 4091 36231 4097
rect 37918 4088 37924 4100
rect 37976 4088 37982 4140
rect 38013 4131 38071 4137
rect 38013 4097 38025 4131
rect 38059 4097 38071 4131
rect 41690 4128 41696 4140
rect 41651 4100 41696 4128
rect 38013 4091 38071 4097
rect 28960 4032 31754 4060
rect 28960 4020 28966 4032
rect 35434 4020 35440 4072
rect 35492 4060 35498 4072
rect 37366 4060 37372 4072
rect 35492 4032 37372 4060
rect 35492 4020 35498 4032
rect 37366 4020 37372 4032
rect 37424 4020 37430 4072
rect 37458 4020 37464 4072
rect 37516 4060 37522 4072
rect 38028 4060 38056 4091
rect 41690 4088 41696 4100
rect 41748 4088 41754 4140
rect 45830 4128 45836 4140
rect 45791 4100 45836 4128
rect 45830 4088 45836 4100
rect 45888 4088 45894 4140
rect 45922 4088 45928 4140
rect 45980 4128 45986 4140
rect 46845 4131 46903 4137
rect 46845 4128 46857 4131
rect 45980 4100 46857 4128
rect 45980 4088 45986 4100
rect 46845 4097 46857 4100
rect 46891 4097 46903 4131
rect 46845 4091 46903 4097
rect 46934 4088 46940 4140
rect 46992 4128 46998 4140
rect 47857 4131 47915 4137
rect 46992 4100 47037 4128
rect 46992 4088 46998 4100
rect 47857 4097 47869 4131
rect 47903 4097 47915 4131
rect 47857 4091 47915 4097
rect 38746 4060 38752 4072
rect 37516 4032 38056 4060
rect 38707 4032 38752 4060
rect 37516 4020 37522 4032
rect 38746 4020 38752 4032
rect 38804 4020 38810 4072
rect 38933 4063 38991 4069
rect 38933 4029 38945 4063
rect 38979 4029 38991 4063
rect 39758 4060 39764 4072
rect 39719 4032 39764 4060
rect 38933 4023 38991 4029
rect 2700 3964 9674 3992
rect 1578 3924 1584 3936
rect 1539 3896 1584 3924
rect 1578 3884 1584 3896
rect 1636 3884 1642 3936
rect 1670 3884 1676 3936
rect 1728 3924 1734 3936
rect 2133 3927 2191 3933
rect 2133 3924 2145 3927
rect 1728 3896 2145 3924
rect 1728 3884 1734 3896
rect 2133 3893 2145 3896
rect 2179 3893 2191 3927
rect 2133 3887 2191 3893
rect 2777 3927 2835 3933
rect 2777 3893 2789 3927
rect 2823 3924 2835 3927
rect 2866 3924 2872 3936
rect 2823 3896 2872 3924
rect 2823 3893 2835 3896
rect 2777 3887 2835 3893
rect 2866 3884 2872 3896
rect 2924 3884 2930 3936
rect 3510 3924 3516 3936
rect 3471 3896 3516 3924
rect 3510 3884 3516 3896
rect 3568 3884 3574 3936
rect 4433 3927 4491 3933
rect 4433 3893 4445 3927
rect 4479 3924 4491 3927
rect 4614 3924 4620 3936
rect 4479 3896 4620 3924
rect 4479 3893 4491 3896
rect 4433 3887 4491 3893
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 4982 3924 4988 3936
rect 4943 3896 4988 3924
rect 4982 3884 4988 3896
rect 5040 3884 5046 3936
rect 6546 3884 6552 3936
rect 6604 3924 6610 3936
rect 6825 3927 6883 3933
rect 6825 3924 6837 3927
rect 6604 3896 6837 3924
rect 6604 3884 6610 3896
rect 6825 3893 6837 3896
rect 6871 3893 6883 3927
rect 7558 3924 7564 3936
rect 7519 3896 7564 3924
rect 6825 3887 6883 3893
rect 7558 3884 7564 3896
rect 7616 3884 7622 3936
rect 9646 3924 9674 3964
rect 11532 3964 12434 3992
rect 11532 3924 11560 3964
rect 17494 3952 17500 4004
rect 17552 3992 17558 4004
rect 32030 3992 32036 4004
rect 17552 3964 32036 3992
rect 17552 3952 17558 3964
rect 32030 3952 32036 3964
rect 32088 3952 32094 4004
rect 32122 3952 32128 4004
rect 32180 3992 32186 4004
rect 32953 3995 33011 4001
rect 32953 3992 32965 3995
rect 32180 3964 32965 3992
rect 32180 3952 32186 3964
rect 32953 3961 32965 3964
rect 32999 3961 33011 3995
rect 32953 3955 33011 3961
rect 36170 3952 36176 4004
rect 36228 3992 36234 4004
rect 38105 3995 38163 4001
rect 36228 3964 36676 3992
rect 36228 3952 36234 3964
rect 9646 3896 11560 3924
rect 11698 3884 11704 3936
rect 11756 3924 11762 3936
rect 11977 3927 12035 3933
rect 11977 3924 11989 3927
rect 11756 3896 11989 3924
rect 11756 3884 11762 3896
rect 11977 3893 11989 3896
rect 12023 3893 12035 3927
rect 11977 3887 12035 3893
rect 12158 3884 12164 3936
rect 12216 3924 12222 3936
rect 12713 3927 12771 3933
rect 12713 3924 12725 3927
rect 12216 3896 12725 3924
rect 12216 3884 12222 3896
rect 12713 3893 12725 3896
rect 12759 3893 12771 3927
rect 12713 3887 12771 3893
rect 14182 3884 14188 3936
rect 14240 3924 14246 3936
rect 19334 3924 19340 3936
rect 14240 3896 19340 3924
rect 14240 3884 14246 3896
rect 19334 3884 19340 3896
rect 19392 3884 19398 3936
rect 19978 3884 19984 3936
rect 20036 3924 20042 3936
rect 20165 3927 20223 3933
rect 20165 3924 20177 3927
rect 20036 3896 20177 3924
rect 20036 3884 20042 3896
rect 20165 3893 20177 3896
rect 20211 3893 20223 3927
rect 29546 3924 29552 3936
rect 29507 3896 29552 3924
rect 20165 3887 20223 3893
rect 29546 3884 29552 3896
rect 29604 3884 29610 3936
rect 29730 3884 29736 3936
rect 29788 3924 29794 3936
rect 30193 3927 30251 3933
rect 30193 3924 30205 3927
rect 29788 3896 30205 3924
rect 29788 3884 29794 3896
rect 30193 3893 30205 3896
rect 30239 3893 30251 3927
rect 30193 3887 30251 3893
rect 30837 3927 30895 3933
rect 30837 3893 30849 3927
rect 30883 3924 30895 3927
rect 31294 3924 31300 3936
rect 30883 3896 31300 3924
rect 30883 3893 30895 3896
rect 30837 3887 30895 3893
rect 31294 3884 31300 3896
rect 31352 3884 31358 3936
rect 32217 3927 32275 3933
rect 32217 3893 32229 3927
rect 32263 3924 32275 3927
rect 32306 3924 32312 3936
rect 32263 3896 32312 3924
rect 32263 3893 32275 3896
rect 32217 3887 32275 3893
rect 32306 3884 32312 3896
rect 32364 3884 32370 3936
rect 36265 3927 36323 3933
rect 36265 3893 36277 3927
rect 36311 3924 36323 3927
rect 36538 3924 36544 3936
rect 36311 3896 36544 3924
rect 36311 3893 36323 3896
rect 36265 3887 36323 3893
rect 36538 3884 36544 3896
rect 36596 3884 36602 3936
rect 36648 3924 36676 3964
rect 38105 3961 38117 3995
rect 38151 3992 38163 3995
rect 38948 3992 38976 4023
rect 39758 4020 39764 4032
rect 39816 4020 39822 4072
rect 42426 4060 42432 4072
rect 42387 4032 42432 4060
rect 42426 4020 42432 4032
rect 42484 4020 42490 4072
rect 42613 4063 42671 4069
rect 42613 4029 42625 4063
rect 42659 4029 42671 4063
rect 42613 4023 42671 4029
rect 41785 3995 41843 4001
rect 38151 3964 38976 3992
rect 39040 3964 41644 3992
rect 38151 3961 38163 3964
rect 38105 3955 38163 3961
rect 39040 3924 39068 3964
rect 36648 3896 39068 3924
rect 41233 3927 41291 3933
rect 41233 3893 41245 3927
rect 41279 3924 41291 3927
rect 41506 3924 41512 3936
rect 41279 3896 41512 3924
rect 41279 3893 41291 3896
rect 41233 3887 41291 3893
rect 41506 3884 41512 3896
rect 41564 3884 41570 3936
rect 41616 3924 41644 3964
rect 41785 3961 41797 3995
rect 41831 3992 41843 3995
rect 42628 3992 42656 4023
rect 42702 4020 42708 4072
rect 42760 4060 42766 4072
rect 42889 4063 42947 4069
rect 42889 4060 42901 4063
rect 42760 4032 42901 4060
rect 42760 4020 42766 4032
rect 42889 4029 42901 4032
rect 42935 4029 42947 4063
rect 42889 4023 42947 4029
rect 46750 4020 46756 4072
rect 46808 4060 46814 4072
rect 47872 4060 47900 4091
rect 46808 4032 47900 4060
rect 46808 4020 46814 4032
rect 47578 3992 47584 4004
rect 41831 3964 42656 3992
rect 42720 3964 47584 3992
rect 41831 3961 41843 3964
rect 41785 3955 41843 3961
rect 42720 3924 42748 3964
rect 47578 3952 47584 3964
rect 47636 3952 47642 4004
rect 45370 3924 45376 3936
rect 41616 3896 42748 3924
rect 45331 3896 45376 3924
rect 45370 3884 45376 3896
rect 45428 3884 45434 3936
rect 45925 3927 45983 3933
rect 45925 3893 45937 3927
rect 45971 3924 45983 3927
rect 46198 3924 46204 3936
rect 45971 3896 46204 3924
rect 45971 3893 45983 3896
rect 45925 3887 45983 3893
rect 46198 3884 46204 3896
rect 46256 3884 46262 3936
rect 48038 3924 48044 3936
rect 47999 3896 48044 3924
rect 48038 3884 48044 3896
rect 48096 3884 48102 3936
rect 1104 3834 48852 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 48852 3834
rect 1104 3760 48852 3782
rect 1946 3680 1952 3732
rect 2004 3720 2010 3732
rect 6270 3720 6276 3732
rect 2004 3692 6276 3720
rect 2004 3680 2010 3692
rect 6270 3680 6276 3692
rect 6328 3680 6334 3732
rect 6730 3680 6736 3732
rect 6788 3720 6794 3732
rect 10502 3720 10508 3732
rect 6788 3692 10508 3720
rect 6788 3680 6794 3692
rect 10502 3680 10508 3692
rect 10560 3720 10566 3732
rect 20346 3720 20352 3732
rect 10560 3692 20352 3720
rect 10560 3680 10566 3692
rect 20346 3680 20352 3692
rect 20404 3680 20410 3732
rect 20806 3680 20812 3732
rect 20864 3720 20870 3732
rect 20864 3692 36308 3720
rect 20864 3680 20870 3692
rect 3510 3652 3516 3664
rect 1412 3624 3516 3652
rect 1412 3593 1440 3624
rect 3510 3612 3516 3624
rect 3568 3612 3574 3664
rect 3878 3612 3884 3664
rect 3936 3652 3942 3664
rect 13078 3652 13084 3664
rect 3936 3624 13084 3652
rect 3936 3612 3942 3624
rect 13078 3612 13084 3624
rect 13136 3612 13142 3664
rect 19426 3652 19432 3664
rect 13464 3624 19432 3652
rect 1397 3587 1455 3593
rect 1397 3553 1409 3587
rect 1443 3553 1455 3587
rect 1397 3547 1455 3553
rect 1581 3587 1639 3593
rect 1581 3553 1593 3587
rect 1627 3584 1639 3587
rect 1670 3584 1676 3596
rect 1627 3556 1676 3584
rect 1627 3553 1639 3556
rect 1581 3547 1639 3553
rect 1670 3544 1676 3556
rect 1728 3544 1734 3596
rect 1854 3584 1860 3596
rect 1815 3556 1860 3584
rect 1854 3544 1860 3556
rect 1912 3544 1918 3596
rect 4433 3587 4491 3593
rect 4433 3553 4445 3587
rect 4479 3584 4491 3587
rect 4614 3584 4620 3596
rect 4479 3556 4620 3584
rect 4479 3553 4491 3556
rect 4433 3547 4491 3553
rect 4614 3544 4620 3556
rect 4672 3544 4678 3596
rect 5166 3584 5172 3596
rect 5127 3556 5172 3584
rect 5166 3544 5172 3556
rect 5224 3544 5230 3596
rect 7374 3544 7380 3596
rect 7432 3584 7438 3596
rect 9950 3584 9956 3596
rect 7432 3556 9956 3584
rect 7432 3544 7438 3556
rect 9950 3544 9956 3556
rect 10008 3544 10014 3596
rect 11606 3544 11612 3596
rect 11664 3584 11670 3596
rect 13354 3584 13360 3596
rect 11664 3556 13360 3584
rect 11664 3544 11670 3556
rect 13354 3544 13360 3556
rect 13412 3544 13418 3596
rect 3786 3516 3792 3528
rect 3747 3488 3792 3516
rect 3786 3476 3792 3488
rect 3844 3476 3850 3528
rect 6638 3476 6644 3528
rect 6696 3516 6702 3528
rect 8113 3519 8171 3525
rect 8113 3516 8125 3519
rect 6696 3488 8125 3516
rect 6696 3476 6702 3488
rect 8113 3485 8125 3488
rect 8159 3485 8171 3519
rect 11790 3516 11796 3528
rect 11751 3488 11796 3516
rect 8113 3479 8171 3485
rect 11790 3476 11796 3488
rect 11848 3476 11854 3528
rect 11974 3476 11980 3528
rect 12032 3516 12038 3528
rect 12437 3519 12495 3525
rect 12437 3516 12449 3519
rect 12032 3488 12449 3516
rect 12032 3476 12038 3488
rect 12437 3485 12449 3488
rect 12483 3485 12495 3519
rect 12437 3479 12495 3485
rect 12618 3476 12624 3528
rect 12676 3516 12682 3528
rect 13464 3516 13492 3624
rect 19426 3612 19432 3624
rect 19484 3612 19490 3664
rect 27982 3612 27988 3664
rect 28040 3652 28046 3664
rect 36170 3652 36176 3664
rect 28040 3624 36176 3652
rect 28040 3612 28046 3624
rect 36170 3612 36176 3624
rect 36228 3612 36234 3664
rect 36280 3652 36308 3692
rect 38746 3680 38752 3732
rect 38804 3720 38810 3732
rect 38933 3723 38991 3729
rect 38933 3720 38945 3723
rect 38804 3692 38945 3720
rect 38804 3680 38810 3692
rect 38933 3689 38945 3692
rect 38979 3689 38991 3723
rect 38933 3683 38991 3689
rect 41690 3680 41696 3732
rect 41748 3720 41754 3732
rect 47118 3720 47124 3732
rect 41748 3692 47124 3720
rect 41748 3680 41754 3692
rect 47118 3680 47124 3692
rect 47176 3680 47182 3732
rect 38838 3652 38844 3664
rect 36280 3624 38844 3652
rect 38838 3612 38844 3624
rect 38896 3612 38902 3664
rect 45646 3652 45652 3664
rect 44744 3624 45652 3652
rect 17034 3544 17040 3596
rect 17092 3584 17098 3596
rect 17221 3587 17279 3593
rect 17221 3584 17233 3587
rect 17092 3556 17233 3584
rect 17092 3544 17098 3556
rect 17221 3553 17233 3556
rect 17267 3553 17279 3587
rect 19978 3584 19984 3596
rect 19939 3556 19984 3584
rect 17221 3547 17279 3553
rect 19978 3544 19984 3556
rect 20036 3544 20042 3596
rect 20622 3584 20628 3596
rect 20583 3556 20628 3584
rect 20622 3544 20628 3556
rect 20680 3544 20686 3596
rect 27706 3584 27712 3596
rect 23584 3556 27712 3584
rect 23584 3528 23612 3556
rect 12676 3488 13492 3516
rect 12676 3476 12682 3488
rect 14274 3476 14280 3528
rect 14332 3516 14338 3528
rect 14553 3519 14611 3525
rect 14553 3516 14565 3519
rect 14332 3488 14565 3516
rect 14332 3476 14338 3488
rect 14553 3485 14565 3488
rect 14599 3485 14611 3519
rect 14553 3479 14611 3485
rect 15013 3519 15071 3525
rect 15013 3485 15025 3519
rect 15059 3516 15071 3519
rect 17126 3516 17132 3528
rect 15059 3488 17132 3516
rect 15059 3485 15071 3488
rect 15013 3479 15071 3485
rect 17126 3476 17132 3488
rect 17184 3476 17190 3528
rect 17402 3476 17408 3528
rect 17460 3516 17466 3528
rect 17681 3519 17739 3525
rect 17681 3516 17693 3519
rect 17460 3488 17693 3516
rect 17460 3476 17466 3488
rect 17681 3485 17693 3488
rect 17727 3516 17739 3519
rect 18322 3516 18328 3528
rect 17727 3488 18328 3516
rect 17727 3485 17739 3488
rect 17681 3479 17739 3485
rect 18322 3476 18328 3488
rect 18380 3516 18386 3528
rect 19886 3516 19892 3528
rect 18380 3488 19892 3516
rect 18380 3476 18386 3488
rect 19886 3476 19892 3488
rect 19944 3476 19950 3528
rect 23109 3519 23167 3525
rect 23109 3485 23121 3519
rect 23155 3516 23167 3519
rect 23198 3516 23204 3528
rect 23155 3488 23204 3516
rect 23155 3485 23167 3488
rect 23109 3479 23167 3485
rect 23198 3476 23204 3488
rect 23256 3476 23262 3528
rect 23566 3516 23572 3528
rect 23527 3488 23572 3516
rect 23566 3476 23572 3488
rect 23624 3476 23630 3528
rect 25332 3525 25360 3556
rect 27706 3544 27712 3556
rect 27764 3544 27770 3596
rect 31294 3584 31300 3596
rect 31255 3556 31300 3584
rect 31294 3544 31300 3556
rect 31352 3544 31358 3596
rect 31570 3584 31576 3596
rect 31531 3556 31576 3584
rect 31570 3544 31576 3556
rect 31628 3544 31634 3596
rect 36538 3584 36544 3596
rect 36499 3556 36544 3584
rect 36538 3544 36544 3556
rect 36596 3544 36602 3596
rect 36722 3544 36728 3596
rect 36780 3584 36786 3596
rect 36817 3587 36875 3593
rect 36817 3584 36829 3587
rect 36780 3556 36829 3584
rect 36780 3544 36786 3556
rect 36817 3553 36829 3556
rect 36863 3553 36875 3587
rect 36817 3547 36875 3553
rect 38102 3544 38108 3596
rect 38160 3584 38166 3596
rect 39022 3584 39028 3596
rect 38160 3556 39028 3584
rect 38160 3544 38166 3556
rect 39022 3544 39028 3556
rect 39080 3544 39086 3596
rect 41506 3584 41512 3596
rect 39132 3556 40908 3584
rect 41467 3556 41512 3584
rect 25317 3519 25375 3525
rect 25317 3485 25329 3519
rect 25363 3485 25375 3519
rect 25958 3516 25964 3528
rect 25919 3488 25964 3516
rect 25317 3479 25375 3485
rect 25958 3476 25964 3488
rect 26016 3476 26022 3528
rect 27430 3476 27436 3528
rect 27488 3516 27494 3528
rect 27801 3519 27859 3525
rect 27801 3516 27813 3519
rect 27488 3488 27813 3516
rect 27488 3476 27494 3488
rect 27801 3485 27813 3488
rect 27847 3485 27859 3519
rect 27801 3479 27859 3485
rect 27982 3476 27988 3528
rect 28040 3516 28046 3528
rect 28721 3519 28779 3525
rect 28721 3516 28733 3519
rect 28040 3488 28733 3516
rect 28040 3476 28046 3488
rect 28721 3485 28733 3488
rect 28767 3485 28779 3519
rect 28721 3479 28779 3485
rect 28810 3476 28816 3528
rect 28868 3516 28874 3528
rect 29733 3519 29791 3525
rect 29733 3516 29745 3519
rect 28868 3488 29745 3516
rect 28868 3476 28874 3488
rect 29733 3485 29745 3488
rect 29779 3485 29791 3519
rect 29733 3479 29791 3485
rect 30653 3519 30711 3525
rect 30653 3485 30665 3519
rect 30699 3516 30711 3519
rect 31113 3519 31171 3525
rect 31113 3516 31125 3519
rect 30699 3488 31125 3516
rect 30699 3485 30711 3488
rect 30653 3479 30711 3485
rect 31113 3485 31125 3488
rect 31159 3485 31171 3519
rect 36354 3516 36360 3528
rect 36315 3488 36360 3516
rect 31113 3479 31171 3485
rect 36354 3476 36360 3488
rect 36412 3476 36418 3528
rect 38838 3476 38844 3528
rect 38896 3516 38902 3528
rect 39132 3516 39160 3556
rect 39850 3516 39856 3528
rect 38896 3488 39160 3516
rect 39811 3488 39856 3516
rect 38896 3476 38902 3488
rect 39850 3476 39856 3488
rect 39908 3476 39914 3528
rect 40880 3525 40908 3556
rect 41506 3544 41512 3556
rect 41564 3544 41570 3596
rect 41874 3544 41880 3596
rect 41932 3584 41938 3596
rect 41969 3587 42027 3593
rect 41969 3584 41981 3587
rect 41932 3556 41981 3584
rect 41932 3544 41938 3556
rect 41969 3553 41981 3556
rect 42015 3553 42027 3587
rect 41969 3547 42027 3553
rect 40865 3519 40923 3525
rect 40865 3485 40877 3519
rect 40911 3485 40923 3519
rect 40865 3479 40923 3485
rect 43809 3519 43867 3525
rect 43809 3485 43821 3519
rect 43855 3516 43867 3519
rect 44744 3516 44772 3624
rect 45646 3612 45652 3624
rect 45704 3612 45710 3664
rect 45370 3544 45376 3596
rect 45428 3584 45434 3596
rect 46017 3587 46075 3593
rect 46017 3584 46029 3587
rect 45428 3556 46029 3584
rect 45428 3544 45434 3556
rect 46017 3553 46029 3556
rect 46063 3553 46075 3587
rect 46198 3584 46204 3596
rect 46159 3556 46204 3584
rect 46017 3547 46075 3553
rect 46198 3544 46204 3556
rect 46256 3544 46262 3596
rect 46382 3544 46388 3596
rect 46440 3584 46446 3596
rect 46477 3587 46535 3593
rect 46477 3584 46489 3587
rect 46440 3556 46489 3584
rect 46440 3544 46446 3556
rect 46477 3553 46489 3556
rect 46523 3553 46535 3587
rect 46477 3547 46535 3553
rect 43855 3488 44772 3516
rect 45005 3519 45063 3525
rect 43855 3485 43867 3488
rect 43809 3479 43867 3485
rect 45005 3485 45017 3519
rect 45051 3516 45063 3519
rect 45922 3516 45928 3528
rect 45051 3488 45928 3516
rect 45051 3485 45063 3488
rect 45005 3479 45063 3485
rect 2038 3408 2044 3460
rect 2096 3448 2102 3460
rect 4617 3451 4675 3457
rect 2096 3420 4568 3448
rect 2096 3408 2102 3420
rect 3510 3340 3516 3392
rect 3568 3380 3574 3392
rect 3881 3383 3939 3389
rect 3881 3380 3893 3383
rect 3568 3352 3893 3380
rect 3568 3340 3574 3352
rect 3881 3349 3893 3352
rect 3927 3349 3939 3383
rect 4540 3380 4568 3420
rect 4617 3417 4629 3451
rect 4663 3448 4675 3451
rect 4982 3448 4988 3460
rect 4663 3420 4988 3448
rect 4663 3417 4675 3420
rect 4617 3411 4675 3417
rect 4982 3408 4988 3420
rect 5040 3408 5046 3460
rect 7098 3408 7104 3460
rect 7156 3448 7162 3460
rect 7285 3451 7343 3457
rect 7285 3448 7297 3451
rect 7156 3420 7297 3448
rect 7156 3408 7162 3420
rect 7285 3417 7297 3420
rect 7331 3417 7343 3451
rect 7285 3411 7343 3417
rect 7469 3451 7527 3457
rect 7469 3417 7481 3451
rect 7515 3448 7527 3451
rect 20165 3451 20223 3457
rect 7515 3420 17954 3448
rect 7515 3417 7527 3420
rect 7469 3411 7527 3417
rect 11882 3380 11888 3392
rect 4540 3352 11888 3380
rect 3881 3343 3939 3349
rect 11882 3340 11888 3352
rect 11940 3340 11946 3392
rect 14458 3340 14464 3392
rect 14516 3380 14522 3392
rect 15105 3383 15163 3389
rect 15105 3380 15117 3383
rect 14516 3352 15117 3380
rect 14516 3340 14522 3352
rect 15105 3349 15117 3352
rect 15151 3349 15163 3383
rect 15105 3343 15163 3349
rect 17494 3340 17500 3392
rect 17552 3380 17558 3392
rect 17773 3383 17831 3389
rect 17773 3380 17785 3383
rect 17552 3352 17785 3380
rect 17552 3340 17558 3352
rect 17773 3349 17785 3352
rect 17819 3349 17831 3383
rect 17926 3380 17954 3420
rect 20165 3417 20177 3451
rect 20211 3448 20223 3451
rect 20346 3448 20352 3460
rect 20211 3420 20352 3448
rect 20211 3417 20223 3420
rect 20165 3411 20223 3417
rect 20346 3408 20352 3420
rect 20404 3408 20410 3460
rect 25409 3451 25467 3457
rect 25409 3417 25421 3451
rect 25455 3448 25467 3451
rect 26145 3451 26203 3457
rect 26145 3448 26157 3451
rect 25455 3420 26157 3448
rect 25455 3417 25467 3420
rect 25409 3411 25467 3417
rect 26145 3417 26157 3420
rect 26191 3417 26203 3451
rect 26145 3411 26203 3417
rect 26234 3408 26240 3460
rect 26292 3448 26298 3460
rect 40957 3451 41015 3457
rect 26292 3420 40264 3448
rect 26292 3408 26298 3420
rect 23014 3380 23020 3392
rect 17926 3352 23020 3380
rect 17773 3343 17831 3349
rect 23014 3340 23020 3352
rect 23072 3340 23078 3392
rect 23382 3340 23388 3392
rect 23440 3380 23446 3392
rect 23661 3383 23719 3389
rect 23661 3380 23673 3383
rect 23440 3352 23673 3380
rect 23440 3340 23446 3352
rect 23661 3349 23673 3352
rect 23707 3349 23719 3383
rect 23661 3343 23719 3349
rect 26418 3340 26424 3392
rect 26476 3380 26482 3392
rect 27430 3380 27436 3392
rect 26476 3352 27436 3380
rect 26476 3340 26482 3352
rect 27430 3340 27436 3352
rect 27488 3340 27494 3392
rect 28813 3383 28871 3389
rect 28813 3349 28825 3383
rect 28859 3380 28871 3383
rect 29638 3380 29644 3392
rect 28859 3352 29644 3380
rect 28859 3349 28871 3352
rect 28813 3343 28871 3349
rect 29638 3340 29644 3352
rect 29696 3340 29702 3392
rect 29825 3383 29883 3389
rect 29825 3349 29837 3383
rect 29871 3380 29883 3383
rect 29914 3380 29920 3392
rect 29871 3352 29920 3380
rect 29871 3349 29883 3352
rect 29825 3343 29883 3349
rect 29914 3340 29920 3352
rect 29972 3340 29978 3392
rect 39945 3383 40003 3389
rect 39945 3349 39957 3383
rect 39991 3380 40003 3383
rect 40126 3380 40132 3392
rect 39991 3352 40132 3380
rect 39991 3349 40003 3352
rect 39945 3343 40003 3349
rect 40126 3340 40132 3352
rect 40184 3340 40190 3392
rect 40236 3380 40264 3420
rect 40957 3417 40969 3451
rect 41003 3448 41015 3451
rect 41693 3451 41751 3457
rect 41693 3448 41705 3451
rect 41003 3420 41705 3448
rect 41003 3417 41015 3420
rect 40957 3411 41015 3417
rect 41693 3417 41705 3420
rect 41739 3417 41751 3451
rect 45020 3448 45048 3479
rect 45922 3476 45928 3488
rect 45980 3476 45986 3528
rect 41693 3411 41751 3417
rect 43824 3420 45048 3448
rect 43824 3380 43852 3420
rect 40236 3352 43852 3380
rect 43901 3383 43959 3389
rect 43901 3349 43913 3383
rect 43947 3380 43959 3383
rect 44174 3380 44180 3392
rect 43947 3352 44180 3380
rect 43947 3349 43959 3352
rect 43901 3343 43959 3349
rect 44174 3340 44180 3352
rect 44232 3340 44238 3392
rect 45097 3383 45155 3389
rect 45097 3349 45109 3383
rect 45143 3380 45155 3383
rect 45186 3380 45192 3392
rect 45143 3352 45192 3380
rect 45143 3349 45155 3352
rect 45097 3343 45155 3349
rect 45186 3340 45192 3352
rect 45244 3340 45250 3392
rect 1104 3290 48852 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 48852 3290
rect 1104 3216 48852 3238
rect 1946 3176 1952 3188
rect 1907 3148 1952 3176
rect 1946 3136 1952 3148
rect 2004 3136 2010 3188
rect 2590 3136 2596 3188
rect 2648 3176 2654 3188
rect 20346 3176 20352 3188
rect 2648 3148 17632 3176
rect 20307 3148 20352 3176
rect 2648 3136 2654 3148
rect 1857 3111 1915 3117
rect 1857 3077 1869 3111
rect 1903 3108 1915 3111
rect 2774 3108 2780 3120
rect 1903 3080 2780 3108
rect 1903 3077 1915 3080
rect 1857 3071 1915 3077
rect 2774 3068 2780 3080
rect 2832 3068 2838 3120
rect 3510 3108 3516 3120
rect 3471 3080 3516 3108
rect 3510 3068 3516 3080
rect 3568 3068 3574 3120
rect 6825 3111 6883 3117
rect 6825 3077 6837 3111
rect 6871 3108 6883 3111
rect 7558 3108 7564 3120
rect 6871 3080 7564 3108
rect 6871 3077 6883 3080
rect 6825 3071 6883 3077
rect 7558 3068 7564 3080
rect 7616 3068 7622 3120
rect 12158 3108 12164 3120
rect 12119 3080 12164 3108
rect 12158 3068 12164 3080
rect 12216 3068 12222 3120
rect 12250 3068 12256 3120
rect 12308 3108 12314 3120
rect 14182 3108 14188 3120
rect 12308 3080 14188 3108
rect 12308 3068 12314 3080
rect 14182 3068 14188 3080
rect 14240 3068 14246 3120
rect 14458 3108 14464 3120
rect 14419 3080 14464 3108
rect 14458 3068 14464 3080
rect 14516 3068 14522 3120
rect 17494 3108 17500 3120
rect 17455 3080 17500 3108
rect 17494 3068 17500 3080
rect 17552 3068 17558 3120
rect 17604 3108 17632 3148
rect 20346 3136 20352 3148
rect 20404 3136 20410 3188
rect 20438 3136 20444 3188
rect 20496 3176 20502 3188
rect 20496 3148 28304 3176
rect 20496 3136 20502 3148
rect 23382 3108 23388 3120
rect 17604 3080 23060 3108
rect 23343 3080 23388 3108
rect 1946 3000 1952 3052
rect 2004 3040 2010 3052
rect 2501 3043 2559 3049
rect 2501 3040 2513 3043
rect 2004 3012 2513 3040
rect 2004 3000 2010 3012
rect 2501 3009 2513 3012
rect 2547 3009 2559 3043
rect 6638 3040 6644 3052
rect 6599 3012 6644 3040
rect 2501 3003 2559 3009
rect 6638 3000 6644 3012
rect 6696 3000 6702 3052
rect 8386 3000 8392 3052
rect 8444 3040 8450 3052
rect 8941 3043 8999 3049
rect 8941 3040 8953 3043
rect 8444 3012 8953 3040
rect 8444 3000 8450 3012
rect 8941 3009 8953 3012
rect 8987 3009 8999 3043
rect 11974 3040 11980 3052
rect 8941 3003 8999 3009
rect 9048 3012 10088 3040
rect 11935 3012 11980 3040
rect 3326 2972 3332 2984
rect 3287 2944 3332 2972
rect 3326 2932 3332 2944
rect 3384 2932 3390 2984
rect 3789 2975 3847 2981
rect 3789 2941 3801 2975
rect 3835 2941 3847 2975
rect 3789 2935 3847 2941
rect 658 2864 664 2916
rect 716 2904 722 2916
rect 716 2876 3188 2904
rect 716 2864 722 2876
rect 2682 2836 2688 2848
rect 2643 2808 2688 2836
rect 2682 2796 2688 2808
rect 2740 2796 2746 2848
rect 3160 2836 3188 2876
rect 3234 2864 3240 2916
rect 3292 2904 3298 2916
rect 3804 2904 3832 2935
rect 6454 2932 6460 2984
rect 6512 2972 6518 2984
rect 7101 2975 7159 2981
rect 7101 2972 7113 2975
rect 6512 2944 7113 2972
rect 6512 2932 6518 2944
rect 7101 2941 7113 2944
rect 7147 2941 7159 2975
rect 7101 2935 7159 2941
rect 9048 2904 9076 3012
rect 3292 2876 3832 2904
rect 3896 2876 9076 2904
rect 10060 2904 10088 3012
rect 11974 3000 11980 3012
rect 12032 3000 12038 3052
rect 14274 3040 14280 3052
rect 14235 3012 14280 3040
rect 14274 3000 14280 3012
rect 14332 3000 14338 3052
rect 17034 3000 17040 3052
rect 17092 3040 17098 3052
rect 17313 3043 17371 3049
rect 17313 3040 17325 3043
rect 17092 3012 17325 3040
rect 17092 3000 17098 3012
rect 17313 3009 17325 3012
rect 17359 3009 17371 3043
rect 17313 3003 17371 3009
rect 20257 3043 20315 3049
rect 20257 3009 20269 3043
rect 20303 3040 20315 3043
rect 20530 3040 20536 3052
rect 20303 3012 20536 3040
rect 20303 3009 20315 3012
rect 20257 3003 20315 3009
rect 20530 3000 20536 3012
rect 20588 3000 20594 3052
rect 10962 2932 10968 2984
rect 11020 2972 11026 2984
rect 12250 2972 12256 2984
rect 11020 2944 12256 2972
rect 11020 2932 11026 2944
rect 12250 2932 12256 2944
rect 12308 2932 12314 2984
rect 12710 2972 12716 2984
rect 12360 2944 12716 2972
rect 12360 2904 12388 2944
rect 12710 2932 12716 2944
rect 12768 2932 12774 2984
rect 12894 2972 12900 2984
rect 12855 2944 12900 2972
rect 12894 2932 12900 2944
rect 12952 2932 12958 2984
rect 15470 2972 15476 2984
rect 15431 2944 15476 2972
rect 15470 2932 15476 2944
rect 15528 2932 15534 2984
rect 18046 2972 18052 2984
rect 18007 2944 18052 2972
rect 18046 2932 18052 2944
rect 18104 2932 18110 2984
rect 10060 2876 12388 2904
rect 3292 2864 3298 2876
rect 3896 2836 3924 2876
rect 12434 2864 12440 2916
rect 12492 2904 12498 2916
rect 23032 2904 23060 3080
rect 23382 3068 23388 3080
rect 23440 3068 23446 3120
rect 23198 3040 23204 3052
rect 23159 3012 23204 3040
rect 23198 3000 23204 3012
rect 23256 3000 23262 3052
rect 25958 3000 25964 3052
rect 26016 3040 26022 3052
rect 26237 3043 26295 3049
rect 26237 3040 26249 3043
rect 26016 3012 26249 3040
rect 26016 3000 26022 3012
rect 26237 3009 26249 3012
rect 26283 3009 26295 3043
rect 26237 3003 26295 3009
rect 23842 2972 23848 2984
rect 23803 2944 23848 2972
rect 23842 2932 23848 2944
rect 23900 2932 23906 2984
rect 28166 2972 28172 2984
rect 23952 2944 28172 2972
rect 23952 2904 23980 2944
rect 28166 2932 28172 2944
rect 28224 2932 28230 2984
rect 12492 2876 22094 2904
rect 23032 2876 23980 2904
rect 28276 2904 28304 3148
rect 28718 3136 28724 3188
rect 28776 3176 28782 3188
rect 48038 3176 48044 3188
rect 28776 3148 48044 3176
rect 28776 3136 28782 3148
rect 48038 3136 48044 3148
rect 48096 3136 48102 3188
rect 29914 3108 29920 3120
rect 29875 3080 29920 3108
rect 29914 3068 29920 3080
rect 29972 3068 29978 3120
rect 32306 3108 32312 3120
rect 32267 3080 32312 3108
rect 32306 3068 32312 3080
rect 32364 3068 32370 3120
rect 40126 3108 40132 3120
rect 40087 3080 40132 3108
rect 40126 3068 40132 3080
rect 40184 3068 40190 3120
rect 44174 3108 44180 3120
rect 44135 3080 44180 3108
rect 44174 3068 44180 3080
rect 44232 3068 44238 3120
rect 44358 3068 44364 3120
rect 44416 3108 44422 3120
rect 46658 3108 46664 3120
rect 44416 3080 46664 3108
rect 44416 3068 44422 3080
rect 46658 3068 46664 3080
rect 46716 3068 46722 3120
rect 29730 3040 29736 3052
rect 29691 3012 29736 3040
rect 29730 3000 29736 3012
rect 29788 3000 29794 3052
rect 32122 3040 32128 3052
rect 32083 3012 32128 3040
rect 32122 3000 32128 3012
rect 32180 3000 32186 3052
rect 36354 3000 36360 3052
rect 36412 3040 36418 3052
rect 36541 3043 36599 3049
rect 36541 3040 36553 3043
rect 36412 3012 36553 3040
rect 36412 3000 36418 3012
rect 36541 3009 36553 3012
rect 36587 3009 36599 3043
rect 36541 3003 36599 3009
rect 42426 3000 42432 3052
rect 42484 3040 42490 3052
rect 42613 3043 42671 3049
rect 42613 3040 42625 3043
rect 42484 3012 42625 3040
rect 42484 3000 42490 3012
rect 42613 3009 42625 3012
rect 42659 3009 42671 3043
rect 42613 3003 42671 3009
rect 45738 3000 45744 3052
rect 45796 3040 45802 3052
rect 46385 3043 46443 3049
rect 46385 3040 46397 3043
rect 45796 3012 46397 3040
rect 45796 3000 45802 3012
rect 46385 3009 46397 3012
rect 46431 3009 46443 3043
rect 46566 3040 46572 3052
rect 46527 3012 46572 3040
rect 46385 3003 46443 3009
rect 46566 3000 46572 3012
rect 46624 3000 46630 3052
rect 47857 3043 47915 3049
rect 47857 3009 47869 3043
rect 47903 3040 47915 3043
rect 49602 3040 49608 3052
rect 47903 3012 49608 3040
rect 47903 3009 47915 3012
rect 47857 3003 47915 3009
rect 49602 3000 49608 3012
rect 49660 3000 49666 3052
rect 30282 2972 30288 2984
rect 30243 2944 30288 2972
rect 30282 2932 30288 2944
rect 30340 2932 30346 2984
rect 33502 2972 33508 2984
rect 33463 2944 33508 2972
rect 33502 2932 33508 2944
rect 33560 2932 33566 2984
rect 39942 2972 39948 2984
rect 39903 2944 39948 2972
rect 39942 2932 39948 2944
rect 40000 2932 40006 2984
rect 41138 2972 41144 2984
rect 41099 2944 41144 2972
rect 41138 2932 41144 2944
rect 41196 2932 41202 2984
rect 43993 2975 44051 2981
rect 43993 2941 44005 2975
rect 44039 2972 44051 2975
rect 44266 2972 44272 2984
rect 44039 2944 44272 2972
rect 44039 2941 44051 2944
rect 43993 2935 44051 2941
rect 44266 2932 44272 2944
rect 44324 2932 44330 2984
rect 44450 2972 44456 2984
rect 44411 2944 44456 2972
rect 44450 2932 44456 2944
rect 44508 2932 44514 2984
rect 28276 2876 31754 2904
rect 12492 2864 12498 2876
rect 5810 2836 5816 2848
rect 3160 2808 3924 2836
rect 5771 2808 5816 2836
rect 5810 2796 5816 2808
rect 5868 2796 5874 2848
rect 9122 2836 9128 2848
rect 9083 2808 9128 2836
rect 9122 2796 9128 2808
rect 9180 2796 9186 2848
rect 9950 2796 9956 2848
rect 10008 2836 10014 2848
rect 12618 2836 12624 2848
rect 10008 2808 12624 2836
rect 10008 2796 10014 2808
rect 12618 2796 12624 2808
rect 12676 2796 12682 2848
rect 12710 2796 12716 2848
rect 12768 2836 12774 2848
rect 20438 2836 20444 2848
rect 12768 2808 20444 2836
rect 12768 2796 12774 2808
rect 20438 2796 20444 2808
rect 20496 2796 20502 2848
rect 22066 2836 22094 2876
rect 28902 2836 28908 2848
rect 22066 2808 28908 2836
rect 28902 2796 28908 2808
rect 28960 2796 28966 2848
rect 29638 2796 29644 2848
rect 29696 2836 29702 2848
rect 29822 2836 29828 2848
rect 29696 2808 29828 2836
rect 29696 2796 29702 2808
rect 29822 2796 29828 2808
rect 29880 2796 29886 2848
rect 31726 2836 31754 2876
rect 32030 2864 32036 2916
rect 32088 2904 32094 2916
rect 48041 2907 48099 2913
rect 48041 2904 48053 2907
rect 32088 2876 48053 2904
rect 32088 2864 32094 2876
rect 48041 2873 48053 2876
rect 48087 2873 48099 2907
rect 48041 2867 48099 2873
rect 33042 2836 33048 2848
rect 31726 2808 33048 2836
rect 33042 2796 33048 2808
rect 33100 2796 33106 2848
rect 37918 2796 37924 2848
rect 37976 2836 37982 2848
rect 44358 2836 44364 2848
rect 37976 2808 44364 2836
rect 37976 2796 37982 2808
rect 44358 2796 44364 2808
rect 44416 2796 44422 2848
rect 1104 2746 48852 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 48852 2746
rect 1104 2672 48852 2694
rect 3326 2592 3332 2644
rect 3384 2632 3390 2644
rect 3973 2635 4031 2641
rect 3973 2632 3985 2635
rect 3384 2604 3985 2632
rect 3384 2592 3390 2604
rect 3973 2601 3985 2604
rect 4019 2601 4031 2635
rect 3973 2595 4031 2601
rect 10413 2635 10471 2641
rect 10413 2601 10425 2635
rect 10459 2632 10471 2635
rect 18230 2632 18236 2644
rect 10459 2604 18236 2632
rect 10459 2601 10471 2604
rect 10413 2595 10471 2601
rect 18230 2592 18236 2604
rect 18288 2592 18294 2644
rect 21358 2592 21364 2644
rect 21416 2632 21422 2644
rect 46842 2632 46848 2644
rect 21416 2604 46848 2632
rect 21416 2592 21422 2604
rect 46842 2592 46848 2604
rect 46900 2592 46906 2644
rect 1302 2524 1308 2576
rect 1360 2564 1366 2576
rect 1360 2536 1900 2564
rect 1360 2524 1366 2536
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2496 1455 2499
rect 1578 2496 1584 2508
rect 1443 2468 1584 2496
rect 1443 2465 1455 2468
rect 1397 2459 1455 2465
rect 1578 2456 1584 2468
rect 1636 2456 1642 2508
rect 1872 2505 1900 2536
rect 6178 2524 6184 2576
rect 6236 2564 6242 2576
rect 17770 2564 17776 2576
rect 6236 2536 6960 2564
rect 6236 2524 6242 2536
rect 1857 2499 1915 2505
rect 1857 2465 1869 2499
rect 1903 2465 1915 2499
rect 1857 2459 1915 2465
rect 5810 2456 5816 2508
rect 5868 2496 5874 2508
rect 6365 2499 6423 2505
rect 6365 2496 6377 2499
rect 5868 2468 6377 2496
rect 5868 2456 5874 2468
rect 6365 2465 6377 2468
rect 6411 2465 6423 2499
rect 6546 2496 6552 2508
rect 6507 2468 6552 2496
rect 6365 2459 6423 2465
rect 6546 2456 6552 2468
rect 6604 2456 6610 2508
rect 6932 2505 6960 2536
rect 9232 2536 16574 2564
rect 17731 2536 17776 2564
rect 9232 2505 9260 2536
rect 6917 2499 6975 2505
rect 6917 2465 6929 2499
rect 6963 2465 6975 2499
rect 6917 2459 6975 2465
rect 9217 2499 9275 2505
rect 9217 2465 9229 2499
rect 9263 2465 9275 2499
rect 9217 2459 9275 2465
rect 11517 2499 11575 2505
rect 11517 2465 11529 2499
rect 11563 2496 11575 2499
rect 11790 2496 11796 2508
rect 11563 2468 11796 2496
rect 11563 2465 11575 2468
rect 11517 2459 11575 2465
rect 11790 2456 11796 2468
rect 11848 2456 11854 2508
rect 12250 2496 12256 2508
rect 12211 2468 12256 2496
rect 12250 2456 12256 2468
rect 12308 2456 12314 2508
rect 14734 2496 14740 2508
rect 14695 2468 14740 2496
rect 14734 2456 14740 2468
rect 14792 2456 14798 2508
rect 16546 2496 16574 2536
rect 17770 2524 17776 2536
rect 17828 2524 17834 2576
rect 23385 2567 23443 2573
rect 23385 2533 23397 2567
rect 23431 2564 23443 2567
rect 23658 2564 23664 2576
rect 23431 2536 23664 2564
rect 23431 2533 23443 2536
rect 23385 2527 23443 2533
rect 23658 2524 23664 2536
rect 23716 2524 23722 2576
rect 25866 2564 25872 2576
rect 25827 2536 25872 2564
rect 25866 2524 25872 2536
rect 25924 2524 25930 2576
rect 35069 2567 35127 2573
rect 35069 2564 35081 2567
rect 26206 2536 35081 2564
rect 22738 2496 22744 2508
rect 16546 2468 22744 2496
rect 22738 2456 22744 2468
rect 22796 2456 22802 2508
rect 23750 2456 23756 2508
rect 23808 2496 23814 2508
rect 24857 2499 24915 2505
rect 24857 2496 24869 2499
rect 23808 2468 24869 2496
rect 23808 2456 23814 2468
rect 24857 2465 24869 2468
rect 24903 2465 24915 2499
rect 26206 2496 26234 2536
rect 35069 2533 35081 2536
rect 35115 2533 35127 2567
rect 47949 2567 48007 2573
rect 47949 2564 47961 2567
rect 35069 2527 35127 2533
rect 35176 2536 47961 2564
rect 24857 2459 24915 2465
rect 24964 2468 26234 2496
rect 26436 2468 27200 2496
rect 4522 2388 4528 2440
rect 4580 2428 4586 2440
rect 4617 2431 4675 2437
rect 4617 2428 4629 2431
rect 4580 2400 4629 2428
rect 4580 2388 4586 2400
rect 4617 2397 4629 2400
rect 4663 2397 4675 2431
rect 4617 2391 4675 2397
rect 7742 2388 7748 2440
rect 7800 2428 7806 2440
rect 8941 2431 8999 2437
rect 8941 2428 8953 2431
rect 7800 2400 8953 2428
rect 7800 2388 7806 2400
rect 8941 2397 8953 2400
rect 8987 2397 8999 2431
rect 8941 2391 8999 2397
rect 19978 2388 19984 2440
rect 20036 2428 20042 2440
rect 20073 2431 20131 2437
rect 20073 2428 20085 2431
rect 20036 2400 20085 2428
rect 20036 2388 20042 2400
rect 20073 2397 20085 2400
rect 20119 2397 20131 2431
rect 20073 2391 20131 2397
rect 22554 2388 22560 2440
rect 22612 2428 22618 2440
rect 22649 2431 22707 2437
rect 22649 2428 22661 2431
rect 22612 2400 22661 2428
rect 22612 2388 22618 2400
rect 22649 2397 22661 2400
rect 22695 2397 22707 2431
rect 22649 2391 22707 2397
rect 23198 2388 23204 2440
rect 23256 2428 23262 2440
rect 23569 2431 23627 2437
rect 23569 2428 23581 2431
rect 23256 2400 23581 2428
rect 23256 2388 23262 2400
rect 23569 2397 23581 2400
rect 23615 2397 23627 2431
rect 23569 2391 23627 2397
rect 24486 2388 24492 2440
rect 24544 2428 24550 2440
rect 24581 2431 24639 2437
rect 24581 2428 24593 2431
rect 24544 2400 24593 2428
rect 24544 2388 24550 2400
rect 24581 2397 24593 2400
rect 24627 2397 24639 2431
rect 24581 2391 24639 2397
rect 24670 2388 24676 2440
rect 24728 2428 24734 2440
rect 24964 2428 24992 2468
rect 24728 2400 24992 2428
rect 24728 2388 24734 2400
rect 25130 2388 25136 2440
rect 25188 2428 25194 2440
rect 26053 2431 26111 2437
rect 26053 2428 26065 2431
rect 25188 2400 26065 2428
rect 25188 2388 25194 2400
rect 26053 2397 26065 2400
rect 26099 2397 26111 2431
rect 26053 2391 26111 2397
rect 1581 2363 1639 2369
rect 1581 2329 1593 2363
rect 1627 2360 1639 2363
rect 2866 2360 2872 2372
rect 1627 2332 2872 2360
rect 1627 2329 1639 2332
rect 1581 2323 1639 2329
rect 2866 2320 2872 2332
rect 2924 2320 2930 2372
rect 3418 2320 3424 2372
rect 3476 2360 3482 2372
rect 8662 2360 8668 2372
rect 3476 2332 8668 2360
rect 3476 2320 3482 2332
rect 8662 2320 8668 2332
rect 8720 2320 8726 2372
rect 9674 2320 9680 2372
rect 9732 2360 9738 2372
rect 10321 2363 10379 2369
rect 10321 2360 10333 2363
rect 9732 2332 10333 2360
rect 9732 2320 9738 2332
rect 10321 2329 10333 2332
rect 10367 2329 10379 2363
rect 11698 2360 11704 2372
rect 11659 2332 11704 2360
rect 10321 2323 10379 2329
rect 11698 2320 11704 2332
rect 11756 2320 11762 2372
rect 14182 2320 14188 2372
rect 14240 2360 14246 2372
rect 14553 2363 14611 2369
rect 14553 2360 14565 2363
rect 14240 2332 14565 2360
rect 14240 2320 14246 2332
rect 14553 2329 14565 2332
rect 14599 2329 14611 2363
rect 14553 2323 14611 2329
rect 17402 2320 17408 2372
rect 17460 2360 17466 2372
rect 17589 2363 17647 2369
rect 17589 2360 17601 2363
rect 17460 2332 17601 2360
rect 17460 2320 17466 2332
rect 17589 2329 17601 2332
rect 17635 2329 17647 2363
rect 26436 2360 26464 2468
rect 27062 2428 27068 2440
rect 27023 2400 27068 2428
rect 27062 2388 27068 2400
rect 27120 2388 27126 2440
rect 27172 2428 27200 2468
rect 27338 2456 27344 2508
rect 27396 2496 27402 2508
rect 28077 2499 28135 2505
rect 28077 2496 28089 2499
rect 27396 2468 28089 2496
rect 27396 2456 27402 2468
rect 28077 2465 28089 2468
rect 28123 2465 28135 2499
rect 29546 2496 29552 2508
rect 29507 2468 29552 2496
rect 28077 2459 28135 2465
rect 29546 2456 29552 2468
rect 29604 2456 29610 2508
rect 29730 2496 29736 2508
rect 29691 2468 29736 2496
rect 29730 2456 29736 2468
rect 29788 2456 29794 2508
rect 30926 2496 30932 2508
rect 30887 2468 30932 2496
rect 30926 2456 30932 2468
rect 30984 2456 30990 2508
rect 33870 2456 33876 2508
rect 33928 2496 33934 2508
rect 35176 2496 35204 2536
rect 47949 2533 47961 2536
rect 47995 2533 48007 2567
rect 47949 2527 48007 2533
rect 33928 2468 35204 2496
rect 33928 2456 33934 2468
rect 35894 2456 35900 2508
rect 35952 2496 35958 2508
rect 38749 2499 38807 2505
rect 38749 2496 38761 2499
rect 35952 2468 38761 2496
rect 35952 2456 35958 2468
rect 38749 2465 38761 2468
rect 38795 2465 38807 2499
rect 39942 2496 39948 2508
rect 39903 2468 39948 2496
rect 38749 2459 38807 2465
rect 39942 2456 39948 2468
rect 40000 2456 40006 2508
rect 44266 2496 44272 2508
rect 44227 2468 44272 2496
rect 44266 2456 44272 2468
rect 44324 2456 44330 2508
rect 45002 2496 45008 2508
rect 44963 2468 45008 2496
rect 45002 2456 45008 2468
rect 45060 2456 45066 2508
rect 45186 2496 45192 2508
rect 45147 2468 45192 2496
rect 45186 2456 45192 2468
rect 45244 2456 45250 2508
rect 45370 2456 45376 2508
rect 45428 2496 45434 2508
rect 45557 2499 45615 2505
rect 45557 2496 45569 2499
rect 45428 2468 45569 2496
rect 45428 2456 45434 2468
rect 45557 2465 45569 2468
rect 45603 2465 45615 2499
rect 45557 2459 45615 2465
rect 27172 2400 27384 2428
rect 17589 2323 17647 2329
rect 20272 2332 26464 2360
rect 4798 2292 4804 2304
rect 4759 2264 4804 2292
rect 4798 2252 4804 2264
rect 4856 2252 4862 2304
rect 20272 2301 20300 2332
rect 26510 2320 26516 2372
rect 26568 2360 26574 2372
rect 27154 2360 27160 2372
rect 26568 2332 27160 2360
rect 26568 2320 26574 2332
rect 27154 2320 27160 2332
rect 27212 2320 27218 2372
rect 20257 2295 20315 2301
rect 20257 2261 20269 2295
rect 20303 2261 20315 2295
rect 22830 2292 22836 2304
rect 22791 2264 22836 2292
rect 20257 2255 20315 2261
rect 22830 2252 22836 2264
rect 22888 2252 22894 2304
rect 24026 2252 24032 2304
rect 24084 2292 24090 2304
rect 24670 2292 24676 2304
rect 24084 2264 24676 2292
rect 24084 2252 24090 2264
rect 24670 2252 24676 2264
rect 24728 2252 24734 2304
rect 25314 2252 25320 2304
rect 25372 2292 25378 2304
rect 27249 2295 27307 2301
rect 27249 2292 27261 2295
rect 25372 2264 27261 2292
rect 25372 2252 25378 2264
rect 27249 2261 27261 2264
rect 27295 2261 27307 2295
rect 27356 2292 27384 2400
rect 27706 2388 27712 2440
rect 27764 2428 27770 2440
rect 27801 2431 27859 2437
rect 27801 2428 27813 2431
rect 27764 2400 27813 2428
rect 27764 2388 27770 2400
rect 27801 2397 27813 2400
rect 27847 2397 27859 2431
rect 27801 2391 27859 2397
rect 32858 2388 32864 2440
rect 32916 2428 32922 2440
rect 32953 2431 33011 2437
rect 32953 2428 32965 2431
rect 32916 2400 32965 2428
rect 32916 2388 32922 2400
rect 32953 2397 32965 2400
rect 32999 2397 33011 2431
rect 32953 2391 33011 2397
rect 34790 2388 34796 2440
rect 34848 2428 34854 2440
rect 34885 2431 34943 2437
rect 34885 2428 34897 2431
rect 34848 2400 34897 2428
rect 34848 2388 34854 2400
rect 34885 2397 34897 2400
rect 34931 2397 34943 2431
rect 34885 2391 34943 2397
rect 36078 2388 36084 2440
rect 36136 2428 36142 2440
rect 36357 2431 36415 2437
rect 36357 2428 36369 2431
rect 36136 2400 36369 2428
rect 36136 2388 36142 2400
rect 36357 2397 36369 2400
rect 36403 2397 36415 2431
rect 36357 2391 36415 2397
rect 38473 2431 38531 2437
rect 38473 2397 38485 2431
rect 38519 2428 38531 2431
rect 38654 2428 38660 2440
rect 38519 2400 38660 2428
rect 38519 2397 38531 2400
rect 38473 2391 38531 2397
rect 38654 2388 38660 2400
rect 38712 2388 38718 2440
rect 27522 2320 27528 2372
rect 27580 2360 27586 2372
rect 33965 2363 34023 2369
rect 27580 2332 33180 2360
rect 27580 2320 27586 2332
rect 31386 2292 31392 2304
rect 27356 2264 31392 2292
rect 27249 2255 27307 2261
rect 31386 2252 31392 2264
rect 31444 2252 31450 2304
rect 33152 2301 33180 2332
rect 33965 2329 33977 2363
rect 34011 2360 34023 2363
rect 34146 2360 34152 2372
rect 34011 2332 34152 2360
rect 34011 2329 34023 2332
rect 33965 2323 34023 2329
rect 34146 2320 34152 2332
rect 34204 2320 34210 2372
rect 43162 2320 43168 2372
rect 43220 2360 43226 2372
rect 43349 2363 43407 2369
rect 43349 2360 43361 2363
rect 43220 2332 43361 2360
rect 43220 2320 43226 2332
rect 43349 2329 43361 2332
rect 43395 2329 43407 2363
rect 47762 2360 47768 2372
rect 47723 2332 47768 2360
rect 43349 2323 43407 2329
rect 47762 2320 47768 2332
rect 47820 2320 47826 2372
rect 33137 2295 33195 2301
rect 33137 2261 33149 2295
rect 33183 2261 33195 2295
rect 34054 2292 34060 2304
rect 34015 2264 34060 2292
rect 33137 2255 33195 2261
rect 34054 2252 34060 2264
rect 34112 2252 34118 2304
rect 34514 2252 34520 2304
rect 34572 2292 34578 2304
rect 36173 2295 36231 2301
rect 36173 2292 36185 2295
rect 34572 2264 36185 2292
rect 34572 2252 34578 2264
rect 36173 2261 36185 2264
rect 36219 2261 36231 2295
rect 43438 2292 43444 2304
rect 43399 2264 43444 2292
rect 36173 2255 36231 2261
rect 43438 2252 43444 2264
rect 43496 2252 43502 2304
rect 1104 2202 48852 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 48852 2202
rect 1104 2128 48852 2150
rect 23934 2048 23940 2100
rect 23992 2088 23998 2100
rect 34054 2088 34060 2100
rect 23992 2060 34060 2088
rect 23992 2048 23998 2060
rect 34054 2048 34060 2060
rect 34112 2048 34118 2100
rect 22830 1980 22836 2032
rect 22888 2020 22894 2032
rect 30650 2020 30656 2032
rect 22888 1992 30656 2020
rect 22888 1980 22894 1992
rect 30650 1980 30656 1992
rect 30708 1980 30714 2032
rect 24302 1912 24308 1964
rect 24360 1952 24366 1964
rect 43438 1952 43444 1964
rect 24360 1924 43444 1952
rect 24360 1912 24366 1924
rect 43438 1912 43444 1924
rect 43496 1912 43502 1964
<< via1 >>
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 14188 49240 14240 49292
rect 20444 49376 20496 49428
rect 18052 49240 18104 49292
rect 24216 49308 24268 49360
rect 29092 49308 29144 49360
rect 664 49172 716 49224
rect 3608 49172 3660 49224
rect 4896 49172 4948 49224
rect 6460 49172 6512 49224
rect 7104 49172 7156 49224
rect 10324 49215 10376 49224
rect 10324 49181 10333 49215
rect 10333 49181 10367 49215
rect 10367 49181 10376 49215
rect 10324 49172 10376 49181
rect 11520 49172 11572 49224
rect 11612 49172 11664 49224
rect 13268 49215 13320 49224
rect 13268 49181 13277 49215
rect 13277 49181 13311 49215
rect 13311 49181 13320 49215
rect 13268 49172 13320 49181
rect 16580 49172 16632 49224
rect 16672 49172 16724 49224
rect 21364 49240 21416 49292
rect 22376 49240 22428 49292
rect 22560 49283 22612 49292
rect 22560 49249 22569 49283
rect 22569 49249 22603 49283
rect 22603 49249 22612 49283
rect 22560 49240 22612 49249
rect 24768 49240 24820 49292
rect 30656 49240 30708 49292
rect 30932 49283 30984 49292
rect 30932 49249 30941 49283
rect 30941 49249 30975 49283
rect 30975 49249 30984 49283
rect 30932 49240 30984 49249
rect 40684 49283 40736 49292
rect 40684 49249 40693 49283
rect 40693 49249 40727 49283
rect 40727 49249 40736 49283
rect 40684 49240 40736 49249
rect 46204 49308 46256 49360
rect 46664 49240 46716 49292
rect 46848 49283 46900 49292
rect 46848 49249 46857 49283
rect 46857 49249 46891 49283
rect 46891 49249 46900 49283
rect 46848 49240 46900 49249
rect 19432 49215 19484 49224
rect 19432 49181 19441 49215
rect 19441 49181 19475 49215
rect 19475 49181 19484 49215
rect 19432 49172 19484 49181
rect 20076 49215 20128 49224
rect 20076 49181 20085 49215
rect 20085 49181 20119 49215
rect 20119 49181 20128 49215
rect 20076 49172 20128 49181
rect 20996 49215 21048 49224
rect 20996 49181 21005 49215
rect 21005 49181 21039 49215
rect 21039 49181 21048 49215
rect 20996 49172 21048 49181
rect 2780 49147 2832 49156
rect 2780 49113 2789 49147
rect 2789 49113 2823 49147
rect 2823 49113 2832 49147
rect 2780 49104 2832 49113
rect 2964 49147 3016 49156
rect 2964 49113 2973 49147
rect 2973 49113 3007 49147
rect 3007 49113 3016 49147
rect 2964 49104 3016 49113
rect 4712 49104 4764 49156
rect 21088 49104 21140 49156
rect 22192 49147 22244 49156
rect 22192 49113 22201 49147
rect 22201 49113 22235 49147
rect 22235 49113 22244 49147
rect 22192 49104 22244 49113
rect 1768 49036 1820 49088
rect 5264 49079 5316 49088
rect 5264 49045 5273 49079
rect 5273 49045 5307 49079
rect 5307 49045 5316 49079
rect 5264 49036 5316 49045
rect 6460 49036 6512 49088
rect 8944 49079 8996 49088
rect 8944 49045 8953 49079
rect 8953 49045 8987 49079
rect 8987 49045 8996 49079
rect 8944 49036 8996 49045
rect 11888 49036 11940 49088
rect 13452 49079 13504 49088
rect 13452 49045 13461 49079
rect 13461 49045 13495 49079
rect 13495 49045 13504 49079
rect 13452 49036 13504 49045
rect 20536 49036 20588 49088
rect 26424 49172 26476 49224
rect 27988 49172 28040 49224
rect 24584 49147 24636 49156
rect 24584 49113 24593 49147
rect 24593 49113 24627 49147
rect 24627 49113 24636 49147
rect 24584 49104 24636 49113
rect 27344 49104 27396 49156
rect 29000 49172 29052 49224
rect 33324 49172 33376 49224
rect 35808 49215 35860 49224
rect 35808 49181 35817 49215
rect 35817 49181 35851 49215
rect 35851 49181 35860 49215
rect 35808 49172 35860 49181
rect 38200 49215 38252 49224
rect 29920 49147 29972 49156
rect 29920 49113 29929 49147
rect 29929 49113 29963 49147
rect 29963 49113 29972 49147
rect 29920 49104 29972 49113
rect 25228 49036 25280 49088
rect 25320 49036 25372 49088
rect 26608 49036 26660 49088
rect 27528 49036 27580 49088
rect 29644 49036 29696 49088
rect 32128 49079 32180 49088
rect 32128 49045 32137 49079
rect 32137 49045 32171 49079
rect 32171 49045 32180 49079
rect 32128 49036 32180 49045
rect 34888 49104 34940 49156
rect 38200 49181 38209 49215
rect 38209 49181 38243 49215
rect 38243 49181 38252 49215
rect 38200 49172 38252 49181
rect 39304 49172 39356 49224
rect 42340 49172 42392 49224
rect 44088 49172 44140 49224
rect 47768 49215 47820 49224
rect 47768 49181 47777 49215
rect 47777 49181 47811 49215
rect 47811 49181 47820 49215
rect 47768 49172 47820 49181
rect 38016 49036 38068 49088
rect 44640 49104 44692 49156
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 1952 48764 2004 48816
rect 1676 48696 1728 48748
rect 8944 48739 8996 48748
rect 8944 48705 8953 48739
rect 8953 48705 8987 48739
rect 8987 48705 8996 48739
rect 8944 48696 8996 48705
rect 11520 48739 11572 48748
rect 11520 48705 11529 48739
rect 11529 48705 11563 48739
rect 11563 48705 11572 48739
rect 11520 48696 11572 48705
rect 25320 48832 25372 48884
rect 39672 48832 39724 48884
rect 22008 48807 22060 48816
rect 22008 48773 22017 48807
rect 22017 48773 22051 48807
rect 22051 48773 22060 48807
rect 22008 48764 22060 48773
rect 25964 48807 26016 48816
rect 25964 48773 25973 48807
rect 25973 48773 26007 48807
rect 26007 48773 26016 48807
rect 25964 48764 26016 48773
rect 27528 48764 27580 48816
rect 47768 48807 47820 48816
rect 27344 48739 27396 48748
rect 27344 48705 27353 48739
rect 27353 48705 27387 48739
rect 27387 48705 27396 48739
rect 27344 48696 27396 48705
rect 47768 48773 47777 48807
rect 47777 48773 47811 48807
rect 47811 48773 47820 48807
rect 47768 48764 47820 48773
rect 32128 48739 32180 48748
rect 32128 48705 32137 48739
rect 32137 48705 32171 48739
rect 32171 48705 32180 48739
rect 32128 48696 32180 48705
rect 34888 48739 34940 48748
rect 34888 48705 34897 48739
rect 34897 48705 34931 48739
rect 34931 48705 34940 48739
rect 34888 48696 34940 48705
rect 2228 48671 2280 48680
rect 2228 48637 2237 48671
rect 2237 48637 2271 48671
rect 2271 48637 2280 48671
rect 2228 48628 2280 48637
rect 2872 48671 2924 48680
rect 2872 48637 2881 48671
rect 2881 48637 2915 48671
rect 2915 48637 2924 48671
rect 2872 48628 2924 48637
rect 6552 48671 6604 48680
rect 6552 48637 6561 48671
rect 6561 48637 6595 48671
rect 6595 48637 6604 48671
rect 6552 48628 6604 48637
rect 7196 48671 7248 48680
rect 7196 48637 7205 48671
rect 7205 48637 7239 48671
rect 7239 48637 7248 48671
rect 7196 48628 7248 48637
rect 9128 48671 9180 48680
rect 9128 48637 9137 48671
rect 9137 48637 9171 48671
rect 9171 48637 9180 48671
rect 9128 48628 9180 48637
rect 9680 48671 9732 48680
rect 9680 48637 9689 48671
rect 9689 48637 9723 48671
rect 9723 48637 9732 48671
rect 9680 48628 9732 48637
rect 11704 48671 11756 48680
rect 11704 48637 11713 48671
rect 11713 48637 11747 48671
rect 11747 48637 11756 48671
rect 11704 48628 11756 48637
rect 12440 48671 12492 48680
rect 12440 48637 12449 48671
rect 12449 48637 12483 48671
rect 12483 48637 12492 48671
rect 14188 48671 14240 48680
rect 12440 48628 12492 48637
rect 14188 48637 14197 48671
rect 14197 48637 14231 48671
rect 14231 48637 14240 48671
rect 14188 48628 14240 48637
rect 14372 48671 14424 48680
rect 14372 48637 14381 48671
rect 14381 48637 14415 48671
rect 14415 48637 14424 48671
rect 14372 48628 14424 48637
rect 15200 48671 15252 48680
rect 15200 48637 15209 48671
rect 15209 48637 15243 48671
rect 15243 48637 15252 48671
rect 15200 48628 15252 48637
rect 16948 48671 17000 48680
rect 16948 48637 16957 48671
rect 16957 48637 16991 48671
rect 16991 48637 17000 48671
rect 16948 48628 17000 48637
rect 7564 48560 7616 48612
rect 17224 48628 17276 48680
rect 19432 48671 19484 48680
rect 19432 48637 19441 48671
rect 19441 48637 19475 48671
rect 19475 48637 19484 48671
rect 19432 48628 19484 48637
rect 22652 48671 22704 48680
rect 19340 48560 19392 48612
rect 2136 48492 2188 48544
rect 4620 48492 4672 48544
rect 9036 48492 9088 48544
rect 15108 48492 15160 48544
rect 17960 48492 18012 48544
rect 22652 48637 22661 48671
rect 22661 48637 22695 48671
rect 22695 48637 22704 48671
rect 22652 48628 22704 48637
rect 22836 48671 22888 48680
rect 22836 48637 22845 48671
rect 22845 48637 22879 48671
rect 22879 48637 22888 48671
rect 22836 48628 22888 48637
rect 23480 48671 23532 48680
rect 23480 48637 23489 48671
rect 23489 48637 23523 48671
rect 23523 48637 23532 48671
rect 23480 48628 23532 48637
rect 28724 48628 28776 48680
rect 29828 48671 29880 48680
rect 27620 48560 27672 48612
rect 27712 48560 27764 48612
rect 29828 48637 29837 48671
rect 29837 48637 29871 48671
rect 29871 48637 29880 48671
rect 29828 48628 29880 48637
rect 30012 48628 30064 48680
rect 32312 48671 32364 48680
rect 32312 48637 32321 48671
rect 32321 48637 32355 48671
rect 32355 48637 32364 48671
rect 32312 48628 32364 48637
rect 33140 48671 33192 48680
rect 33140 48637 33149 48671
rect 33149 48637 33183 48671
rect 33183 48637 33192 48671
rect 33140 48628 33192 48637
rect 35900 48628 35952 48680
rect 36084 48671 36136 48680
rect 36084 48637 36093 48671
rect 36093 48637 36127 48671
rect 36127 48637 36136 48671
rect 36084 48628 36136 48637
rect 39764 48671 39816 48680
rect 39764 48637 39773 48671
rect 39773 48637 39807 48671
rect 39807 48637 39816 48671
rect 39764 48628 39816 48637
rect 40040 48671 40092 48680
rect 40040 48637 40049 48671
rect 40049 48637 40083 48671
rect 40083 48637 40092 48671
rect 40040 48628 40092 48637
rect 42432 48671 42484 48680
rect 42432 48637 42441 48671
rect 42441 48637 42475 48671
rect 42475 48637 42484 48671
rect 42432 48628 42484 48637
rect 42616 48671 42668 48680
rect 42616 48637 42625 48671
rect 42625 48637 42659 48671
rect 42659 48637 42668 48671
rect 42616 48628 42668 48637
rect 42800 48628 42852 48680
rect 45376 48671 45428 48680
rect 33416 48560 33468 48612
rect 33876 48560 33928 48612
rect 45376 48637 45385 48671
rect 45385 48637 45419 48671
rect 45419 48637 45428 48671
rect 45376 48628 45428 48637
rect 45744 48671 45796 48680
rect 45744 48637 45753 48671
rect 45753 48637 45787 48671
rect 45787 48637 45796 48671
rect 45744 48628 45796 48637
rect 45468 48560 45520 48612
rect 22100 48535 22152 48544
rect 22100 48501 22109 48535
rect 22109 48501 22143 48535
rect 22143 48501 22152 48535
rect 22100 48492 22152 48501
rect 24952 48492 25004 48544
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 3424 48288 3476 48340
rect 9036 48288 9088 48340
rect 9128 48288 9180 48340
rect 14372 48288 14424 48340
rect 16212 48288 16264 48340
rect 39672 48288 39724 48340
rect 39764 48288 39816 48340
rect 20 48220 72 48272
rect 2780 48220 2832 48272
rect 7564 48263 7616 48272
rect 7564 48229 7573 48263
rect 7573 48229 7607 48263
rect 7607 48229 7616 48263
rect 7564 48220 7616 48229
rect 4068 48152 4120 48204
rect 3608 48084 3660 48136
rect 4436 48127 4488 48136
rect 4436 48093 4445 48127
rect 4445 48093 4479 48127
rect 4479 48093 4488 48127
rect 4436 48084 4488 48093
rect 10324 48152 10376 48204
rect 10692 48152 10744 48204
rect 12900 48127 12952 48136
rect 3148 48016 3200 48068
rect 3240 48059 3292 48068
rect 3240 48025 3249 48059
rect 3249 48025 3283 48059
rect 3283 48025 3292 48059
rect 3240 48016 3292 48025
rect 5356 48016 5408 48068
rect 1952 47948 2004 48000
rect 12900 48093 12909 48127
rect 12909 48093 12943 48127
rect 12943 48093 12952 48127
rect 12900 48084 12952 48093
rect 14464 48127 14516 48136
rect 14464 48093 14473 48127
rect 14473 48093 14507 48127
rect 14507 48093 14516 48127
rect 14464 48084 14516 48093
rect 11612 48016 11664 48068
rect 13728 48016 13780 48068
rect 10968 47948 11020 48000
rect 13360 47948 13412 48000
rect 16948 48220 17000 48272
rect 19340 48263 19392 48272
rect 19340 48229 19349 48263
rect 19349 48229 19383 48263
rect 19383 48229 19392 48263
rect 19340 48220 19392 48229
rect 16580 48195 16632 48204
rect 16580 48161 16589 48195
rect 16589 48161 16623 48195
rect 16623 48161 16632 48195
rect 16580 48152 16632 48161
rect 17408 48195 17460 48204
rect 17408 48161 17417 48195
rect 17417 48161 17451 48195
rect 17451 48161 17460 48195
rect 17408 48152 17460 48161
rect 20996 48220 21048 48272
rect 22836 48220 22888 48272
rect 24584 48220 24636 48272
rect 25228 48263 25280 48272
rect 25228 48229 25237 48263
rect 25237 48229 25271 48263
rect 25271 48229 25280 48263
rect 25228 48220 25280 48229
rect 20628 48152 20680 48204
rect 27068 48195 27120 48204
rect 20076 48084 20128 48136
rect 16028 48016 16080 48068
rect 20168 48016 20220 48068
rect 20260 47948 20312 48000
rect 20352 47948 20404 48000
rect 27068 48161 27077 48195
rect 27077 48161 27111 48195
rect 27111 48161 27120 48195
rect 27068 48152 27120 48161
rect 22652 48084 22704 48136
rect 24400 48127 24452 48136
rect 24400 48093 24409 48127
rect 24409 48093 24443 48127
rect 24443 48093 24452 48127
rect 24400 48084 24452 48093
rect 28724 48263 28776 48272
rect 28724 48229 28733 48263
rect 28733 48229 28767 48263
rect 28767 48229 28776 48263
rect 28724 48220 28776 48229
rect 29920 48220 29972 48272
rect 32220 48195 32272 48204
rect 32220 48161 32229 48195
rect 32229 48161 32263 48195
rect 32263 48161 32272 48195
rect 32220 48152 32272 48161
rect 29736 48127 29788 48136
rect 29736 48093 29745 48127
rect 29745 48093 29779 48127
rect 29779 48093 29788 48127
rect 29736 48084 29788 48093
rect 31024 48127 31076 48136
rect 31024 48093 31033 48127
rect 31033 48093 31067 48127
rect 31067 48093 31076 48127
rect 31024 48084 31076 48093
rect 22928 48016 22980 48068
rect 27068 48016 27120 48068
rect 24400 47948 24452 48000
rect 35808 48152 35860 48204
rect 36728 48195 36780 48204
rect 36728 48161 36737 48195
rect 36737 48161 36771 48195
rect 36771 48161 36780 48195
rect 36728 48152 36780 48161
rect 42616 48220 42668 48272
rect 47032 48220 47084 48272
rect 49608 48220 49660 48272
rect 42524 48152 42576 48204
rect 32496 48084 32548 48136
rect 34796 48084 34848 48136
rect 41052 48127 41104 48136
rect 41052 48093 41061 48127
rect 41061 48093 41095 48127
rect 41095 48093 41104 48127
rect 41052 48084 41104 48093
rect 41788 48127 41840 48136
rect 41788 48093 41797 48127
rect 41797 48093 41831 48127
rect 41831 48093 41840 48127
rect 41788 48084 41840 48093
rect 42800 48152 42852 48204
rect 43168 48195 43220 48204
rect 43168 48161 43177 48195
rect 43177 48161 43211 48195
rect 43211 48161 43220 48195
rect 43168 48152 43220 48161
rect 46756 48195 46808 48204
rect 46756 48161 46765 48195
rect 46765 48161 46799 48195
rect 46799 48161 46808 48195
rect 46756 48152 46808 48161
rect 44732 48084 44784 48136
rect 46296 48127 46348 48136
rect 46296 48093 46305 48127
rect 46305 48093 46339 48127
rect 46339 48093 46348 48127
rect 46296 48084 46348 48093
rect 33508 47948 33560 48000
rect 41880 47991 41932 48000
rect 41880 47957 41889 47991
rect 41889 47957 41923 47991
rect 41923 47957 41932 47991
rect 41880 47948 41932 47957
rect 42064 48016 42116 48068
rect 47676 48016 47728 48068
rect 44180 47948 44232 48000
rect 45100 47948 45152 48000
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 1308 47744 1360 47796
rect 3240 47744 3292 47796
rect 5356 47787 5408 47796
rect 5356 47753 5365 47787
rect 5365 47753 5399 47787
rect 5399 47753 5408 47787
rect 5356 47744 5408 47753
rect 6552 47787 6604 47796
rect 6552 47753 6561 47787
rect 6561 47753 6595 47787
rect 6595 47753 6604 47787
rect 6552 47744 6604 47753
rect 11612 47787 11664 47796
rect 11612 47753 11621 47787
rect 11621 47753 11655 47787
rect 11655 47753 11664 47787
rect 11612 47744 11664 47753
rect 11704 47744 11756 47796
rect 16028 47787 16080 47796
rect 16028 47753 16037 47787
rect 16037 47753 16071 47787
rect 16071 47753 16080 47787
rect 16028 47744 16080 47753
rect 2136 47719 2188 47728
rect 2136 47685 2145 47719
rect 2145 47685 2179 47719
rect 2179 47685 2188 47719
rect 2136 47676 2188 47685
rect 5172 47676 5224 47728
rect 17960 47744 18012 47796
rect 19432 47744 19484 47796
rect 20168 47787 20220 47796
rect 20168 47753 20177 47787
rect 20177 47753 20211 47787
rect 20211 47753 20220 47787
rect 20168 47744 20220 47753
rect 20260 47744 20312 47796
rect 27068 47787 27120 47796
rect 1952 47651 2004 47660
rect 1952 47617 1961 47651
rect 1961 47617 1995 47651
rect 1995 47617 2004 47651
rect 1952 47608 2004 47617
rect 4436 47608 4488 47660
rect 3056 47583 3108 47592
rect 3056 47549 3065 47583
rect 3065 47549 3099 47583
rect 3099 47549 3108 47583
rect 3056 47540 3108 47549
rect 6920 47608 6972 47660
rect 7104 47651 7156 47660
rect 7104 47617 7113 47651
rect 7113 47617 7147 47651
rect 7147 47617 7156 47651
rect 7104 47608 7156 47617
rect 11520 47651 11572 47660
rect 11520 47617 11529 47651
rect 11529 47617 11563 47651
rect 11563 47617 11572 47651
rect 11520 47608 11572 47617
rect 12072 47608 12124 47660
rect 14188 47608 14240 47660
rect 15568 47608 15620 47660
rect 18420 47676 18472 47728
rect 22192 47676 22244 47728
rect 27068 47753 27077 47787
rect 27077 47753 27111 47787
rect 27111 47753 27120 47787
rect 27068 47744 27120 47753
rect 29828 47744 29880 47796
rect 32312 47744 32364 47796
rect 35900 47787 35952 47796
rect 35900 47753 35909 47787
rect 35909 47753 35943 47787
rect 35943 47753 35952 47787
rect 35900 47744 35952 47753
rect 42064 47744 42116 47796
rect 42524 47744 42576 47796
rect 31852 47676 31904 47728
rect 33508 47719 33560 47728
rect 19064 47651 19116 47660
rect 19064 47617 19073 47651
rect 19073 47617 19107 47651
rect 19107 47617 19116 47651
rect 19064 47608 19116 47617
rect 19340 47608 19392 47660
rect 21732 47608 21784 47660
rect 22376 47608 22428 47660
rect 24124 47651 24176 47660
rect 24124 47617 24133 47651
rect 24133 47617 24167 47651
rect 24167 47617 24176 47651
rect 24124 47608 24176 47617
rect 7656 47540 7708 47592
rect 7748 47583 7800 47592
rect 7748 47549 7757 47583
rect 7757 47549 7791 47583
rect 7791 47549 7800 47583
rect 16948 47583 17000 47592
rect 7748 47540 7800 47549
rect 16948 47549 16957 47583
rect 16957 47549 16991 47583
rect 16991 47549 17000 47583
rect 16948 47540 17000 47549
rect 15108 47472 15160 47524
rect 27620 47608 27672 47660
rect 30012 47651 30064 47660
rect 30012 47617 30021 47651
rect 30021 47617 30055 47651
rect 30055 47617 30064 47651
rect 30012 47608 30064 47617
rect 31024 47608 31076 47660
rect 33508 47685 33517 47719
rect 33517 47685 33551 47719
rect 33551 47685 33560 47719
rect 33508 47676 33560 47685
rect 33324 47651 33376 47660
rect 33324 47617 33333 47651
rect 33333 47617 33367 47651
rect 33367 47617 33376 47651
rect 33324 47608 33376 47617
rect 41696 47651 41748 47660
rect 28172 47540 28224 47592
rect 28356 47583 28408 47592
rect 28356 47549 28365 47583
rect 28365 47549 28399 47583
rect 28399 47549 28408 47583
rect 28356 47540 28408 47549
rect 29828 47540 29880 47592
rect 32496 47540 32548 47592
rect 34704 47583 34756 47592
rect 34704 47549 34713 47583
rect 34713 47549 34747 47583
rect 34747 47549 34756 47583
rect 34704 47540 34756 47549
rect 26976 47472 27028 47524
rect 30748 47472 30800 47524
rect 13268 47404 13320 47456
rect 19064 47404 19116 47456
rect 20076 47404 20128 47456
rect 23940 47447 23992 47456
rect 23940 47413 23949 47447
rect 23949 47413 23983 47447
rect 23983 47413 23992 47447
rect 23940 47404 23992 47413
rect 34520 47404 34572 47456
rect 41696 47617 41705 47651
rect 41705 47617 41739 47651
rect 41739 47617 41748 47651
rect 41696 47608 41748 47617
rect 46204 47744 46256 47796
rect 48320 47744 48372 47796
rect 47768 47719 47820 47728
rect 47768 47685 47777 47719
rect 47777 47685 47811 47719
rect 47811 47685 47820 47719
rect 47768 47676 47820 47685
rect 43444 47540 43496 47592
rect 46020 47540 46072 47592
rect 40684 47472 40736 47524
rect 44548 47404 44600 47456
rect 45192 47404 45244 47456
rect 46388 47404 46440 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 2228 47200 2280 47252
rect 3148 47200 3200 47252
rect 7656 47243 7708 47252
rect 7656 47209 7665 47243
rect 7665 47209 7699 47243
rect 7699 47209 7708 47243
rect 7656 47200 7708 47209
rect 16948 47243 17000 47252
rect 16948 47209 16957 47243
rect 16957 47209 16991 47243
rect 16991 47209 17000 47243
rect 16948 47200 17000 47209
rect 18052 47200 18104 47252
rect 40684 47200 40736 47252
rect 42432 47200 42484 47252
rect 43444 47243 43496 47252
rect 43444 47209 43453 47243
rect 43453 47209 43487 47243
rect 43487 47209 43496 47243
rect 43444 47200 43496 47209
rect 6920 47132 6972 47184
rect 17868 47132 17920 47184
rect 18236 47132 18288 47184
rect 26976 47132 27028 47184
rect 14464 47064 14516 47116
rect 29828 47132 29880 47184
rect 30656 47175 30708 47184
rect 30656 47141 30665 47175
rect 30665 47141 30699 47175
rect 30699 47141 30708 47175
rect 30656 47132 30708 47141
rect 30748 47132 30800 47184
rect 41696 47132 41748 47184
rect 43996 47132 44048 47184
rect 1400 47039 1452 47048
rect 1400 47005 1409 47039
rect 1409 47005 1443 47039
rect 1443 47005 1452 47039
rect 1400 46996 1452 47005
rect 2412 47039 2464 47048
rect 2412 47005 2421 47039
rect 2421 47005 2455 47039
rect 2455 47005 2464 47039
rect 2412 46996 2464 47005
rect 2780 46996 2832 47048
rect 7932 46996 7984 47048
rect 19248 47039 19300 47048
rect 19248 47005 19257 47039
rect 19257 47005 19291 47039
rect 19291 47005 19300 47039
rect 19248 46996 19300 47005
rect 30012 47064 30064 47116
rect 39856 47064 39908 47116
rect 45192 47107 45244 47116
rect 45192 47073 45201 47107
rect 45201 47073 45235 47107
rect 45235 47073 45244 47107
rect 45192 47064 45244 47073
rect 45284 47064 45336 47116
rect 28080 47039 28132 47048
rect 28080 47005 28089 47039
rect 28089 47005 28123 47039
rect 28123 47005 28132 47039
rect 28080 46996 28132 47005
rect 28172 47039 28224 47048
rect 28172 47005 28181 47039
rect 28181 47005 28215 47039
rect 28215 47005 28224 47039
rect 43904 47039 43956 47048
rect 28172 46996 28224 47005
rect 43904 47005 43913 47039
rect 43913 47005 43947 47039
rect 43947 47005 43956 47039
rect 43904 46996 43956 47005
rect 45008 47039 45060 47048
rect 45008 47005 45017 47039
rect 45017 47005 45051 47039
rect 45051 47005 45060 47039
rect 45008 46996 45060 47005
rect 48964 46996 49016 47048
rect 20076 46971 20128 46980
rect 20076 46937 20085 46971
rect 20085 46937 20119 46971
rect 20119 46937 20128 46971
rect 20076 46928 20128 46937
rect 31024 46928 31076 46980
rect 47952 46860 48004 46912
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 44640 46699 44692 46708
rect 44640 46665 44649 46699
rect 44649 46665 44683 46699
rect 44683 46665 44692 46699
rect 44640 46656 44692 46665
rect 47676 46699 47728 46708
rect 47676 46665 47685 46699
rect 47685 46665 47719 46699
rect 47719 46665 47728 46699
rect 47676 46656 47728 46665
rect 2780 46588 2832 46640
rect 3792 46631 3844 46640
rect 3792 46597 3801 46631
rect 3801 46597 3835 46631
rect 3835 46597 3844 46631
rect 3792 46588 3844 46597
rect 18236 46631 18288 46640
rect 18236 46597 18245 46631
rect 18245 46597 18279 46631
rect 18279 46597 18288 46631
rect 18236 46588 18288 46597
rect 22928 46588 22980 46640
rect 19248 46520 19300 46572
rect 42800 46563 42852 46572
rect 42800 46529 42809 46563
rect 42809 46529 42843 46563
rect 42843 46529 42852 46563
rect 42800 46520 42852 46529
rect 44088 46563 44140 46572
rect 44088 46529 44097 46563
rect 44097 46529 44131 46563
rect 44131 46529 44140 46563
rect 44088 46520 44140 46529
rect 44548 46563 44600 46572
rect 44548 46529 44557 46563
rect 44557 46529 44591 46563
rect 44591 46529 44600 46563
rect 44548 46520 44600 46529
rect 47032 46563 47084 46572
rect 47032 46529 47041 46563
rect 47041 46529 47075 46563
rect 47075 46529 47084 46563
rect 47032 46520 47084 46529
rect 2504 46452 2556 46504
rect 20076 46495 20128 46504
rect 20076 46461 20085 46495
rect 20085 46461 20119 46495
rect 20119 46461 20128 46495
rect 20076 46452 20128 46461
rect 46388 46452 46440 46504
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 2504 46155 2556 46164
rect 2504 46121 2513 46155
rect 2513 46121 2547 46155
rect 2547 46121 2556 46155
rect 2504 46112 2556 46121
rect 19248 46112 19300 46164
rect 45008 46112 45060 46164
rect 45376 46112 45428 46164
rect 47768 45976 47820 46028
rect 48136 46019 48188 46028
rect 48136 45985 48145 46019
rect 48145 45985 48179 46019
rect 48179 45985 48188 46019
rect 48136 45976 48188 45985
rect 1400 45951 1452 45960
rect 1400 45917 1409 45951
rect 1409 45917 1443 45951
rect 1443 45917 1452 45951
rect 1400 45908 1452 45917
rect 2504 45908 2556 45960
rect 3240 45951 3292 45960
rect 3240 45917 3249 45951
rect 3249 45917 3283 45951
rect 3283 45917 3292 45951
rect 3240 45908 3292 45917
rect 3976 45951 4028 45960
rect 3976 45917 3985 45951
rect 3985 45917 4019 45951
rect 4019 45917 4028 45951
rect 3976 45908 4028 45917
rect 13268 45951 13320 45960
rect 13268 45917 13277 45951
rect 13277 45917 13311 45951
rect 13311 45917 13320 45951
rect 13268 45908 13320 45917
rect 18236 45908 18288 45960
rect 18420 45951 18472 45960
rect 18420 45917 18429 45951
rect 18429 45917 18463 45951
rect 18463 45917 18472 45951
rect 19248 45951 19300 45960
rect 18420 45908 18472 45917
rect 19248 45917 19257 45951
rect 19257 45917 19291 45951
rect 19291 45917 19300 45951
rect 19248 45908 19300 45917
rect 44180 45908 44232 45960
rect 45928 45908 45980 45960
rect 13084 45772 13136 45824
rect 19156 45840 19208 45892
rect 19984 45840 20036 45892
rect 34520 45840 34572 45892
rect 47676 45840 47728 45892
rect 22836 45772 22888 45824
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 2504 45568 2556 45620
rect 3240 45500 3292 45552
rect 20076 45568 20128 45620
rect 28080 45568 28132 45620
rect 28816 45568 28868 45620
rect 13084 45543 13136 45552
rect 3884 45364 3936 45416
rect 4068 45407 4120 45416
rect 4068 45373 4077 45407
rect 4077 45373 4111 45407
rect 4111 45373 4120 45407
rect 4068 45364 4120 45373
rect 13084 45509 13093 45543
rect 13093 45509 13127 45543
rect 13127 45509 13136 45543
rect 13084 45500 13136 45509
rect 47676 45543 47728 45552
rect 19248 45432 19300 45484
rect 13176 45364 13228 45416
rect 13820 45407 13872 45416
rect 13820 45373 13829 45407
rect 13829 45373 13863 45407
rect 13863 45373 13872 45407
rect 13820 45364 13872 45373
rect 21548 45364 21600 45416
rect 28816 45364 28868 45416
rect 42340 45432 42392 45484
rect 45468 45475 45520 45484
rect 45468 45441 45477 45475
rect 45477 45441 45511 45475
rect 45511 45441 45520 45475
rect 45468 45432 45520 45441
rect 46296 45432 46348 45484
rect 47676 45509 47685 45543
rect 47685 45509 47719 45543
rect 47719 45509 47728 45543
rect 47676 45500 47728 45509
rect 46756 45364 46808 45416
rect 47124 45432 47176 45484
rect 1400 45228 1452 45280
rect 2044 45228 2096 45280
rect 46480 45228 46532 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 3884 45067 3936 45076
rect 3884 45033 3893 45067
rect 3893 45033 3927 45067
rect 3927 45033 3936 45067
rect 3884 45024 3936 45033
rect 13176 45067 13228 45076
rect 13176 45033 13185 45067
rect 13185 45033 13219 45067
rect 13219 45033 13228 45067
rect 13176 45024 13228 45033
rect 1400 44931 1452 44940
rect 1400 44897 1409 44931
rect 1409 44897 1443 44931
rect 1443 44897 1452 44931
rect 1400 44888 1452 44897
rect 2780 44931 2832 44940
rect 2780 44897 2789 44931
rect 2789 44897 2823 44931
rect 2823 44897 2832 44931
rect 2780 44888 2832 44897
rect 46480 44931 46532 44940
rect 46480 44897 46489 44931
rect 46489 44897 46523 44931
rect 46523 44897 46532 44931
rect 46480 44888 46532 44897
rect 48136 44931 48188 44940
rect 48136 44897 48145 44931
rect 48145 44897 48179 44931
rect 48179 44897 48188 44931
rect 48136 44888 48188 44897
rect 3792 44863 3844 44872
rect 3792 44829 3801 44863
rect 3801 44829 3835 44863
rect 3835 44829 3844 44863
rect 3792 44820 3844 44829
rect 45192 44863 45244 44872
rect 45192 44829 45201 44863
rect 45201 44829 45235 44863
rect 45235 44829 45244 44863
rect 45192 44820 45244 44829
rect 2780 44752 2832 44804
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 3976 44480 4028 44532
rect 2044 44455 2096 44464
rect 2044 44421 2053 44455
rect 2053 44421 2087 44455
rect 2087 44421 2096 44455
rect 2044 44412 2096 44421
rect 47308 44412 47360 44464
rect 45192 44387 45244 44396
rect 45192 44353 45201 44387
rect 45201 44353 45235 44387
rect 45235 44353 45244 44387
rect 45192 44344 45244 44353
rect 47768 44387 47820 44396
rect 47768 44353 47777 44387
rect 47777 44353 47811 44387
rect 47811 44353 47820 44387
rect 47768 44344 47820 44353
rect 2872 44319 2924 44328
rect 2872 44285 2881 44319
rect 2881 44285 2915 44319
rect 2915 44285 2924 44319
rect 2872 44276 2924 44285
rect 46848 44319 46900 44328
rect 46848 44285 46857 44319
rect 46857 44285 46891 44319
rect 46891 44285 46900 44319
rect 46848 44276 46900 44285
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 2780 43979 2832 43988
rect 2780 43945 2789 43979
rect 2789 43945 2823 43979
rect 2823 43945 2832 43979
rect 2780 43936 2832 43945
rect 1860 43775 1912 43784
rect 1860 43741 1869 43775
rect 1869 43741 1903 43775
rect 1903 43741 1912 43775
rect 1860 43732 1912 43741
rect 2136 43732 2188 43784
rect 46940 43664 46992 43716
rect 48136 43707 48188 43716
rect 48136 43673 48145 43707
rect 48145 43673 48179 43707
rect 48179 43673 48188 43707
rect 48136 43664 48188 43673
rect 1952 43639 2004 43648
rect 1952 43605 1961 43639
rect 1961 43605 1995 43639
rect 1995 43605 2004 43639
rect 1952 43596 2004 43605
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 46940 43435 46992 43444
rect 46940 43401 46949 43435
rect 46949 43401 46983 43435
rect 46983 43401 46992 43435
rect 46940 43392 46992 43401
rect 1860 43367 1912 43376
rect 1860 43333 1869 43367
rect 1869 43333 1903 43367
rect 1903 43333 1912 43367
rect 1860 43324 1912 43333
rect 7932 43256 7984 43308
rect 47860 43299 47912 43308
rect 47860 43265 47869 43299
rect 47869 43265 47903 43299
rect 47903 43265 47912 43299
rect 47860 43256 47912 43265
rect 2228 43052 2280 43104
rect 48228 43052 48280 43104
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 47308 42755 47360 42764
rect 47308 42721 47317 42755
rect 47317 42721 47351 42755
rect 47351 42721 47360 42755
rect 47308 42712 47360 42721
rect 47216 42687 47268 42696
rect 47216 42653 47225 42687
rect 47225 42653 47259 42687
rect 47259 42653 47268 42687
rect 47216 42644 47268 42653
rect 47952 42619 48004 42628
rect 22652 42508 22704 42560
rect 47952 42585 47961 42619
rect 47961 42585 47995 42619
rect 47995 42585 48004 42619
rect 47952 42576 48004 42585
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 46756 42211 46808 42220
rect 46756 42177 46765 42211
rect 46765 42177 46799 42211
rect 46799 42177 46808 42211
rect 46756 42168 46808 42177
rect 20444 42032 20496 42084
rect 20628 42032 20680 42084
rect 1400 41964 1452 42016
rect 46480 41964 46532 42016
rect 47768 42007 47820 42016
rect 47768 41973 47777 42007
rect 47777 41973 47811 42007
rect 47811 41973 47820 42007
rect 47768 41964 47820 41973
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 1400 41667 1452 41676
rect 1400 41633 1409 41667
rect 1409 41633 1443 41667
rect 1443 41633 1452 41667
rect 1400 41624 1452 41633
rect 1860 41667 1912 41676
rect 1860 41633 1869 41667
rect 1869 41633 1903 41667
rect 1903 41633 1912 41667
rect 1860 41624 1912 41633
rect 47768 41692 47820 41744
rect 46480 41667 46532 41676
rect 46480 41633 46489 41667
rect 46489 41633 46523 41667
rect 46523 41633 46532 41667
rect 46480 41624 46532 41633
rect 21088 41556 21140 41608
rect 24124 41556 24176 41608
rect 1584 41531 1636 41540
rect 1584 41497 1593 41531
rect 1593 41497 1627 41531
rect 1627 41497 1636 41531
rect 1584 41488 1636 41497
rect 48136 41531 48188 41540
rect 48136 41497 48145 41531
rect 48145 41497 48179 41531
rect 48179 41497 48188 41531
rect 48136 41488 48188 41497
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 1584 41216 1636 41268
rect 1860 41123 1912 41132
rect 1860 41089 1869 41123
rect 1869 41089 1903 41123
rect 1903 41089 1912 41123
rect 1860 41080 1912 41089
rect 1492 41012 1544 41064
rect 45744 41080 45796 41132
rect 46204 41055 46256 41064
rect 46204 41021 46213 41055
rect 46213 41021 46247 41055
rect 46247 41021 46256 41055
rect 46204 41012 46256 41021
rect 2320 40944 2372 40996
rect 46296 40876 46348 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 21824 40536 21876 40588
rect 1400 40511 1452 40520
rect 1400 40477 1409 40511
rect 1409 40477 1443 40511
rect 1443 40477 1452 40511
rect 1400 40468 1452 40477
rect 22652 40511 22704 40520
rect 22652 40477 22661 40511
rect 22661 40477 22695 40511
rect 22695 40477 22704 40511
rect 22652 40468 22704 40477
rect 23388 40536 23440 40588
rect 46296 40579 46348 40588
rect 46296 40545 46305 40579
rect 46305 40545 46339 40579
rect 46339 40545 46348 40579
rect 46296 40536 46348 40545
rect 22468 40400 22520 40452
rect 23848 40468 23900 40520
rect 47676 40400 47728 40452
rect 48136 40443 48188 40452
rect 48136 40409 48145 40443
rect 48145 40409 48179 40443
rect 48179 40409 48188 40443
rect 48136 40400 48188 40409
rect 1584 40375 1636 40384
rect 1584 40341 1593 40375
rect 1593 40341 1627 40375
rect 1627 40341 1636 40375
rect 1584 40332 1636 40341
rect 22376 40375 22428 40384
rect 22376 40341 22385 40375
rect 22385 40341 22419 40375
rect 22419 40341 22428 40375
rect 22376 40332 22428 40341
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 22652 40128 22704 40180
rect 24032 40128 24084 40180
rect 22376 40060 22428 40112
rect 20996 40035 21048 40044
rect 20996 40001 21005 40035
rect 21005 40001 21039 40035
rect 21039 40001 21048 40035
rect 20996 39992 21048 40001
rect 21272 40035 21324 40044
rect 21272 40001 21281 40035
rect 21281 40001 21315 40035
rect 21315 40001 21324 40035
rect 21272 39992 21324 40001
rect 23112 39992 23164 40044
rect 44548 39992 44600 40044
rect 47308 39992 47360 40044
rect 47676 40035 47728 40044
rect 47676 40001 47685 40035
rect 47685 40001 47719 40035
rect 47719 40001 47728 40035
rect 47676 39992 47728 40001
rect 20444 39924 20496 39976
rect 23664 39967 23716 39976
rect 23664 39933 23673 39967
rect 23673 39933 23707 39967
rect 23707 39933 23716 39967
rect 23664 39924 23716 39933
rect 18880 39856 18932 39908
rect 20904 39788 20956 39840
rect 24400 39788 24452 39840
rect 25044 39831 25096 39840
rect 25044 39797 25053 39831
rect 25053 39797 25087 39831
rect 25087 39797 25096 39831
rect 25044 39788 25096 39797
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 23112 39627 23164 39636
rect 23112 39593 23121 39627
rect 23121 39593 23155 39627
rect 23155 39593 23164 39627
rect 23112 39584 23164 39593
rect 23940 39584 23992 39636
rect 20444 39491 20496 39500
rect 20444 39457 20453 39491
rect 20453 39457 20487 39491
rect 20487 39457 20496 39491
rect 20444 39448 20496 39457
rect 2044 39380 2096 39432
rect 18236 39380 18288 39432
rect 18328 39423 18380 39432
rect 18328 39389 18337 39423
rect 18337 39389 18371 39423
rect 18371 39389 18380 39423
rect 18328 39380 18380 39389
rect 20720 39355 20772 39364
rect 20720 39321 20754 39355
rect 20754 39321 20772 39355
rect 23388 39516 23440 39568
rect 23756 39516 23808 39568
rect 23664 39448 23716 39500
rect 23572 39423 23624 39432
rect 23572 39389 23581 39423
rect 23581 39389 23615 39423
rect 23615 39389 23624 39423
rect 23572 39380 23624 39389
rect 23848 39380 23900 39432
rect 26700 39380 26752 39432
rect 47676 39423 47728 39432
rect 47676 39389 47685 39423
rect 47685 39389 47719 39423
rect 47719 39389 47728 39423
rect 47676 39380 47728 39389
rect 20720 39312 20772 39321
rect 23664 39312 23716 39364
rect 26976 39312 27028 39364
rect 17224 39244 17276 39296
rect 19432 39244 19484 39296
rect 21272 39244 21324 39296
rect 22008 39244 22060 39296
rect 23020 39244 23072 39296
rect 25044 39244 25096 39296
rect 25780 39287 25832 39296
rect 25780 39253 25789 39287
rect 25789 39253 25823 39287
rect 25823 39253 25832 39287
rect 25780 39244 25832 39253
rect 29276 39244 29328 39296
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 20720 39040 20772 39092
rect 22652 39083 22704 39092
rect 22652 39049 22661 39083
rect 22661 39049 22695 39083
rect 22695 39049 22704 39083
rect 22652 39040 22704 39049
rect 23296 39040 23348 39092
rect 23480 39040 23532 39092
rect 26976 39083 27028 39092
rect 26976 39049 26985 39083
rect 26985 39049 27019 39083
rect 27019 39049 27028 39083
rect 26976 39040 27028 39049
rect 2964 38972 3016 39024
rect 2044 38947 2096 38956
rect 2044 38913 2053 38947
rect 2053 38913 2087 38947
rect 2087 38913 2096 38947
rect 2044 38904 2096 38913
rect 17224 38947 17276 38956
rect 17224 38913 17233 38947
rect 17233 38913 17267 38947
rect 17267 38913 17276 38947
rect 17224 38904 17276 38913
rect 18604 38947 18656 38956
rect 18604 38913 18613 38947
rect 18613 38913 18647 38947
rect 18647 38913 18656 38947
rect 18604 38904 18656 38913
rect 21824 38972 21876 39024
rect 20904 38947 20956 38956
rect 20904 38913 20913 38947
rect 20913 38913 20947 38947
rect 20947 38913 20956 38947
rect 20904 38904 20956 38913
rect 21088 38947 21140 38956
rect 21088 38913 21097 38947
rect 21097 38913 21131 38947
rect 21131 38913 21140 38947
rect 21088 38904 21140 38913
rect 22560 38904 22612 38956
rect 23020 38904 23072 38956
rect 23940 38972 23992 39024
rect 26700 38972 26752 39024
rect 26792 38972 26844 39024
rect 2964 38836 3016 38888
rect 3056 38879 3108 38888
rect 3056 38845 3065 38879
rect 3065 38845 3099 38879
rect 3099 38845 3108 38879
rect 18880 38879 18932 38888
rect 3056 38836 3108 38845
rect 18880 38845 18889 38879
rect 18889 38845 18923 38879
rect 18923 38845 18932 38879
rect 18880 38836 18932 38845
rect 23204 38836 23256 38888
rect 23756 38836 23808 38888
rect 25136 38904 25188 38956
rect 13728 38768 13780 38820
rect 18328 38700 18380 38752
rect 19984 38743 20036 38752
rect 19984 38709 19993 38743
rect 19993 38709 20027 38743
rect 20027 38709 20036 38743
rect 19984 38700 20036 38709
rect 21088 38768 21140 38820
rect 23848 38768 23900 38820
rect 26240 38836 26292 38888
rect 27528 38904 27580 38956
rect 26148 38768 26200 38820
rect 30196 38904 30248 38956
rect 30932 38904 30984 38956
rect 47952 38947 48004 38956
rect 47952 38913 47961 38947
rect 47961 38913 47995 38947
rect 47995 38913 48004 38947
rect 47952 38904 48004 38913
rect 26424 38743 26476 38752
rect 26424 38709 26433 38743
rect 26433 38709 26467 38743
rect 26467 38709 26476 38743
rect 26424 38700 26476 38709
rect 31116 38700 31168 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 2964 38539 3016 38548
rect 2964 38505 2973 38539
rect 2973 38505 3007 38539
rect 3007 38505 3016 38539
rect 2964 38496 3016 38505
rect 21824 38539 21876 38548
rect 21824 38505 21833 38539
rect 21833 38505 21867 38539
rect 21867 38505 21876 38539
rect 21824 38496 21876 38505
rect 22468 38496 22520 38548
rect 38752 38496 38804 38548
rect 23940 38428 23992 38480
rect 25136 38428 25188 38480
rect 35164 38428 35216 38480
rect 39304 38428 39356 38480
rect 19432 38403 19484 38412
rect 19432 38369 19441 38403
rect 19441 38369 19475 38403
rect 19475 38369 19484 38403
rect 19432 38360 19484 38369
rect 20996 38360 21048 38412
rect 21640 38360 21692 38412
rect 8944 38292 8996 38344
rect 6920 38224 6972 38276
rect 15568 38224 15620 38276
rect 16120 38292 16172 38344
rect 19248 38335 19300 38344
rect 19248 38301 19257 38335
rect 19257 38301 19291 38335
rect 19291 38301 19300 38335
rect 19248 38292 19300 38301
rect 22652 38360 22704 38412
rect 22928 38360 22980 38412
rect 17408 38224 17460 38276
rect 18328 38156 18380 38208
rect 22376 38224 22428 38276
rect 22744 38335 22796 38344
rect 22744 38301 22753 38335
rect 22753 38301 22787 38335
rect 22787 38301 22796 38335
rect 22744 38292 22796 38301
rect 24032 38360 24084 38412
rect 23480 38335 23532 38344
rect 23480 38301 23489 38335
rect 23489 38301 23523 38335
rect 23523 38301 23532 38335
rect 23480 38292 23532 38301
rect 25780 38360 25832 38412
rect 31300 38360 31352 38412
rect 24216 38292 24268 38344
rect 25228 38335 25280 38344
rect 25228 38301 25237 38335
rect 25237 38301 25271 38335
rect 25271 38301 25280 38335
rect 25228 38292 25280 38301
rect 26148 38292 26200 38344
rect 26424 38292 26476 38344
rect 29460 38292 29512 38344
rect 31484 38292 31536 38344
rect 31668 38335 31720 38344
rect 31668 38301 31677 38335
rect 31677 38301 31711 38335
rect 31711 38301 31720 38335
rect 31668 38292 31720 38301
rect 47676 38360 47728 38412
rect 48136 38403 48188 38412
rect 48136 38369 48145 38403
rect 48145 38369 48179 38403
rect 48179 38369 48188 38403
rect 48136 38360 48188 38369
rect 31944 38292 31996 38344
rect 32128 38292 32180 38344
rect 22652 38156 22704 38208
rect 22744 38156 22796 38208
rect 25872 38224 25924 38276
rect 27896 38224 27948 38276
rect 31392 38267 31444 38276
rect 31392 38233 31401 38267
rect 31401 38233 31435 38267
rect 31435 38233 31444 38267
rect 31392 38224 31444 38233
rect 38936 38224 38988 38276
rect 29920 38156 29972 38208
rect 30012 38156 30064 38208
rect 32036 38156 32088 38208
rect 46664 38156 46716 38208
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 5264 37952 5316 38004
rect 1492 37884 1544 37936
rect 19708 37927 19760 37936
rect 19708 37893 19717 37927
rect 19717 37893 19751 37927
rect 19751 37893 19760 37927
rect 19708 37884 19760 37893
rect 21824 37884 21876 37936
rect 1860 37859 1912 37868
rect 1860 37825 1869 37859
rect 1869 37825 1903 37859
rect 1903 37825 1912 37859
rect 1860 37816 1912 37825
rect 8944 37859 8996 37868
rect 8944 37825 8953 37859
rect 8953 37825 8987 37859
rect 8987 37825 8996 37859
rect 8944 37816 8996 37825
rect 17224 37859 17276 37868
rect 17224 37825 17233 37859
rect 17233 37825 17267 37859
rect 17267 37825 17276 37859
rect 17224 37816 17276 37825
rect 18604 37859 18656 37868
rect 1676 37748 1728 37800
rect 15568 37748 15620 37800
rect 9128 37612 9180 37664
rect 14004 37680 14056 37732
rect 14096 37680 14148 37732
rect 17408 37791 17460 37800
rect 17408 37757 17417 37791
rect 17417 37757 17451 37791
rect 17451 37757 17460 37791
rect 18604 37825 18613 37859
rect 18613 37825 18647 37859
rect 18647 37825 18656 37859
rect 18604 37816 18656 37825
rect 22284 37859 22336 37868
rect 22284 37825 22293 37859
rect 22293 37825 22327 37859
rect 22327 37825 22336 37859
rect 22284 37816 22336 37825
rect 22468 37859 22520 37868
rect 22468 37825 22477 37859
rect 22477 37825 22511 37859
rect 22511 37825 22520 37859
rect 23020 37859 23072 37868
rect 22468 37816 22520 37825
rect 23020 37825 23029 37859
rect 23029 37825 23063 37859
rect 23063 37825 23072 37859
rect 23020 37816 23072 37825
rect 23204 37859 23256 37868
rect 23204 37825 23213 37859
rect 23213 37825 23247 37859
rect 23247 37825 23256 37859
rect 23204 37816 23256 37825
rect 24860 37816 24912 37868
rect 25412 37859 25464 37868
rect 25412 37825 25421 37859
rect 25421 37825 25455 37859
rect 25455 37825 25464 37859
rect 25412 37816 25464 37825
rect 26332 37952 26384 38004
rect 27896 37927 27948 37936
rect 27896 37893 27905 37927
rect 27905 37893 27939 37927
rect 27939 37893 27948 37927
rect 27896 37884 27948 37893
rect 20720 37791 20772 37800
rect 17408 37748 17460 37757
rect 20720 37757 20729 37791
rect 20729 37757 20763 37791
rect 20763 37757 20772 37791
rect 20720 37748 20772 37757
rect 22560 37748 22612 37800
rect 23388 37748 23440 37800
rect 26056 37748 26108 37800
rect 21824 37655 21876 37664
rect 21824 37621 21833 37655
rect 21833 37621 21867 37655
rect 21867 37621 21876 37655
rect 21824 37612 21876 37621
rect 28908 37816 28960 37868
rect 29368 37859 29420 37868
rect 29368 37825 29377 37859
rect 29377 37825 29411 37859
rect 29411 37825 29420 37859
rect 29368 37816 29420 37825
rect 29184 37748 29236 37800
rect 29460 37791 29512 37800
rect 29460 37757 29469 37791
rect 29469 37757 29503 37791
rect 29503 37757 29512 37791
rect 29460 37748 29512 37757
rect 30288 37748 30340 37800
rect 31116 37859 31168 37868
rect 31116 37825 31125 37859
rect 31125 37825 31159 37859
rect 31159 37825 31168 37859
rect 31116 37816 31168 37825
rect 47032 37884 47084 37936
rect 47216 37884 47268 37936
rect 47860 37859 47912 37868
rect 31208 37748 31260 37800
rect 28356 37680 28408 37732
rect 28908 37680 28960 37732
rect 47860 37825 47869 37859
rect 47869 37825 47903 37859
rect 47903 37825 47912 37859
rect 47860 37816 47912 37825
rect 31484 37748 31536 37800
rect 31576 37680 31628 37732
rect 32036 37680 32088 37732
rect 23388 37655 23440 37664
rect 23388 37621 23397 37655
rect 23397 37621 23431 37655
rect 23431 37621 23440 37655
rect 23388 37612 23440 37621
rect 26792 37612 26844 37664
rect 29000 37655 29052 37664
rect 29000 37621 29009 37655
rect 29009 37621 29043 37655
rect 29043 37621 29052 37655
rect 29000 37612 29052 37621
rect 29368 37612 29420 37664
rect 30012 37612 30064 37664
rect 30564 37612 30616 37664
rect 35624 37612 35676 37664
rect 47492 37612 47544 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 8944 37408 8996 37460
rect 20720 37408 20772 37460
rect 21456 37408 21508 37460
rect 23020 37408 23072 37460
rect 4068 37340 4120 37392
rect 1400 37315 1452 37324
rect 1400 37281 1409 37315
rect 1409 37281 1443 37315
rect 1443 37281 1452 37315
rect 1400 37272 1452 37281
rect 9128 37315 9180 37324
rect 9128 37281 9137 37315
rect 9137 37281 9171 37315
rect 9171 37281 9180 37315
rect 9128 37272 9180 37281
rect 14004 37340 14056 37392
rect 17408 37340 17460 37392
rect 22376 37340 22428 37392
rect 25228 37408 25280 37460
rect 27436 37408 27488 37460
rect 29184 37408 29236 37460
rect 26148 37340 26200 37392
rect 28356 37340 28408 37392
rect 31300 37340 31352 37392
rect 15292 37272 15344 37324
rect 23572 37315 23624 37324
rect 23572 37281 23581 37315
rect 23581 37281 23615 37315
rect 23615 37281 23624 37315
rect 23572 37272 23624 37281
rect 25688 37272 25740 37324
rect 25872 37272 25924 37324
rect 1676 37247 1728 37256
rect 1676 37213 1685 37247
rect 1685 37213 1719 37247
rect 1719 37213 1728 37247
rect 1676 37204 1728 37213
rect 8944 37247 8996 37256
rect 8944 37213 8953 37247
rect 8953 37213 8987 37247
rect 8987 37213 8996 37247
rect 8944 37204 8996 37213
rect 15108 37247 15160 37256
rect 15108 37213 15117 37247
rect 15117 37213 15151 37247
rect 15151 37213 15160 37247
rect 15108 37204 15160 37213
rect 17224 37204 17276 37256
rect 15292 37179 15344 37188
rect 15292 37145 15301 37179
rect 15301 37145 15335 37179
rect 15335 37145 15344 37179
rect 15292 37136 15344 37145
rect 3608 37068 3660 37120
rect 18144 37136 18196 37188
rect 18604 37204 18656 37256
rect 20444 37204 20496 37256
rect 21824 37204 21876 37256
rect 21916 37204 21968 37256
rect 22468 37204 22520 37256
rect 24860 37247 24912 37256
rect 24860 37213 24869 37247
rect 24869 37213 24903 37247
rect 24903 37213 24912 37247
rect 24860 37204 24912 37213
rect 25228 37204 25280 37256
rect 26240 37204 26292 37256
rect 30288 37272 30340 37324
rect 31392 37272 31444 37324
rect 26700 37204 26752 37256
rect 29000 37204 29052 37256
rect 29920 37204 29972 37256
rect 31484 37247 31536 37256
rect 31484 37213 31493 37247
rect 31493 37213 31527 37247
rect 31527 37213 31536 37247
rect 31484 37204 31536 37213
rect 20352 37179 20404 37188
rect 20352 37145 20361 37179
rect 20361 37145 20395 37179
rect 20395 37145 20404 37179
rect 20352 37136 20404 37145
rect 22376 37136 22428 37188
rect 23572 37136 23624 37188
rect 24676 37179 24728 37188
rect 24676 37145 24685 37179
rect 24685 37145 24719 37179
rect 24719 37145 24728 37179
rect 24676 37136 24728 37145
rect 28816 37179 28868 37188
rect 28816 37145 28825 37179
rect 28825 37145 28859 37179
rect 28859 37145 28868 37179
rect 30564 37179 30616 37188
rect 28816 37136 28868 37145
rect 22468 37111 22520 37120
rect 22468 37077 22477 37111
rect 22477 37077 22511 37111
rect 22511 37077 22520 37111
rect 22468 37068 22520 37077
rect 24860 37068 24912 37120
rect 25504 37068 25556 37120
rect 30012 37068 30064 37120
rect 30196 37111 30248 37120
rect 30196 37077 30205 37111
rect 30205 37077 30239 37111
rect 30239 37077 30248 37111
rect 30196 37068 30248 37077
rect 30564 37145 30573 37179
rect 30573 37145 30607 37179
rect 30607 37145 30616 37179
rect 30564 37136 30616 37145
rect 31208 37136 31260 37188
rect 46848 37204 46900 37256
rect 47952 37247 48004 37256
rect 47952 37213 47961 37247
rect 47961 37213 47995 37247
rect 47995 37213 48004 37247
rect 47952 37204 48004 37213
rect 30932 37068 30984 37120
rect 46480 37068 46532 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 8944 36864 8996 36916
rect 1676 36796 1728 36848
rect 8300 36728 8352 36780
rect 9036 36728 9088 36780
rect 1676 36660 1728 36712
rect 1952 36660 2004 36712
rect 13360 36839 13412 36848
rect 13360 36805 13369 36839
rect 13369 36805 13403 36839
rect 13403 36805 13412 36839
rect 13360 36796 13412 36805
rect 15108 36864 15160 36916
rect 16488 36796 16540 36848
rect 18788 36796 18840 36848
rect 21732 36864 21784 36916
rect 22284 36864 22336 36916
rect 22376 36864 22428 36916
rect 24676 36907 24728 36916
rect 20444 36796 20496 36848
rect 24676 36873 24685 36907
rect 24685 36873 24719 36907
rect 24719 36873 24728 36907
rect 24676 36864 24728 36873
rect 26240 36907 26292 36916
rect 26240 36873 26249 36907
rect 26249 36873 26283 36907
rect 26283 36873 26292 36907
rect 26240 36864 26292 36873
rect 31944 36864 31996 36916
rect 14464 36771 14516 36780
rect 14464 36737 14498 36771
rect 14498 36737 14516 36771
rect 17224 36771 17276 36780
rect 14464 36728 14516 36737
rect 17224 36737 17233 36771
rect 17233 36737 17267 36771
rect 17267 36737 17276 36771
rect 17224 36728 17276 36737
rect 18604 36771 18656 36780
rect 18604 36737 18613 36771
rect 18613 36737 18647 36771
rect 18647 36737 18656 36771
rect 18604 36728 18656 36737
rect 21088 36728 21140 36780
rect 21916 36728 21968 36780
rect 11704 36703 11756 36712
rect 11704 36669 11713 36703
rect 11713 36669 11747 36703
rect 11747 36669 11756 36703
rect 11704 36660 11756 36669
rect 14096 36592 14148 36644
rect 2504 36524 2556 36576
rect 12716 36524 12768 36576
rect 13820 36524 13872 36576
rect 16856 36660 16908 36712
rect 17868 36660 17920 36712
rect 20352 36660 20404 36712
rect 22468 36728 22520 36780
rect 23020 36771 23072 36780
rect 23020 36737 23054 36771
rect 23054 36737 23072 36771
rect 23020 36728 23072 36737
rect 25872 36771 25924 36780
rect 22652 36660 22704 36712
rect 24308 36660 24360 36712
rect 22376 36592 22428 36644
rect 25872 36737 25881 36771
rect 25881 36737 25915 36771
rect 25915 36737 25924 36771
rect 25872 36728 25924 36737
rect 26056 36771 26108 36780
rect 26056 36737 26065 36771
rect 26065 36737 26099 36771
rect 26099 36737 26108 36771
rect 26056 36728 26108 36737
rect 26332 36728 26384 36780
rect 27804 36728 27856 36780
rect 25688 36660 25740 36712
rect 26700 36660 26752 36712
rect 26424 36592 26476 36644
rect 45836 36796 45888 36848
rect 46756 36796 46808 36848
rect 30932 36771 30984 36780
rect 30932 36737 30941 36771
rect 30941 36737 30975 36771
rect 30975 36737 30984 36771
rect 30932 36728 30984 36737
rect 30012 36703 30064 36712
rect 30012 36669 30021 36703
rect 30021 36669 30055 36703
rect 30055 36669 30064 36703
rect 30012 36660 30064 36669
rect 30288 36660 30340 36712
rect 31208 36592 31260 36644
rect 15200 36524 15252 36576
rect 24860 36524 24912 36576
rect 25964 36524 26016 36576
rect 28908 36524 28960 36576
rect 46848 36524 46900 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 11704 36320 11756 36372
rect 16488 36363 16540 36372
rect 2136 36184 2188 36236
rect 2504 36184 2556 36236
rect 3700 36116 3752 36168
rect 3792 36116 3844 36168
rect 16488 36329 16497 36363
rect 16497 36329 16531 36363
rect 16531 36329 16540 36363
rect 16488 36320 16540 36329
rect 18604 36363 18656 36372
rect 18604 36329 18613 36363
rect 18613 36329 18647 36363
rect 18647 36329 18656 36363
rect 18604 36320 18656 36329
rect 25872 36320 25924 36372
rect 26332 36363 26384 36372
rect 26332 36329 26341 36363
rect 26341 36329 26375 36363
rect 26375 36329 26384 36363
rect 26332 36320 26384 36329
rect 18144 36252 18196 36304
rect 24860 36252 24912 36304
rect 26148 36252 26200 36304
rect 19984 36184 20036 36236
rect 22652 36227 22704 36236
rect 22652 36193 22661 36227
rect 22661 36193 22695 36227
rect 22695 36193 22704 36227
rect 22652 36184 22704 36193
rect 25688 36227 25740 36236
rect 25688 36193 25697 36227
rect 25697 36193 25731 36227
rect 25731 36193 25740 36227
rect 25688 36184 25740 36193
rect 15200 36116 15252 36168
rect 15844 36048 15896 36100
rect 16028 36048 16080 36100
rect 3056 36023 3108 36032
rect 3056 35989 3065 36023
rect 3065 35989 3099 36023
rect 3099 35989 3108 36023
rect 3056 35980 3108 35989
rect 15016 35980 15068 36032
rect 17040 36048 17092 36100
rect 17408 36159 17460 36168
rect 17408 36125 17417 36159
rect 17417 36125 17451 36159
rect 17451 36125 17460 36159
rect 17408 36116 17460 36125
rect 17592 36159 17644 36168
rect 17592 36125 17601 36159
rect 17601 36125 17635 36159
rect 17635 36125 17644 36159
rect 17592 36116 17644 36125
rect 18144 36116 18196 36168
rect 19156 36116 19208 36168
rect 22192 36116 22244 36168
rect 23296 36116 23348 36168
rect 25504 36159 25556 36168
rect 18236 36048 18288 36100
rect 16948 36023 17000 36032
rect 16948 35989 16957 36023
rect 16957 35989 16991 36023
rect 16991 35989 17000 36023
rect 16948 35980 17000 35989
rect 19156 35980 19208 36032
rect 21732 36048 21784 36100
rect 21916 36091 21968 36100
rect 21916 36057 21925 36091
rect 21925 36057 21959 36091
rect 21959 36057 21968 36091
rect 21916 36048 21968 36057
rect 25504 36125 25513 36159
rect 25513 36125 25547 36159
rect 25547 36125 25556 36159
rect 25504 36116 25556 36125
rect 25780 36116 25832 36168
rect 26240 36116 26292 36168
rect 21272 35980 21324 36032
rect 26056 36048 26108 36100
rect 26792 36159 26844 36168
rect 26792 36125 26801 36159
rect 26801 36125 26835 36159
rect 26835 36125 26844 36159
rect 26792 36116 26844 36125
rect 31116 36159 31168 36168
rect 31116 36125 31125 36159
rect 31125 36125 31159 36159
rect 31159 36125 31168 36159
rect 31116 36116 31168 36125
rect 31300 36252 31352 36304
rect 31852 36184 31904 36236
rect 47952 36252 48004 36304
rect 46480 36227 46532 36236
rect 46480 36193 46489 36227
rect 46489 36193 46523 36227
rect 46523 36193 46532 36227
rect 46480 36184 46532 36193
rect 48136 36227 48188 36236
rect 48136 36193 48145 36227
rect 48145 36193 48179 36227
rect 48179 36193 48188 36227
rect 48136 36184 48188 36193
rect 27160 36048 27212 36100
rect 27436 36048 27488 36100
rect 29184 36048 29236 36100
rect 29736 36048 29788 36100
rect 31576 36116 31628 36168
rect 31668 36048 31720 36100
rect 27896 35980 27948 36032
rect 32036 35980 32088 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 9036 35819 9088 35828
rect 9036 35785 9045 35819
rect 9045 35785 9079 35819
rect 9079 35785 9088 35819
rect 9036 35776 9088 35785
rect 15292 35776 15344 35828
rect 3056 35708 3108 35760
rect 3700 35708 3752 35760
rect 12072 35708 12124 35760
rect 16488 35708 16540 35760
rect 16948 35708 17000 35760
rect 17960 35776 18012 35828
rect 19248 35776 19300 35828
rect 21088 35776 21140 35828
rect 20260 35708 20312 35760
rect 21732 35776 21784 35828
rect 23020 35776 23072 35828
rect 2044 35683 2096 35692
rect 2044 35649 2053 35683
rect 2053 35649 2087 35683
rect 2087 35649 2096 35683
rect 2044 35640 2096 35649
rect 9404 35640 9456 35692
rect 14832 35640 14884 35692
rect 16764 35640 16816 35692
rect 19248 35683 19300 35692
rect 19248 35649 19257 35683
rect 19257 35649 19291 35683
rect 19291 35649 19300 35683
rect 19248 35640 19300 35649
rect 20628 35640 20680 35692
rect 20996 35683 21048 35692
rect 20996 35649 21005 35683
rect 21005 35649 21039 35683
rect 21039 35649 21048 35683
rect 20996 35640 21048 35649
rect 2780 35615 2832 35624
rect 2780 35581 2789 35615
rect 2789 35581 2823 35615
rect 2823 35581 2832 35615
rect 2780 35572 2832 35581
rect 16028 35572 16080 35624
rect 20720 35572 20772 35624
rect 22284 35708 22336 35760
rect 21548 35640 21600 35692
rect 21732 35572 21784 35624
rect 23296 35683 23348 35692
rect 23296 35649 23305 35683
rect 23305 35649 23339 35683
rect 23339 35649 23348 35683
rect 23296 35640 23348 35649
rect 23388 35683 23440 35692
rect 23388 35649 23397 35683
rect 23397 35649 23431 35683
rect 23431 35649 23440 35683
rect 24860 35776 24912 35828
rect 25412 35776 25464 35828
rect 28356 35819 28408 35828
rect 28356 35785 28365 35819
rect 28365 35785 28399 35819
rect 28399 35785 28408 35819
rect 28356 35776 28408 35785
rect 29000 35776 29052 35828
rect 23388 35640 23440 35649
rect 24032 35683 24084 35692
rect 24032 35649 24041 35683
rect 24041 35649 24075 35683
rect 24075 35649 24084 35683
rect 24032 35640 24084 35649
rect 24308 35683 24360 35692
rect 23756 35572 23808 35624
rect 24308 35649 24317 35683
rect 24317 35649 24351 35683
rect 24351 35649 24360 35683
rect 28908 35708 28960 35760
rect 32864 35776 32916 35828
rect 31852 35708 31904 35760
rect 32036 35708 32088 35760
rect 24308 35640 24360 35649
rect 25596 35640 25648 35692
rect 25044 35572 25096 35624
rect 25688 35615 25740 35624
rect 25688 35581 25697 35615
rect 25697 35581 25731 35615
rect 25731 35581 25740 35615
rect 25688 35572 25740 35581
rect 26332 35683 26384 35692
rect 26332 35649 26341 35683
rect 26341 35649 26375 35683
rect 26375 35649 26384 35683
rect 26332 35640 26384 35649
rect 27712 35640 27764 35692
rect 28724 35640 28776 35692
rect 28356 35572 28408 35624
rect 28816 35572 28868 35624
rect 1952 35436 2004 35488
rect 16304 35436 16356 35488
rect 22284 35504 22336 35556
rect 34796 35640 34848 35692
rect 45928 35640 45980 35692
rect 46664 35640 46716 35692
rect 47860 35683 47912 35692
rect 47860 35649 47869 35683
rect 47869 35649 47903 35683
rect 47903 35649 47912 35683
rect 47860 35640 47912 35649
rect 20628 35479 20680 35488
rect 20628 35445 20637 35479
rect 20637 35445 20671 35479
rect 20671 35445 20680 35479
rect 20628 35436 20680 35445
rect 23572 35436 23624 35488
rect 24492 35479 24544 35488
rect 24492 35445 24501 35479
rect 24501 35445 24535 35479
rect 24535 35445 24544 35479
rect 24492 35436 24544 35445
rect 24584 35436 24636 35488
rect 29184 35436 29236 35488
rect 29276 35436 29328 35488
rect 30288 35504 30340 35556
rect 31484 35436 31536 35488
rect 32496 35436 32548 35488
rect 32864 35436 32916 35488
rect 46940 35479 46992 35488
rect 46940 35445 46949 35479
rect 46949 35445 46983 35479
rect 46983 35445 46992 35479
rect 46940 35436 46992 35445
rect 47584 35436 47636 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 1952 35275 2004 35284
rect 1952 35241 1961 35275
rect 1961 35241 1995 35275
rect 1995 35241 2004 35275
rect 1952 35232 2004 35241
rect 15844 35275 15896 35284
rect 15844 35241 15853 35275
rect 15853 35241 15887 35275
rect 15887 35241 15896 35275
rect 15844 35232 15896 35241
rect 17408 35232 17460 35284
rect 11520 35096 11572 35148
rect 12164 35071 12216 35080
rect 12164 35037 12173 35071
rect 12173 35037 12207 35071
rect 12207 35037 12216 35071
rect 12164 35028 12216 35037
rect 1860 35003 1912 35012
rect 1860 34969 1869 35003
rect 1869 34969 1903 35003
rect 1903 34969 1912 35003
rect 1860 34960 1912 34969
rect 12256 34960 12308 35012
rect 15108 34960 15160 35012
rect 14188 34892 14240 34944
rect 16304 35071 16356 35080
rect 16304 35037 16313 35071
rect 16313 35037 16347 35071
rect 16347 35037 16356 35071
rect 16304 35028 16356 35037
rect 16764 35028 16816 35080
rect 17960 35028 18012 35080
rect 17592 34960 17644 35012
rect 17040 34892 17092 34944
rect 19984 35096 20036 35148
rect 20444 35232 20496 35284
rect 45928 35232 45980 35284
rect 27620 35207 27672 35216
rect 18420 35028 18472 35080
rect 19156 35028 19208 35080
rect 20628 35028 20680 35080
rect 27620 35173 27629 35207
rect 27629 35173 27663 35207
rect 27663 35173 27672 35207
rect 27620 35164 27672 35173
rect 28816 35164 28868 35216
rect 30288 35164 30340 35216
rect 22560 35139 22612 35148
rect 22560 35105 22569 35139
rect 22569 35105 22603 35139
rect 22603 35105 22612 35139
rect 22560 35096 22612 35105
rect 24584 35096 24636 35148
rect 31024 35164 31076 35216
rect 19248 34892 19300 34944
rect 20812 34892 20864 34944
rect 23296 35028 23348 35080
rect 23940 34960 23992 35012
rect 25596 35003 25648 35012
rect 25596 34969 25605 35003
rect 25605 34969 25639 35003
rect 25639 34969 25648 35003
rect 25596 34960 25648 34969
rect 26792 35028 26844 35080
rect 28356 35028 28408 35080
rect 29736 35028 29788 35080
rect 30748 35028 30800 35080
rect 31576 35164 31628 35216
rect 31668 35096 31720 35148
rect 27252 35003 27304 35012
rect 27252 34969 27261 35003
rect 27261 34969 27295 35003
rect 27295 34969 27304 35003
rect 27252 34960 27304 34969
rect 27344 34960 27396 35012
rect 27896 34960 27948 35012
rect 28724 34960 28776 35012
rect 28908 34960 28960 35012
rect 31576 35003 31628 35012
rect 31576 34969 31585 35003
rect 31585 34969 31619 35003
rect 31619 34969 31628 35003
rect 31576 34960 31628 34969
rect 31668 34960 31720 35012
rect 32496 35028 32548 35080
rect 33048 35003 33100 35012
rect 33048 34969 33082 35003
rect 33082 34969 33100 35003
rect 33048 34960 33100 34969
rect 47676 34960 47728 35012
rect 48136 35003 48188 35012
rect 48136 34969 48145 35003
rect 48145 34969 48179 35003
rect 48179 34969 48188 35003
rect 48136 34960 48188 34969
rect 22284 34892 22336 34944
rect 22928 34892 22980 34944
rect 23204 34935 23256 34944
rect 23204 34901 23213 34935
rect 23213 34901 23247 34935
rect 23247 34901 23256 34935
rect 23204 34892 23256 34901
rect 24400 34892 24452 34944
rect 25688 34935 25740 34944
rect 25688 34901 25697 34935
rect 25697 34901 25731 34935
rect 25731 34901 25740 34935
rect 25688 34892 25740 34901
rect 26700 34935 26752 34944
rect 26700 34901 26709 34935
rect 26709 34901 26743 34935
rect 26743 34901 26752 34935
rect 26700 34892 26752 34901
rect 29828 34935 29880 34944
rect 29828 34901 29837 34935
rect 29837 34901 29871 34935
rect 29871 34901 29880 34935
rect 29828 34892 29880 34901
rect 30196 34935 30248 34944
rect 30196 34901 30205 34935
rect 30205 34901 30239 34935
rect 30239 34901 30248 34935
rect 30196 34892 30248 34901
rect 34244 34892 34296 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 12256 34688 12308 34740
rect 12532 34688 12584 34740
rect 2044 34595 2096 34604
rect 2044 34561 2053 34595
rect 2053 34561 2087 34595
rect 2087 34561 2096 34595
rect 2044 34552 2096 34561
rect 2504 34552 2556 34604
rect 18972 34620 19024 34672
rect 21732 34688 21784 34740
rect 27252 34688 27304 34740
rect 29276 34688 29328 34740
rect 23848 34620 23900 34672
rect 30012 34688 30064 34740
rect 41052 34688 41104 34740
rect 47676 34731 47728 34740
rect 1860 34484 1912 34536
rect 12992 34552 13044 34604
rect 13636 34595 13688 34604
rect 13636 34561 13645 34595
rect 13645 34561 13679 34595
rect 13679 34561 13688 34595
rect 13636 34552 13688 34561
rect 13820 34595 13872 34604
rect 13820 34561 13829 34595
rect 13829 34561 13863 34595
rect 13863 34561 13872 34595
rect 13820 34552 13872 34561
rect 14464 34595 14516 34604
rect 14464 34561 14473 34595
rect 14473 34561 14507 34595
rect 14507 34561 14516 34595
rect 14464 34552 14516 34561
rect 14648 34595 14700 34604
rect 14648 34561 14657 34595
rect 14657 34561 14691 34595
rect 14691 34561 14700 34595
rect 14648 34552 14700 34561
rect 12900 34484 12952 34536
rect 13912 34484 13964 34536
rect 14188 34484 14240 34536
rect 17040 34595 17092 34604
rect 17040 34561 17046 34595
rect 17046 34561 17080 34595
rect 17080 34561 17092 34595
rect 17040 34552 17092 34561
rect 17224 34552 17276 34604
rect 17960 34595 18012 34604
rect 16028 34527 16080 34536
rect 16028 34493 16037 34527
rect 16037 34493 16071 34527
rect 16071 34493 16080 34527
rect 16028 34484 16080 34493
rect 17960 34561 17969 34595
rect 17969 34561 18003 34595
rect 18003 34561 18012 34595
rect 17960 34552 18012 34561
rect 20812 34595 20864 34604
rect 20812 34561 20821 34595
rect 20821 34561 20855 34595
rect 20855 34561 20864 34595
rect 20812 34552 20864 34561
rect 21180 34595 21232 34604
rect 21180 34561 21189 34595
rect 21189 34561 21223 34595
rect 21223 34561 21232 34595
rect 21180 34552 21232 34561
rect 21640 34552 21692 34604
rect 22192 34595 22244 34604
rect 22192 34561 22201 34595
rect 22201 34561 22235 34595
rect 22235 34561 22244 34595
rect 22192 34552 22244 34561
rect 22284 34595 22336 34604
rect 22284 34561 22293 34595
rect 22293 34561 22327 34595
rect 22327 34561 22336 34595
rect 22284 34552 22336 34561
rect 17592 34484 17644 34536
rect 19708 34484 19760 34536
rect 21088 34484 21140 34536
rect 12440 34416 12492 34468
rect 1400 34348 1452 34400
rect 2136 34391 2188 34400
rect 2136 34357 2145 34391
rect 2145 34357 2179 34391
rect 2179 34357 2188 34391
rect 2136 34348 2188 34357
rect 8484 34348 8536 34400
rect 15660 34348 15712 34400
rect 17316 34348 17368 34400
rect 23020 34391 23072 34400
rect 23020 34357 23029 34391
rect 23029 34357 23063 34391
rect 23063 34357 23072 34391
rect 23020 34348 23072 34357
rect 23572 34552 23624 34604
rect 24216 34595 24268 34604
rect 24216 34561 24225 34595
rect 24225 34561 24259 34595
rect 24259 34561 24268 34595
rect 24216 34552 24268 34561
rect 24584 34552 24636 34604
rect 23480 34527 23532 34536
rect 23480 34493 23489 34527
rect 23489 34493 23523 34527
rect 23523 34493 23532 34527
rect 23480 34484 23532 34493
rect 25044 34595 25096 34604
rect 25044 34561 25053 34595
rect 25053 34561 25087 34595
rect 25087 34561 25096 34595
rect 25044 34552 25096 34561
rect 24400 34416 24452 34468
rect 24860 34484 24912 34536
rect 29828 34620 29880 34672
rect 30932 34620 30984 34672
rect 25964 34595 26016 34604
rect 25964 34561 25973 34595
rect 25973 34561 26007 34595
rect 26007 34561 26016 34595
rect 25964 34552 26016 34561
rect 26424 34552 26476 34604
rect 28908 34552 28960 34604
rect 30104 34552 30156 34604
rect 47400 34620 47452 34672
rect 47676 34697 47685 34731
rect 47685 34697 47719 34731
rect 47719 34697 47728 34731
rect 47676 34688 47728 34697
rect 47860 34552 47912 34604
rect 25872 34416 25924 34468
rect 29920 34484 29972 34536
rect 46388 34484 46440 34536
rect 24308 34391 24360 34400
rect 24308 34357 24317 34391
rect 24317 34357 24351 34391
rect 24351 34357 24360 34391
rect 24308 34348 24360 34357
rect 24492 34348 24544 34400
rect 25504 34348 25556 34400
rect 26148 34391 26200 34400
rect 26148 34357 26157 34391
rect 26157 34357 26191 34391
rect 26191 34357 26200 34391
rect 26148 34348 26200 34357
rect 26424 34391 26476 34400
rect 26424 34357 26433 34391
rect 26433 34357 26467 34391
rect 26467 34357 26476 34391
rect 26424 34348 26476 34357
rect 28448 34416 28500 34468
rect 29276 34348 29328 34400
rect 30840 34348 30892 34400
rect 46848 34348 46900 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 8300 34076 8352 34128
rect 12164 34144 12216 34196
rect 1400 34051 1452 34060
rect 1400 34017 1409 34051
rect 1409 34017 1443 34051
rect 1443 34017 1452 34051
rect 1400 34008 1452 34017
rect 2136 34008 2188 34060
rect 2780 34051 2832 34060
rect 2780 34017 2789 34051
rect 2789 34017 2823 34051
rect 2823 34017 2832 34051
rect 2780 34008 2832 34017
rect 10232 34008 10284 34060
rect 9220 33940 9272 33992
rect 10324 33872 10376 33924
rect 10876 33940 10928 33992
rect 14648 34144 14700 34196
rect 21272 34144 21324 34196
rect 21824 34144 21876 34196
rect 22008 34144 22060 34196
rect 23480 34144 23532 34196
rect 24584 34144 24636 34196
rect 24860 34144 24912 34196
rect 25044 34187 25096 34196
rect 25044 34153 25053 34187
rect 25053 34153 25087 34187
rect 25087 34153 25096 34187
rect 25044 34144 25096 34153
rect 26608 34187 26660 34196
rect 26608 34153 26617 34187
rect 26617 34153 26651 34187
rect 26651 34153 26660 34187
rect 26608 34144 26660 34153
rect 23848 34076 23900 34128
rect 27068 34119 27120 34128
rect 27068 34085 27077 34119
rect 27077 34085 27111 34119
rect 27111 34085 27120 34119
rect 27068 34076 27120 34085
rect 12992 34051 13044 34060
rect 12992 34017 13001 34051
rect 13001 34017 13035 34051
rect 13035 34017 13044 34051
rect 12992 34008 13044 34017
rect 14188 34051 14240 34060
rect 14188 34017 14197 34051
rect 14197 34017 14231 34051
rect 14231 34017 14240 34051
rect 14188 34008 14240 34017
rect 13820 33940 13872 33992
rect 15108 34008 15160 34060
rect 16028 34008 16080 34060
rect 17316 34051 17368 34060
rect 17316 34017 17325 34051
rect 17325 34017 17359 34051
rect 17359 34017 17368 34051
rect 17316 34008 17368 34017
rect 20352 34008 20404 34060
rect 26056 34008 26108 34060
rect 27436 34008 27488 34060
rect 28448 34051 28500 34060
rect 28448 34017 28457 34051
rect 28457 34017 28491 34051
rect 28491 34017 28500 34051
rect 28448 34008 28500 34017
rect 29000 34008 29052 34060
rect 30288 34008 30340 34060
rect 37648 34051 37700 34060
rect 37648 34017 37657 34051
rect 37657 34017 37691 34051
rect 37691 34017 37700 34051
rect 37648 34008 37700 34017
rect 46756 34076 46808 34128
rect 46940 34008 46992 34060
rect 48228 34008 48280 34060
rect 10784 33804 10836 33856
rect 15384 33940 15436 33992
rect 19708 33983 19760 33992
rect 19708 33949 19717 33983
rect 19717 33949 19751 33983
rect 19751 33949 19760 33983
rect 19708 33940 19760 33949
rect 20628 33940 20680 33992
rect 23020 33940 23072 33992
rect 24768 33983 24820 33992
rect 24768 33949 24777 33983
rect 24777 33949 24811 33983
rect 24811 33949 24820 33983
rect 24768 33940 24820 33949
rect 25044 33940 25096 33992
rect 25504 33983 25556 33992
rect 25504 33949 25513 33983
rect 25513 33949 25547 33983
rect 25547 33949 25556 33983
rect 25504 33940 25556 33949
rect 25872 33983 25924 33992
rect 25872 33949 25881 33983
rect 25881 33949 25915 33983
rect 25915 33949 25924 33983
rect 25872 33940 25924 33949
rect 26424 33940 26476 33992
rect 26884 33983 26936 33992
rect 26884 33949 26893 33983
rect 26893 33949 26927 33983
rect 26927 33949 26936 33983
rect 26884 33940 26936 33949
rect 29828 33940 29880 33992
rect 30748 33983 30800 33992
rect 30748 33949 30757 33983
rect 30757 33949 30791 33983
rect 30791 33949 30800 33983
rect 30748 33940 30800 33949
rect 22928 33915 22980 33924
rect 22928 33881 22937 33915
rect 22937 33881 22971 33915
rect 22971 33881 22980 33915
rect 22928 33872 22980 33881
rect 25780 33872 25832 33924
rect 28356 33915 28408 33924
rect 28356 33881 28365 33915
rect 28365 33881 28399 33915
rect 28399 33881 28408 33915
rect 28356 33872 28408 33881
rect 30012 33915 30064 33924
rect 30012 33881 30021 33915
rect 30021 33881 30055 33915
rect 30055 33881 30064 33915
rect 35992 33915 36044 33924
rect 30012 33872 30064 33881
rect 35992 33881 36001 33915
rect 36001 33881 36035 33915
rect 36035 33881 36044 33915
rect 35992 33872 36044 33881
rect 18604 33847 18656 33856
rect 18604 33813 18613 33847
rect 18613 33813 18647 33847
rect 18647 33813 18656 33847
rect 18604 33804 18656 33813
rect 22468 33804 22520 33856
rect 25596 33847 25648 33856
rect 25596 33813 25605 33847
rect 25605 33813 25639 33847
rect 25639 33813 25648 33847
rect 25596 33804 25648 33813
rect 27528 33804 27580 33856
rect 30564 33804 30616 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 10324 33643 10376 33652
rect 10324 33609 10333 33643
rect 10333 33609 10367 33643
rect 10367 33609 10376 33643
rect 10324 33600 10376 33609
rect 10232 33532 10284 33584
rect 11244 33532 11296 33584
rect 1860 33507 1912 33516
rect 1860 33473 1869 33507
rect 1869 33473 1903 33507
rect 1903 33473 1912 33507
rect 1860 33464 1912 33473
rect 8300 33464 8352 33516
rect 2780 33439 2832 33448
rect 2780 33405 2789 33439
rect 2789 33405 2823 33439
rect 2823 33405 2832 33439
rect 2780 33396 2832 33405
rect 10508 33464 10560 33516
rect 10692 33507 10744 33516
rect 10692 33473 10701 33507
rect 10701 33473 10735 33507
rect 10735 33473 10744 33507
rect 10692 33464 10744 33473
rect 10784 33507 10836 33516
rect 10784 33473 10798 33507
rect 10798 33473 10832 33507
rect 10832 33473 10836 33507
rect 10968 33507 11020 33516
rect 10784 33464 10836 33473
rect 10968 33473 10977 33507
rect 10977 33473 11011 33507
rect 11011 33473 11020 33507
rect 10968 33464 11020 33473
rect 11980 33464 12032 33516
rect 12808 33600 12860 33652
rect 12900 33600 12952 33652
rect 17224 33600 17276 33652
rect 26608 33600 26660 33652
rect 27252 33600 27304 33652
rect 27804 33600 27856 33652
rect 29828 33600 29880 33652
rect 30104 33600 30156 33652
rect 32956 33600 33008 33652
rect 35992 33600 36044 33652
rect 46388 33600 46440 33652
rect 12164 33532 12216 33584
rect 12348 33464 12400 33516
rect 13084 33464 13136 33516
rect 16028 33532 16080 33584
rect 18972 33575 19024 33584
rect 18972 33541 18981 33575
rect 18981 33541 19015 33575
rect 19015 33541 19024 33575
rect 18972 33532 19024 33541
rect 22192 33575 22244 33584
rect 22192 33541 22201 33575
rect 22201 33541 22235 33575
rect 22235 33541 22244 33575
rect 22192 33532 22244 33541
rect 14556 33507 14608 33516
rect 14556 33473 14590 33507
rect 14590 33473 14608 33507
rect 14556 33464 14608 33473
rect 16764 33464 16816 33516
rect 18604 33464 18656 33516
rect 19984 33464 20036 33516
rect 20444 33464 20496 33516
rect 21640 33464 21692 33516
rect 12256 33439 12308 33448
rect 12256 33405 12265 33439
rect 12265 33405 12299 33439
rect 12299 33405 12308 33439
rect 12992 33439 13044 33448
rect 12256 33396 12308 33405
rect 12992 33405 13001 33439
rect 13001 33405 13035 33439
rect 13035 33405 13044 33439
rect 12992 33396 13044 33405
rect 13820 33396 13872 33448
rect 22652 33464 22704 33516
rect 26332 33532 26384 33584
rect 26884 33532 26936 33584
rect 27528 33575 27580 33584
rect 27528 33541 27537 33575
rect 27537 33541 27571 33575
rect 27571 33541 27580 33575
rect 27528 33532 27580 33541
rect 30564 33532 30616 33584
rect 24216 33396 24268 33448
rect 23848 33371 23900 33380
rect 23848 33337 23857 33371
rect 23857 33337 23891 33371
rect 23891 33337 23900 33371
rect 23848 33328 23900 33337
rect 26056 33328 26108 33380
rect 27344 33396 27396 33448
rect 27528 33396 27580 33448
rect 28448 33464 28500 33516
rect 30656 33507 30708 33516
rect 30656 33473 30665 33507
rect 30665 33473 30699 33507
rect 30699 33473 30708 33507
rect 30656 33464 30708 33473
rect 30840 33507 30892 33516
rect 30840 33473 30849 33507
rect 30849 33473 30883 33507
rect 30883 33473 30892 33507
rect 30840 33464 30892 33473
rect 31024 33507 31076 33516
rect 31024 33473 31033 33507
rect 31033 33473 31067 33507
rect 31067 33473 31076 33507
rect 31024 33464 31076 33473
rect 33048 33464 33100 33516
rect 35900 33464 35952 33516
rect 46664 33464 46716 33516
rect 47952 33507 48004 33516
rect 47952 33473 47961 33507
rect 47961 33473 47995 33507
rect 47995 33473 48004 33507
rect 47952 33464 48004 33473
rect 26608 33328 26660 33380
rect 28264 33328 28316 33380
rect 32312 33396 32364 33448
rect 32496 33439 32548 33448
rect 32496 33405 32505 33439
rect 32505 33405 32539 33439
rect 32539 33405 32548 33439
rect 32496 33396 32548 33405
rect 2780 33260 2832 33312
rect 9772 33303 9824 33312
rect 9772 33269 9781 33303
rect 9781 33269 9815 33303
rect 9815 33269 9824 33303
rect 9772 33260 9824 33269
rect 10876 33260 10928 33312
rect 12808 33303 12860 33312
rect 12808 33269 12817 33303
rect 12817 33269 12851 33303
rect 12851 33269 12860 33303
rect 12808 33260 12860 33269
rect 13636 33260 13688 33312
rect 14280 33260 14332 33312
rect 15384 33260 15436 33312
rect 18880 33260 18932 33312
rect 19064 33260 19116 33312
rect 20996 33260 21048 33312
rect 26240 33260 26292 33312
rect 26516 33260 26568 33312
rect 28172 33260 28224 33312
rect 30380 33303 30432 33312
rect 30380 33269 30389 33303
rect 30389 33269 30423 33303
rect 30423 33269 30432 33303
rect 30380 33260 30432 33269
rect 46940 33260 46992 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 2780 33099 2832 33108
rect 2780 33065 2789 33099
rect 2789 33065 2823 33099
rect 2823 33065 2832 33099
rect 2780 33056 2832 33065
rect 10232 33056 10284 33108
rect 11244 33099 11296 33108
rect 11244 33065 11253 33099
rect 11253 33065 11287 33099
rect 11287 33065 11296 33099
rect 11244 33056 11296 33065
rect 12164 33056 12216 33108
rect 12532 33056 12584 33108
rect 20444 33099 20496 33108
rect 20444 33065 20453 33099
rect 20453 33065 20487 33099
rect 20487 33065 20496 33099
rect 20444 33056 20496 33065
rect 12348 32988 12400 33040
rect 13728 32988 13780 33040
rect 19984 32988 20036 33040
rect 20628 32988 20680 33040
rect 2044 32852 2096 32904
rect 2688 32895 2740 32904
rect 2688 32861 2697 32895
rect 2697 32861 2731 32895
rect 2731 32861 2740 32895
rect 2688 32852 2740 32861
rect 11060 32920 11112 32972
rect 12440 32920 12492 32972
rect 13176 32852 13228 32904
rect 13544 32852 13596 32904
rect 14188 32852 14240 32904
rect 14740 32852 14792 32904
rect 15384 32852 15436 32904
rect 20809 32895 20861 32904
rect 20809 32861 20836 32895
rect 20836 32861 20861 32895
rect 10784 32784 10836 32836
rect 12256 32784 12308 32836
rect 13084 32784 13136 32836
rect 7656 32716 7708 32768
rect 18328 32784 18380 32836
rect 13728 32716 13780 32768
rect 18880 32716 18932 32768
rect 19432 32716 19484 32768
rect 20809 32852 20861 32861
rect 20996 32920 21048 32972
rect 22008 32852 22060 32904
rect 28448 33056 28500 33108
rect 30656 33056 30708 33108
rect 30932 33056 30984 33108
rect 31024 33056 31076 33108
rect 32404 33056 32456 33108
rect 33048 33099 33100 33108
rect 33048 33065 33057 33099
rect 33057 33065 33091 33099
rect 33091 33065 33100 33099
rect 33048 33056 33100 33065
rect 47400 33056 47452 33108
rect 27528 32988 27580 33040
rect 26792 32852 26844 32904
rect 22284 32784 22336 32836
rect 28172 32895 28224 32904
rect 28172 32861 28181 32895
rect 28181 32861 28215 32895
rect 28215 32861 28224 32895
rect 28172 32852 28224 32861
rect 28264 32895 28316 32904
rect 28632 32988 28684 33040
rect 30288 32963 30340 32972
rect 30288 32929 30297 32963
rect 30297 32929 30331 32963
rect 30331 32929 30340 32963
rect 30288 32920 30340 32929
rect 30564 32920 30616 32972
rect 28264 32861 28278 32895
rect 28278 32861 28312 32895
rect 28312 32861 28316 32895
rect 28264 32852 28316 32861
rect 30104 32895 30156 32904
rect 30104 32861 30113 32895
rect 30113 32861 30147 32895
rect 30147 32861 30156 32895
rect 30104 32852 30156 32861
rect 30196 32852 30248 32904
rect 30380 32852 30432 32904
rect 33324 32895 33376 32904
rect 33324 32861 33333 32895
rect 33333 32861 33367 32895
rect 33367 32861 33376 32895
rect 33324 32852 33376 32861
rect 21732 32716 21784 32768
rect 22100 32716 22152 32768
rect 27160 32784 27212 32836
rect 23572 32759 23624 32768
rect 23572 32725 23581 32759
rect 23581 32725 23615 32759
rect 23615 32725 23624 32759
rect 23572 32716 23624 32725
rect 25044 32716 25096 32768
rect 29736 32759 29788 32768
rect 29736 32725 29745 32759
rect 29745 32725 29779 32759
rect 29779 32725 29788 32759
rect 29736 32716 29788 32725
rect 32312 32784 32364 32836
rect 33508 32895 33560 32904
rect 33508 32861 33517 32895
rect 33517 32861 33551 32895
rect 33551 32861 33560 32895
rect 33508 32852 33560 32861
rect 32588 32759 32640 32768
rect 32588 32725 32597 32759
rect 32597 32725 32631 32759
rect 32631 32725 32640 32759
rect 32588 32716 32640 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 12992 32512 13044 32564
rect 14556 32512 14608 32564
rect 17960 32512 18012 32564
rect 2044 32419 2096 32428
rect 2044 32385 2053 32419
rect 2053 32385 2087 32419
rect 2087 32385 2096 32419
rect 2044 32376 2096 32385
rect 10324 32376 10376 32428
rect 10692 32444 10744 32496
rect 12164 32444 12216 32496
rect 13544 32444 13596 32496
rect 10600 32419 10652 32428
rect 10600 32385 10614 32419
rect 10614 32385 10648 32419
rect 10648 32385 10652 32419
rect 10600 32376 10652 32385
rect 10968 32376 11020 32428
rect 11796 32376 11848 32428
rect 12256 32419 12308 32428
rect 2780 32308 2832 32360
rect 2872 32351 2924 32360
rect 2872 32317 2881 32351
rect 2881 32317 2915 32351
rect 2915 32317 2924 32351
rect 12256 32385 12265 32419
rect 12265 32385 12299 32419
rect 12299 32385 12308 32419
rect 12256 32376 12308 32385
rect 13084 32419 13136 32428
rect 13084 32385 13093 32419
rect 13093 32385 13127 32419
rect 13127 32385 13136 32419
rect 13084 32376 13136 32385
rect 13820 32376 13872 32428
rect 2872 32308 2924 32317
rect 13544 32308 13596 32360
rect 13636 32308 13688 32360
rect 11612 32240 11664 32292
rect 12992 32240 13044 32292
rect 14280 32240 14332 32292
rect 8300 32172 8352 32224
rect 10232 32172 10284 32224
rect 11060 32172 11112 32224
rect 12808 32172 12860 32224
rect 13176 32172 13228 32224
rect 14740 32376 14792 32428
rect 15108 32419 15160 32428
rect 15108 32385 15117 32419
rect 15117 32385 15151 32419
rect 15151 32385 15160 32419
rect 15108 32376 15160 32385
rect 16028 32376 16080 32428
rect 17224 32419 17276 32428
rect 17224 32385 17258 32419
rect 17258 32385 17276 32419
rect 17224 32376 17276 32385
rect 15108 32172 15160 32224
rect 18696 32172 18748 32224
rect 23848 32444 23900 32496
rect 20168 32376 20220 32428
rect 20352 32376 20404 32428
rect 22008 32419 22060 32428
rect 22008 32385 22017 32419
rect 22017 32385 22051 32419
rect 22051 32385 22060 32419
rect 22008 32376 22060 32385
rect 23112 32376 23164 32428
rect 24860 32512 24912 32564
rect 25412 32555 25464 32564
rect 25412 32521 25421 32555
rect 25421 32521 25455 32555
rect 25455 32521 25464 32555
rect 25412 32512 25464 32521
rect 24308 32444 24360 32496
rect 33508 32512 33560 32564
rect 25964 32376 26016 32428
rect 27528 32376 27580 32428
rect 29184 32444 29236 32496
rect 29736 32444 29788 32496
rect 29920 32376 29972 32428
rect 30012 32376 30064 32428
rect 24032 32308 24084 32360
rect 24768 32240 24820 32292
rect 26148 32308 26200 32360
rect 29000 32308 29052 32360
rect 30288 32351 30340 32360
rect 30288 32317 30297 32351
rect 30297 32317 30331 32351
rect 30331 32317 30340 32351
rect 30656 32376 30708 32428
rect 32496 32376 32548 32428
rect 32772 32376 32824 32428
rect 33324 32376 33376 32428
rect 33876 32376 33928 32428
rect 47676 32419 47728 32428
rect 47676 32385 47685 32419
rect 47685 32385 47719 32419
rect 47719 32385 47728 32419
rect 47676 32376 47728 32385
rect 30288 32308 30340 32317
rect 29184 32240 29236 32292
rect 30656 32240 30708 32292
rect 20352 32172 20404 32224
rect 21364 32172 21416 32224
rect 23388 32172 23440 32224
rect 23480 32172 23532 32224
rect 24492 32172 24544 32224
rect 28540 32172 28592 32224
rect 30472 32172 30524 32224
rect 46848 32308 46900 32360
rect 34060 32215 34112 32224
rect 34060 32181 34069 32215
rect 34069 32181 34103 32215
rect 34103 32181 34112 32215
rect 34060 32172 34112 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 2780 31968 2832 32020
rect 10600 31968 10652 32020
rect 10508 31900 10560 31952
rect 12532 31968 12584 32020
rect 17224 31968 17276 32020
rect 17316 31968 17368 32020
rect 11520 31943 11572 31952
rect 1860 31807 1912 31816
rect 1860 31773 1869 31807
rect 1869 31773 1903 31807
rect 1903 31773 1912 31807
rect 1860 31764 1912 31773
rect 2044 31807 2096 31816
rect 2044 31773 2053 31807
rect 2053 31773 2087 31807
rect 2087 31773 2096 31807
rect 2044 31764 2096 31773
rect 7656 31764 7708 31816
rect 9680 31807 9732 31816
rect 9680 31773 9689 31807
rect 9689 31773 9723 31807
rect 9723 31773 9732 31807
rect 9680 31764 9732 31773
rect 10232 31764 10284 31816
rect 11520 31909 11529 31943
rect 11529 31909 11563 31943
rect 11563 31909 11572 31943
rect 11520 31900 11572 31909
rect 11704 31900 11756 31952
rect 12900 31900 12952 31952
rect 12992 31900 13044 31952
rect 12440 31832 12492 31884
rect 10876 31764 10928 31816
rect 10968 31807 11020 31816
rect 10968 31773 10977 31807
rect 10977 31773 11011 31807
rect 11011 31773 11020 31807
rect 10968 31764 11020 31773
rect 11704 31764 11756 31816
rect 11796 31807 11848 31816
rect 11796 31773 11805 31807
rect 11805 31773 11839 31807
rect 11839 31773 11848 31807
rect 12532 31807 12584 31816
rect 11796 31764 11848 31773
rect 12532 31773 12541 31807
rect 12541 31773 12575 31807
rect 12575 31773 12584 31807
rect 12532 31764 12584 31773
rect 15292 31900 15344 31952
rect 18328 31943 18380 31952
rect 18328 31909 18337 31943
rect 18337 31909 18371 31943
rect 18371 31909 18380 31943
rect 18328 31900 18380 31909
rect 19432 31875 19484 31884
rect 19432 31841 19441 31875
rect 19441 31841 19475 31875
rect 19475 31841 19484 31875
rect 19432 31832 19484 31841
rect 22284 31968 22336 32020
rect 23112 32011 23164 32020
rect 23112 31977 23121 32011
rect 23121 31977 23155 32011
rect 23155 31977 23164 32011
rect 23112 31968 23164 31977
rect 25412 31968 25464 32020
rect 29920 31968 29972 32020
rect 31668 31968 31720 32020
rect 32772 31968 32824 32020
rect 27436 31900 27488 31952
rect 12900 31807 12952 31816
rect 11612 31696 11664 31748
rect 12164 31696 12216 31748
rect 12900 31773 12909 31807
rect 12909 31773 12943 31807
rect 12943 31773 12952 31807
rect 12900 31764 12952 31773
rect 13544 31807 13596 31816
rect 13544 31773 13553 31807
rect 13553 31773 13587 31807
rect 13587 31773 13596 31807
rect 13544 31764 13596 31773
rect 14280 31764 14332 31816
rect 14924 31696 14976 31748
rect 10324 31671 10376 31680
rect 10324 31637 10333 31671
rect 10333 31637 10367 31671
rect 10367 31637 10376 31671
rect 10324 31628 10376 31637
rect 10692 31628 10744 31680
rect 12256 31628 12308 31680
rect 14832 31628 14884 31680
rect 15016 31628 15068 31680
rect 21088 31807 21140 31816
rect 21088 31773 21097 31807
rect 21097 31773 21131 31807
rect 21131 31773 21140 31807
rect 21088 31764 21140 31773
rect 22928 31832 22980 31884
rect 22468 31807 22520 31816
rect 22468 31773 22477 31807
rect 22477 31773 22511 31807
rect 22511 31773 22520 31807
rect 22468 31764 22520 31773
rect 23388 31807 23440 31816
rect 16580 31696 16632 31748
rect 16672 31696 16724 31748
rect 17316 31696 17368 31748
rect 22100 31696 22152 31748
rect 23388 31773 23397 31807
rect 23397 31773 23431 31807
rect 23431 31773 23440 31807
rect 23388 31764 23440 31773
rect 28172 31832 28224 31884
rect 23572 31807 23624 31816
rect 23572 31773 23581 31807
rect 23581 31773 23615 31807
rect 23615 31773 23624 31807
rect 23572 31764 23624 31773
rect 24492 31807 24544 31816
rect 24492 31773 24501 31807
rect 24501 31773 24535 31807
rect 24535 31773 24544 31807
rect 24492 31764 24544 31773
rect 26700 31764 26752 31816
rect 28540 31832 28592 31884
rect 29368 31900 29420 31952
rect 29552 31900 29604 31952
rect 30196 31875 30248 31884
rect 24032 31696 24084 31748
rect 24584 31696 24636 31748
rect 25320 31696 25372 31748
rect 28632 31807 28684 31816
rect 28632 31773 28641 31807
rect 28641 31773 28675 31807
rect 28675 31773 28684 31807
rect 28632 31764 28684 31773
rect 30196 31841 30205 31875
rect 30205 31841 30239 31875
rect 30239 31841 30248 31875
rect 30196 31832 30248 31841
rect 30012 31807 30064 31816
rect 30012 31773 30021 31807
rect 30021 31773 30055 31807
rect 30055 31773 30064 31807
rect 30012 31764 30064 31773
rect 31208 31764 31260 31816
rect 31852 31764 31904 31816
rect 32312 31832 32364 31884
rect 33508 31875 33560 31884
rect 33508 31841 33517 31875
rect 33517 31841 33551 31875
rect 33551 31841 33560 31875
rect 33508 31832 33560 31841
rect 46112 31832 46164 31884
rect 32220 31807 32272 31816
rect 32220 31773 32234 31807
rect 32234 31773 32268 31807
rect 32268 31773 32272 31807
rect 32220 31764 32272 31773
rect 32404 31807 32456 31816
rect 32404 31773 32413 31807
rect 32413 31773 32447 31807
rect 32447 31773 32456 31807
rect 32404 31764 32456 31773
rect 34060 31764 34112 31816
rect 35992 31807 36044 31816
rect 35992 31773 36001 31807
rect 36001 31773 36035 31807
rect 36035 31773 36044 31807
rect 35992 31764 36044 31773
rect 47952 31807 48004 31816
rect 47952 31773 47961 31807
rect 47961 31773 47995 31807
rect 47995 31773 48004 31807
rect 47952 31764 48004 31773
rect 36176 31739 36228 31748
rect 36176 31705 36185 31739
rect 36185 31705 36219 31739
rect 36219 31705 36228 31739
rect 36176 31696 36228 31705
rect 17040 31628 17092 31680
rect 25780 31628 25832 31680
rect 27988 31671 28040 31680
rect 27988 31637 27997 31671
rect 27997 31637 28031 31671
rect 28031 31637 28040 31671
rect 27988 31628 28040 31637
rect 28264 31628 28316 31680
rect 34244 31628 34296 31680
rect 48044 31671 48096 31680
rect 48044 31637 48053 31671
rect 48053 31637 48087 31671
rect 48087 31637 48096 31671
rect 48044 31628 48096 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 1584 31424 1636 31476
rect 1952 31263 2004 31272
rect 1952 31229 1961 31263
rect 1961 31229 1995 31263
rect 1995 31229 2004 31263
rect 1952 31220 2004 31229
rect 2872 31220 2924 31272
rect 3056 31263 3108 31272
rect 3056 31229 3065 31263
rect 3065 31229 3099 31263
rect 3099 31229 3108 31263
rect 3056 31220 3108 31229
rect 10324 31356 10376 31408
rect 10876 31399 10928 31408
rect 10876 31365 10885 31399
rect 10885 31365 10919 31399
rect 10919 31365 10928 31399
rect 10876 31356 10928 31365
rect 12992 31424 13044 31476
rect 13268 31424 13320 31476
rect 13636 31424 13688 31476
rect 14464 31467 14516 31476
rect 14464 31433 14473 31467
rect 14473 31433 14507 31467
rect 14507 31433 14516 31467
rect 14464 31424 14516 31433
rect 16672 31399 16724 31408
rect 10968 31331 11020 31340
rect 8208 31220 8260 31272
rect 10968 31297 10977 31331
rect 10977 31297 11011 31331
rect 11011 31297 11020 31331
rect 10968 31288 11020 31297
rect 11796 31288 11848 31340
rect 11980 31331 12032 31340
rect 11980 31297 11989 31331
rect 11989 31297 12023 31331
rect 12023 31297 12032 31331
rect 11980 31288 12032 31297
rect 11520 31220 11572 31272
rect 13084 31288 13136 31340
rect 13360 31331 13412 31340
rect 13360 31297 13369 31331
rect 13369 31297 13403 31331
rect 13403 31297 13412 31331
rect 13360 31288 13412 31297
rect 8300 31152 8352 31204
rect 10416 31152 10468 31204
rect 13268 31220 13320 31272
rect 14464 31288 14516 31340
rect 14832 31288 14884 31340
rect 15016 31288 15068 31340
rect 15200 31331 15252 31340
rect 15200 31297 15209 31331
rect 15209 31297 15243 31331
rect 15243 31297 15252 31331
rect 15200 31288 15252 31297
rect 10140 31084 10192 31136
rect 10784 31084 10836 31136
rect 11704 31084 11756 31136
rect 14464 31152 14516 31204
rect 14924 31195 14976 31204
rect 14924 31161 14933 31195
rect 14933 31161 14967 31195
rect 14967 31161 14976 31195
rect 14924 31152 14976 31161
rect 16672 31365 16681 31399
rect 16681 31365 16715 31399
rect 16715 31365 16724 31399
rect 16672 31356 16724 31365
rect 16764 31356 16816 31408
rect 18328 31356 18380 31408
rect 18880 31399 18932 31408
rect 18880 31365 18889 31399
rect 18889 31365 18923 31399
rect 18923 31365 18932 31399
rect 18880 31356 18932 31365
rect 20168 31356 20220 31408
rect 16028 31288 16080 31340
rect 17040 31331 17092 31340
rect 17040 31297 17049 31331
rect 17049 31297 17083 31331
rect 17083 31297 17092 31331
rect 17040 31288 17092 31297
rect 17224 31288 17276 31340
rect 23572 31424 23624 31476
rect 24400 31424 24452 31476
rect 25320 31467 25372 31476
rect 25320 31433 25329 31467
rect 25329 31433 25363 31467
rect 25363 31433 25372 31467
rect 25320 31424 25372 31433
rect 28632 31424 28684 31476
rect 32220 31424 32272 31476
rect 36176 31424 36228 31476
rect 25044 31356 25096 31408
rect 18696 31263 18748 31272
rect 18696 31229 18705 31263
rect 18705 31229 18739 31263
rect 18739 31229 18748 31263
rect 18696 31220 18748 31229
rect 20536 31263 20588 31272
rect 20536 31229 20545 31263
rect 20545 31229 20579 31263
rect 20579 31229 20588 31263
rect 20536 31220 20588 31229
rect 17684 31152 17736 31204
rect 22100 31263 22152 31272
rect 22100 31229 22109 31263
rect 22109 31229 22143 31263
rect 22143 31229 22152 31263
rect 23388 31288 23440 31340
rect 23480 31288 23532 31340
rect 24676 31288 24728 31340
rect 26056 31356 26108 31408
rect 30748 31356 30800 31408
rect 24768 31263 24820 31272
rect 22100 31220 22152 31229
rect 22744 31152 22796 31204
rect 23296 31152 23348 31204
rect 24768 31229 24777 31263
rect 24777 31229 24811 31263
rect 24811 31229 24820 31263
rect 24768 31220 24820 31229
rect 25780 31331 25832 31340
rect 25780 31297 25794 31331
rect 25794 31297 25828 31331
rect 25828 31297 25832 31331
rect 25780 31288 25832 31297
rect 25964 31331 26016 31340
rect 25964 31297 25973 31331
rect 25973 31297 26007 31331
rect 26007 31297 26016 31331
rect 25964 31288 26016 31297
rect 27896 31288 27948 31340
rect 28816 31288 28868 31340
rect 30472 31331 30524 31340
rect 30472 31297 30481 31331
rect 30481 31297 30515 31331
rect 30515 31297 30524 31331
rect 30472 31288 30524 31297
rect 30656 31331 30708 31340
rect 30656 31297 30665 31331
rect 30665 31297 30699 31331
rect 30699 31297 30708 31331
rect 30656 31288 30708 31297
rect 48044 31356 48096 31408
rect 32128 31331 32180 31340
rect 32128 31297 32137 31331
rect 32137 31297 32171 31331
rect 32171 31297 32180 31331
rect 32128 31288 32180 31297
rect 31208 31220 31260 31272
rect 35900 31288 35952 31340
rect 12716 31084 12768 31136
rect 14280 31127 14332 31136
rect 14280 31093 14289 31127
rect 14289 31093 14323 31127
rect 14323 31093 14332 31127
rect 14280 31084 14332 31093
rect 21640 31084 21692 31136
rect 23388 31084 23440 31136
rect 24400 31084 24452 31136
rect 30472 31152 30524 31204
rect 27160 31084 27212 31136
rect 28816 31127 28868 31136
rect 28816 31093 28825 31127
rect 28825 31093 28859 31127
rect 28859 31093 28868 31127
rect 28816 31084 28868 31093
rect 31300 31084 31352 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 1952 30880 2004 30932
rect 2872 30923 2924 30932
rect 2872 30889 2881 30923
rect 2881 30889 2915 30923
rect 2915 30889 2924 30923
rect 2872 30880 2924 30889
rect 10416 30923 10468 30932
rect 10416 30889 10425 30923
rect 10425 30889 10459 30923
rect 10459 30889 10468 30923
rect 10416 30880 10468 30889
rect 10508 30880 10560 30932
rect 10968 30880 11020 30932
rect 13636 30880 13688 30932
rect 15200 30880 15252 30932
rect 16764 30880 16816 30932
rect 24676 30880 24728 30932
rect 30472 30923 30524 30932
rect 30472 30889 30481 30923
rect 30481 30889 30515 30923
rect 30515 30889 30524 30923
rect 30472 30880 30524 30889
rect 35992 30880 36044 30932
rect 11060 30812 11112 30864
rect 12072 30812 12124 30864
rect 14372 30812 14424 30864
rect 14924 30812 14976 30864
rect 15292 30855 15344 30864
rect 15292 30821 15301 30855
rect 15301 30821 15335 30855
rect 15335 30821 15344 30855
rect 15292 30812 15344 30821
rect 16580 30812 16632 30864
rect 31300 30812 31352 30864
rect 7656 30676 7708 30728
rect 10784 30676 10836 30728
rect 12164 30676 12216 30728
rect 11612 30608 11664 30660
rect 11796 30608 11848 30660
rect 11980 30540 12032 30592
rect 12348 30583 12400 30592
rect 12348 30549 12357 30583
rect 12357 30549 12391 30583
rect 12391 30549 12400 30583
rect 12348 30540 12400 30549
rect 12808 30719 12860 30728
rect 12808 30685 12817 30719
rect 12817 30685 12851 30719
rect 12851 30685 12860 30719
rect 12808 30676 12860 30685
rect 13084 30719 13136 30728
rect 13084 30685 13093 30719
rect 13093 30685 13127 30719
rect 13127 30685 13136 30719
rect 13084 30676 13136 30685
rect 13360 30676 13412 30728
rect 14372 30676 14424 30728
rect 18420 30744 18472 30796
rect 22928 30787 22980 30796
rect 22928 30753 22937 30787
rect 22937 30753 22971 30787
rect 22971 30753 22980 30787
rect 22928 30744 22980 30753
rect 24032 30744 24084 30796
rect 16672 30719 16724 30728
rect 16672 30685 16681 30719
rect 16681 30685 16715 30719
rect 16715 30685 16724 30719
rect 16672 30676 16724 30685
rect 16764 30676 16816 30728
rect 17960 30676 18012 30728
rect 20168 30676 20220 30728
rect 21916 30676 21968 30728
rect 22468 30676 22520 30728
rect 23388 30676 23440 30728
rect 24400 30719 24452 30728
rect 24400 30685 24409 30719
rect 24409 30685 24443 30719
rect 24443 30685 24452 30719
rect 24400 30676 24452 30685
rect 25412 30719 25464 30728
rect 25412 30685 25421 30719
rect 25421 30685 25455 30719
rect 25455 30685 25464 30719
rect 25412 30676 25464 30685
rect 25504 30676 25556 30728
rect 25964 30676 26016 30728
rect 27712 30744 27764 30796
rect 27896 30676 27948 30728
rect 12716 30651 12768 30660
rect 12716 30617 12725 30651
rect 12725 30617 12759 30651
rect 12759 30617 12768 30651
rect 12716 30608 12768 30617
rect 18696 30608 18748 30660
rect 23480 30608 23532 30660
rect 24584 30651 24636 30660
rect 24584 30617 24593 30651
rect 24593 30617 24627 30651
rect 24627 30617 24636 30651
rect 24584 30608 24636 30617
rect 24860 30608 24912 30660
rect 31024 30744 31076 30796
rect 30472 30676 30524 30728
rect 13176 30540 13228 30592
rect 17224 30540 17276 30592
rect 25320 30540 25372 30592
rect 26700 30540 26752 30592
rect 27528 30540 27580 30592
rect 28172 30540 28224 30592
rect 31944 30719 31996 30728
rect 31944 30685 31953 30719
rect 31953 30685 31987 30719
rect 31987 30685 31996 30719
rect 31944 30676 31996 30685
rect 35348 30676 35400 30728
rect 34520 30608 34572 30660
rect 32312 30540 32364 30592
rect 33324 30583 33376 30592
rect 33324 30549 33333 30583
rect 33333 30549 33367 30583
rect 33367 30549 33376 30583
rect 33324 30540 33376 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 11796 30379 11848 30388
rect 11796 30345 11805 30379
rect 11805 30345 11839 30379
rect 11839 30345 11848 30379
rect 11796 30336 11848 30345
rect 12256 30336 12308 30388
rect 14372 30379 14424 30388
rect 9680 30268 9732 30320
rect 10508 30243 10560 30252
rect 10508 30209 10517 30243
rect 10517 30209 10551 30243
rect 10551 30209 10560 30243
rect 10508 30200 10560 30209
rect 11704 30268 11756 30320
rect 12072 30268 12124 30320
rect 13268 30311 13320 30320
rect 13268 30277 13277 30311
rect 13277 30277 13311 30311
rect 13311 30277 13320 30311
rect 13268 30268 13320 30277
rect 14372 30345 14381 30379
rect 14381 30345 14415 30379
rect 14415 30345 14424 30379
rect 14372 30336 14424 30345
rect 19340 30336 19392 30388
rect 20444 30336 20496 30388
rect 20904 30336 20956 30388
rect 22928 30336 22980 30388
rect 24032 30336 24084 30388
rect 24308 30336 24360 30388
rect 24860 30379 24912 30388
rect 24860 30345 24869 30379
rect 24869 30345 24903 30379
rect 24903 30345 24912 30379
rect 24860 30336 24912 30345
rect 27988 30336 28040 30388
rect 32128 30379 32180 30388
rect 32128 30345 32137 30379
rect 32137 30345 32171 30379
rect 32171 30345 32180 30379
rect 32128 30336 32180 30345
rect 1952 30175 2004 30184
rect 1952 30141 1961 30175
rect 1961 30141 1995 30175
rect 1995 30141 2004 30175
rect 1952 30132 2004 30141
rect 2780 30132 2832 30184
rect 2872 30175 2924 30184
rect 2872 30141 2881 30175
rect 2881 30141 2915 30175
rect 2915 30141 2924 30175
rect 2872 30132 2924 30141
rect 10232 30132 10284 30184
rect 12532 30200 12584 30252
rect 14372 30243 14424 30252
rect 14372 30209 14381 30243
rect 14381 30209 14415 30243
rect 14415 30209 14424 30243
rect 14372 30200 14424 30209
rect 19524 30268 19576 30320
rect 16028 30200 16080 30252
rect 17040 30200 17092 30252
rect 19708 30243 19760 30252
rect 19708 30209 19717 30243
rect 19717 30209 19751 30243
rect 19751 30209 19760 30243
rect 19708 30200 19760 30209
rect 20168 30200 20220 30252
rect 12256 30132 12308 30184
rect 14188 30175 14240 30184
rect 14188 30141 14197 30175
rect 14197 30141 14231 30175
rect 14231 30141 14240 30175
rect 14188 30132 14240 30141
rect 8944 29996 8996 30048
rect 16672 30132 16724 30184
rect 17500 30132 17552 30184
rect 19984 30175 20036 30184
rect 19984 30141 19993 30175
rect 19993 30141 20027 30175
rect 20027 30141 20036 30175
rect 19984 30132 20036 30141
rect 20904 30132 20956 30184
rect 21916 30200 21968 30252
rect 23204 30200 23256 30252
rect 23480 30200 23532 30252
rect 25044 30268 25096 30320
rect 26056 30311 26108 30320
rect 22468 30132 22520 30184
rect 24124 30243 24176 30252
rect 24124 30209 24133 30243
rect 24133 30209 24167 30243
rect 24167 30209 24176 30243
rect 24124 30200 24176 30209
rect 24308 30243 24360 30252
rect 24308 30209 24317 30243
rect 24317 30209 24351 30243
rect 24351 30209 24360 30243
rect 26056 30277 26065 30311
rect 26065 30277 26099 30311
rect 26099 30277 26108 30311
rect 26056 30268 26108 30277
rect 29828 30268 29880 30320
rect 32588 30311 32640 30320
rect 32588 30277 32597 30311
rect 32597 30277 32631 30311
rect 32631 30277 32640 30311
rect 32588 30268 32640 30277
rect 33048 30268 33100 30320
rect 24308 30200 24360 30209
rect 25044 30132 25096 30184
rect 25320 30243 25372 30252
rect 25320 30209 25329 30243
rect 25329 30209 25363 30243
rect 25363 30209 25372 30243
rect 25320 30200 25372 30209
rect 25504 30243 25556 30252
rect 25504 30209 25513 30243
rect 25513 30209 25547 30243
rect 25547 30209 25556 30243
rect 25504 30200 25556 30209
rect 27620 30200 27672 30252
rect 25780 30132 25832 30184
rect 26332 30132 26384 30184
rect 27528 30132 27580 30184
rect 21824 30064 21876 30116
rect 27804 30064 27856 30116
rect 28172 30200 28224 30252
rect 33324 30200 33376 30252
rect 35992 30268 36044 30320
rect 28540 30175 28592 30184
rect 28540 30141 28549 30175
rect 28549 30141 28583 30175
rect 28583 30141 28592 30175
rect 28540 30132 28592 30141
rect 33508 30132 33560 30184
rect 29920 30107 29972 30116
rect 29920 30073 29929 30107
rect 29929 30073 29963 30107
rect 29963 30073 29972 30107
rect 29920 30064 29972 30073
rect 30104 30064 30156 30116
rect 34612 30200 34664 30252
rect 35808 30064 35860 30116
rect 46020 30064 46072 30116
rect 15200 29996 15252 30048
rect 16764 29996 16816 30048
rect 17132 29996 17184 30048
rect 20444 30039 20496 30048
rect 20444 30005 20453 30039
rect 20453 30005 20487 30039
rect 20487 30005 20496 30039
rect 20444 29996 20496 30005
rect 20536 29996 20588 30048
rect 22376 29996 22428 30048
rect 23112 30039 23164 30048
rect 23112 30005 23121 30039
rect 23121 30005 23155 30039
rect 23155 30005 23164 30039
rect 23112 29996 23164 30005
rect 23664 30039 23716 30048
rect 23664 30005 23673 30039
rect 23673 30005 23707 30039
rect 23707 30005 23716 30039
rect 23664 29996 23716 30005
rect 23756 29996 23808 30048
rect 25688 29996 25740 30048
rect 27436 30039 27488 30048
rect 27436 30005 27445 30039
rect 27445 30005 27479 30039
rect 27479 30005 27488 30039
rect 27436 29996 27488 30005
rect 30196 29996 30248 30048
rect 33324 29996 33376 30048
rect 34520 29996 34572 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 1952 29792 2004 29844
rect 2780 29792 2832 29844
rect 14188 29792 14240 29844
rect 15108 29792 15160 29844
rect 15936 29792 15988 29844
rect 16580 29792 16632 29844
rect 17224 29792 17276 29844
rect 2872 29588 2924 29640
rect 8944 29724 8996 29776
rect 12532 29724 12584 29776
rect 8208 29656 8260 29708
rect 9312 29656 9364 29708
rect 13268 29656 13320 29708
rect 17776 29724 17828 29776
rect 15108 29656 15160 29708
rect 12164 29588 12216 29640
rect 8300 29520 8352 29572
rect 8944 29563 8996 29572
rect 8944 29529 8953 29563
rect 8953 29529 8987 29563
rect 8987 29529 8996 29563
rect 8944 29520 8996 29529
rect 8484 29452 8536 29504
rect 12348 29520 12400 29572
rect 9496 29452 9548 29504
rect 12256 29495 12308 29504
rect 12256 29461 12265 29495
rect 12265 29461 12299 29495
rect 12299 29461 12308 29495
rect 14280 29588 14332 29640
rect 14832 29588 14884 29640
rect 15016 29631 15068 29640
rect 15016 29597 15025 29631
rect 15025 29597 15059 29631
rect 15059 29597 15068 29631
rect 15016 29588 15068 29597
rect 15568 29588 15620 29640
rect 16028 29631 16080 29640
rect 16028 29597 16037 29631
rect 16037 29597 16071 29631
rect 16071 29597 16080 29631
rect 16028 29588 16080 29597
rect 16488 29656 16540 29708
rect 17132 29631 17184 29640
rect 17132 29597 17141 29631
rect 17141 29597 17175 29631
rect 17175 29597 17184 29631
rect 17132 29588 17184 29597
rect 17592 29588 17644 29640
rect 17684 29588 17736 29640
rect 18328 29631 18380 29640
rect 18328 29597 18337 29631
rect 18337 29597 18371 29631
rect 18371 29597 18380 29631
rect 19524 29792 19576 29844
rect 19984 29792 20036 29844
rect 21548 29835 21600 29844
rect 21548 29801 21557 29835
rect 21557 29801 21591 29835
rect 21591 29801 21600 29835
rect 21548 29792 21600 29801
rect 22744 29792 22796 29844
rect 24124 29792 24176 29844
rect 25688 29792 25740 29844
rect 27712 29792 27764 29844
rect 27804 29835 27856 29844
rect 27804 29801 27813 29835
rect 27813 29801 27847 29835
rect 27847 29801 27856 29835
rect 27804 29792 27856 29801
rect 27988 29792 28040 29844
rect 46940 29792 46992 29844
rect 20444 29699 20496 29708
rect 18328 29588 18380 29597
rect 12992 29520 13044 29572
rect 12256 29452 12308 29461
rect 15476 29452 15528 29504
rect 17224 29452 17276 29504
rect 17408 29495 17460 29504
rect 17408 29461 17417 29495
rect 17417 29461 17451 29495
rect 17451 29461 17460 29495
rect 17408 29452 17460 29461
rect 17868 29495 17920 29504
rect 17868 29461 17877 29495
rect 17877 29461 17911 29495
rect 17911 29461 17920 29495
rect 17868 29452 17920 29461
rect 17960 29452 18012 29504
rect 19340 29588 19392 29640
rect 20444 29665 20453 29699
rect 20453 29665 20487 29699
rect 20487 29665 20496 29699
rect 20444 29656 20496 29665
rect 21640 29656 21692 29708
rect 24032 29724 24084 29776
rect 25872 29724 25924 29776
rect 35808 29724 35860 29776
rect 25504 29656 25556 29708
rect 26608 29656 26660 29708
rect 26792 29656 26844 29708
rect 28540 29656 28592 29708
rect 29552 29656 29604 29708
rect 30196 29699 30248 29708
rect 30196 29665 30205 29699
rect 30205 29665 30239 29699
rect 30239 29665 30248 29699
rect 30196 29656 30248 29665
rect 20536 29588 20588 29640
rect 22376 29631 22428 29640
rect 22376 29597 22385 29631
rect 22385 29597 22419 29631
rect 22419 29597 22428 29631
rect 22376 29588 22428 29597
rect 21824 29520 21876 29572
rect 23112 29588 23164 29640
rect 23756 29588 23808 29640
rect 25412 29588 25464 29640
rect 26976 29588 27028 29640
rect 23664 29520 23716 29572
rect 26792 29563 26844 29572
rect 21548 29452 21600 29504
rect 23388 29452 23440 29504
rect 23756 29495 23808 29504
rect 23756 29461 23765 29495
rect 23765 29461 23799 29495
rect 23799 29461 23808 29495
rect 23756 29452 23808 29461
rect 24032 29452 24084 29504
rect 24860 29452 24912 29504
rect 26424 29452 26476 29504
rect 26792 29529 26801 29563
rect 26801 29529 26835 29563
rect 26835 29529 26844 29563
rect 26792 29520 26844 29529
rect 28816 29631 28868 29640
rect 28816 29597 28825 29631
rect 28825 29597 28859 29631
rect 28859 29597 28868 29631
rect 28816 29588 28868 29597
rect 34796 29656 34848 29708
rect 27528 29520 27580 29572
rect 30380 29520 30432 29572
rect 31024 29520 31076 29572
rect 32036 29631 32088 29640
rect 32036 29597 32045 29631
rect 32045 29597 32079 29631
rect 32079 29597 32088 29631
rect 32036 29588 32088 29597
rect 32312 29588 32364 29640
rect 32772 29588 32824 29640
rect 35072 29631 35124 29640
rect 35072 29597 35095 29631
rect 35095 29597 35124 29631
rect 35072 29588 35124 29597
rect 32404 29520 32456 29572
rect 29920 29495 29972 29504
rect 29920 29461 29929 29495
rect 29929 29461 29963 29495
rect 29963 29461 29972 29495
rect 29920 29452 29972 29461
rect 31576 29495 31628 29504
rect 31576 29461 31585 29495
rect 31585 29461 31619 29495
rect 31619 29461 31628 29495
rect 31576 29452 31628 29461
rect 31760 29452 31812 29504
rect 32128 29452 32180 29504
rect 34796 29495 34848 29504
rect 34796 29461 34805 29495
rect 34805 29461 34839 29495
rect 34839 29461 34848 29495
rect 34796 29452 34848 29461
rect 35532 29656 35584 29708
rect 35716 29588 35768 29640
rect 47308 29631 47360 29640
rect 47308 29597 47317 29631
rect 47317 29597 47351 29631
rect 47351 29597 47360 29631
rect 47308 29588 47360 29597
rect 35624 29520 35676 29572
rect 35440 29452 35492 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 7012 29112 7064 29164
rect 8208 29180 8260 29232
rect 16580 29248 16632 29300
rect 16672 29248 16724 29300
rect 17224 29291 17276 29300
rect 17224 29257 17233 29291
rect 17233 29257 17267 29291
rect 17267 29257 17276 29291
rect 17224 29248 17276 29257
rect 17316 29248 17368 29300
rect 12164 29180 12216 29232
rect 9404 29155 9456 29164
rect 9404 29121 9413 29155
rect 9413 29121 9447 29155
rect 9447 29121 9456 29155
rect 9404 29112 9456 29121
rect 9496 29155 9548 29164
rect 9496 29121 9505 29155
rect 9505 29121 9539 29155
rect 9539 29121 9548 29155
rect 9496 29112 9548 29121
rect 9680 29155 9732 29164
rect 9680 29121 9689 29155
rect 9689 29121 9723 29155
rect 9723 29121 9732 29155
rect 12532 29155 12584 29164
rect 9680 29112 9732 29121
rect 12532 29121 12541 29155
rect 12541 29121 12575 29155
rect 12575 29121 12584 29155
rect 12532 29112 12584 29121
rect 9772 29044 9824 29096
rect 10324 29044 10376 29096
rect 13268 29112 13320 29164
rect 15292 29180 15344 29232
rect 15476 29180 15528 29232
rect 17500 29180 17552 29232
rect 17868 29180 17920 29232
rect 20168 29248 20220 29300
rect 23204 29291 23256 29300
rect 23204 29257 23213 29291
rect 23213 29257 23247 29291
rect 23247 29257 23256 29291
rect 23204 29248 23256 29257
rect 27068 29248 27120 29300
rect 14096 29155 14148 29164
rect 14096 29121 14130 29155
rect 14130 29121 14148 29155
rect 14096 29112 14148 29121
rect 15752 29112 15804 29164
rect 15936 29155 15988 29164
rect 15936 29121 15945 29155
rect 15945 29121 15979 29155
rect 15979 29121 15988 29155
rect 15936 29112 15988 29121
rect 17132 29112 17184 29164
rect 17684 29155 17736 29164
rect 17684 29121 17693 29155
rect 17693 29121 17727 29155
rect 17727 29121 17736 29155
rect 17684 29112 17736 29121
rect 17776 29112 17828 29164
rect 19892 29112 19944 29164
rect 8484 28976 8536 29028
rect 11980 28976 12032 29028
rect 2044 28951 2096 28960
rect 2044 28917 2053 28951
rect 2053 28917 2087 28951
rect 2087 28917 2096 28951
rect 2044 28908 2096 28917
rect 12992 28908 13044 28960
rect 15568 29044 15620 29096
rect 16488 29044 16540 29096
rect 17500 29044 17552 29096
rect 17960 29044 18012 29096
rect 20628 29180 20680 29232
rect 20904 29112 20956 29164
rect 21824 29155 21876 29164
rect 21824 29121 21833 29155
rect 21833 29121 21867 29155
rect 21867 29121 21876 29155
rect 21824 29112 21876 29121
rect 22376 29180 22428 29232
rect 25504 29180 25556 29232
rect 27528 29223 27580 29232
rect 27528 29189 27537 29223
rect 27537 29189 27571 29223
rect 27571 29189 27580 29223
rect 27528 29180 27580 29189
rect 22744 29112 22796 29164
rect 23756 29112 23808 29164
rect 24768 29112 24820 29164
rect 24860 29112 24912 29164
rect 27436 29112 27488 29164
rect 29920 29248 29972 29300
rect 30012 29248 30064 29300
rect 31576 29248 31628 29300
rect 31760 29248 31812 29300
rect 32956 29248 33008 29300
rect 34704 29291 34756 29300
rect 34704 29257 34713 29291
rect 34713 29257 34747 29291
rect 34747 29257 34756 29291
rect 34704 29248 34756 29257
rect 33232 29180 33284 29232
rect 33324 29180 33376 29232
rect 15108 28976 15160 29028
rect 17592 29019 17644 29028
rect 17592 28985 17601 29019
rect 17601 28985 17635 29019
rect 17635 28985 17644 29019
rect 17592 28976 17644 28985
rect 14464 28908 14516 28960
rect 15016 28908 15068 28960
rect 16488 28908 16540 28960
rect 22468 29044 22520 29096
rect 27620 29044 27672 29096
rect 33968 29112 34020 29164
rect 36636 29248 36688 29300
rect 34704 29112 34756 29164
rect 34796 29112 34848 29164
rect 46020 29180 46072 29232
rect 35256 29112 35308 29164
rect 46756 29112 46808 29164
rect 19340 28908 19392 28960
rect 19616 28908 19668 28960
rect 26976 28976 27028 29028
rect 33508 29044 33560 29096
rect 31024 28908 31076 28960
rect 33692 28976 33744 29028
rect 46664 28976 46716 29028
rect 46296 28908 46348 28960
rect 46480 28908 46532 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 2044 28568 2096 28620
rect 2780 28611 2832 28620
rect 2780 28577 2789 28611
rect 2789 28577 2823 28611
rect 2823 28577 2832 28611
rect 7012 28611 7064 28620
rect 2780 28568 2832 28577
rect 7012 28577 7021 28611
rect 7021 28577 7055 28611
rect 7055 28577 7064 28611
rect 7012 28568 7064 28577
rect 9220 28543 9272 28552
rect 9220 28509 9229 28543
rect 9229 28509 9263 28543
rect 9263 28509 9272 28543
rect 9220 28500 9272 28509
rect 9404 28704 9456 28756
rect 14096 28704 14148 28756
rect 15660 28704 15712 28756
rect 23480 28704 23532 28756
rect 26332 28704 26384 28756
rect 31208 28704 31260 28756
rect 32036 28704 32088 28756
rect 33232 28747 33284 28756
rect 33232 28713 33241 28747
rect 33241 28713 33275 28747
rect 33275 28713 33284 28747
rect 33232 28704 33284 28713
rect 18328 28636 18380 28688
rect 20168 28679 20220 28688
rect 20168 28645 20177 28679
rect 20177 28645 20211 28679
rect 20211 28645 20220 28679
rect 20168 28636 20220 28645
rect 22836 28636 22888 28688
rect 24308 28636 24360 28688
rect 14464 28568 14516 28620
rect 27068 28611 27120 28620
rect 9404 28543 9456 28552
rect 9404 28509 9413 28543
rect 9413 28509 9447 28543
rect 9447 28509 9456 28543
rect 9404 28500 9456 28509
rect 9680 28500 9732 28552
rect 10140 28543 10192 28552
rect 10140 28509 10149 28543
rect 10149 28509 10183 28543
rect 10183 28509 10192 28543
rect 10140 28500 10192 28509
rect 2136 28432 2188 28484
rect 8392 28407 8444 28416
rect 8392 28373 8401 28407
rect 8401 28373 8435 28407
rect 8435 28373 8444 28407
rect 8392 28364 8444 28373
rect 10232 28407 10284 28416
rect 10232 28373 10241 28407
rect 10241 28373 10275 28407
rect 10275 28373 10284 28407
rect 10232 28364 10284 28373
rect 15016 28500 15068 28552
rect 15200 28432 15252 28484
rect 15844 28500 15896 28552
rect 16028 28543 16080 28552
rect 16028 28509 16037 28543
rect 16037 28509 16071 28543
rect 16071 28509 16080 28543
rect 16028 28500 16080 28509
rect 16488 28543 16540 28552
rect 16488 28509 16497 28543
rect 16497 28509 16531 28543
rect 16531 28509 16540 28543
rect 16488 28500 16540 28509
rect 19892 28500 19944 28552
rect 20720 28500 20772 28552
rect 21180 28500 21232 28552
rect 17224 28432 17276 28484
rect 19616 28432 19668 28484
rect 20536 28432 20588 28484
rect 26332 28432 26384 28484
rect 17592 28364 17644 28416
rect 23204 28364 23256 28416
rect 26240 28364 26292 28416
rect 27068 28577 27077 28611
rect 27077 28577 27111 28611
rect 27111 28577 27120 28611
rect 27068 28568 27120 28577
rect 27344 28568 27396 28620
rect 27252 28500 27304 28552
rect 27712 28500 27764 28552
rect 29552 28636 29604 28688
rect 30104 28636 30156 28688
rect 34704 28611 34756 28620
rect 34704 28577 34713 28611
rect 34713 28577 34747 28611
rect 34747 28577 34756 28611
rect 34704 28568 34756 28577
rect 36636 28611 36688 28620
rect 36636 28577 36645 28611
rect 36645 28577 36679 28611
rect 36679 28577 36688 28611
rect 36636 28568 36688 28577
rect 46296 28611 46348 28620
rect 46296 28577 46305 28611
rect 46305 28577 46339 28611
rect 46339 28577 46348 28611
rect 46296 28568 46348 28577
rect 46480 28611 46532 28620
rect 46480 28577 46489 28611
rect 46489 28577 46523 28611
rect 46523 28577 46532 28611
rect 46480 28568 46532 28577
rect 47492 28568 47544 28620
rect 47676 28568 47728 28620
rect 48136 28611 48188 28620
rect 48136 28577 48145 28611
rect 48145 28577 48179 28611
rect 48179 28577 48188 28611
rect 48136 28568 48188 28577
rect 28356 28543 28408 28552
rect 27344 28432 27396 28484
rect 28356 28509 28365 28543
rect 28365 28509 28399 28543
rect 28399 28509 28408 28543
rect 28356 28500 28408 28509
rect 30380 28543 30432 28552
rect 30380 28509 30389 28543
rect 30389 28509 30423 28543
rect 30423 28509 30432 28543
rect 30380 28500 30432 28509
rect 31944 28500 31996 28552
rect 32588 28500 32640 28552
rect 33692 28543 33744 28552
rect 33692 28509 33701 28543
rect 33701 28509 33735 28543
rect 33735 28509 33744 28543
rect 33692 28500 33744 28509
rect 34520 28500 34572 28552
rect 35900 28500 35952 28552
rect 31024 28475 31076 28484
rect 31024 28441 31033 28475
rect 31033 28441 31067 28475
rect 31067 28441 31076 28475
rect 31024 28432 31076 28441
rect 31208 28475 31260 28484
rect 31208 28441 31217 28475
rect 31217 28441 31251 28475
rect 31251 28441 31260 28475
rect 31208 28432 31260 28441
rect 31760 28432 31812 28484
rect 27436 28364 27488 28416
rect 27712 28407 27764 28416
rect 27712 28373 27721 28407
rect 27721 28373 27755 28407
rect 27755 28373 27764 28407
rect 27712 28364 27764 28373
rect 38476 28475 38528 28484
rect 38476 28441 38485 28475
rect 38485 28441 38519 28475
rect 38519 28441 38528 28475
rect 38476 28432 38528 28441
rect 34060 28407 34112 28416
rect 34060 28373 34069 28407
rect 34069 28373 34103 28407
rect 34103 28373 34112 28407
rect 34060 28364 34112 28373
rect 47584 28364 47636 28416
rect 47860 28364 47912 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 2136 28203 2188 28212
rect 2136 28169 2145 28203
rect 2145 28169 2179 28203
rect 2179 28169 2188 28203
rect 2136 28160 2188 28169
rect 6368 28160 6420 28212
rect 13084 28160 13136 28212
rect 16028 28160 16080 28212
rect 17500 28203 17552 28212
rect 17500 28169 17509 28203
rect 17509 28169 17543 28203
rect 17543 28169 17552 28203
rect 17500 28160 17552 28169
rect 18420 28135 18472 28144
rect 2044 28067 2096 28076
rect 2044 28033 2053 28067
rect 2053 28033 2087 28067
rect 2087 28033 2096 28067
rect 2044 28024 2096 28033
rect 9772 28024 9824 28076
rect 9956 28067 10008 28076
rect 9956 28033 9965 28067
rect 9965 28033 9999 28067
rect 9999 28033 10008 28067
rect 9956 28024 10008 28033
rect 10324 28024 10376 28076
rect 18420 28101 18429 28135
rect 18429 28101 18463 28135
rect 18463 28101 18472 28135
rect 18420 28092 18472 28101
rect 20168 28135 20220 28144
rect 20168 28101 20202 28135
rect 20202 28101 20220 28135
rect 20168 28092 20220 28101
rect 23204 28135 23256 28144
rect 23204 28101 23213 28135
rect 23213 28101 23247 28135
rect 23247 28101 23256 28135
rect 23204 28092 23256 28101
rect 27712 28092 27764 28144
rect 27804 28092 27856 28144
rect 12992 28067 13044 28076
rect 12992 28033 13001 28067
rect 13001 28033 13035 28067
rect 13035 28033 13044 28067
rect 12992 28024 13044 28033
rect 15568 28067 15620 28076
rect 15568 28033 15577 28067
rect 15577 28033 15611 28067
rect 15611 28033 15620 28067
rect 15568 28024 15620 28033
rect 19340 28024 19392 28076
rect 19984 28024 20036 28076
rect 26056 28067 26108 28076
rect 26056 28033 26065 28067
rect 26065 28033 26099 28067
rect 26099 28033 26108 28067
rect 26056 28024 26108 28033
rect 9772 27820 9824 27872
rect 11152 27956 11204 28008
rect 15200 27956 15252 28008
rect 17684 27999 17736 28008
rect 17684 27965 17693 27999
rect 17693 27965 17727 27999
rect 17727 27965 17736 27999
rect 17684 27956 17736 27965
rect 23480 27999 23532 28008
rect 12900 27931 12952 27940
rect 12900 27897 12909 27931
rect 12909 27897 12943 27931
rect 12943 27897 12952 27931
rect 23480 27965 23489 27999
rect 23489 27965 23523 27999
rect 23523 27965 23532 27999
rect 23480 27956 23532 27965
rect 26240 28067 26292 28076
rect 26240 28033 26254 28067
rect 26254 28033 26288 28067
rect 26288 28033 26292 28067
rect 26240 28024 26292 28033
rect 28172 28024 28224 28076
rect 33048 28092 33100 28144
rect 26700 27956 26752 28008
rect 26976 27999 27028 28008
rect 26976 27965 26985 27999
rect 26985 27965 27019 27999
rect 27019 27965 27028 27999
rect 26976 27956 27028 27965
rect 29552 28067 29604 28076
rect 29552 28033 29561 28067
rect 29561 28033 29595 28067
rect 29595 28033 29604 28067
rect 29736 28067 29788 28076
rect 29552 28024 29604 28033
rect 29736 28033 29745 28067
rect 29745 28033 29779 28067
rect 29779 28033 29788 28067
rect 29736 28024 29788 28033
rect 32036 28024 32088 28076
rect 34796 28024 34848 28076
rect 29920 27956 29972 28008
rect 32588 27999 32640 28008
rect 32588 27965 32597 27999
rect 32597 27965 32631 27999
rect 32631 27965 32640 27999
rect 32588 27956 32640 27965
rect 35440 28067 35492 28076
rect 35440 28033 35449 28067
rect 35449 28033 35483 28067
rect 35483 28033 35492 28067
rect 35624 28067 35676 28076
rect 35440 28024 35492 28033
rect 35624 28033 35633 28067
rect 35633 28033 35667 28067
rect 35667 28033 35676 28067
rect 35624 28024 35676 28033
rect 47124 28024 47176 28076
rect 47860 28067 47912 28076
rect 47860 28033 47869 28067
rect 47869 28033 47903 28067
rect 47903 28033 47912 28067
rect 47860 28024 47912 28033
rect 12900 27888 12952 27897
rect 9956 27820 10008 27872
rect 17592 27820 17644 27872
rect 20628 27820 20680 27872
rect 26240 27820 26292 27872
rect 28080 27888 28132 27940
rect 33968 27931 34020 27940
rect 27712 27820 27764 27872
rect 29644 27820 29696 27872
rect 33968 27897 33977 27931
rect 33977 27897 34011 27931
rect 34011 27897 34020 27931
rect 33968 27888 34020 27897
rect 35900 27888 35952 27940
rect 35992 27820 36044 27872
rect 47032 27863 47084 27872
rect 47032 27829 47041 27863
rect 47041 27829 47075 27863
rect 47075 27829 47084 27863
rect 47032 27820 47084 27829
rect 47124 27820 47176 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 2044 27616 2096 27668
rect 2596 27616 2648 27668
rect 17040 27616 17092 27668
rect 20904 27616 20956 27668
rect 27344 27659 27396 27668
rect 27344 27625 27353 27659
rect 27353 27625 27387 27659
rect 27387 27625 27396 27659
rect 27344 27616 27396 27625
rect 27436 27616 27488 27668
rect 28080 27616 28132 27668
rect 28356 27616 28408 27668
rect 29736 27616 29788 27668
rect 32036 27659 32088 27668
rect 32036 27625 32045 27659
rect 32045 27625 32079 27659
rect 32079 27625 32088 27659
rect 32036 27616 32088 27625
rect 9680 27548 9732 27600
rect 11152 27591 11204 27600
rect 11152 27557 11161 27591
rect 11161 27557 11195 27591
rect 11195 27557 11204 27591
rect 11152 27548 11204 27557
rect 17776 27548 17828 27600
rect 20720 27591 20772 27600
rect 20720 27557 20729 27591
rect 20729 27557 20763 27591
rect 20763 27557 20772 27591
rect 20720 27548 20772 27557
rect 24860 27548 24912 27600
rect 25596 27548 25648 27600
rect 30564 27548 30616 27600
rect 33140 27616 33192 27668
rect 35624 27616 35676 27668
rect 34796 27548 34848 27600
rect 35072 27548 35124 27600
rect 1860 27523 1912 27532
rect 1860 27489 1869 27523
rect 1869 27489 1903 27523
rect 1903 27489 1912 27523
rect 1860 27480 1912 27489
rect 9312 27480 9364 27532
rect 12164 27523 12216 27532
rect 1400 27455 1452 27464
rect 1400 27421 1409 27455
rect 1409 27421 1443 27455
rect 1443 27421 1452 27455
rect 1400 27412 1452 27421
rect 9036 27412 9088 27464
rect 10324 27412 10376 27464
rect 12164 27489 12173 27523
rect 12173 27489 12207 27523
rect 12207 27489 12216 27523
rect 12164 27480 12216 27489
rect 24584 27480 24636 27532
rect 12440 27455 12492 27464
rect 12440 27421 12474 27455
rect 12474 27421 12492 27455
rect 2136 27344 2188 27396
rect 10232 27344 10284 27396
rect 10508 27344 10560 27396
rect 12440 27412 12492 27421
rect 16488 27412 16540 27464
rect 17408 27455 17460 27464
rect 17408 27421 17417 27455
rect 17417 27421 17451 27455
rect 17451 27421 17460 27455
rect 17408 27412 17460 27421
rect 20628 27412 20680 27464
rect 15108 27387 15160 27396
rect 15108 27353 15142 27387
rect 15142 27353 15160 27387
rect 15108 27344 15160 27353
rect 22928 27344 22980 27396
rect 24768 27412 24820 27464
rect 26792 27412 26844 27464
rect 26976 27412 27028 27464
rect 27068 27412 27120 27464
rect 28632 27455 28684 27464
rect 28632 27421 28641 27455
rect 28641 27421 28675 27455
rect 28675 27421 28684 27455
rect 28632 27412 28684 27421
rect 29644 27412 29696 27464
rect 26240 27387 26292 27396
rect 26240 27353 26274 27387
rect 26274 27353 26292 27387
rect 26240 27344 26292 27353
rect 27712 27344 27764 27396
rect 31208 27344 31260 27396
rect 9220 27276 9272 27328
rect 10876 27276 10928 27328
rect 14188 27276 14240 27328
rect 15200 27276 15252 27328
rect 17684 27276 17736 27328
rect 23204 27276 23256 27328
rect 24676 27319 24728 27328
rect 24676 27285 24685 27319
rect 24685 27285 24719 27319
rect 24719 27285 24728 27319
rect 24676 27276 24728 27285
rect 28632 27276 28684 27328
rect 32404 27415 32410 27442
rect 32410 27415 32444 27442
rect 32444 27415 32456 27442
rect 32404 27390 32456 27415
rect 34060 27480 34112 27532
rect 34520 27480 34572 27532
rect 32772 27412 32824 27464
rect 33324 27387 33376 27396
rect 33324 27353 33333 27387
rect 33333 27353 33367 27387
rect 33367 27353 33376 27387
rect 33324 27344 33376 27353
rect 34704 27276 34756 27328
rect 35348 27412 35400 27464
rect 35992 27412 36044 27464
rect 38108 27548 38160 27600
rect 47032 27480 47084 27532
rect 48228 27480 48280 27532
rect 46664 27344 46716 27396
rect 46940 27276 46992 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 2136 27115 2188 27124
rect 2136 27081 2145 27115
rect 2145 27081 2179 27115
rect 2179 27081 2188 27115
rect 2136 27072 2188 27081
rect 9496 27072 9548 27124
rect 1400 27004 1452 27056
rect 10324 27072 10376 27124
rect 10416 27004 10468 27056
rect 14188 27047 14240 27056
rect 14188 27013 14197 27047
rect 14197 27013 14231 27047
rect 14231 27013 14240 27047
rect 14188 27004 14240 27013
rect 8668 26979 8720 26988
rect 8668 26945 8677 26979
rect 8677 26945 8711 26979
rect 8711 26945 8720 26979
rect 8668 26936 8720 26945
rect 8852 26979 8904 26988
rect 8852 26945 8861 26979
rect 8861 26945 8895 26979
rect 8895 26945 8904 26979
rect 8852 26936 8904 26945
rect 9036 26979 9088 26988
rect 9036 26945 9045 26979
rect 9045 26945 9079 26979
rect 9079 26945 9088 26979
rect 9036 26936 9088 26945
rect 10692 26979 10744 26988
rect 2504 26868 2556 26920
rect 2320 26800 2372 26852
rect 9128 26868 9180 26920
rect 10692 26945 10701 26979
rect 10701 26945 10735 26979
rect 10735 26945 10744 26979
rect 10692 26936 10744 26945
rect 10876 26979 10928 26988
rect 10876 26945 10885 26979
rect 10885 26945 10919 26979
rect 10919 26945 10928 26979
rect 10876 26936 10928 26945
rect 15384 27072 15436 27124
rect 22928 27115 22980 27124
rect 22928 27081 22937 27115
rect 22937 27081 22971 27115
rect 22971 27081 22980 27115
rect 22928 27072 22980 27081
rect 14556 27004 14608 27056
rect 1400 26732 1452 26784
rect 9680 26800 9732 26852
rect 10600 26868 10652 26920
rect 19524 26936 19576 26988
rect 23204 26979 23256 26988
rect 23204 26945 23213 26979
rect 23213 26945 23247 26979
rect 23247 26945 23256 26979
rect 23204 26936 23256 26945
rect 24860 27072 24912 27124
rect 24676 27004 24728 27056
rect 24768 27004 24820 27056
rect 30564 27072 30616 27124
rect 34704 27072 34756 27124
rect 36084 27072 36136 27124
rect 33692 27004 33744 27056
rect 46388 27004 46440 27056
rect 27068 26979 27120 26988
rect 15016 26868 15068 26920
rect 20996 26868 21048 26920
rect 27068 26945 27077 26979
rect 27077 26945 27111 26979
rect 27111 26945 27120 26979
rect 27068 26936 27120 26945
rect 32680 26979 32732 26988
rect 32680 26945 32689 26979
rect 32689 26945 32723 26979
rect 32723 26945 32732 26979
rect 32680 26936 32732 26945
rect 27252 26911 27304 26920
rect 27252 26877 27261 26911
rect 27261 26877 27295 26911
rect 27295 26877 27304 26911
rect 27252 26868 27304 26877
rect 28080 26911 28132 26920
rect 28080 26877 28089 26911
rect 28089 26877 28123 26911
rect 28123 26877 28132 26911
rect 28080 26868 28132 26877
rect 29920 26911 29972 26920
rect 7564 26732 7616 26784
rect 9864 26732 9916 26784
rect 10048 26800 10100 26852
rect 26332 26800 26384 26852
rect 26424 26800 26476 26852
rect 29920 26877 29929 26911
rect 29929 26877 29963 26911
rect 29963 26877 29972 26911
rect 29920 26868 29972 26877
rect 32864 26979 32916 26988
rect 32864 26945 32873 26979
rect 32873 26945 32907 26979
rect 32907 26945 32916 26979
rect 32864 26936 32916 26945
rect 33140 26936 33192 26988
rect 10508 26732 10560 26784
rect 14096 26732 14148 26784
rect 14280 26775 14332 26784
rect 14280 26741 14289 26775
rect 14289 26741 14323 26775
rect 14323 26741 14332 26775
rect 14280 26732 14332 26741
rect 15108 26732 15160 26784
rect 21088 26732 21140 26784
rect 32220 26732 32272 26784
rect 32404 26775 32456 26784
rect 32404 26741 32413 26775
rect 32413 26741 32447 26775
rect 32447 26741 32456 26775
rect 32404 26732 32456 26741
rect 32956 26868 33008 26920
rect 34336 26979 34388 26988
rect 33232 26800 33284 26852
rect 34336 26945 34345 26979
rect 34345 26945 34379 26979
rect 34379 26945 34388 26979
rect 34336 26936 34388 26945
rect 35072 26979 35124 26988
rect 35072 26945 35081 26979
rect 35081 26945 35115 26979
rect 35115 26945 35124 26979
rect 35072 26936 35124 26945
rect 34244 26868 34296 26920
rect 35992 26936 36044 26988
rect 36084 26979 36136 26988
rect 36084 26945 36093 26979
rect 36093 26945 36127 26979
rect 36127 26945 36136 26979
rect 36084 26936 36136 26945
rect 32772 26732 32824 26784
rect 32864 26732 32916 26784
rect 35532 26800 35584 26852
rect 34612 26732 34664 26784
rect 35440 26732 35492 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 6184 26571 6236 26580
rect 6184 26537 6193 26571
rect 6193 26537 6227 26571
rect 6227 26537 6236 26571
rect 6184 26528 6236 26537
rect 9772 26571 9824 26580
rect 9312 26460 9364 26512
rect 9772 26537 9781 26571
rect 9781 26537 9815 26571
rect 9815 26537 9824 26571
rect 9772 26528 9824 26537
rect 10600 26503 10652 26512
rect 10600 26469 10609 26503
rect 10609 26469 10643 26503
rect 10643 26469 10652 26503
rect 10600 26460 10652 26469
rect 12072 26503 12124 26512
rect 12072 26469 12081 26503
rect 12081 26469 12115 26503
rect 12115 26469 12124 26503
rect 12072 26460 12124 26469
rect 14832 26460 14884 26512
rect 18144 26460 18196 26512
rect 1400 26435 1452 26444
rect 1400 26401 1409 26435
rect 1409 26401 1443 26435
rect 1443 26401 1452 26435
rect 1400 26392 1452 26401
rect 2780 26435 2832 26444
rect 2780 26401 2789 26435
rect 2789 26401 2823 26435
rect 2823 26401 2832 26435
rect 6276 26435 6328 26444
rect 2780 26392 2832 26401
rect 6276 26401 6285 26435
rect 6285 26401 6319 26435
rect 6319 26401 6328 26435
rect 6276 26392 6328 26401
rect 7564 26392 7616 26444
rect 9220 26392 9272 26444
rect 6460 26367 6512 26376
rect 6460 26333 6469 26367
rect 6469 26333 6503 26367
rect 6503 26333 6512 26367
rect 6460 26324 6512 26333
rect 1584 26299 1636 26308
rect 1584 26265 1593 26299
rect 1593 26265 1627 26299
rect 1627 26265 1636 26299
rect 1584 26256 1636 26265
rect 6368 26256 6420 26308
rect 9220 26256 9272 26308
rect 10324 26324 10376 26376
rect 10876 26324 10928 26376
rect 12348 26367 12400 26376
rect 12348 26333 12357 26367
rect 12357 26333 12391 26367
rect 12391 26333 12400 26367
rect 12348 26324 12400 26333
rect 14096 26367 14148 26376
rect 14096 26333 14105 26367
rect 14105 26333 14139 26367
rect 14139 26333 14148 26367
rect 14096 26324 14148 26333
rect 14372 26367 14424 26376
rect 14372 26333 14381 26367
rect 14381 26333 14415 26367
rect 14415 26333 14424 26367
rect 14372 26324 14424 26333
rect 15200 26324 15252 26376
rect 15292 26367 15344 26376
rect 15292 26333 15301 26367
rect 15301 26333 15335 26367
rect 15335 26333 15344 26367
rect 15292 26324 15344 26333
rect 17592 26324 17644 26376
rect 19524 26528 19576 26580
rect 27252 26528 27304 26580
rect 29920 26571 29972 26580
rect 29920 26537 29929 26571
rect 29929 26537 29963 26571
rect 29963 26537 29972 26571
rect 29920 26528 29972 26537
rect 34336 26528 34388 26580
rect 35992 26528 36044 26580
rect 38936 26571 38988 26580
rect 38936 26537 38945 26571
rect 38945 26537 38979 26571
rect 38979 26537 38988 26571
rect 38936 26528 38988 26537
rect 37280 26460 37332 26512
rect 19524 26367 19576 26376
rect 10140 26256 10192 26308
rect 1952 26188 2004 26240
rect 5724 26188 5776 26240
rect 10692 26256 10744 26308
rect 12164 26256 12216 26308
rect 15016 26256 15068 26308
rect 12256 26231 12308 26240
rect 12256 26197 12265 26231
rect 12265 26197 12299 26231
rect 12299 26197 12308 26231
rect 12256 26188 12308 26197
rect 14280 26231 14332 26240
rect 14280 26197 14289 26231
rect 14289 26197 14323 26231
rect 14323 26197 14332 26231
rect 14280 26188 14332 26197
rect 15384 26256 15436 26308
rect 16948 26188 17000 26240
rect 18144 26188 18196 26240
rect 19524 26333 19533 26367
rect 19533 26333 19567 26367
rect 19567 26333 19576 26367
rect 19524 26324 19576 26333
rect 20076 26324 20128 26376
rect 23572 26392 23624 26444
rect 32864 26392 32916 26444
rect 24768 26324 24820 26376
rect 27436 26324 27488 26376
rect 29828 26367 29880 26376
rect 29828 26333 29837 26367
rect 29837 26333 29871 26367
rect 29871 26333 29880 26367
rect 29828 26324 29880 26333
rect 30748 26367 30800 26376
rect 30748 26333 30757 26367
rect 30757 26333 30791 26367
rect 30791 26333 30800 26367
rect 30748 26324 30800 26333
rect 19156 26256 19208 26308
rect 20260 26256 20312 26308
rect 26332 26256 26384 26308
rect 31116 26299 31168 26308
rect 31116 26265 31125 26299
rect 31125 26265 31159 26299
rect 31159 26265 31168 26299
rect 31116 26256 31168 26265
rect 31208 26256 31260 26308
rect 34336 26256 34388 26308
rect 34520 26324 34572 26376
rect 35348 26367 35400 26376
rect 35348 26333 35357 26367
rect 35357 26333 35391 26367
rect 35391 26333 35400 26367
rect 35348 26324 35400 26333
rect 35440 26324 35492 26376
rect 37372 26324 37424 26376
rect 35256 26256 35308 26308
rect 47952 26299 48004 26308
rect 47952 26265 47961 26299
rect 47961 26265 47995 26299
rect 47995 26265 48004 26299
rect 47952 26256 48004 26265
rect 48044 26256 48096 26308
rect 19432 26188 19484 26240
rect 20536 26188 20588 26240
rect 20812 26188 20864 26240
rect 30196 26188 30248 26240
rect 30380 26188 30432 26240
rect 36544 26188 36596 26240
rect 38292 26188 38344 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 1584 25984 1636 26036
rect 1584 25891 1636 25900
rect 1584 25857 1593 25891
rect 1593 25857 1627 25891
rect 1627 25857 1636 25891
rect 1584 25848 1636 25857
rect 2504 25848 2556 25900
rect 12900 25984 12952 26036
rect 13268 25984 13320 26036
rect 17960 25984 18012 26036
rect 18052 25984 18104 26036
rect 19064 25984 19116 26036
rect 20260 25984 20312 26036
rect 5724 25916 5776 25968
rect 19892 25916 19944 25968
rect 22928 25959 22980 25968
rect 22928 25925 22937 25959
rect 22937 25925 22971 25959
rect 22971 25925 22980 25959
rect 22928 25916 22980 25925
rect 23940 25984 23992 26036
rect 24400 25984 24452 26036
rect 24676 25984 24728 26036
rect 30380 25984 30432 26036
rect 31760 25984 31812 26036
rect 32128 25984 32180 26036
rect 32588 25984 32640 26036
rect 33324 25984 33376 26036
rect 6184 25712 6236 25764
rect 10324 25848 10376 25900
rect 7012 25823 7064 25832
rect 7012 25789 7021 25823
rect 7021 25789 7055 25823
rect 7055 25789 7064 25823
rect 7012 25780 7064 25789
rect 8668 25823 8720 25832
rect 8668 25789 8677 25823
rect 8677 25789 8711 25823
rect 8711 25789 8720 25823
rect 8668 25780 8720 25789
rect 10140 25780 10192 25832
rect 11060 25780 11112 25832
rect 12532 25848 12584 25900
rect 13544 25848 13596 25900
rect 14556 25891 14608 25900
rect 14556 25857 14565 25891
rect 14565 25857 14599 25891
rect 14599 25857 14608 25891
rect 14556 25848 14608 25857
rect 14832 25891 14884 25900
rect 14832 25857 14841 25891
rect 14841 25857 14875 25891
rect 14875 25857 14884 25891
rect 14832 25848 14884 25857
rect 16948 25891 17000 25900
rect 16948 25857 16982 25891
rect 16982 25857 17000 25891
rect 16948 25848 17000 25857
rect 17960 25848 18012 25900
rect 18880 25848 18932 25900
rect 19064 25891 19116 25900
rect 19064 25857 19073 25891
rect 19073 25857 19107 25891
rect 19107 25857 19116 25891
rect 19064 25848 19116 25857
rect 13636 25823 13688 25832
rect 8392 25712 8444 25764
rect 9588 25644 9640 25696
rect 10876 25644 10928 25696
rect 12072 25644 12124 25696
rect 13268 25644 13320 25696
rect 13636 25789 13645 25823
rect 13645 25789 13679 25823
rect 13679 25789 13688 25823
rect 13636 25780 13688 25789
rect 16672 25823 16724 25832
rect 16672 25789 16681 25823
rect 16681 25789 16715 25823
rect 16715 25789 16724 25823
rect 16672 25780 16724 25789
rect 18144 25780 18196 25832
rect 19248 25891 19300 25900
rect 19248 25857 19257 25891
rect 19257 25857 19291 25891
rect 19291 25857 19300 25891
rect 19248 25848 19300 25857
rect 19432 25891 19484 25900
rect 19432 25857 19441 25891
rect 19441 25857 19475 25891
rect 19475 25857 19484 25891
rect 19432 25848 19484 25857
rect 20260 25848 20312 25900
rect 20536 25891 20588 25900
rect 20536 25857 20545 25891
rect 20545 25857 20579 25891
rect 20579 25857 20588 25891
rect 20536 25848 20588 25857
rect 20720 25891 20772 25900
rect 20720 25857 20729 25891
rect 20729 25857 20763 25891
rect 20763 25857 20772 25891
rect 20720 25848 20772 25857
rect 23848 25891 23900 25900
rect 20812 25780 20864 25832
rect 23112 25823 23164 25832
rect 23112 25789 23121 25823
rect 23121 25789 23155 25823
rect 23155 25789 23164 25823
rect 23112 25780 23164 25789
rect 14464 25644 14516 25696
rect 17040 25644 17092 25696
rect 19984 25712 20036 25764
rect 18052 25687 18104 25696
rect 18052 25653 18061 25687
rect 18061 25653 18095 25687
rect 18095 25653 18104 25687
rect 18052 25644 18104 25653
rect 18788 25687 18840 25696
rect 18788 25653 18797 25687
rect 18797 25653 18831 25687
rect 18831 25653 18840 25687
rect 18788 25644 18840 25653
rect 19892 25644 19944 25696
rect 23848 25857 23857 25891
rect 23857 25857 23891 25891
rect 23891 25857 23900 25891
rect 23848 25848 23900 25857
rect 24032 25848 24084 25900
rect 24308 25848 24360 25900
rect 25964 25848 26016 25900
rect 27988 25916 28040 25968
rect 29828 25916 29880 25968
rect 34520 25984 34572 26036
rect 35256 25984 35308 26036
rect 35624 26027 35676 26036
rect 35624 25993 35633 26027
rect 35633 25993 35667 26027
rect 35667 25993 35676 26027
rect 35624 25984 35676 25993
rect 36544 25984 36596 26036
rect 46848 25984 46900 26036
rect 23940 25644 23992 25696
rect 24124 25687 24176 25696
rect 24124 25653 24133 25687
rect 24133 25653 24167 25687
rect 24167 25653 24176 25687
rect 24124 25644 24176 25653
rect 24768 25687 24820 25696
rect 24768 25653 24777 25687
rect 24777 25653 24811 25687
rect 24811 25653 24820 25687
rect 24768 25644 24820 25653
rect 24860 25644 24912 25696
rect 25228 25687 25280 25696
rect 25228 25653 25237 25687
rect 25237 25653 25271 25687
rect 25271 25653 25280 25687
rect 25228 25644 25280 25653
rect 30748 25848 30800 25900
rect 30104 25823 30156 25832
rect 30104 25789 30113 25823
rect 30113 25789 30147 25823
rect 30147 25789 30156 25823
rect 32220 25848 32272 25900
rect 30104 25780 30156 25789
rect 32128 25780 32180 25832
rect 32404 25848 32456 25900
rect 34612 25916 34664 25968
rect 38292 25959 38344 25968
rect 38292 25925 38301 25959
rect 38301 25925 38335 25959
rect 38335 25925 38344 25959
rect 38292 25916 38344 25925
rect 38108 25891 38160 25900
rect 38108 25857 38117 25891
rect 38117 25857 38151 25891
rect 38151 25857 38160 25891
rect 38108 25848 38160 25857
rect 46480 25916 46532 25968
rect 46848 25891 46900 25900
rect 46848 25857 46857 25891
rect 46857 25857 46891 25891
rect 46891 25857 46900 25891
rect 46848 25848 46900 25857
rect 48504 25780 48556 25832
rect 36544 25644 36596 25696
rect 45192 25644 45244 25696
rect 47768 25687 47820 25696
rect 47768 25653 47777 25687
rect 47777 25653 47811 25687
rect 47811 25653 47820 25687
rect 47768 25644 47820 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 7012 25483 7064 25492
rect 7012 25449 7021 25483
rect 7021 25449 7055 25483
rect 7055 25449 7064 25483
rect 7012 25440 7064 25449
rect 9312 25440 9364 25492
rect 9956 25483 10008 25492
rect 9956 25449 9965 25483
rect 9965 25449 9999 25483
rect 9999 25449 10008 25483
rect 9956 25440 10008 25449
rect 10140 25483 10192 25492
rect 10140 25449 10149 25483
rect 10149 25449 10183 25483
rect 10183 25449 10192 25483
rect 10140 25440 10192 25449
rect 11060 25483 11112 25492
rect 11060 25449 11069 25483
rect 11069 25449 11103 25483
rect 11103 25449 11112 25483
rect 11060 25440 11112 25449
rect 12256 25440 12308 25492
rect 12532 25483 12584 25492
rect 12532 25449 12541 25483
rect 12541 25449 12575 25483
rect 12575 25449 12584 25483
rect 12532 25440 12584 25449
rect 14280 25483 14332 25492
rect 14280 25449 14289 25483
rect 14289 25449 14323 25483
rect 14323 25449 14332 25483
rect 14280 25440 14332 25449
rect 14464 25483 14516 25492
rect 14464 25449 14473 25483
rect 14473 25449 14507 25483
rect 14507 25449 14516 25483
rect 14464 25440 14516 25449
rect 14556 25440 14608 25492
rect 19524 25440 19576 25492
rect 23572 25483 23624 25492
rect 23572 25449 23581 25483
rect 23581 25449 23615 25483
rect 23615 25449 23624 25483
rect 23572 25440 23624 25449
rect 23756 25483 23808 25492
rect 23756 25449 23765 25483
rect 23765 25449 23799 25483
rect 23799 25449 23808 25483
rect 23756 25440 23808 25449
rect 6644 25236 6696 25288
rect 6920 25279 6972 25288
rect 6920 25245 6929 25279
rect 6929 25245 6963 25279
rect 6963 25245 6972 25279
rect 6920 25236 6972 25245
rect 9312 25347 9364 25356
rect 9312 25313 9321 25347
rect 9321 25313 9355 25347
rect 9355 25313 9364 25347
rect 9312 25304 9364 25313
rect 21180 25372 21232 25424
rect 10692 25347 10744 25356
rect 10692 25313 10701 25347
rect 10701 25313 10735 25347
rect 10735 25313 10744 25347
rect 10692 25304 10744 25313
rect 10876 25304 10928 25356
rect 17040 25304 17092 25356
rect 18236 25304 18288 25356
rect 30104 25440 30156 25492
rect 30196 25440 30248 25492
rect 38108 25483 38160 25492
rect 23940 25372 23992 25424
rect 36544 25372 36596 25424
rect 9312 25168 9364 25220
rect 9496 25168 9548 25220
rect 10048 25236 10100 25288
rect 10784 25279 10836 25288
rect 10784 25245 10793 25279
rect 10793 25245 10827 25279
rect 10827 25245 10836 25279
rect 10784 25236 10836 25245
rect 16580 25236 16632 25288
rect 16672 25236 16724 25288
rect 20076 25279 20128 25288
rect 20076 25245 20085 25279
rect 20085 25245 20119 25279
rect 20119 25245 20128 25279
rect 20076 25236 20128 25245
rect 24952 25304 25004 25356
rect 12164 25211 12216 25220
rect 12164 25177 12173 25211
rect 12173 25177 12207 25211
rect 12207 25177 12216 25211
rect 12164 25168 12216 25177
rect 12348 25211 12400 25220
rect 12348 25177 12373 25211
rect 12373 25177 12400 25211
rect 12348 25168 12400 25177
rect 14188 25168 14240 25220
rect 14372 25168 14424 25220
rect 18788 25168 18840 25220
rect 19156 25168 19208 25220
rect 19524 25168 19576 25220
rect 20168 25168 20220 25220
rect 21272 25236 21324 25288
rect 21916 25236 21968 25288
rect 23388 25211 23440 25220
rect 23388 25177 23397 25211
rect 23397 25177 23431 25211
rect 23431 25177 23440 25211
rect 23388 25168 23440 25177
rect 24124 25236 24176 25288
rect 24400 25279 24452 25288
rect 24400 25245 24409 25279
rect 24409 25245 24443 25279
rect 24443 25245 24452 25279
rect 24400 25236 24452 25245
rect 25320 25279 25372 25288
rect 25320 25245 25329 25279
rect 25329 25245 25363 25279
rect 25363 25245 25372 25279
rect 25320 25236 25372 25245
rect 25964 25304 26016 25356
rect 38108 25449 38117 25483
rect 38117 25449 38151 25483
rect 38151 25449 38160 25483
rect 38108 25440 38160 25449
rect 25596 25236 25648 25288
rect 30748 25236 30800 25288
rect 31484 25236 31536 25288
rect 24676 25168 24728 25220
rect 31668 25168 31720 25220
rect 47768 25304 47820 25356
rect 38016 25279 38068 25288
rect 38016 25245 38025 25279
rect 38025 25245 38059 25279
rect 38059 25245 38068 25279
rect 38016 25236 38068 25245
rect 38292 25279 38344 25288
rect 38292 25245 38301 25279
rect 38301 25245 38335 25279
rect 38335 25245 38344 25279
rect 38292 25236 38344 25245
rect 46480 25211 46532 25220
rect 13084 25143 13136 25152
rect 13084 25109 13093 25143
rect 13093 25109 13127 25143
rect 13127 25109 13136 25143
rect 13084 25100 13136 25109
rect 14832 25100 14884 25152
rect 17960 25100 18012 25152
rect 18236 25100 18288 25152
rect 20536 25100 20588 25152
rect 22468 25100 22520 25152
rect 22928 25100 22980 25152
rect 23572 25143 23624 25152
rect 23572 25109 23581 25143
rect 23581 25109 23615 25143
rect 23615 25109 23624 25143
rect 23572 25100 23624 25109
rect 24400 25100 24452 25152
rect 25136 25100 25188 25152
rect 29828 25100 29880 25152
rect 32772 25143 32824 25152
rect 32772 25109 32781 25143
rect 32781 25109 32815 25143
rect 32815 25109 32824 25143
rect 32772 25100 32824 25109
rect 46480 25177 46489 25211
rect 46489 25177 46523 25211
rect 46523 25177 46532 25211
rect 46480 25168 46532 25177
rect 48136 25211 48188 25220
rect 48136 25177 48145 25211
rect 48145 25177 48179 25211
rect 48179 25177 48188 25211
rect 48136 25168 48188 25177
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 7656 24803 7708 24812
rect 7656 24769 7665 24803
rect 7665 24769 7699 24803
rect 7699 24769 7708 24803
rect 7656 24760 7708 24769
rect 2228 24692 2280 24744
rect 11520 24896 11572 24948
rect 14372 24896 14424 24948
rect 16580 24896 16632 24948
rect 8484 24828 8536 24880
rect 10048 24828 10100 24880
rect 18236 24871 18288 24880
rect 18236 24837 18245 24871
rect 18245 24837 18279 24871
rect 18279 24837 18288 24871
rect 18236 24828 18288 24837
rect 19248 24896 19300 24948
rect 20168 24896 20220 24948
rect 23572 24896 23624 24948
rect 24676 24896 24728 24948
rect 25504 24896 25556 24948
rect 25688 24896 25740 24948
rect 47492 24896 47544 24948
rect 19892 24828 19944 24880
rect 13268 24760 13320 24812
rect 8760 24735 8812 24744
rect 8760 24701 8769 24735
rect 8769 24701 8803 24735
rect 8803 24701 8812 24735
rect 11520 24735 11572 24744
rect 8760 24692 8812 24701
rect 11520 24701 11529 24735
rect 11529 24701 11563 24735
rect 11563 24701 11572 24735
rect 11520 24692 11572 24701
rect 13084 24692 13136 24744
rect 13360 24735 13412 24744
rect 13360 24701 13369 24735
rect 13369 24701 13403 24735
rect 13403 24701 13412 24735
rect 13360 24692 13412 24701
rect 13728 24760 13780 24812
rect 17408 24803 17460 24812
rect 14188 24692 14240 24744
rect 17408 24769 17417 24803
rect 17417 24769 17451 24803
rect 17451 24769 17460 24803
rect 17408 24760 17460 24769
rect 17684 24760 17736 24812
rect 19156 24760 19208 24812
rect 19432 24760 19484 24812
rect 18420 24692 18472 24744
rect 18788 24692 18840 24744
rect 1584 24556 1636 24608
rect 12256 24556 12308 24608
rect 13452 24556 13504 24608
rect 13544 24556 13596 24608
rect 15108 24556 15160 24608
rect 17408 24624 17460 24676
rect 18052 24624 18104 24676
rect 20536 24803 20588 24812
rect 20536 24769 20545 24803
rect 20545 24769 20579 24803
rect 20579 24769 20588 24803
rect 20536 24760 20588 24769
rect 20720 24803 20772 24812
rect 20720 24769 20729 24803
rect 20729 24769 20763 24803
rect 20763 24769 20772 24803
rect 20720 24760 20772 24769
rect 21824 24760 21876 24812
rect 24860 24828 24912 24880
rect 20812 24692 20864 24744
rect 21916 24624 21968 24676
rect 23940 24803 23992 24812
rect 22744 24692 22796 24744
rect 23940 24769 23949 24803
rect 23949 24769 23983 24803
rect 23983 24769 23992 24803
rect 23940 24760 23992 24769
rect 24952 24760 25004 24812
rect 27160 24760 27212 24812
rect 25228 24692 25280 24744
rect 21548 24556 21600 24608
rect 21824 24599 21876 24608
rect 21824 24565 21833 24599
rect 21833 24565 21867 24599
rect 21867 24565 21876 24599
rect 21824 24556 21876 24565
rect 23480 24556 23532 24608
rect 24584 24624 24636 24676
rect 26700 24624 26752 24676
rect 27436 24803 27488 24812
rect 27436 24769 27445 24803
rect 27445 24769 27479 24803
rect 27479 24769 27488 24803
rect 27436 24760 27488 24769
rect 27620 24803 27672 24812
rect 27620 24769 27629 24803
rect 27629 24769 27663 24803
rect 27663 24769 27672 24803
rect 27620 24760 27672 24769
rect 28908 24760 28960 24812
rect 29276 24828 29328 24880
rect 31484 24871 31536 24880
rect 31484 24837 31493 24871
rect 31493 24837 31527 24871
rect 31527 24837 31536 24871
rect 31484 24828 31536 24837
rect 29368 24760 29420 24812
rect 30196 24760 30248 24812
rect 30380 24760 30432 24812
rect 32220 24760 32272 24812
rect 33140 24760 33192 24812
rect 33324 24760 33376 24812
rect 36544 24803 36596 24812
rect 36544 24769 36553 24803
rect 36553 24769 36587 24803
rect 36587 24769 36596 24803
rect 36544 24760 36596 24769
rect 39120 24803 39172 24812
rect 39120 24769 39129 24803
rect 39129 24769 39163 24803
rect 39163 24769 39172 24803
rect 39120 24760 39172 24769
rect 47952 24803 48004 24812
rect 47952 24769 47961 24803
rect 47961 24769 47995 24803
rect 47995 24769 48004 24803
rect 47952 24760 48004 24769
rect 29276 24624 29328 24676
rect 29552 24692 29604 24744
rect 34796 24692 34848 24744
rect 35440 24735 35492 24744
rect 35440 24701 35449 24735
rect 35449 24701 35483 24735
rect 35483 24701 35492 24735
rect 35440 24692 35492 24701
rect 35624 24692 35676 24744
rect 25320 24556 25372 24608
rect 27068 24556 27120 24608
rect 29828 24556 29880 24608
rect 32496 24556 32548 24608
rect 32772 24556 32824 24608
rect 36544 24556 36596 24608
rect 37372 24556 37424 24608
rect 38568 24556 38620 24608
rect 39120 24556 39172 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 1584 24395 1636 24404
rect 1584 24361 1593 24395
rect 1593 24361 1627 24395
rect 1627 24361 1636 24395
rect 1584 24352 1636 24361
rect 1768 24352 1820 24404
rect 10692 24352 10744 24404
rect 12348 24352 12400 24404
rect 13268 24395 13320 24404
rect 13268 24361 13277 24395
rect 13277 24361 13311 24395
rect 13311 24361 13320 24395
rect 13268 24352 13320 24361
rect 13452 24395 13504 24404
rect 13452 24361 13461 24395
rect 13461 24361 13495 24395
rect 13495 24361 13504 24395
rect 13452 24352 13504 24361
rect 13728 24352 13780 24404
rect 14648 24352 14700 24404
rect 22652 24395 22704 24404
rect 22652 24361 22661 24395
rect 22661 24361 22695 24395
rect 22695 24361 22704 24395
rect 22652 24352 22704 24361
rect 32772 24352 32824 24404
rect 34796 24395 34848 24404
rect 34796 24361 34805 24395
rect 34805 24361 34839 24395
rect 34839 24361 34848 24395
rect 34796 24352 34848 24361
rect 8208 24216 8260 24268
rect 12256 24216 12308 24268
rect 13912 24216 13964 24268
rect 18144 24259 18196 24268
rect 18144 24225 18153 24259
rect 18153 24225 18187 24259
rect 18187 24225 18196 24259
rect 18144 24216 18196 24225
rect 23296 24284 23348 24336
rect 23940 24284 23992 24336
rect 29184 24284 29236 24336
rect 32680 24284 32732 24336
rect 43996 24284 44048 24336
rect 1400 24191 1452 24200
rect 1400 24157 1409 24191
rect 1409 24157 1443 24191
rect 1443 24157 1452 24191
rect 1400 24148 1452 24157
rect 8852 24148 8904 24200
rect 9956 24148 10008 24200
rect 4068 24080 4120 24132
rect 3056 24012 3108 24064
rect 12256 24080 12308 24132
rect 12900 24148 12952 24200
rect 12992 24123 13044 24132
rect 12992 24089 13001 24123
rect 13001 24089 13035 24123
rect 13035 24089 13044 24123
rect 14188 24148 14240 24200
rect 16948 24148 17000 24200
rect 17868 24191 17920 24200
rect 17868 24157 17877 24191
rect 17877 24157 17911 24191
rect 17911 24157 17920 24191
rect 17868 24148 17920 24157
rect 19156 24148 19208 24200
rect 22192 24148 22244 24200
rect 22744 24148 22796 24200
rect 23664 24148 23716 24200
rect 24584 24191 24636 24200
rect 24584 24157 24593 24191
rect 24593 24157 24627 24191
rect 24627 24157 24636 24191
rect 24584 24148 24636 24157
rect 24676 24191 24728 24200
rect 24676 24157 24685 24191
rect 24685 24157 24719 24191
rect 24719 24157 24728 24191
rect 25136 24191 25188 24200
rect 24676 24148 24728 24157
rect 25136 24157 25145 24191
rect 25145 24157 25179 24191
rect 25179 24157 25188 24191
rect 25136 24148 25188 24157
rect 25596 24148 25648 24200
rect 26608 24216 26660 24268
rect 26792 24259 26844 24268
rect 26792 24225 26801 24259
rect 26801 24225 26835 24259
rect 26835 24225 26844 24259
rect 26792 24216 26844 24225
rect 32496 24259 32548 24268
rect 32496 24225 32505 24259
rect 32505 24225 32539 24259
rect 32539 24225 32548 24259
rect 32496 24216 32548 24225
rect 33140 24216 33192 24268
rect 37280 24259 37332 24268
rect 26240 24148 26292 24200
rect 26332 24191 26384 24200
rect 26332 24157 26341 24191
rect 26341 24157 26375 24191
rect 26375 24157 26384 24191
rect 29552 24191 29604 24200
rect 26332 24148 26384 24157
rect 29552 24157 29561 24191
rect 29561 24157 29595 24191
rect 29595 24157 29604 24191
rect 29552 24148 29604 24157
rect 29828 24191 29880 24200
rect 29828 24157 29862 24191
rect 29862 24157 29880 24191
rect 32312 24191 32364 24200
rect 29828 24148 29880 24157
rect 32312 24157 32321 24191
rect 32321 24157 32355 24191
rect 32355 24157 32364 24191
rect 32312 24148 32364 24157
rect 37280 24225 37289 24259
rect 37289 24225 37323 24259
rect 37323 24225 37332 24259
rect 37280 24216 37332 24225
rect 46940 24216 46992 24268
rect 47308 24191 47360 24200
rect 47308 24157 47317 24191
rect 47317 24157 47351 24191
rect 47351 24157 47360 24191
rect 47308 24148 47360 24157
rect 21364 24123 21416 24132
rect 12992 24080 13044 24089
rect 21364 24089 21373 24123
rect 21373 24089 21407 24123
rect 21407 24089 21416 24123
rect 21364 24080 21416 24089
rect 21548 24080 21600 24132
rect 23848 24080 23900 24132
rect 14280 24012 14332 24064
rect 17592 24012 17644 24064
rect 20168 24012 20220 24064
rect 28448 24080 28500 24132
rect 37464 24123 37516 24132
rect 27988 24012 28040 24064
rect 28172 24055 28224 24064
rect 28172 24021 28181 24055
rect 28181 24021 28215 24055
rect 28215 24021 28224 24055
rect 28172 24012 28224 24021
rect 28540 24012 28592 24064
rect 37464 24089 37473 24123
rect 37473 24089 37507 24123
rect 37507 24089 37516 24123
rect 37464 24080 37516 24089
rect 39120 24123 39172 24132
rect 39120 24089 39129 24123
rect 39129 24089 39163 24123
rect 39163 24089 39172 24123
rect 39120 24080 39172 24089
rect 38660 24012 38712 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 4712 23808 4764 23860
rect 8300 23740 8352 23792
rect 17592 23740 17644 23792
rect 19156 23808 19208 23860
rect 27160 23808 27212 23860
rect 27988 23808 28040 23860
rect 30472 23808 30524 23860
rect 37464 23851 37516 23860
rect 8944 23672 8996 23724
rect 12992 23672 13044 23724
rect 13912 23715 13964 23724
rect 13912 23681 13921 23715
rect 13921 23681 13955 23715
rect 13955 23681 13964 23715
rect 14648 23715 14700 23724
rect 13912 23672 13964 23681
rect 14648 23681 14657 23715
rect 14657 23681 14691 23715
rect 14691 23681 14700 23715
rect 14648 23672 14700 23681
rect 15108 23604 15160 23656
rect 11520 23536 11572 23588
rect 17592 23604 17644 23656
rect 17960 23536 18012 23588
rect 19248 23672 19300 23724
rect 19432 23604 19484 23656
rect 2044 23511 2096 23520
rect 2044 23477 2053 23511
rect 2053 23477 2087 23511
rect 2087 23477 2096 23511
rect 2044 23468 2096 23477
rect 8208 23468 8260 23520
rect 13544 23468 13596 23520
rect 13728 23468 13780 23520
rect 14740 23511 14792 23520
rect 14740 23477 14749 23511
rect 14749 23477 14783 23511
rect 14783 23477 14792 23511
rect 14740 23468 14792 23477
rect 16856 23468 16908 23520
rect 17684 23468 17736 23520
rect 20168 23536 20220 23588
rect 23112 23536 23164 23588
rect 23480 23740 23532 23792
rect 25964 23740 26016 23792
rect 29000 23740 29052 23792
rect 31024 23740 31076 23792
rect 37464 23817 37473 23851
rect 37473 23817 37507 23851
rect 37507 23817 37516 23851
rect 37464 23808 37516 23817
rect 32404 23740 32456 23792
rect 48044 23740 48096 23792
rect 23664 23715 23716 23724
rect 23664 23681 23673 23715
rect 23673 23681 23707 23715
rect 23707 23681 23716 23715
rect 23664 23672 23716 23681
rect 24952 23672 25004 23724
rect 26700 23672 26752 23724
rect 26792 23672 26844 23724
rect 27068 23672 27120 23724
rect 28448 23672 28500 23724
rect 29552 23672 29604 23724
rect 37372 23715 37424 23724
rect 37372 23681 37381 23715
rect 37381 23681 37415 23715
rect 37415 23681 37424 23715
rect 37372 23672 37424 23681
rect 25136 23604 25188 23656
rect 25228 23536 25280 23588
rect 23388 23511 23440 23520
rect 23388 23477 23397 23511
rect 23397 23477 23431 23511
rect 23431 23477 23440 23511
rect 23388 23468 23440 23477
rect 23480 23468 23532 23520
rect 24676 23511 24728 23520
rect 24676 23477 24685 23511
rect 24685 23477 24719 23511
rect 24719 23477 24728 23511
rect 24676 23468 24728 23477
rect 24860 23511 24912 23520
rect 24860 23477 24869 23511
rect 24869 23477 24903 23511
rect 24903 23477 24912 23511
rect 24860 23468 24912 23477
rect 25044 23468 25096 23520
rect 27988 23604 28040 23656
rect 29092 23604 29144 23656
rect 29736 23647 29788 23656
rect 29736 23613 29745 23647
rect 29745 23613 29779 23647
rect 29779 23613 29788 23647
rect 29736 23604 29788 23613
rect 33232 23647 33284 23656
rect 33232 23613 33241 23647
rect 33241 23613 33275 23647
rect 33275 23613 33284 23647
rect 33232 23604 33284 23613
rect 33416 23647 33468 23656
rect 33416 23613 33425 23647
rect 33425 23613 33459 23647
rect 33459 23613 33468 23647
rect 33416 23604 33468 23613
rect 40040 23604 40092 23656
rect 28632 23536 28684 23588
rect 27896 23468 27948 23520
rect 29644 23468 29696 23520
rect 47676 23468 47728 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 1584 23196 1636 23248
rect 23020 23264 23072 23316
rect 23112 23264 23164 23316
rect 8944 23239 8996 23248
rect 8944 23205 8953 23239
rect 8953 23205 8987 23239
rect 8987 23205 8996 23239
rect 8944 23196 8996 23205
rect 9312 23196 9364 23248
rect 12072 23196 12124 23248
rect 2044 23128 2096 23180
rect 2780 23171 2832 23180
rect 2780 23137 2789 23171
rect 2789 23137 2823 23171
rect 2823 23137 2832 23171
rect 15108 23196 15160 23248
rect 16948 23196 17000 23248
rect 19984 23196 20036 23248
rect 20260 23196 20312 23248
rect 22192 23239 22244 23248
rect 22192 23205 22201 23239
rect 22201 23205 22235 23239
rect 22235 23205 22244 23239
rect 22192 23196 22244 23205
rect 23204 23196 23256 23248
rect 23572 23264 23624 23316
rect 25044 23264 25096 23316
rect 26240 23264 26292 23316
rect 27712 23264 27764 23316
rect 28264 23264 28316 23316
rect 29552 23307 29604 23316
rect 29552 23273 29561 23307
rect 29561 23273 29595 23307
rect 29595 23273 29604 23307
rect 29552 23264 29604 23273
rect 29736 23264 29788 23316
rect 32128 23264 32180 23316
rect 33416 23264 33468 23316
rect 47860 23307 47912 23316
rect 47860 23273 47869 23307
rect 47869 23273 47903 23307
rect 47903 23273 47912 23307
rect 47860 23264 47912 23273
rect 24768 23196 24820 23248
rect 2780 23128 2832 23137
rect 8208 23103 8260 23112
rect 8208 23069 8217 23103
rect 8217 23069 8251 23103
rect 8251 23069 8260 23103
rect 8208 23060 8260 23069
rect 8852 23060 8904 23112
rect 2320 22992 2372 23044
rect 8024 23035 8076 23044
rect 8024 23001 8033 23035
rect 8033 23001 8067 23035
rect 8067 23001 8076 23035
rect 8024 22992 8076 23001
rect 8392 23035 8444 23044
rect 8392 23001 8401 23035
rect 8401 23001 8435 23035
rect 8435 23001 8444 23035
rect 8392 22992 8444 23001
rect 9772 23060 9824 23112
rect 11796 23060 11848 23112
rect 11980 23103 12032 23112
rect 11980 23069 11989 23103
rect 11989 23069 12023 23103
rect 12023 23069 12032 23103
rect 11980 23060 12032 23069
rect 12072 23103 12124 23112
rect 12072 23069 12081 23103
rect 12081 23069 12115 23103
rect 12115 23069 12124 23103
rect 12072 23060 12124 23069
rect 12348 23060 12400 23112
rect 13452 23060 13504 23112
rect 17040 23060 17092 23112
rect 19156 23128 19208 23180
rect 9864 22992 9916 23044
rect 12900 23035 12952 23044
rect 4620 22924 4672 22976
rect 11612 22967 11664 22976
rect 11612 22933 11621 22967
rect 11621 22933 11655 22967
rect 11655 22933 11664 22967
rect 11612 22924 11664 22933
rect 12900 23001 12909 23035
rect 12909 23001 12943 23035
rect 12943 23001 12952 23035
rect 12900 22992 12952 23001
rect 14188 22992 14240 23044
rect 15568 22992 15620 23044
rect 18236 23103 18288 23112
rect 18236 23069 18245 23103
rect 18245 23069 18279 23103
rect 18279 23069 18288 23103
rect 18236 23060 18288 23069
rect 17960 22992 18012 23044
rect 18696 23060 18748 23112
rect 19892 23128 19944 23180
rect 19432 23103 19484 23112
rect 19432 23069 19449 23103
rect 19449 23069 19483 23103
rect 19483 23069 19484 23103
rect 19432 23060 19484 23069
rect 20168 23060 20220 23112
rect 20904 23060 20956 23112
rect 21824 23060 21876 23112
rect 23480 23103 23532 23112
rect 23480 23069 23489 23103
rect 23489 23069 23523 23103
rect 23523 23069 23532 23103
rect 23480 23060 23532 23069
rect 24860 23060 24912 23112
rect 26424 23196 26476 23248
rect 27988 23196 28040 23248
rect 26332 23128 26384 23180
rect 28172 23060 28224 23112
rect 28632 23060 28684 23112
rect 17776 22967 17828 22976
rect 17776 22933 17785 22967
rect 17785 22933 17819 22967
rect 17819 22933 17828 22967
rect 17776 22924 17828 22933
rect 19248 22967 19300 22976
rect 19248 22933 19257 22967
rect 19257 22933 19291 22967
rect 19291 22933 19300 22967
rect 19248 22924 19300 22933
rect 20076 22924 20128 22976
rect 20444 22924 20496 22976
rect 25688 22992 25740 23044
rect 26976 22992 27028 23044
rect 28816 23100 28868 23112
rect 28816 23066 28825 23100
rect 28825 23066 28859 23100
rect 28859 23066 28868 23100
rect 28816 23060 28868 23066
rect 29000 23103 29052 23112
rect 29000 23069 29009 23103
rect 29009 23069 29043 23103
rect 29043 23069 29052 23103
rect 48228 23196 48280 23248
rect 45744 23128 45796 23180
rect 29000 23060 29052 23069
rect 29460 22992 29512 23044
rect 29368 22924 29420 22976
rect 29644 22924 29696 22976
rect 30196 23103 30248 23112
rect 30196 23069 30205 23103
rect 30205 23069 30239 23103
rect 30239 23069 30248 23103
rect 33140 23103 33192 23112
rect 30196 23060 30248 23069
rect 33140 23069 33149 23103
rect 33149 23069 33183 23103
rect 33183 23069 33192 23103
rect 33140 23060 33192 23069
rect 47492 23103 47544 23112
rect 47492 23069 47501 23103
rect 47501 23069 47535 23103
rect 47535 23069 47544 23103
rect 47492 23060 47544 23069
rect 46664 22992 46716 23044
rect 48044 22967 48096 22976
rect 48044 22933 48053 22967
rect 48053 22933 48087 22967
rect 48087 22933 48096 22967
rect 48044 22924 48096 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 1584 22763 1636 22772
rect 1584 22729 1593 22763
rect 1593 22729 1627 22763
rect 1627 22729 1636 22763
rect 1584 22720 1636 22729
rect 2320 22763 2372 22772
rect 2320 22729 2329 22763
rect 2329 22729 2363 22763
rect 2363 22729 2372 22763
rect 2320 22720 2372 22729
rect 8024 22720 8076 22772
rect 1400 22627 1452 22636
rect 1400 22593 1409 22627
rect 1409 22593 1443 22627
rect 1443 22593 1452 22627
rect 1400 22584 1452 22593
rect 2136 22584 2188 22636
rect 8300 22652 8352 22704
rect 8944 22652 8996 22704
rect 11980 22720 12032 22772
rect 14188 22763 14240 22772
rect 8852 22584 8904 22636
rect 11612 22652 11664 22704
rect 13728 22652 13780 22704
rect 14188 22729 14197 22763
rect 14197 22729 14231 22763
rect 14231 22729 14240 22763
rect 14188 22720 14240 22729
rect 14464 22720 14516 22772
rect 14280 22652 14332 22704
rect 15568 22720 15620 22772
rect 15752 22720 15804 22772
rect 16212 22720 16264 22772
rect 11520 22627 11572 22636
rect 11520 22593 11529 22627
rect 11529 22593 11563 22627
rect 11563 22593 11572 22627
rect 11520 22584 11572 22593
rect 13452 22584 13504 22636
rect 14464 22627 14516 22636
rect 14464 22593 14473 22627
rect 14473 22593 14507 22627
rect 14507 22593 14516 22627
rect 14464 22584 14516 22593
rect 8208 22380 8260 22432
rect 9404 22423 9456 22432
rect 9404 22389 9413 22423
rect 9413 22389 9447 22423
rect 9447 22389 9456 22423
rect 9404 22380 9456 22389
rect 10784 22516 10836 22568
rect 15016 22584 15068 22636
rect 15752 22627 15804 22636
rect 15752 22593 15761 22627
rect 15761 22593 15795 22627
rect 15795 22593 15804 22627
rect 15752 22584 15804 22593
rect 15936 22627 15988 22636
rect 15936 22593 15945 22627
rect 15945 22593 15979 22627
rect 15979 22593 15988 22627
rect 15936 22584 15988 22593
rect 16212 22584 16264 22636
rect 17040 22584 17092 22636
rect 17776 22627 17828 22636
rect 17776 22593 17810 22627
rect 17810 22593 17828 22627
rect 17776 22584 17828 22593
rect 19432 22584 19484 22636
rect 21916 22652 21968 22704
rect 23480 22584 23532 22636
rect 24124 22627 24176 22636
rect 24124 22593 24133 22627
rect 24133 22593 24167 22627
rect 24167 22593 24176 22627
rect 24124 22584 24176 22593
rect 26424 22652 26476 22704
rect 27436 22720 27488 22772
rect 28816 22763 28868 22772
rect 28816 22729 28825 22763
rect 28825 22729 28859 22763
rect 28859 22729 28868 22763
rect 28816 22720 28868 22729
rect 41880 22720 41932 22772
rect 47492 22720 47544 22772
rect 25044 22627 25096 22636
rect 12716 22380 12768 22432
rect 12900 22423 12952 22432
rect 12900 22389 12909 22423
rect 12909 22389 12943 22423
rect 12943 22389 12952 22423
rect 12900 22380 12952 22389
rect 17868 22380 17920 22432
rect 18880 22423 18932 22432
rect 18880 22389 18889 22423
rect 18889 22389 18923 22423
rect 18923 22389 18932 22423
rect 18880 22380 18932 22389
rect 23572 22448 23624 22500
rect 25044 22593 25053 22627
rect 25053 22593 25087 22627
rect 25087 22593 25096 22627
rect 25044 22584 25096 22593
rect 26148 22627 26200 22636
rect 26148 22593 26157 22627
rect 26157 22593 26191 22627
rect 26191 22593 26200 22627
rect 26148 22584 26200 22593
rect 26976 22627 27028 22636
rect 26976 22593 26985 22627
rect 26985 22593 27019 22627
rect 27019 22593 27028 22627
rect 26976 22584 27028 22593
rect 27804 22584 27856 22636
rect 28448 22627 28500 22636
rect 28448 22593 28457 22627
rect 28457 22593 28491 22627
rect 28491 22593 28500 22627
rect 29736 22652 29788 22704
rect 30380 22652 30432 22704
rect 28448 22584 28500 22593
rect 25504 22516 25556 22568
rect 24676 22448 24728 22500
rect 20720 22423 20772 22432
rect 20720 22389 20729 22423
rect 20729 22389 20763 22423
rect 20763 22389 20772 22423
rect 20720 22380 20772 22389
rect 22192 22380 22244 22432
rect 24216 22423 24268 22432
rect 24216 22389 24225 22423
rect 24225 22389 24259 22423
rect 24259 22389 24268 22423
rect 24216 22380 24268 22389
rect 25320 22423 25372 22432
rect 25320 22389 25329 22423
rect 25329 22389 25363 22423
rect 25363 22389 25372 22423
rect 25320 22380 25372 22389
rect 28080 22380 28132 22432
rect 29368 22584 29420 22636
rect 32128 22627 32180 22636
rect 32128 22593 32137 22627
rect 32137 22593 32171 22627
rect 32171 22593 32180 22627
rect 32128 22584 32180 22593
rect 48136 22627 48188 22636
rect 48136 22593 48145 22627
rect 48145 22593 48179 22627
rect 48179 22593 48188 22627
rect 48136 22584 48188 22593
rect 33232 22448 33284 22500
rect 33508 22491 33560 22500
rect 33508 22457 33517 22491
rect 33517 22457 33551 22491
rect 33551 22457 33560 22491
rect 33508 22448 33560 22457
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 12992 22219 13044 22228
rect 2136 22108 2188 22160
rect 9036 22108 9088 22160
rect 11520 22108 11572 22160
rect 12992 22185 13001 22219
rect 13001 22185 13035 22219
rect 13035 22185 13044 22219
rect 12992 22176 13044 22185
rect 15936 22219 15988 22228
rect 15936 22185 15945 22219
rect 15945 22185 15979 22219
rect 15979 22185 15988 22219
rect 15936 22176 15988 22185
rect 16212 22176 16264 22228
rect 18236 22176 18288 22228
rect 19800 22176 19852 22228
rect 21916 22176 21968 22228
rect 23020 22176 23072 22228
rect 27712 22176 27764 22228
rect 30380 22219 30432 22228
rect 30380 22185 30389 22219
rect 30389 22185 30423 22219
rect 30423 22185 30432 22219
rect 30380 22176 30432 22185
rect 8208 22040 8260 22092
rect 8852 22040 8904 22092
rect 18696 22108 18748 22160
rect 19892 22108 19944 22160
rect 21180 22108 21232 22160
rect 19432 22040 19484 22092
rect 25320 22108 25372 22160
rect 30656 22108 30708 22160
rect 9220 22015 9272 22024
rect 9220 21981 9229 22015
rect 9229 21981 9263 22015
rect 9263 21981 9272 22015
rect 9220 21972 9272 21981
rect 6736 21904 6788 21956
rect 4068 21836 4120 21888
rect 9312 21836 9364 21888
rect 9404 21836 9456 21888
rect 9772 21972 9824 22024
rect 17592 21972 17644 22024
rect 10140 21836 10192 21888
rect 11612 21904 11664 21956
rect 13452 21904 13504 21956
rect 12808 21836 12860 21888
rect 16948 21904 17000 21956
rect 18052 21904 18104 21956
rect 18880 21904 18932 21956
rect 17500 21836 17552 21888
rect 19156 21836 19208 21888
rect 19892 22015 19944 22024
rect 19892 21981 19901 22015
rect 19901 21981 19935 22015
rect 19935 21981 19944 22015
rect 19892 21972 19944 21981
rect 20904 21972 20956 22024
rect 23296 22040 23348 22092
rect 20352 21904 20404 21956
rect 22192 21904 22244 21956
rect 22744 21904 22796 21956
rect 24124 21904 24176 21956
rect 25136 21972 25188 22024
rect 30745 22015 30797 22024
rect 30745 21981 30772 22015
rect 30772 21981 30797 22015
rect 30745 21972 30797 21981
rect 31484 22108 31536 22160
rect 31576 22108 31628 22160
rect 48044 22108 48096 22160
rect 30380 21904 30432 21956
rect 32036 22040 32088 22092
rect 32128 22015 32180 22024
rect 32128 21981 32137 22015
rect 32137 21981 32171 22015
rect 32171 21981 32180 22015
rect 32128 21972 32180 21981
rect 32588 22015 32640 22024
rect 32588 21981 32597 22015
rect 32597 21981 32631 22015
rect 32631 21981 32640 22015
rect 32588 21972 32640 21981
rect 33508 21972 33560 22024
rect 21548 21836 21600 21888
rect 23388 21836 23440 21888
rect 24676 21836 24728 21888
rect 24860 21836 24912 21888
rect 25964 21836 26016 21888
rect 28264 21836 28316 21888
rect 31484 21879 31536 21888
rect 31484 21845 31493 21879
rect 31493 21845 31527 21879
rect 31527 21845 31536 21879
rect 31484 21836 31536 21845
rect 33324 21904 33376 21956
rect 45468 21972 45520 22024
rect 47952 21947 48004 21956
rect 34796 21836 34848 21888
rect 47952 21913 47961 21947
rect 47961 21913 47995 21947
rect 47995 21913 48004 21947
rect 47952 21904 48004 21913
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 6736 21675 6788 21684
rect 6736 21641 6745 21675
rect 6745 21641 6779 21675
rect 6779 21641 6788 21675
rect 6736 21632 6788 21641
rect 8484 21632 8536 21684
rect 11612 21675 11664 21684
rect 9312 21564 9364 21616
rect 10140 21564 10192 21616
rect 6644 21539 6696 21548
rect 6644 21505 6653 21539
rect 6653 21505 6687 21539
rect 6687 21505 6696 21539
rect 6644 21496 6696 21505
rect 9404 21496 9456 21548
rect 9864 21539 9916 21548
rect 9864 21505 9873 21539
rect 9873 21505 9907 21539
rect 9907 21505 9916 21539
rect 11612 21641 11621 21675
rect 11621 21641 11655 21675
rect 11655 21641 11664 21675
rect 11612 21632 11664 21641
rect 11980 21632 12032 21684
rect 20352 21632 20404 21684
rect 13452 21564 13504 21616
rect 14740 21564 14792 21616
rect 18052 21564 18104 21616
rect 19064 21564 19116 21616
rect 19248 21564 19300 21616
rect 9864 21496 9916 21505
rect 11152 21428 11204 21480
rect 12348 21496 12400 21548
rect 13544 21496 13596 21548
rect 18420 21496 18472 21548
rect 13820 21471 13872 21480
rect 13820 21437 13829 21471
rect 13829 21437 13863 21471
rect 13863 21437 13872 21471
rect 13820 21428 13872 21437
rect 18880 21496 18932 21548
rect 25596 21632 25648 21684
rect 33324 21632 33376 21684
rect 22744 21607 22796 21616
rect 22744 21573 22753 21607
rect 22753 21573 22787 21607
rect 22787 21573 22796 21607
rect 22744 21564 22796 21573
rect 23112 21564 23164 21616
rect 22376 21496 22428 21548
rect 3976 21360 4028 21412
rect 18972 21428 19024 21480
rect 24860 21496 24912 21548
rect 27620 21564 27672 21616
rect 31484 21564 31536 21616
rect 25228 21539 25280 21548
rect 25228 21505 25262 21539
rect 25262 21505 25280 21539
rect 25228 21496 25280 21505
rect 25596 21496 25648 21548
rect 24216 21471 24268 21480
rect 24216 21437 24225 21471
rect 24225 21437 24259 21471
rect 24259 21437 24268 21471
rect 24216 21428 24268 21437
rect 30748 21428 30800 21480
rect 31392 21539 31444 21548
rect 31392 21505 31401 21539
rect 31401 21505 31435 21539
rect 31435 21505 31444 21539
rect 31392 21496 31444 21505
rect 31576 21539 31628 21548
rect 31576 21505 31585 21539
rect 31585 21505 31619 21539
rect 31619 21505 31628 21539
rect 31576 21496 31628 21505
rect 32128 21496 32180 21548
rect 31484 21428 31536 21480
rect 34520 21471 34572 21480
rect 34520 21437 34529 21471
rect 34529 21437 34563 21471
rect 34563 21437 34572 21471
rect 34520 21428 34572 21437
rect 34704 21471 34756 21480
rect 34704 21437 34713 21471
rect 34713 21437 34747 21471
rect 34747 21437 34756 21471
rect 34704 21428 34756 21437
rect 46572 21428 46624 21480
rect 9220 21335 9272 21344
rect 9220 21301 9229 21335
rect 9229 21301 9263 21335
rect 9263 21301 9272 21335
rect 9220 21292 9272 21301
rect 12808 21292 12860 21344
rect 18144 21335 18196 21344
rect 18144 21301 18153 21335
rect 18153 21301 18187 21335
rect 18187 21301 18196 21335
rect 18144 21292 18196 21301
rect 20720 21360 20772 21412
rect 21824 21360 21876 21412
rect 23112 21360 23164 21412
rect 24952 21360 25004 21412
rect 22100 21292 22152 21344
rect 22284 21335 22336 21344
rect 22284 21301 22293 21335
rect 22293 21301 22327 21335
rect 22327 21301 22336 21335
rect 22284 21292 22336 21301
rect 23296 21292 23348 21344
rect 24676 21292 24728 21344
rect 24860 21292 24912 21344
rect 32772 21292 32824 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 11152 21131 11204 21140
rect 11152 21097 11161 21131
rect 11161 21097 11195 21131
rect 11195 21097 11204 21131
rect 11152 21088 11204 21097
rect 15568 21088 15620 21140
rect 18972 21088 19024 21140
rect 21548 21088 21600 21140
rect 18420 21063 18472 21072
rect 18420 21029 18429 21063
rect 18429 21029 18463 21063
rect 18463 21029 18472 21063
rect 22376 21088 22428 21140
rect 18420 21020 18472 21029
rect 17040 20995 17092 21004
rect 17040 20961 17049 20995
rect 17049 20961 17083 20995
rect 17083 20961 17092 20995
rect 17040 20952 17092 20961
rect 21548 20952 21600 21004
rect 23296 21088 23348 21140
rect 25228 21088 25280 21140
rect 25688 21088 25740 21140
rect 5632 20884 5684 20936
rect 6644 20927 6696 20936
rect 6644 20893 6653 20927
rect 6653 20893 6687 20927
rect 6687 20893 6696 20927
rect 6644 20884 6696 20893
rect 8024 20927 8076 20936
rect 8024 20893 8033 20927
rect 8033 20893 8067 20927
rect 8067 20893 8076 20927
rect 8024 20884 8076 20893
rect 8944 20927 8996 20936
rect 8944 20893 8953 20927
rect 8953 20893 8987 20927
rect 8987 20893 8996 20927
rect 8944 20884 8996 20893
rect 9220 20927 9272 20936
rect 9220 20893 9254 20927
rect 9254 20893 9272 20927
rect 9220 20884 9272 20893
rect 10784 20927 10836 20936
rect 10784 20893 10793 20927
rect 10793 20893 10827 20927
rect 10827 20893 10836 20927
rect 10784 20884 10836 20893
rect 12992 20884 13044 20936
rect 15936 20884 15988 20936
rect 20996 20927 21048 20936
rect 20996 20893 21005 20927
rect 21005 20893 21039 20927
rect 21039 20893 21048 20927
rect 20996 20884 21048 20893
rect 21088 20927 21140 20936
rect 21088 20893 21097 20927
rect 21097 20893 21131 20927
rect 21131 20893 21140 20927
rect 22192 20995 22244 21004
rect 22192 20961 22201 20995
rect 22201 20961 22235 20995
rect 22235 20961 22244 20995
rect 22192 20952 22244 20961
rect 21088 20884 21140 20893
rect 8208 20859 8260 20868
rect 8208 20825 8217 20859
rect 8217 20825 8251 20859
rect 8251 20825 8260 20859
rect 8208 20816 8260 20825
rect 9128 20816 9180 20868
rect 6644 20748 6696 20800
rect 9404 20748 9456 20800
rect 10324 20791 10376 20800
rect 10324 20757 10333 20791
rect 10333 20757 10367 20791
rect 10367 20757 10376 20791
rect 13912 20816 13964 20868
rect 16856 20816 16908 20868
rect 22376 20884 22428 20936
rect 25136 21020 25188 21072
rect 23480 20952 23532 21004
rect 24400 20952 24452 21004
rect 24952 20995 25004 21004
rect 24952 20961 24961 20995
rect 24961 20961 24995 20995
rect 24995 20961 25004 20995
rect 24952 20952 25004 20961
rect 25320 20952 25372 21004
rect 23112 20884 23164 20936
rect 24676 20927 24728 20936
rect 24676 20893 24685 20927
rect 24685 20893 24719 20927
rect 24719 20893 24728 20927
rect 24676 20884 24728 20893
rect 25136 20884 25188 20936
rect 25596 20884 25648 20936
rect 24952 20816 25004 20868
rect 26148 20995 26200 21004
rect 26148 20961 26157 20995
rect 26157 20961 26191 20995
rect 26191 20961 26200 20995
rect 26148 20952 26200 20961
rect 25872 20927 25924 20936
rect 25872 20893 25881 20927
rect 25881 20893 25915 20927
rect 25915 20893 25924 20927
rect 25872 20884 25924 20893
rect 25964 20927 26016 20936
rect 25964 20893 25973 20927
rect 25973 20893 26007 20927
rect 26007 20893 26016 20927
rect 31392 21088 31444 21140
rect 34796 21131 34848 21140
rect 34796 21097 34805 21131
rect 34805 21097 34839 21131
rect 34839 21097 34848 21131
rect 34796 21088 34848 21097
rect 30748 20995 30800 21004
rect 30748 20961 30757 20995
rect 30757 20961 30791 20995
rect 30791 20961 30800 20995
rect 30748 20952 30800 20961
rect 25964 20884 26016 20893
rect 27620 20927 27672 20936
rect 27620 20893 27629 20927
rect 27629 20893 27663 20927
rect 27663 20893 27672 20927
rect 27620 20884 27672 20893
rect 28632 20884 28684 20936
rect 31484 20884 31536 20936
rect 32128 20884 32180 20936
rect 32772 20884 32824 20936
rect 34244 20884 34296 20936
rect 27712 20816 27764 20868
rect 15568 20791 15620 20800
rect 10324 20748 10376 20757
rect 15568 20757 15577 20791
rect 15577 20757 15611 20791
rect 15611 20757 15620 20791
rect 15568 20748 15620 20757
rect 21548 20748 21600 20800
rect 23480 20748 23532 20800
rect 23664 20791 23716 20800
rect 23664 20757 23673 20791
rect 23673 20757 23707 20791
rect 23707 20757 23716 20791
rect 23664 20748 23716 20757
rect 23756 20748 23808 20800
rect 26424 20748 26476 20800
rect 29000 20791 29052 20800
rect 29000 20757 29009 20791
rect 29009 20757 29043 20791
rect 29043 20757 29052 20791
rect 29000 20748 29052 20757
rect 32220 20748 32272 20800
rect 32588 20748 32640 20800
rect 34520 20816 34572 20868
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 5632 20451 5684 20460
rect 5632 20417 5641 20451
rect 5641 20417 5675 20451
rect 5675 20417 5684 20451
rect 5632 20408 5684 20417
rect 10324 20544 10376 20596
rect 13912 20587 13964 20596
rect 13912 20553 13921 20587
rect 13921 20553 13955 20587
rect 13955 20553 13964 20587
rect 13912 20544 13964 20553
rect 9128 20476 9180 20528
rect 10784 20476 10836 20528
rect 14832 20544 14884 20596
rect 16856 20587 16908 20596
rect 16856 20553 16865 20587
rect 16865 20553 16899 20587
rect 16899 20553 16908 20587
rect 16856 20544 16908 20553
rect 8944 20451 8996 20460
rect 8944 20417 8978 20451
rect 8978 20417 8996 20451
rect 10692 20451 10744 20460
rect 8944 20408 8996 20417
rect 10692 20417 10701 20451
rect 10701 20417 10735 20451
rect 10735 20417 10744 20451
rect 10692 20408 10744 20417
rect 14188 20451 14240 20460
rect 14188 20417 14211 20451
rect 14211 20417 14240 20451
rect 14188 20408 14240 20417
rect 8024 20383 8076 20392
rect 8024 20349 8033 20383
rect 8033 20349 8067 20383
rect 8067 20349 8076 20383
rect 8024 20340 8076 20349
rect 14556 20451 14608 20460
rect 14556 20417 14565 20451
rect 14565 20417 14599 20451
rect 14599 20417 14608 20451
rect 14556 20408 14608 20417
rect 16580 20408 16632 20460
rect 17132 20451 17184 20460
rect 17132 20417 17141 20451
rect 17141 20417 17175 20451
rect 17175 20417 17184 20451
rect 17132 20408 17184 20417
rect 18144 20476 18196 20528
rect 18236 20451 18288 20460
rect 18236 20417 18245 20451
rect 18245 20417 18279 20451
rect 18279 20417 18288 20451
rect 18236 20408 18288 20417
rect 19156 20544 19208 20596
rect 20076 20544 20128 20596
rect 23296 20544 23348 20596
rect 24124 20544 24176 20596
rect 24492 20544 24544 20596
rect 25872 20544 25924 20596
rect 32864 20544 32916 20596
rect 34704 20544 34756 20596
rect 18696 20408 18748 20460
rect 19064 20451 19116 20460
rect 19064 20417 19073 20451
rect 19073 20417 19107 20451
rect 19107 20417 19116 20451
rect 19064 20408 19116 20417
rect 19248 20451 19300 20460
rect 19248 20417 19257 20451
rect 19257 20417 19291 20451
rect 19291 20417 19300 20451
rect 19248 20408 19300 20417
rect 19156 20340 19208 20392
rect 22284 20476 22336 20528
rect 20076 20408 20128 20460
rect 20536 20408 20588 20460
rect 20996 20408 21048 20460
rect 21548 20408 21600 20460
rect 24216 20476 24268 20528
rect 23664 20408 23716 20460
rect 25964 20451 26016 20460
rect 25964 20417 25973 20451
rect 25973 20417 26007 20451
rect 26007 20417 26016 20451
rect 25964 20408 26016 20417
rect 21272 20340 21324 20392
rect 21640 20340 21692 20392
rect 29000 20476 29052 20528
rect 27804 20451 27856 20460
rect 27804 20417 27813 20451
rect 27813 20417 27847 20451
rect 27847 20417 27856 20451
rect 27804 20408 27856 20417
rect 27988 20383 28040 20392
rect 27988 20349 27997 20383
rect 27997 20349 28031 20383
rect 28031 20349 28040 20383
rect 27988 20340 28040 20349
rect 29184 20408 29236 20460
rect 30472 20408 30524 20460
rect 30380 20340 30432 20392
rect 32220 20408 32272 20460
rect 32588 20408 32640 20460
rect 34244 20408 34296 20460
rect 14280 20272 14332 20324
rect 27804 20272 27856 20324
rect 28724 20272 28776 20324
rect 31760 20272 31812 20324
rect 8208 20204 8260 20256
rect 10140 20204 10192 20256
rect 12532 20204 12584 20256
rect 17592 20204 17644 20256
rect 20352 20247 20404 20256
rect 20352 20213 20361 20247
rect 20361 20213 20395 20247
rect 20395 20213 20404 20247
rect 20996 20247 21048 20256
rect 20352 20204 20404 20213
rect 20996 20213 21005 20247
rect 21005 20213 21039 20247
rect 21039 20213 21048 20247
rect 20996 20204 21048 20213
rect 22284 20204 22336 20256
rect 24492 20247 24544 20256
rect 24492 20213 24501 20247
rect 24501 20213 24535 20247
rect 24535 20213 24544 20247
rect 24492 20204 24544 20213
rect 24768 20204 24820 20256
rect 25320 20204 25372 20256
rect 25688 20204 25740 20256
rect 26700 20204 26752 20256
rect 27528 20204 27580 20256
rect 29092 20204 29144 20256
rect 33140 20204 33192 20256
rect 46296 20204 46348 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 8944 20043 8996 20052
rect 8944 20009 8953 20043
rect 8953 20009 8987 20043
rect 8987 20009 8996 20043
rect 8944 20000 8996 20009
rect 8208 19932 8260 19984
rect 18604 20000 18656 20052
rect 19248 20000 19300 20052
rect 21456 20000 21508 20052
rect 27712 20043 27764 20052
rect 27712 20009 27721 20043
rect 27721 20009 27755 20043
rect 27755 20009 27764 20043
rect 27712 20000 27764 20009
rect 6644 19907 6696 19916
rect 6644 19873 6653 19907
rect 6653 19873 6687 19907
rect 6687 19873 6696 19907
rect 6644 19864 6696 19873
rect 6920 19907 6972 19916
rect 6920 19873 6929 19907
rect 6929 19873 6963 19907
rect 6963 19873 6972 19907
rect 6920 19864 6972 19873
rect 20536 19932 20588 19984
rect 21180 19932 21232 19984
rect 22192 19932 22244 19984
rect 30748 19932 30800 19984
rect 21640 19907 21692 19916
rect 3976 19728 4028 19780
rect 9036 19796 9088 19848
rect 9312 19839 9364 19848
rect 9312 19805 9321 19839
rect 9321 19805 9355 19839
rect 9355 19805 9364 19839
rect 9312 19796 9364 19805
rect 9404 19836 9456 19848
rect 9404 19802 9413 19836
rect 9413 19802 9447 19836
rect 9447 19802 9456 19836
rect 9404 19796 9456 19802
rect 9772 19796 9824 19848
rect 10232 19796 10284 19848
rect 21640 19873 21649 19907
rect 21649 19873 21683 19907
rect 21683 19873 21692 19907
rect 21640 19864 21692 19873
rect 22284 19864 22336 19916
rect 23756 19864 23808 19916
rect 24584 19864 24636 19916
rect 27436 19864 27488 19916
rect 13636 19796 13688 19848
rect 13820 19796 13872 19848
rect 17316 19839 17368 19848
rect 17316 19805 17325 19839
rect 17325 19805 17359 19839
rect 17359 19805 17368 19839
rect 17316 19796 17368 19805
rect 17592 19839 17644 19848
rect 17592 19805 17626 19839
rect 17626 19805 17644 19839
rect 17592 19796 17644 19805
rect 17868 19796 17920 19848
rect 20352 19796 20404 19848
rect 23020 19796 23072 19848
rect 23480 19796 23532 19848
rect 26424 19839 26476 19848
rect 26424 19805 26433 19839
rect 26433 19805 26467 19839
rect 26467 19805 26476 19839
rect 26424 19796 26476 19805
rect 26700 19839 26752 19848
rect 26700 19805 26709 19839
rect 26709 19805 26743 19839
rect 26743 19805 26752 19839
rect 26700 19796 26752 19805
rect 27620 19796 27672 19848
rect 28724 19796 28776 19848
rect 30380 19796 30432 19848
rect 32312 19864 32364 19916
rect 46296 19907 46348 19916
rect 46296 19873 46305 19907
rect 46305 19873 46339 19907
rect 46339 19873 46348 19907
rect 46296 19864 46348 19873
rect 14372 19728 14424 19780
rect 20904 19728 20956 19780
rect 15108 19660 15160 19712
rect 20628 19703 20680 19712
rect 20628 19669 20637 19703
rect 20637 19669 20671 19703
rect 20671 19669 20680 19703
rect 21456 19703 21508 19712
rect 20628 19660 20680 19669
rect 21456 19669 21465 19703
rect 21465 19669 21499 19703
rect 21499 19669 21508 19703
rect 25872 19728 25924 19780
rect 29000 19728 29052 19780
rect 22284 19703 22336 19712
rect 21456 19660 21508 19669
rect 22284 19669 22293 19703
rect 22293 19669 22327 19703
rect 22327 19669 22336 19703
rect 22284 19660 22336 19669
rect 27528 19660 27580 19712
rect 31484 19728 31536 19780
rect 31576 19703 31628 19712
rect 31576 19669 31585 19703
rect 31585 19669 31619 19703
rect 31619 19669 31628 19703
rect 31576 19660 31628 19669
rect 32680 19703 32732 19712
rect 32680 19669 32689 19703
rect 32689 19669 32723 19703
rect 32723 19669 32732 19703
rect 32680 19660 32732 19669
rect 32864 19728 32916 19780
rect 33140 19839 33192 19848
rect 33140 19805 33149 19839
rect 33149 19805 33183 19839
rect 33183 19805 33192 19839
rect 33140 19796 33192 19805
rect 48136 19839 48188 19848
rect 48136 19805 48145 19839
rect 48145 19805 48179 19839
rect 48179 19805 48188 19839
rect 48136 19796 48188 19805
rect 46940 19728 46992 19780
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 2320 19456 2372 19508
rect 3976 19456 4028 19508
rect 4068 19456 4120 19508
rect 15936 19499 15988 19508
rect 12532 19431 12584 19440
rect 12532 19397 12541 19431
rect 12541 19397 12575 19431
rect 12575 19397 12584 19431
rect 12532 19388 12584 19397
rect 15936 19465 15945 19499
rect 15945 19465 15979 19499
rect 15979 19465 15988 19499
rect 15936 19456 15988 19465
rect 17040 19456 17092 19508
rect 17868 19456 17920 19508
rect 22284 19456 22336 19508
rect 24676 19456 24728 19508
rect 25596 19456 25648 19508
rect 16764 19388 16816 19440
rect 9404 19363 9456 19372
rect 9404 19329 9438 19363
rect 9438 19329 9456 19363
rect 9404 19320 9456 19329
rect 9864 19320 9916 19372
rect 9128 19295 9180 19304
rect 9128 19261 9137 19295
rect 9137 19261 9171 19295
rect 9171 19261 9180 19295
rect 9128 19252 9180 19261
rect 10692 19320 10744 19372
rect 13728 19320 13780 19372
rect 12624 19252 12676 19304
rect 14464 19252 14516 19304
rect 15108 19363 15160 19372
rect 15108 19329 15117 19363
rect 15117 19329 15151 19363
rect 15151 19329 15160 19363
rect 15108 19320 15160 19329
rect 15292 19363 15344 19372
rect 15292 19329 15301 19363
rect 15301 19329 15335 19363
rect 15335 19329 15344 19363
rect 16672 19363 16724 19372
rect 15292 19320 15344 19329
rect 1400 19116 1452 19168
rect 2228 19159 2280 19168
rect 2228 19125 2237 19159
rect 2237 19125 2271 19159
rect 2271 19125 2280 19159
rect 2228 19116 2280 19125
rect 9772 19116 9824 19168
rect 15568 19184 15620 19236
rect 16672 19329 16681 19363
rect 16681 19329 16715 19363
rect 16715 19329 16724 19363
rect 16672 19320 16724 19329
rect 20628 19363 20680 19372
rect 20628 19329 20637 19363
rect 20637 19329 20671 19363
rect 20671 19329 20680 19363
rect 20628 19320 20680 19329
rect 16580 19252 16632 19304
rect 20904 19295 20956 19304
rect 20904 19261 20913 19295
rect 20913 19261 20947 19295
rect 20947 19261 20956 19295
rect 20904 19252 20956 19261
rect 21088 19184 21140 19236
rect 22744 19320 22796 19372
rect 23296 19320 23348 19372
rect 23480 19388 23532 19440
rect 24216 19388 24268 19440
rect 24768 19388 24820 19440
rect 26700 19388 26752 19440
rect 28356 19456 28408 19508
rect 29184 19388 29236 19440
rect 31760 19456 31812 19508
rect 32312 19456 32364 19508
rect 32588 19456 32640 19508
rect 46940 19499 46992 19508
rect 46940 19465 46949 19499
rect 46949 19465 46983 19499
rect 46983 19465 46992 19499
rect 46940 19456 46992 19465
rect 32680 19388 32732 19440
rect 24860 19363 24912 19372
rect 24860 19329 24869 19363
rect 24869 19329 24903 19363
rect 24903 19329 24912 19363
rect 24860 19320 24912 19329
rect 27344 19320 27396 19372
rect 28264 19320 28316 19372
rect 28632 19363 28684 19372
rect 28632 19329 28641 19363
rect 28641 19329 28675 19363
rect 28675 19329 28684 19363
rect 28632 19320 28684 19329
rect 28908 19363 28960 19372
rect 28908 19329 28942 19363
rect 28942 19329 28960 19363
rect 28908 19320 28960 19329
rect 31760 19320 31812 19372
rect 32128 19363 32180 19372
rect 32128 19329 32137 19363
rect 32137 19329 32171 19363
rect 32171 19329 32180 19363
rect 32128 19320 32180 19329
rect 46756 19320 46808 19372
rect 47952 19363 48004 19372
rect 47952 19329 47961 19363
rect 47961 19329 47995 19363
rect 47995 19329 48004 19363
rect 47952 19320 48004 19329
rect 14648 19159 14700 19168
rect 14648 19125 14657 19159
rect 14657 19125 14691 19159
rect 14691 19125 14700 19159
rect 14648 19116 14700 19125
rect 20076 19116 20128 19168
rect 21916 19252 21968 19304
rect 23388 19295 23440 19304
rect 23388 19261 23397 19295
rect 23397 19261 23431 19295
rect 23431 19261 23440 19295
rect 23388 19252 23440 19261
rect 26424 19252 26476 19304
rect 27988 19295 28040 19304
rect 27988 19261 27997 19295
rect 27997 19261 28031 19295
rect 28031 19261 28040 19295
rect 27988 19252 28040 19261
rect 23020 19184 23072 19236
rect 24860 19184 24912 19236
rect 21824 19116 21876 19168
rect 22376 19159 22428 19168
rect 22376 19125 22385 19159
rect 22385 19125 22419 19159
rect 22419 19125 22428 19159
rect 22376 19116 22428 19125
rect 25964 19116 26016 19168
rect 27344 19116 27396 19168
rect 48044 19159 48096 19168
rect 48044 19125 48053 19159
rect 48053 19125 48087 19159
rect 48087 19125 48096 19159
rect 48044 19116 48096 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 9404 18912 9456 18964
rect 12624 18955 12676 18964
rect 12624 18921 12633 18955
rect 12633 18921 12667 18955
rect 12667 18921 12676 18955
rect 12624 18912 12676 18921
rect 20996 18912 21048 18964
rect 14372 18844 14424 18896
rect 20812 18844 20864 18896
rect 21456 18844 21508 18896
rect 25596 18912 25648 18964
rect 25872 18912 25924 18964
rect 26700 18912 26752 18964
rect 26792 18912 26844 18964
rect 27528 18955 27580 18964
rect 27528 18921 27537 18955
rect 27537 18921 27571 18955
rect 27571 18921 27580 18955
rect 27528 18912 27580 18921
rect 28264 18912 28316 18964
rect 21640 18844 21692 18896
rect 21824 18844 21876 18896
rect 1400 18819 1452 18828
rect 1400 18785 1409 18819
rect 1409 18785 1443 18819
rect 1443 18785 1452 18819
rect 1400 18776 1452 18785
rect 2228 18776 2280 18828
rect 2780 18819 2832 18828
rect 2780 18785 2789 18819
rect 2789 18785 2823 18819
rect 2823 18785 2832 18819
rect 2780 18776 2832 18785
rect 9312 18776 9364 18828
rect 9772 18708 9824 18760
rect 10140 18708 10192 18760
rect 10232 18751 10284 18760
rect 10232 18717 10241 18751
rect 10241 18717 10275 18751
rect 10275 18717 10284 18751
rect 11244 18751 11296 18760
rect 10232 18708 10284 18717
rect 11244 18717 11253 18751
rect 11253 18717 11287 18751
rect 11287 18717 11296 18751
rect 12992 18776 13044 18828
rect 11244 18708 11296 18717
rect 12624 18708 12676 18760
rect 16672 18776 16724 18828
rect 20536 18819 20588 18828
rect 13544 18708 13596 18760
rect 14464 18751 14516 18760
rect 14464 18717 14473 18751
rect 14473 18717 14507 18751
rect 14507 18717 14516 18751
rect 14464 18708 14516 18717
rect 15292 18708 15344 18760
rect 17316 18708 17368 18760
rect 20536 18785 20545 18819
rect 20545 18785 20579 18819
rect 20579 18785 20588 18819
rect 20536 18776 20588 18785
rect 16672 18640 16724 18692
rect 17224 18640 17276 18692
rect 20076 18708 20128 18760
rect 21548 18776 21600 18828
rect 23112 18844 23164 18896
rect 26424 18887 26476 18896
rect 26424 18853 26433 18887
rect 26433 18853 26467 18887
rect 26467 18853 26476 18887
rect 26424 18844 26476 18853
rect 21640 18708 21692 18760
rect 23388 18751 23440 18760
rect 23388 18717 23397 18751
rect 23397 18717 23431 18751
rect 23431 18717 23440 18751
rect 23388 18708 23440 18717
rect 23480 18751 23532 18760
rect 23480 18717 23489 18751
rect 23489 18717 23523 18751
rect 23523 18717 23532 18751
rect 26792 18776 26844 18828
rect 23480 18708 23532 18717
rect 25964 18751 26016 18760
rect 17776 18572 17828 18624
rect 21548 18572 21600 18624
rect 22100 18572 22152 18624
rect 25320 18640 25372 18692
rect 25964 18717 25973 18751
rect 25973 18717 26007 18751
rect 26007 18717 26016 18751
rect 25964 18708 26016 18717
rect 26884 18708 26936 18760
rect 27068 18708 27120 18760
rect 26148 18640 26200 18692
rect 24676 18572 24728 18624
rect 25688 18572 25740 18624
rect 28356 18819 28408 18828
rect 28356 18785 28365 18819
rect 28365 18785 28399 18819
rect 28399 18785 28408 18819
rect 28356 18776 28408 18785
rect 27344 18751 27396 18760
rect 27344 18717 27353 18751
rect 27353 18717 27387 18751
rect 27387 18717 27396 18751
rect 27344 18708 27396 18717
rect 27804 18708 27856 18760
rect 28264 18751 28316 18760
rect 28264 18717 28273 18751
rect 28273 18717 28307 18751
rect 28307 18717 28316 18751
rect 28264 18708 28316 18717
rect 28908 18912 28960 18964
rect 28724 18708 28776 18760
rect 31576 18708 31628 18760
rect 31760 18572 31812 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 13820 18368 13872 18420
rect 16672 18411 16724 18420
rect 16672 18377 16681 18411
rect 16681 18377 16715 18411
rect 16715 18377 16724 18411
rect 16672 18368 16724 18377
rect 17776 18411 17828 18420
rect 17776 18377 17785 18411
rect 17785 18377 17819 18411
rect 17819 18377 17828 18411
rect 17776 18368 17828 18377
rect 21640 18368 21692 18420
rect 21824 18368 21876 18420
rect 12992 18300 13044 18352
rect 14372 18300 14424 18352
rect 16028 18300 16080 18352
rect 16580 18300 16632 18352
rect 20352 18300 20404 18352
rect 20996 18343 21048 18352
rect 20996 18309 21005 18343
rect 21005 18309 21039 18343
rect 21039 18309 21048 18343
rect 20996 18300 21048 18309
rect 21916 18300 21968 18352
rect 14648 18232 14700 18284
rect 14924 18275 14976 18284
rect 14924 18241 14947 18275
rect 14947 18241 14976 18275
rect 14924 18232 14976 18241
rect 15292 18275 15344 18284
rect 1952 18207 2004 18216
rect 1952 18173 1961 18207
rect 1961 18173 1995 18207
rect 1995 18173 2004 18207
rect 1952 18164 2004 18173
rect 2780 18207 2832 18216
rect 2780 18173 2789 18207
rect 2789 18173 2823 18207
rect 2823 18173 2832 18207
rect 2780 18164 2832 18173
rect 14464 18164 14516 18216
rect 15292 18241 15301 18275
rect 15301 18241 15335 18275
rect 15335 18241 15344 18275
rect 15292 18232 15344 18241
rect 15844 18232 15896 18284
rect 17224 18232 17276 18284
rect 18512 18232 18564 18284
rect 18604 18275 18656 18284
rect 18604 18241 18613 18275
rect 18613 18241 18647 18275
rect 18647 18241 18656 18275
rect 18604 18232 18656 18241
rect 17408 18164 17460 18216
rect 20720 18232 20772 18284
rect 20904 18275 20956 18284
rect 20904 18241 20913 18275
rect 20913 18241 20947 18275
rect 20947 18241 20956 18275
rect 20904 18232 20956 18241
rect 21824 18232 21876 18284
rect 22100 18275 22152 18284
rect 22100 18241 22109 18275
rect 22109 18241 22143 18275
rect 22143 18241 22152 18275
rect 23664 18368 23716 18420
rect 24216 18368 24268 18420
rect 25136 18368 25188 18420
rect 27804 18411 27856 18420
rect 23020 18300 23072 18352
rect 24032 18300 24084 18352
rect 26148 18300 26200 18352
rect 22100 18232 22152 18241
rect 24124 18275 24176 18284
rect 24124 18241 24133 18275
rect 24133 18241 24167 18275
rect 24167 18241 24176 18275
rect 24124 18232 24176 18241
rect 25320 18232 25372 18284
rect 27528 18300 27580 18352
rect 27804 18377 27813 18411
rect 27813 18377 27847 18411
rect 27847 18377 27856 18411
rect 27804 18368 27856 18377
rect 28264 18300 28316 18352
rect 28356 18300 28408 18352
rect 28540 18232 28592 18284
rect 34336 18232 34388 18284
rect 21548 18164 21600 18216
rect 4068 18096 4120 18148
rect 8300 18096 8352 18148
rect 17224 18096 17276 18148
rect 22284 18207 22336 18216
rect 22284 18173 22293 18207
rect 22293 18173 22327 18207
rect 22327 18173 22336 18207
rect 22284 18164 22336 18173
rect 24216 18164 24268 18216
rect 24676 18164 24728 18216
rect 26148 18164 26200 18216
rect 29000 18164 29052 18216
rect 32864 18207 32916 18216
rect 32864 18173 32873 18207
rect 32873 18173 32907 18207
rect 32907 18173 32916 18207
rect 32864 18164 32916 18173
rect 34428 18164 34480 18216
rect 23296 18096 23348 18148
rect 25596 18096 25648 18148
rect 14924 18028 14976 18080
rect 17500 18028 17552 18080
rect 18696 18071 18748 18080
rect 18696 18037 18705 18071
rect 18705 18037 18739 18071
rect 18739 18037 18748 18071
rect 18696 18028 18748 18037
rect 20720 18028 20772 18080
rect 22192 18028 22244 18080
rect 23112 18028 23164 18080
rect 23388 18028 23440 18080
rect 23572 18028 23624 18080
rect 24032 18028 24084 18080
rect 27620 18071 27672 18080
rect 27620 18037 27629 18071
rect 27629 18037 27663 18071
rect 27663 18037 27672 18071
rect 27620 18028 27672 18037
rect 28724 18071 28776 18080
rect 28724 18037 28733 18071
rect 28733 18037 28767 18071
rect 28767 18037 28776 18071
rect 28724 18028 28776 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 1952 17824 2004 17876
rect 8300 17799 8352 17808
rect 8300 17765 8309 17799
rect 8309 17765 8343 17799
rect 8343 17765 8352 17799
rect 8300 17756 8352 17765
rect 13728 17824 13780 17876
rect 16028 17867 16080 17876
rect 14648 17756 14700 17808
rect 9128 17688 9180 17740
rect 11244 17688 11296 17740
rect 11336 17731 11388 17740
rect 11336 17697 11345 17731
rect 11345 17697 11379 17731
rect 11379 17697 11388 17731
rect 11336 17688 11388 17697
rect 12808 17688 12860 17740
rect 1768 17620 1820 17672
rect 2044 17663 2096 17672
rect 2044 17629 2053 17663
rect 2053 17629 2087 17663
rect 2087 17629 2096 17663
rect 2044 17620 2096 17629
rect 2596 17620 2648 17672
rect 9864 17663 9916 17672
rect 9864 17629 9873 17663
rect 9873 17629 9907 17663
rect 9907 17629 9916 17663
rect 9864 17620 9916 17629
rect 11980 17620 12032 17672
rect 14464 17688 14516 17740
rect 16028 17833 16037 17867
rect 16037 17833 16071 17867
rect 16071 17833 16080 17867
rect 16028 17824 16080 17833
rect 16120 17824 16172 17876
rect 22284 17824 22336 17876
rect 23480 17824 23532 17876
rect 16764 17799 16816 17808
rect 16764 17765 16773 17799
rect 16773 17765 16807 17799
rect 16807 17765 16816 17799
rect 16764 17756 16816 17765
rect 17040 17688 17092 17740
rect 14372 17620 14424 17672
rect 17316 17620 17368 17672
rect 17500 17663 17552 17672
rect 17500 17629 17534 17663
rect 17534 17629 17552 17663
rect 17500 17620 17552 17629
rect 23020 17756 23072 17808
rect 23112 17756 23164 17808
rect 24768 17824 24820 17876
rect 25136 17824 25188 17876
rect 25320 17867 25372 17876
rect 25320 17833 25329 17867
rect 25329 17833 25363 17867
rect 25363 17833 25372 17867
rect 25320 17824 25372 17833
rect 26700 17824 26752 17876
rect 27620 17824 27672 17876
rect 34428 17824 34480 17876
rect 20076 17688 20128 17740
rect 24124 17688 24176 17740
rect 21640 17663 21692 17672
rect 8852 17552 8904 17604
rect 10048 17595 10100 17604
rect 10048 17561 10057 17595
rect 10057 17561 10091 17595
rect 10091 17561 10100 17595
rect 10048 17552 10100 17561
rect 14924 17595 14976 17604
rect 14924 17561 14958 17595
rect 14958 17561 14976 17595
rect 14924 17552 14976 17561
rect 15016 17552 15068 17604
rect 16120 17552 16172 17604
rect 16580 17595 16632 17604
rect 16580 17561 16589 17595
rect 16589 17561 16623 17595
rect 16623 17561 16632 17595
rect 16580 17552 16632 17561
rect 1952 17484 2004 17536
rect 7564 17484 7616 17536
rect 10416 17484 10468 17536
rect 10508 17484 10560 17536
rect 20628 17552 20680 17604
rect 21640 17629 21649 17663
rect 21649 17629 21683 17663
rect 21683 17629 21692 17663
rect 21640 17620 21692 17629
rect 22100 17663 22152 17672
rect 22100 17629 22109 17663
rect 22109 17629 22143 17663
rect 22143 17629 22152 17663
rect 22100 17620 22152 17629
rect 22376 17620 22428 17672
rect 22928 17620 22980 17672
rect 23112 17552 23164 17604
rect 24216 17620 24268 17672
rect 24032 17552 24084 17604
rect 24584 17688 24636 17740
rect 24952 17688 25004 17740
rect 26148 17595 26200 17604
rect 26148 17561 26157 17595
rect 26157 17561 26191 17595
rect 26191 17561 26200 17595
rect 26148 17552 26200 17561
rect 20904 17484 20956 17536
rect 22284 17527 22336 17536
rect 22284 17493 22293 17527
rect 22293 17493 22327 17527
rect 22327 17493 22336 17527
rect 22284 17484 22336 17493
rect 24768 17527 24820 17536
rect 24768 17493 24777 17527
rect 24777 17493 24811 17527
rect 24811 17493 24820 17527
rect 24768 17484 24820 17493
rect 26792 17663 26844 17672
rect 26792 17629 26801 17663
rect 26801 17629 26835 17663
rect 26835 17629 26844 17663
rect 26792 17620 26844 17629
rect 26976 17663 27028 17672
rect 26976 17629 26985 17663
rect 26985 17629 27019 17663
rect 27019 17629 27028 17663
rect 26976 17620 27028 17629
rect 28356 17688 28408 17740
rect 28632 17688 28684 17740
rect 27344 17620 27396 17672
rect 31760 17688 31812 17740
rect 33048 17731 33100 17740
rect 33048 17697 33057 17731
rect 33057 17697 33091 17731
rect 33091 17697 33100 17731
rect 33048 17688 33100 17697
rect 34244 17620 34296 17672
rect 46296 17620 46348 17672
rect 29644 17552 29696 17604
rect 29828 17484 29880 17536
rect 33508 17484 33560 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 1676 17280 1728 17332
rect 7564 17280 7616 17332
rect 8852 17323 8904 17332
rect 8852 17289 8861 17323
rect 8861 17289 8895 17323
rect 8895 17289 8904 17323
rect 8852 17280 8904 17289
rect 10048 17323 10100 17332
rect 10048 17289 10057 17323
rect 10057 17289 10091 17323
rect 10091 17289 10100 17323
rect 10048 17280 10100 17289
rect 1952 17255 2004 17264
rect 1952 17221 1961 17255
rect 1961 17221 1995 17255
rect 1995 17221 2004 17255
rect 1952 17212 2004 17221
rect 1768 17187 1820 17196
rect 1768 17153 1777 17187
rect 1777 17153 1811 17187
rect 1811 17153 1820 17187
rect 1768 17144 1820 17153
rect 9772 17144 9824 17196
rect 9956 17187 10008 17196
rect 9956 17153 9965 17187
rect 9965 17153 9999 17187
rect 9999 17153 10008 17187
rect 9956 17144 10008 17153
rect 10508 17144 10560 17196
rect 2780 17119 2832 17128
rect 2780 17085 2789 17119
rect 2789 17085 2823 17119
rect 2823 17085 2832 17119
rect 2780 17076 2832 17085
rect 11520 17144 11572 17196
rect 12900 17212 12952 17264
rect 11980 17187 12032 17196
rect 11980 17153 11989 17187
rect 11989 17153 12023 17187
rect 12023 17153 12032 17187
rect 11980 17144 12032 17153
rect 12716 17187 12768 17196
rect 12716 17153 12725 17187
rect 12725 17153 12759 17187
rect 12759 17153 12768 17187
rect 12716 17144 12768 17153
rect 15292 17280 15344 17332
rect 15936 17280 15988 17332
rect 18512 17280 18564 17332
rect 20812 17280 20864 17332
rect 20996 17280 21048 17332
rect 21272 17280 21324 17332
rect 21824 17280 21876 17332
rect 22100 17280 22152 17332
rect 14464 17212 14516 17264
rect 15384 17144 15436 17196
rect 16028 17212 16080 17264
rect 22928 17255 22980 17264
rect 22928 17221 22937 17255
rect 22937 17221 22971 17255
rect 22971 17221 22980 17255
rect 22928 17212 22980 17221
rect 23020 17212 23072 17264
rect 13728 17076 13780 17128
rect 15936 17187 15988 17196
rect 15936 17153 15945 17187
rect 15945 17153 15979 17187
rect 15979 17153 15988 17187
rect 15936 17144 15988 17153
rect 18328 17144 18380 17196
rect 20536 17144 20588 17196
rect 22192 17187 22244 17196
rect 22192 17153 22201 17187
rect 22201 17153 22235 17187
rect 22235 17153 22244 17187
rect 22192 17144 22244 17153
rect 23112 17187 23164 17196
rect 17408 17076 17460 17128
rect 20904 17076 20956 17128
rect 21640 17076 21692 17128
rect 23112 17153 23121 17187
rect 23121 17153 23155 17187
rect 23155 17153 23164 17187
rect 23112 17144 23164 17153
rect 23572 17144 23624 17196
rect 25044 17280 25096 17332
rect 25136 17280 25188 17332
rect 26792 17280 26844 17332
rect 24860 17212 24912 17264
rect 29092 17280 29144 17332
rect 28080 17255 28132 17264
rect 28080 17221 28089 17255
rect 28089 17221 28123 17255
rect 28123 17221 28132 17255
rect 28080 17212 28132 17221
rect 29460 17212 29512 17264
rect 33508 17255 33560 17264
rect 33508 17221 33517 17255
rect 33517 17221 33551 17255
rect 33551 17221 33560 17255
rect 33508 17212 33560 17221
rect 23296 17076 23348 17128
rect 25136 17144 25188 17196
rect 27160 17144 27212 17196
rect 27344 17144 27396 17196
rect 30288 17144 30340 17196
rect 47400 17144 47452 17196
rect 24124 17076 24176 17128
rect 24308 17076 24360 17128
rect 11704 16940 11756 16992
rect 11888 17008 11940 17060
rect 15384 17008 15436 17060
rect 15844 17008 15896 17060
rect 20628 17008 20680 17060
rect 22560 17008 22612 17060
rect 14280 16940 14332 16992
rect 15200 16940 15252 16992
rect 15476 16940 15528 16992
rect 18604 16940 18656 16992
rect 18972 16940 19024 16992
rect 20168 16940 20220 16992
rect 20444 16940 20496 16992
rect 20812 16940 20864 16992
rect 23848 17008 23900 17060
rect 24768 17008 24820 17060
rect 23480 16940 23532 16992
rect 23664 16983 23716 16992
rect 23664 16949 23673 16983
rect 23673 16949 23707 16983
rect 23707 16949 23716 16983
rect 23664 16940 23716 16949
rect 27252 17008 27304 17060
rect 33508 17076 33560 17128
rect 33600 17076 33652 17128
rect 29552 16940 29604 16992
rect 30196 16983 30248 16992
rect 30196 16949 30205 16983
rect 30205 16949 30239 16983
rect 30239 16949 30248 16983
rect 30196 16940 30248 16949
rect 47676 16983 47728 16992
rect 47676 16949 47685 16983
rect 47685 16949 47719 16983
rect 47719 16949 47728 16983
rect 47676 16940 47728 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 2688 16668 2740 16720
rect 1860 16575 1912 16584
rect 1860 16541 1869 16575
rect 1869 16541 1903 16575
rect 1903 16541 1912 16575
rect 1860 16532 1912 16541
rect 11244 16600 11296 16652
rect 14372 16643 14424 16652
rect 14372 16609 14381 16643
rect 14381 16609 14415 16643
rect 14415 16609 14424 16643
rect 14372 16600 14424 16609
rect 16580 16736 16632 16788
rect 17684 16736 17736 16788
rect 20076 16736 20128 16788
rect 20536 16779 20588 16788
rect 20536 16745 20545 16779
rect 20545 16745 20579 16779
rect 20579 16745 20588 16779
rect 20536 16736 20588 16745
rect 17408 16711 17460 16720
rect 17408 16677 17417 16711
rect 17417 16677 17451 16711
rect 17451 16677 17460 16711
rect 17408 16668 17460 16677
rect 23020 16600 23072 16652
rect 28356 16736 28408 16788
rect 28908 16736 28960 16788
rect 30288 16779 30340 16788
rect 27160 16643 27212 16652
rect 27160 16609 27169 16643
rect 27169 16609 27203 16643
rect 27203 16609 27212 16643
rect 28540 16643 28592 16652
rect 27160 16600 27212 16609
rect 11704 16575 11756 16584
rect 11704 16541 11738 16575
rect 11738 16541 11756 16575
rect 11704 16532 11756 16541
rect 15200 16532 15252 16584
rect 11888 16464 11940 16516
rect 17868 16464 17920 16516
rect 18972 16464 19024 16516
rect 20720 16575 20772 16584
rect 20720 16541 20729 16575
rect 20729 16541 20763 16575
rect 20763 16541 20772 16575
rect 20720 16532 20772 16541
rect 20812 16464 20864 16516
rect 20996 16575 21048 16584
rect 20996 16541 21005 16575
rect 21005 16541 21039 16575
rect 21039 16541 21048 16575
rect 20996 16532 21048 16541
rect 21456 16532 21508 16584
rect 23664 16532 23716 16584
rect 27436 16532 27488 16584
rect 11704 16396 11756 16448
rect 11796 16396 11848 16448
rect 16672 16396 16724 16448
rect 20996 16396 21048 16448
rect 25136 16396 25188 16448
rect 28540 16609 28549 16643
rect 28549 16609 28583 16643
rect 28583 16609 28592 16643
rect 28540 16600 28592 16609
rect 28632 16643 28684 16652
rect 28632 16609 28641 16643
rect 28641 16609 28675 16643
rect 28675 16609 28684 16643
rect 28632 16600 28684 16609
rect 28080 16532 28132 16584
rect 29460 16532 29512 16584
rect 30288 16745 30297 16779
rect 30297 16745 30331 16779
rect 30331 16745 30340 16779
rect 30288 16736 30340 16745
rect 46296 16643 46348 16652
rect 46296 16609 46305 16643
rect 46305 16609 46339 16643
rect 46339 16609 46348 16643
rect 46296 16600 46348 16609
rect 48136 16643 48188 16652
rect 48136 16609 48145 16643
rect 48145 16609 48179 16643
rect 48179 16609 48188 16643
rect 48136 16600 48188 16609
rect 29828 16575 29880 16584
rect 29828 16541 29837 16575
rect 29837 16541 29871 16575
rect 29871 16541 29880 16575
rect 29828 16532 29880 16541
rect 30196 16532 30248 16584
rect 32864 16532 32916 16584
rect 30380 16464 30432 16516
rect 31484 16464 31536 16516
rect 31668 16464 31720 16516
rect 47676 16464 47728 16516
rect 30748 16396 30800 16448
rect 31944 16439 31996 16448
rect 31944 16405 31953 16439
rect 31953 16405 31987 16439
rect 31987 16405 31996 16439
rect 31944 16396 31996 16405
rect 36544 16396 36596 16448
rect 47492 16396 47544 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 11520 16192 11572 16244
rect 11796 16192 11848 16244
rect 15844 16192 15896 16244
rect 11704 16167 11756 16176
rect 11704 16133 11713 16167
rect 11713 16133 11747 16167
rect 11747 16133 11756 16167
rect 11704 16124 11756 16133
rect 14280 16124 14332 16176
rect 15384 16124 15436 16176
rect 27160 16192 27212 16244
rect 27436 16235 27488 16244
rect 27436 16201 27445 16235
rect 27445 16201 27479 16235
rect 27479 16201 27488 16235
rect 27436 16192 27488 16201
rect 28264 16192 28316 16244
rect 28908 16192 28960 16244
rect 29644 16235 29696 16244
rect 29644 16201 29653 16235
rect 29653 16201 29687 16235
rect 29687 16201 29696 16235
rect 29644 16192 29696 16201
rect 11520 16099 11572 16108
rect 11520 16065 11529 16099
rect 11529 16065 11563 16099
rect 11563 16065 11572 16099
rect 11520 16056 11572 16065
rect 16672 16099 16724 16108
rect 16672 16065 16681 16099
rect 16681 16065 16715 16099
rect 16715 16065 16724 16099
rect 16672 16056 16724 16065
rect 18328 16056 18380 16108
rect 18972 16099 19024 16108
rect 18972 16065 18981 16099
rect 18981 16065 19015 16099
rect 19015 16065 19024 16099
rect 18972 16056 19024 16065
rect 20720 16056 20772 16108
rect 20904 16099 20956 16108
rect 20904 16065 20913 16099
rect 20913 16065 20947 16099
rect 20947 16065 20956 16099
rect 20904 16056 20956 16065
rect 18512 16031 18564 16040
rect 20 15920 72 15972
rect 18512 15997 18521 16031
rect 18521 15997 18555 16031
rect 18555 15997 18564 16031
rect 18512 15988 18564 15997
rect 19524 16031 19576 16040
rect 19524 15997 19533 16031
rect 19533 15997 19567 16031
rect 19567 15997 19576 16031
rect 19524 15988 19576 15997
rect 20076 15988 20128 16040
rect 25136 16099 25188 16108
rect 25136 16065 25145 16099
rect 25145 16065 25179 16099
rect 25179 16065 25188 16099
rect 25136 16056 25188 16065
rect 25688 16056 25740 16108
rect 28080 16056 28132 16108
rect 26608 15988 26660 16040
rect 20168 15920 20220 15972
rect 20628 15920 20680 15972
rect 13176 15852 13228 15904
rect 23020 15852 23072 15904
rect 25044 15852 25096 15904
rect 25320 15895 25372 15904
rect 25320 15861 25329 15895
rect 25329 15861 25363 15895
rect 25363 15861 25372 15895
rect 25320 15852 25372 15861
rect 27068 15920 27120 15972
rect 27344 15852 27396 15904
rect 29000 16056 29052 16108
rect 36544 16192 36596 16244
rect 30840 16124 30892 16176
rect 31024 16124 31076 16176
rect 30748 16056 30800 16108
rect 31944 16124 31996 16176
rect 31576 16099 31628 16108
rect 28724 16031 28776 16040
rect 28724 15997 28733 16031
rect 28733 15997 28767 16031
rect 28767 15997 28776 16031
rect 28724 15988 28776 15997
rect 28540 15920 28592 15972
rect 29184 15988 29236 16040
rect 30840 15988 30892 16040
rect 31024 15988 31076 16040
rect 31576 16065 31585 16099
rect 31585 16065 31619 16099
rect 31619 16065 31628 16099
rect 31576 16056 31628 16065
rect 32128 16099 32180 16108
rect 32128 16065 32137 16099
rect 32137 16065 32171 16099
rect 32171 16065 32180 16099
rect 32128 16056 32180 16065
rect 32220 16056 32272 16108
rect 31484 15988 31536 16040
rect 29092 15920 29144 15972
rect 29184 15852 29236 15904
rect 29552 15852 29604 15904
rect 31760 15852 31812 15904
rect 46756 15920 46808 15972
rect 33508 15895 33560 15904
rect 33508 15861 33517 15895
rect 33517 15861 33551 15895
rect 33551 15861 33560 15895
rect 33508 15852 33560 15861
rect 46296 15852 46348 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 2412 15580 2464 15632
rect 19524 15648 19576 15700
rect 21180 15648 21232 15700
rect 22560 15691 22612 15700
rect 22560 15657 22569 15691
rect 22569 15657 22603 15691
rect 22603 15657 22612 15691
rect 22560 15648 22612 15657
rect 25044 15648 25096 15700
rect 26700 15648 26752 15700
rect 27436 15691 27488 15700
rect 27436 15657 27445 15691
rect 27445 15657 27479 15691
rect 27479 15657 27488 15691
rect 27436 15648 27488 15657
rect 18696 15580 18748 15632
rect 7656 15512 7708 15564
rect 18420 15512 18472 15564
rect 29092 15580 29144 15632
rect 32864 15623 32916 15632
rect 32864 15589 32873 15623
rect 32873 15589 32907 15623
rect 32907 15589 32916 15623
rect 32864 15580 32916 15589
rect 28080 15512 28132 15564
rect 46296 15555 46348 15564
rect 46296 15521 46305 15555
rect 46305 15521 46339 15555
rect 46339 15521 46348 15555
rect 46296 15512 46348 15521
rect 48136 15555 48188 15564
rect 48136 15521 48145 15555
rect 48145 15521 48179 15555
rect 48179 15521 48188 15555
rect 48136 15512 48188 15521
rect 18328 15444 18380 15496
rect 20720 15487 20772 15496
rect 20720 15453 20729 15487
rect 20729 15453 20763 15487
rect 20763 15453 20772 15487
rect 20720 15444 20772 15453
rect 20904 15444 20956 15496
rect 21088 15487 21140 15496
rect 21088 15453 21097 15487
rect 21097 15453 21131 15487
rect 21131 15453 21140 15487
rect 21088 15444 21140 15453
rect 24860 15444 24912 15496
rect 26608 15487 26660 15496
rect 26608 15453 26617 15487
rect 26617 15453 26651 15487
rect 26651 15453 26660 15487
rect 26608 15444 26660 15453
rect 26884 15487 26936 15496
rect 26884 15453 26893 15487
rect 26893 15453 26927 15487
rect 26927 15453 26936 15487
rect 26884 15444 26936 15453
rect 19432 15308 19484 15360
rect 20536 15351 20588 15360
rect 20536 15317 20545 15351
rect 20545 15317 20579 15351
rect 20579 15317 20588 15351
rect 20536 15308 20588 15317
rect 22192 15308 22244 15360
rect 23572 15308 23624 15360
rect 23664 15308 23716 15360
rect 24952 15308 25004 15360
rect 25872 15308 25924 15360
rect 26148 15308 26200 15360
rect 28356 15444 28408 15496
rect 29184 15444 29236 15496
rect 29552 15487 29604 15496
rect 29552 15453 29561 15487
rect 29561 15453 29595 15487
rect 29595 15453 29604 15487
rect 29552 15444 29604 15453
rect 31116 15444 31168 15496
rect 31484 15487 31536 15496
rect 31484 15453 31493 15487
rect 31493 15453 31527 15487
rect 31527 15453 31536 15487
rect 31484 15444 31536 15453
rect 31760 15487 31812 15496
rect 31760 15453 31794 15487
rect 31794 15453 31812 15487
rect 31760 15444 31812 15453
rect 28724 15308 28776 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 20536 15104 20588 15156
rect 20720 15104 20772 15156
rect 22192 15147 22244 15156
rect 22192 15113 22201 15147
rect 22201 15113 22235 15147
rect 22235 15113 22244 15147
rect 22192 15104 22244 15113
rect 22560 15104 22612 15156
rect 32220 15104 32272 15156
rect 46664 15104 46716 15156
rect 17684 15079 17736 15088
rect 17684 15045 17693 15079
rect 17693 15045 17727 15079
rect 17727 15045 17736 15079
rect 17684 15036 17736 15045
rect 19156 15079 19208 15088
rect 19156 15045 19165 15079
rect 19165 15045 19199 15079
rect 19199 15045 19208 15079
rect 19156 15036 19208 15045
rect 21640 15036 21692 15088
rect 22100 15036 22152 15088
rect 18328 15011 18380 15020
rect 18328 14977 18337 15011
rect 18337 14977 18371 15011
rect 18371 14977 18380 15011
rect 18328 14968 18380 14977
rect 21180 14968 21232 15020
rect 23388 15036 23440 15088
rect 31024 15036 31076 15088
rect 2872 14900 2924 14952
rect 19156 14900 19208 14952
rect 17868 14875 17920 14884
rect 17868 14841 17877 14875
rect 17877 14841 17911 14875
rect 17911 14841 17920 14875
rect 17868 14832 17920 14841
rect 20720 14900 20772 14952
rect 22192 14900 22244 14952
rect 23572 15011 23624 15020
rect 23572 14977 23581 15011
rect 23581 14977 23615 15011
rect 23615 14977 23624 15011
rect 23572 14968 23624 14977
rect 24584 14968 24636 15020
rect 25136 15011 25188 15020
rect 25136 14977 25145 15011
rect 25145 14977 25179 15011
rect 25179 14977 25188 15011
rect 25136 14968 25188 14977
rect 25964 14968 26016 15020
rect 27988 14968 28040 15020
rect 28448 14968 28500 15020
rect 30840 14968 30892 15020
rect 33508 15036 33560 15088
rect 31576 15011 31628 15020
rect 22928 14900 22980 14952
rect 21456 14832 21508 14884
rect 22284 14832 22336 14884
rect 27528 14900 27580 14952
rect 31576 14977 31585 15011
rect 31585 14977 31619 15011
rect 31619 14977 31628 15011
rect 31576 14968 31628 14977
rect 31668 14968 31720 15020
rect 46848 14968 46900 15020
rect 47584 15011 47636 15020
rect 47584 14977 47593 15011
rect 47593 14977 47627 15011
rect 47627 14977 47636 15011
rect 47584 14968 47636 14977
rect 24952 14832 25004 14884
rect 28264 14832 28316 14884
rect 19432 14764 19484 14816
rect 20628 14764 20680 14816
rect 23480 14764 23532 14816
rect 24860 14764 24912 14816
rect 27160 14807 27212 14816
rect 27160 14773 27169 14807
rect 27169 14773 27203 14807
rect 27203 14773 27212 14807
rect 27160 14764 27212 14773
rect 27620 14764 27672 14816
rect 46480 14764 46532 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 20904 14560 20956 14612
rect 17960 14424 18012 14476
rect 20168 14424 20220 14476
rect 19432 14399 19484 14408
rect 19432 14365 19441 14399
rect 19441 14365 19475 14399
rect 19475 14365 19484 14399
rect 19432 14356 19484 14365
rect 19616 14288 19668 14340
rect 17316 14263 17368 14272
rect 17316 14229 17325 14263
rect 17325 14229 17359 14263
rect 17359 14229 17368 14263
rect 17316 14220 17368 14229
rect 17408 14220 17460 14272
rect 17592 14220 17644 14272
rect 19248 14263 19300 14272
rect 19248 14229 19257 14263
rect 19257 14229 19291 14263
rect 19291 14229 19300 14263
rect 19248 14220 19300 14229
rect 20536 14492 20588 14544
rect 21180 14560 21232 14612
rect 21456 14560 21508 14612
rect 23112 14560 23164 14612
rect 24584 14603 24636 14612
rect 21272 14492 21324 14544
rect 22744 14467 22796 14476
rect 22744 14433 22753 14467
rect 22753 14433 22787 14467
rect 22787 14433 22796 14467
rect 22744 14424 22796 14433
rect 23664 14492 23716 14544
rect 23848 14492 23900 14544
rect 24584 14569 24593 14603
rect 24593 14569 24627 14603
rect 24627 14569 24636 14603
rect 24584 14560 24636 14569
rect 24676 14560 24728 14612
rect 26884 14560 26936 14612
rect 27068 14560 27120 14612
rect 27436 14560 27488 14612
rect 25688 14492 25740 14544
rect 26148 14492 26200 14544
rect 28448 14492 28500 14544
rect 28908 14492 28960 14544
rect 20812 14356 20864 14408
rect 21180 14356 21232 14408
rect 23112 14356 23164 14408
rect 20720 14288 20772 14340
rect 21088 14288 21140 14340
rect 22008 14288 22060 14340
rect 22468 14288 22520 14340
rect 20904 14220 20956 14272
rect 21640 14220 21692 14272
rect 22192 14263 22244 14272
rect 22192 14229 22201 14263
rect 22201 14229 22235 14263
rect 22235 14229 22244 14263
rect 22192 14220 22244 14229
rect 23296 14288 23348 14340
rect 24032 14356 24084 14408
rect 24952 14424 25004 14476
rect 26700 14424 26752 14476
rect 46480 14467 46532 14476
rect 27160 14399 27212 14408
rect 27160 14365 27169 14399
rect 27169 14365 27203 14399
rect 27203 14365 27212 14399
rect 27160 14356 27212 14365
rect 27528 14399 27580 14408
rect 27528 14365 27537 14399
rect 27537 14365 27571 14399
rect 27571 14365 27580 14399
rect 27528 14356 27580 14365
rect 46480 14433 46489 14467
rect 46489 14433 46523 14467
rect 46523 14433 46532 14467
rect 46480 14424 46532 14433
rect 28356 14399 28408 14408
rect 28356 14365 28365 14399
rect 28365 14365 28399 14399
rect 28399 14365 28408 14399
rect 28356 14356 28408 14365
rect 31484 14399 31536 14408
rect 31484 14365 31493 14399
rect 31493 14365 31527 14399
rect 31527 14365 31536 14399
rect 31484 14356 31536 14365
rect 22836 14220 22888 14272
rect 25044 14288 25096 14340
rect 24400 14220 24452 14272
rect 24676 14220 24728 14272
rect 27160 14220 27212 14272
rect 47676 14288 47728 14340
rect 48136 14331 48188 14340
rect 48136 14297 48145 14331
rect 48145 14297 48179 14331
rect 48179 14297 48188 14331
rect 48136 14288 48188 14297
rect 27620 14220 27672 14272
rect 28080 14220 28132 14272
rect 32404 14220 32456 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 19248 13948 19300 14000
rect 2044 13923 2096 13932
rect 2044 13889 2053 13923
rect 2053 13889 2087 13923
rect 2087 13889 2096 13923
rect 2044 13880 2096 13889
rect 17408 13923 17460 13932
rect 17408 13889 17417 13923
rect 17417 13889 17451 13923
rect 17451 13889 17460 13923
rect 17408 13880 17460 13889
rect 17500 13923 17552 13932
rect 17500 13889 17509 13923
rect 17509 13889 17543 13923
rect 17543 13889 17552 13923
rect 17500 13880 17552 13889
rect 17960 13880 18012 13932
rect 21272 14016 21324 14068
rect 22468 14016 22520 14068
rect 23388 14016 23440 14068
rect 27160 14016 27212 14068
rect 20628 13991 20680 14000
rect 20628 13957 20637 13991
rect 20637 13957 20671 13991
rect 20671 13957 20680 13991
rect 20628 13948 20680 13957
rect 20536 13923 20588 13932
rect 20536 13889 20543 13923
rect 20543 13889 20588 13923
rect 20536 13880 20588 13889
rect 18144 13812 18196 13864
rect 1584 13676 1636 13728
rect 2872 13719 2924 13728
rect 2872 13685 2881 13719
rect 2881 13685 2915 13719
rect 2915 13685 2924 13719
rect 2872 13676 2924 13685
rect 17224 13719 17276 13728
rect 17224 13685 17233 13719
rect 17233 13685 17267 13719
rect 17267 13685 17276 13719
rect 17224 13676 17276 13685
rect 19248 13676 19300 13728
rect 20628 13812 20680 13864
rect 20904 13880 20956 13932
rect 22008 13948 22060 14000
rect 23296 13948 23348 14000
rect 23664 13948 23716 14000
rect 24032 13948 24084 14000
rect 23480 13923 23532 13932
rect 23480 13889 23514 13923
rect 23514 13889 23532 13923
rect 23480 13880 23532 13889
rect 27160 13923 27212 13932
rect 27160 13889 27169 13923
rect 27169 13889 27203 13923
rect 27203 13889 27212 13923
rect 27160 13880 27212 13889
rect 27620 14016 27672 14068
rect 31024 14016 31076 14068
rect 31852 14016 31904 14068
rect 27436 13923 27488 13932
rect 27436 13889 27445 13923
rect 27445 13889 27479 13923
rect 27479 13889 27488 13923
rect 27436 13880 27488 13889
rect 22284 13855 22336 13864
rect 22284 13821 22293 13855
rect 22293 13821 22327 13855
rect 22327 13821 22336 13855
rect 22284 13812 22336 13821
rect 21640 13744 21692 13796
rect 20996 13719 21048 13728
rect 20996 13685 21005 13719
rect 21005 13685 21039 13719
rect 21039 13685 21048 13719
rect 20996 13676 21048 13685
rect 21548 13676 21600 13728
rect 25596 13812 25648 13864
rect 29552 13948 29604 14000
rect 32404 13991 32456 14000
rect 28080 13880 28132 13932
rect 28632 13880 28684 13932
rect 32404 13957 32413 13991
rect 32413 13957 32447 13991
rect 32447 13957 32456 13991
rect 32404 13948 32456 13957
rect 31576 13880 31628 13932
rect 32036 13812 32088 13864
rect 32220 13855 32272 13864
rect 32220 13821 32229 13855
rect 32229 13821 32263 13855
rect 32263 13821 32272 13855
rect 32220 13812 32272 13821
rect 46204 13880 46256 13932
rect 47860 13923 47912 13932
rect 47860 13889 47869 13923
rect 47869 13889 47903 13923
rect 47903 13889 47912 13923
rect 47860 13880 47912 13889
rect 25320 13676 25372 13728
rect 27896 13676 27948 13728
rect 28908 13676 28960 13728
rect 30748 13719 30800 13728
rect 30748 13685 30757 13719
rect 30757 13685 30791 13719
rect 30791 13685 30800 13719
rect 30748 13676 30800 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 20536 13472 20588 13524
rect 22284 13515 22336 13524
rect 22284 13481 22293 13515
rect 22293 13481 22327 13515
rect 22327 13481 22336 13515
rect 22284 13472 22336 13481
rect 23572 13472 23624 13524
rect 25136 13472 25188 13524
rect 26700 13472 26752 13524
rect 32220 13472 32272 13524
rect 47676 13515 47728 13524
rect 47676 13481 47685 13515
rect 47685 13481 47719 13515
rect 47719 13481 47728 13515
rect 47676 13472 47728 13481
rect 2872 13404 2924 13456
rect 4068 13404 4120 13456
rect 6920 13404 6972 13456
rect 22836 13404 22888 13456
rect 1584 13379 1636 13388
rect 1584 13345 1593 13379
rect 1593 13345 1627 13379
rect 1627 13345 1636 13379
rect 1584 13336 1636 13345
rect 2780 13379 2832 13388
rect 2780 13345 2789 13379
rect 2789 13345 2823 13379
rect 2823 13345 2832 13379
rect 2780 13336 2832 13345
rect 12532 13336 12584 13388
rect 20720 13336 20772 13388
rect 21548 13379 21600 13388
rect 19248 13311 19300 13320
rect 19248 13277 19257 13311
rect 19257 13277 19291 13311
rect 19291 13277 19300 13311
rect 19248 13268 19300 13277
rect 20996 13268 21048 13320
rect 21548 13345 21557 13379
rect 21557 13345 21591 13379
rect 21591 13345 21600 13379
rect 21548 13336 21600 13345
rect 21640 13336 21692 13388
rect 27344 13336 27396 13388
rect 27896 13336 27948 13388
rect 28540 13336 28592 13388
rect 31116 13379 31168 13388
rect 31116 13345 31125 13379
rect 31125 13345 31159 13379
rect 31159 13345 31168 13379
rect 31116 13336 31168 13345
rect 21456 13268 21508 13320
rect 22468 13311 22520 13320
rect 22468 13277 22477 13311
rect 22477 13277 22511 13311
rect 22511 13277 22520 13311
rect 22468 13268 22520 13277
rect 23664 13268 23716 13320
rect 24216 13268 24268 13320
rect 25320 13268 25372 13320
rect 27620 13268 27672 13320
rect 30472 13268 30524 13320
rect 30748 13268 30800 13320
rect 14004 13200 14056 13252
rect 17224 13200 17276 13252
rect 21824 13200 21876 13252
rect 23296 13243 23348 13252
rect 17316 13132 17368 13184
rect 18052 13132 18104 13184
rect 18696 13132 18748 13184
rect 20628 13132 20680 13184
rect 23296 13209 23305 13243
rect 23305 13209 23339 13243
rect 23339 13209 23348 13243
rect 23296 13200 23348 13209
rect 27160 13200 27212 13252
rect 27988 13243 28040 13252
rect 23848 13132 23900 13184
rect 26976 13132 27028 13184
rect 27988 13209 27997 13243
rect 27997 13209 28031 13243
rect 28031 13209 28040 13243
rect 27988 13200 28040 13209
rect 27712 13132 27764 13184
rect 28540 13132 28592 13184
rect 30564 13132 30616 13184
rect 31668 13132 31720 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 14004 12971 14056 12980
rect 14004 12937 14013 12971
rect 14013 12937 14047 12971
rect 14047 12937 14056 12971
rect 14004 12928 14056 12937
rect 18144 12971 18196 12980
rect 18144 12937 18153 12971
rect 18153 12937 18187 12971
rect 18187 12937 18196 12971
rect 18144 12928 18196 12937
rect 21180 12971 21232 12980
rect 21180 12937 21189 12971
rect 21189 12937 21223 12971
rect 21223 12937 21232 12971
rect 21180 12928 21232 12937
rect 8484 12792 8536 12844
rect 9772 12835 9824 12844
rect 9772 12801 9781 12835
rect 9781 12801 9815 12835
rect 9815 12801 9824 12835
rect 9772 12792 9824 12801
rect 11612 12792 11664 12844
rect 15476 12792 15528 12844
rect 18052 12860 18104 12912
rect 19616 12860 19668 12912
rect 20076 12860 20128 12912
rect 22652 12860 22704 12912
rect 1400 12767 1452 12776
rect 1400 12733 1409 12767
rect 1409 12733 1443 12767
rect 1443 12733 1452 12767
rect 1400 12724 1452 12733
rect 7932 12724 7984 12776
rect 10508 12724 10560 12776
rect 21548 12792 21600 12844
rect 22468 12792 22520 12844
rect 22928 12792 22980 12844
rect 23296 12928 23348 12980
rect 27344 12971 27396 12980
rect 27344 12937 27353 12971
rect 27353 12937 27387 12971
rect 27387 12937 27396 12971
rect 28908 12971 28960 12980
rect 27344 12928 27396 12937
rect 23848 12860 23900 12912
rect 24400 12903 24452 12912
rect 24400 12869 24409 12903
rect 24409 12869 24443 12903
rect 24443 12869 24452 12903
rect 24400 12860 24452 12869
rect 25320 12860 25372 12912
rect 27804 12903 27856 12912
rect 27804 12869 27813 12903
rect 27813 12869 27847 12903
rect 27847 12869 27856 12903
rect 27804 12860 27856 12869
rect 28908 12937 28917 12971
rect 28917 12937 28951 12971
rect 28951 12937 28960 12971
rect 28908 12928 28960 12937
rect 32036 12928 32088 12980
rect 31668 12860 31720 12912
rect 32220 12860 32272 12912
rect 21456 12724 21508 12776
rect 23664 12724 23716 12776
rect 25136 12835 25188 12844
rect 25136 12801 25145 12835
rect 25145 12801 25179 12835
rect 25179 12801 25188 12835
rect 25136 12792 25188 12801
rect 26700 12792 26752 12844
rect 27712 12835 27764 12844
rect 27712 12801 27721 12835
rect 27721 12801 27755 12835
rect 27755 12801 27764 12835
rect 27712 12792 27764 12801
rect 28632 12792 28684 12844
rect 25044 12724 25096 12776
rect 27620 12724 27672 12776
rect 27896 12767 27948 12776
rect 27896 12733 27905 12767
rect 27905 12733 27939 12767
rect 27939 12733 27948 12767
rect 27896 12724 27948 12733
rect 22560 12656 22612 12708
rect 18604 12588 18656 12640
rect 19432 12588 19484 12640
rect 22192 12631 22244 12640
rect 22192 12597 22201 12631
rect 22201 12597 22235 12631
rect 22235 12597 22244 12631
rect 22192 12588 22244 12597
rect 23848 12588 23900 12640
rect 25320 12631 25372 12640
rect 25320 12597 25329 12631
rect 25329 12597 25363 12631
rect 25363 12597 25372 12631
rect 25320 12588 25372 12597
rect 25688 12588 25740 12640
rect 25964 12631 26016 12640
rect 25964 12597 25973 12631
rect 25973 12597 26007 12631
rect 26007 12597 26016 12631
rect 25964 12588 26016 12597
rect 26332 12656 26384 12708
rect 27528 12656 27580 12708
rect 30840 12792 30892 12844
rect 31024 12792 31076 12844
rect 42800 12656 42852 12708
rect 46848 12656 46900 12708
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 23388 12384 23440 12436
rect 19248 12316 19300 12368
rect 11612 12223 11664 12232
rect 11612 12189 11621 12223
rect 11621 12189 11655 12223
rect 11655 12189 11664 12223
rect 11612 12180 11664 12189
rect 17868 12180 17920 12232
rect 20076 12316 20128 12368
rect 22560 12316 22612 12368
rect 21088 12248 21140 12300
rect 21548 12223 21600 12232
rect 21548 12189 21557 12223
rect 21557 12189 21591 12223
rect 21591 12189 21600 12223
rect 21548 12180 21600 12189
rect 21824 12291 21876 12300
rect 21824 12257 21833 12291
rect 21833 12257 21867 12291
rect 21867 12257 21876 12291
rect 21824 12248 21876 12257
rect 23020 12248 23072 12300
rect 24124 12316 24176 12368
rect 25320 12384 25372 12436
rect 25596 12384 25648 12436
rect 25872 12384 25924 12436
rect 26608 12384 26660 12436
rect 30472 12384 30524 12436
rect 38476 12384 38528 12436
rect 46848 12384 46900 12436
rect 27068 12316 27120 12368
rect 28540 12316 28592 12368
rect 30380 12316 30432 12368
rect 30840 12316 30892 12368
rect 23848 12291 23900 12300
rect 23848 12257 23853 12291
rect 23853 12257 23887 12291
rect 23887 12257 23900 12291
rect 23848 12248 23900 12257
rect 26148 12248 26200 12300
rect 19616 12112 19668 12164
rect 20076 12112 20128 12164
rect 22192 12180 22244 12232
rect 23204 12180 23256 12232
rect 24952 12223 25004 12232
rect 23480 12112 23532 12164
rect 24952 12189 24961 12223
rect 24961 12189 24995 12223
rect 24995 12189 25004 12223
rect 24952 12180 25004 12189
rect 25136 12180 25188 12232
rect 25688 12223 25740 12232
rect 24400 12112 24452 12164
rect 25688 12189 25697 12223
rect 25697 12189 25731 12223
rect 25731 12189 25740 12223
rect 25688 12180 25740 12189
rect 26332 12180 26384 12232
rect 27160 12223 27212 12232
rect 27160 12189 27169 12223
rect 27169 12189 27203 12223
rect 27203 12189 27212 12223
rect 27160 12180 27212 12189
rect 27896 12248 27948 12300
rect 27988 12248 28040 12300
rect 11704 12087 11756 12096
rect 11704 12053 11713 12087
rect 11713 12053 11747 12087
rect 11747 12053 11756 12087
rect 11704 12044 11756 12053
rect 19340 12044 19392 12096
rect 22284 12087 22336 12096
rect 22284 12053 22293 12087
rect 22293 12053 22327 12087
rect 22327 12053 22336 12087
rect 22284 12044 22336 12053
rect 22652 12044 22704 12096
rect 26240 12087 26292 12096
rect 26240 12053 26249 12087
rect 26249 12053 26283 12087
rect 26283 12053 26292 12087
rect 26240 12044 26292 12053
rect 26424 12112 26476 12164
rect 27712 12223 27764 12232
rect 27712 12189 27721 12223
rect 27721 12189 27755 12223
rect 27755 12189 27764 12223
rect 27712 12180 27764 12189
rect 28264 12180 28316 12232
rect 28448 12223 28500 12232
rect 28448 12189 28457 12223
rect 28457 12189 28491 12223
rect 28491 12189 28500 12223
rect 28448 12180 28500 12189
rect 28540 12180 28592 12232
rect 31852 12223 31904 12232
rect 31852 12189 31861 12223
rect 31861 12189 31895 12223
rect 31895 12189 31904 12223
rect 31852 12180 31904 12189
rect 30656 12112 30708 12164
rect 31576 12112 31628 12164
rect 27068 12044 27120 12096
rect 27528 12044 27580 12096
rect 28080 12044 28132 12096
rect 30748 12044 30800 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 12716 11840 12768 11892
rect 21548 11840 21600 11892
rect 24124 11840 24176 11892
rect 24952 11840 25004 11892
rect 27436 11840 27488 11892
rect 21824 11772 21876 11824
rect 26792 11772 26844 11824
rect 26976 11815 27028 11824
rect 26976 11781 26985 11815
rect 26985 11781 27019 11815
rect 27019 11781 27028 11815
rect 26976 11772 27028 11781
rect 27896 11772 27948 11824
rect 19892 11704 19944 11756
rect 19064 11679 19116 11688
rect 19064 11645 19073 11679
rect 19073 11645 19107 11679
rect 19107 11645 19116 11679
rect 20536 11704 20588 11756
rect 22192 11747 22244 11756
rect 22192 11713 22201 11747
rect 22201 11713 22235 11747
rect 22235 11713 22244 11747
rect 22192 11704 22244 11713
rect 24400 11747 24452 11756
rect 19064 11636 19116 11645
rect 22744 11636 22796 11688
rect 17040 11500 17092 11552
rect 18972 11500 19024 11552
rect 20536 11543 20588 11552
rect 20536 11509 20545 11543
rect 20545 11509 20579 11543
rect 20579 11509 20588 11543
rect 20536 11500 20588 11509
rect 22468 11568 22520 11620
rect 24400 11713 24409 11747
rect 24409 11713 24443 11747
rect 24443 11713 24452 11747
rect 24400 11704 24452 11713
rect 24216 11636 24268 11688
rect 25780 11704 25832 11756
rect 26332 11704 26384 11756
rect 26700 11704 26752 11756
rect 27344 11704 27396 11756
rect 28080 11772 28132 11824
rect 31852 11840 31904 11892
rect 28356 11704 28408 11756
rect 30380 11747 30432 11790
rect 30380 11738 30389 11747
rect 30389 11738 30423 11747
rect 30423 11738 30432 11747
rect 30472 11747 30524 11756
rect 30472 11713 30481 11747
rect 30481 11713 30515 11747
rect 30515 11713 30524 11747
rect 30472 11704 30524 11713
rect 30656 11747 30708 11756
rect 30656 11713 30665 11747
rect 30665 11713 30699 11747
rect 30699 11713 30708 11747
rect 30656 11704 30708 11713
rect 42800 11772 42852 11824
rect 25044 11636 25096 11688
rect 22652 11500 22704 11552
rect 22744 11500 22796 11552
rect 25596 11500 25648 11552
rect 26976 11543 27028 11552
rect 26976 11509 26985 11543
rect 26985 11509 27019 11543
rect 27019 11509 27028 11543
rect 26976 11500 27028 11509
rect 29644 11636 29696 11688
rect 30564 11636 30616 11688
rect 37464 11679 37516 11688
rect 37464 11645 37473 11679
rect 37473 11645 37507 11679
rect 37507 11645 37516 11679
rect 37464 11636 37516 11645
rect 29736 11568 29788 11620
rect 31300 11568 31352 11620
rect 27896 11500 27948 11552
rect 27988 11500 28040 11552
rect 30012 11543 30064 11552
rect 30012 11509 30021 11543
rect 30021 11509 30055 11543
rect 30055 11509 30064 11543
rect 30012 11500 30064 11509
rect 30104 11500 30156 11552
rect 37280 11568 37332 11620
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 18052 11296 18104 11348
rect 21824 11296 21876 11348
rect 23480 11296 23532 11348
rect 2504 11135 2556 11144
rect 2504 11101 2513 11135
rect 2513 11101 2547 11135
rect 2547 11101 2556 11135
rect 2504 11092 2556 11101
rect 1860 11067 1912 11076
rect 1860 11033 1869 11067
rect 1869 11033 1903 11067
rect 1903 11033 1912 11067
rect 1860 11024 1912 11033
rect 11704 11203 11756 11212
rect 11704 11169 11713 11203
rect 11713 11169 11747 11203
rect 11747 11169 11756 11203
rect 11704 11160 11756 11169
rect 13084 11203 13136 11212
rect 13084 11169 13093 11203
rect 13093 11169 13127 11203
rect 13127 11169 13136 11203
rect 13084 11160 13136 11169
rect 18972 11160 19024 11212
rect 20260 11160 20312 11212
rect 20720 11160 20772 11212
rect 14188 11092 14240 11144
rect 17960 11092 18012 11144
rect 19432 11092 19484 11144
rect 22008 11092 22060 11144
rect 18788 11024 18840 11076
rect 19248 11024 19300 11076
rect 22284 11024 22336 11076
rect 24676 11067 24728 11076
rect 24676 11033 24710 11067
rect 24710 11033 24728 11067
rect 24676 11024 24728 11033
rect 25964 11296 26016 11348
rect 27160 11296 27212 11348
rect 30472 11296 30524 11348
rect 37464 11296 37516 11348
rect 26148 11228 26200 11280
rect 30104 11228 30156 11280
rect 26332 11160 26384 11212
rect 27160 11160 27212 11212
rect 27896 11160 27948 11212
rect 29552 11160 29604 11212
rect 26240 11135 26292 11144
rect 26240 11101 26249 11135
rect 26249 11101 26283 11135
rect 26283 11101 26292 11135
rect 26240 11092 26292 11101
rect 26424 11135 26476 11144
rect 26424 11101 26433 11135
rect 26433 11101 26467 11135
rect 26467 11101 26476 11135
rect 26424 11092 26476 11101
rect 26608 11135 26660 11144
rect 26608 11101 26617 11135
rect 26617 11101 26651 11135
rect 26651 11101 26660 11135
rect 26608 11092 26660 11101
rect 26792 11135 26844 11144
rect 26792 11101 26801 11135
rect 26801 11101 26835 11135
rect 26835 11101 26844 11135
rect 26792 11092 26844 11101
rect 26976 11092 27028 11144
rect 28908 11135 28960 11144
rect 28908 11101 28917 11135
rect 28917 11101 28951 11135
rect 28951 11101 28960 11135
rect 28908 11092 28960 11101
rect 30748 11135 30800 11144
rect 30748 11101 30782 11135
rect 30782 11101 30800 11135
rect 30748 11092 30800 11101
rect 37280 11135 37332 11144
rect 37280 11101 37289 11135
rect 37289 11101 37323 11135
rect 37323 11101 37332 11135
rect 37280 11092 37332 11101
rect 47124 11135 47176 11144
rect 47124 11101 47133 11135
rect 47133 11101 47167 11135
rect 47167 11101 47176 11135
rect 47124 11092 47176 11101
rect 47952 11135 48004 11144
rect 47952 11101 47961 11135
rect 47961 11101 47995 11135
rect 47995 11101 48004 11135
rect 47952 11092 48004 11101
rect 2596 10999 2648 11008
rect 2596 10965 2605 10999
rect 2605 10965 2639 10999
rect 2639 10965 2648 10999
rect 2596 10956 2648 10965
rect 18328 10956 18380 11008
rect 19156 10956 19208 11008
rect 25320 10956 25372 11008
rect 26976 10999 27028 11008
rect 26976 10965 26985 10999
rect 26985 10965 27019 10999
rect 27019 10965 27028 10999
rect 26976 10956 27028 10965
rect 27528 11024 27580 11076
rect 29644 11067 29696 11076
rect 29644 11033 29653 11067
rect 29653 11033 29687 11067
rect 29687 11033 29696 11067
rect 29644 11024 29696 11033
rect 30380 11024 30432 11076
rect 31300 11024 31352 11076
rect 28356 10956 28408 11008
rect 47216 10999 47268 11008
rect 47216 10965 47225 10999
rect 47225 10965 47259 10999
rect 47259 10965 47268 10999
rect 47216 10956 47268 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 18788 10795 18840 10804
rect 18788 10761 18797 10795
rect 18797 10761 18831 10795
rect 18831 10761 18840 10795
rect 18788 10752 18840 10761
rect 19248 10752 19300 10804
rect 21272 10795 21324 10804
rect 2596 10684 2648 10736
rect 18052 10684 18104 10736
rect 21272 10761 21281 10795
rect 21281 10761 21315 10795
rect 21315 10761 21324 10795
rect 21272 10752 21324 10761
rect 24676 10795 24728 10804
rect 24676 10761 24685 10795
rect 24685 10761 24719 10795
rect 24719 10761 24728 10795
rect 24676 10752 24728 10761
rect 25320 10795 25372 10804
rect 25320 10761 25329 10795
rect 25329 10761 25363 10795
rect 25363 10761 25372 10795
rect 25320 10752 25372 10761
rect 18972 10616 19024 10668
rect 19432 10659 19484 10668
rect 1584 10548 1636 10600
rect 2964 10591 3016 10600
rect 2964 10557 2973 10591
rect 2973 10557 3007 10591
rect 3007 10557 3016 10591
rect 2964 10548 3016 10557
rect 19432 10625 19441 10659
rect 19441 10625 19475 10659
rect 19475 10625 19484 10659
rect 19432 10616 19484 10625
rect 19800 10616 19852 10668
rect 20076 10684 20128 10736
rect 20904 10684 20956 10736
rect 21732 10684 21784 10736
rect 20168 10659 20220 10668
rect 20168 10625 20202 10659
rect 20202 10625 20220 10659
rect 20168 10616 20220 10625
rect 23388 10616 23440 10668
rect 19340 10548 19392 10600
rect 23480 10548 23532 10600
rect 24216 10659 24268 10668
rect 24216 10625 24225 10659
rect 24225 10625 24259 10659
rect 24259 10625 24268 10659
rect 24216 10616 24268 10625
rect 24400 10616 24452 10668
rect 27528 10684 27580 10736
rect 30012 10727 30064 10736
rect 30012 10693 30046 10727
rect 30046 10693 30064 10727
rect 30012 10684 30064 10693
rect 47768 10659 47820 10668
rect 22192 10480 22244 10532
rect 24216 10480 24268 10532
rect 24400 10480 24452 10532
rect 23020 10412 23072 10464
rect 26608 10548 26660 10600
rect 29552 10548 29604 10600
rect 30380 10412 30432 10464
rect 47768 10625 47777 10659
rect 47777 10625 47811 10659
rect 47811 10625 47820 10659
rect 47768 10616 47820 10625
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 1584 10251 1636 10260
rect 1584 10217 1593 10251
rect 1593 10217 1627 10251
rect 1627 10217 1636 10251
rect 1584 10208 1636 10217
rect 20168 10208 20220 10260
rect 27160 10251 27212 10260
rect 27160 10217 27169 10251
rect 27169 10217 27203 10251
rect 27203 10217 27212 10251
rect 27160 10208 27212 10217
rect 19340 10140 19392 10192
rect 20444 10140 20496 10192
rect 20536 10140 20588 10192
rect 1952 10004 2004 10056
rect 3056 10004 3108 10056
rect 19156 9936 19208 9988
rect 19432 9979 19484 9988
rect 19432 9945 19441 9979
rect 19441 9945 19475 9979
rect 19475 9945 19484 9979
rect 19432 9936 19484 9945
rect 2780 9911 2832 9920
rect 2780 9877 2789 9911
rect 2789 9877 2823 9911
rect 2823 9877 2832 9911
rect 2780 9868 2832 9877
rect 19340 9868 19392 9920
rect 25320 10072 25372 10124
rect 47952 10140 48004 10192
rect 47216 10072 47268 10124
rect 48136 10115 48188 10124
rect 48136 10081 48145 10115
rect 48145 10081 48179 10115
rect 48179 10081 48188 10115
rect 48136 10072 48188 10081
rect 20996 10004 21048 10056
rect 26976 10004 27028 10056
rect 22100 9868 22152 9920
rect 26608 9868 26660 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 18604 9664 18656 9716
rect 2780 9596 2832 9648
rect 4068 9596 4120 9648
rect 12532 9596 12584 9648
rect 1952 9571 2004 9580
rect 1952 9537 1961 9571
rect 1961 9537 1995 9571
rect 1995 9537 2004 9571
rect 1952 9528 2004 9537
rect 17960 9596 18012 9648
rect 19984 9664 20036 9716
rect 20996 9664 21048 9716
rect 2872 9503 2924 9512
rect 2872 9469 2881 9503
rect 2881 9469 2915 9503
rect 2915 9469 2924 9503
rect 2872 9460 2924 9469
rect 18696 9528 18748 9580
rect 19616 9571 19668 9580
rect 19616 9537 19625 9571
rect 19625 9537 19659 9571
rect 19659 9537 19668 9571
rect 19616 9528 19668 9537
rect 19984 9528 20036 9580
rect 20260 9528 20312 9580
rect 23664 9596 23716 9648
rect 26424 9528 26476 9580
rect 27804 9528 27856 9580
rect 27988 9528 28040 9580
rect 38568 9596 38620 9648
rect 46848 9596 46900 9648
rect 31484 9528 31536 9580
rect 20444 9460 20496 9512
rect 23388 9460 23440 9512
rect 26976 9460 27028 9512
rect 27896 9503 27948 9512
rect 27896 9469 27905 9503
rect 27905 9469 27939 9503
rect 27939 9469 27948 9503
rect 27896 9460 27948 9469
rect 17960 9324 18012 9376
rect 19432 9324 19484 9376
rect 23848 9324 23900 9376
rect 24952 9324 25004 9376
rect 27712 9324 27764 9376
rect 27804 9324 27856 9376
rect 28264 9324 28316 9376
rect 30012 9367 30064 9376
rect 30012 9333 30021 9367
rect 30021 9333 30055 9367
rect 30055 9333 30064 9367
rect 30012 9324 30064 9333
rect 30656 9367 30708 9376
rect 30656 9333 30665 9367
rect 30665 9333 30699 9367
rect 30699 9333 30708 9367
rect 30656 9324 30708 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 17776 9120 17828 9172
rect 22376 9120 22428 9172
rect 27988 9120 28040 9172
rect 24952 9052 25004 9104
rect 19248 9027 19300 9036
rect 19248 8993 19257 9027
rect 19257 8993 19291 9027
rect 19291 8993 19300 9027
rect 19248 8984 19300 8993
rect 24492 8984 24544 9036
rect 19156 8916 19208 8968
rect 19432 8780 19484 8832
rect 19984 8848 20036 8900
rect 20996 8848 21048 8900
rect 22928 8916 22980 8968
rect 23296 8916 23348 8968
rect 23664 8916 23716 8968
rect 25044 8916 25096 8968
rect 25136 8959 25188 8968
rect 25136 8925 25145 8959
rect 25145 8925 25179 8959
rect 25179 8925 25188 8959
rect 26424 8959 26476 8968
rect 25136 8916 25188 8925
rect 26424 8925 26433 8959
rect 26433 8925 26467 8959
rect 26467 8925 26476 8959
rect 26424 8916 26476 8925
rect 48044 9052 48096 9104
rect 27804 8984 27856 9036
rect 30012 9027 30064 9036
rect 30012 8993 30021 9027
rect 30021 8993 30055 9027
rect 30055 8993 30064 9027
rect 30012 8984 30064 8993
rect 30288 9027 30340 9036
rect 30288 8993 30297 9027
rect 30297 8993 30331 9027
rect 30331 8993 30340 9027
rect 30288 8984 30340 8993
rect 27712 8959 27764 8968
rect 27712 8925 27721 8959
rect 27721 8925 27755 8959
rect 27755 8925 27764 8959
rect 27712 8916 27764 8925
rect 27896 8959 27948 8968
rect 27896 8925 27905 8959
rect 27905 8925 27939 8959
rect 27939 8925 27948 8959
rect 27896 8916 27948 8925
rect 21180 8848 21232 8900
rect 22192 8891 22244 8900
rect 20628 8823 20680 8832
rect 20628 8789 20637 8823
rect 20637 8789 20671 8823
rect 20671 8789 20680 8823
rect 20628 8780 20680 8789
rect 20812 8780 20864 8832
rect 22192 8857 22201 8891
rect 22201 8857 22235 8891
rect 22235 8857 22244 8891
rect 22192 8848 22244 8857
rect 23388 8848 23440 8900
rect 26608 8891 26660 8900
rect 26608 8857 26617 8891
rect 26617 8857 26651 8891
rect 26651 8857 26660 8891
rect 26608 8848 26660 8857
rect 30380 8848 30432 8900
rect 47952 8891 48004 8900
rect 47952 8857 47961 8891
rect 47961 8857 47995 8891
rect 47995 8857 48004 8891
rect 47952 8848 48004 8857
rect 23204 8780 23256 8832
rect 24952 8780 25004 8832
rect 27068 8780 27120 8832
rect 38292 8780 38344 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 3608 8576 3660 8628
rect 30288 8576 30340 8628
rect 20444 8508 20496 8560
rect 1860 8483 1912 8492
rect 1860 8449 1869 8483
rect 1869 8449 1903 8483
rect 1903 8449 1912 8483
rect 1860 8440 1912 8449
rect 17960 8483 18012 8492
rect 17960 8449 17969 8483
rect 17969 8449 18003 8483
rect 18003 8449 18012 8483
rect 17960 8440 18012 8449
rect 21548 8508 21600 8560
rect 22100 8508 22152 8560
rect 18144 8415 18196 8424
rect 18144 8381 18153 8415
rect 18153 8381 18187 8415
rect 18187 8381 18196 8415
rect 18144 8372 18196 8381
rect 19340 8415 19392 8424
rect 19340 8381 19349 8415
rect 19349 8381 19383 8415
rect 19383 8381 19392 8415
rect 19340 8372 19392 8381
rect 20260 8304 20312 8356
rect 20812 8483 20864 8492
rect 20812 8449 20821 8483
rect 20821 8449 20855 8483
rect 20855 8449 20864 8483
rect 20812 8440 20864 8449
rect 20996 8483 21048 8492
rect 20996 8449 21005 8483
rect 21005 8449 21039 8483
rect 21039 8449 21048 8483
rect 20996 8440 21048 8449
rect 21180 8440 21232 8492
rect 23112 8551 23164 8560
rect 23112 8517 23146 8551
rect 23146 8517 23164 8551
rect 23112 8508 23164 8517
rect 25688 8508 25740 8560
rect 24952 8440 25004 8492
rect 26976 8483 27028 8492
rect 26976 8449 26985 8483
rect 26985 8449 27019 8483
rect 27019 8449 27028 8483
rect 26976 8440 27028 8449
rect 27252 8483 27304 8492
rect 27252 8449 27286 8483
rect 27286 8449 27304 8483
rect 27252 8440 27304 8449
rect 30656 8508 30708 8560
rect 29736 8483 29788 8492
rect 29736 8449 29745 8483
rect 29745 8449 29779 8483
rect 29779 8449 29788 8483
rect 29736 8440 29788 8449
rect 47768 8483 47820 8492
rect 47768 8449 47777 8483
rect 47777 8449 47811 8483
rect 47811 8449 47820 8483
rect 47768 8440 47820 8449
rect 21824 8304 21876 8356
rect 21916 8304 21968 8356
rect 24216 8347 24268 8356
rect 24216 8313 24225 8347
rect 24225 8313 24259 8347
rect 24259 8313 24268 8347
rect 24216 8304 24268 8313
rect 26240 8347 26292 8356
rect 26240 8313 26249 8347
rect 26249 8313 26283 8347
rect 26283 8313 26292 8347
rect 26240 8304 26292 8313
rect 26792 8304 26844 8356
rect 29828 8304 29880 8356
rect 20352 8279 20404 8288
rect 20352 8245 20361 8279
rect 20361 8245 20395 8279
rect 20395 8245 20404 8279
rect 20352 8236 20404 8245
rect 20628 8236 20680 8288
rect 21548 8236 21600 8288
rect 22284 8236 22336 8288
rect 26608 8236 26660 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 18144 8032 18196 8084
rect 20352 8032 20404 8084
rect 22928 8075 22980 8084
rect 2136 7964 2188 8016
rect 7748 7964 7800 8016
rect 18696 7964 18748 8016
rect 20628 7896 20680 7948
rect 22928 8041 22937 8075
rect 22937 8041 22971 8075
rect 22971 8041 22980 8075
rect 22928 8032 22980 8041
rect 25044 8032 25096 8084
rect 27252 8032 27304 8084
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 18604 7828 18656 7880
rect 23848 7896 23900 7948
rect 18880 7760 18932 7812
rect 16672 7692 16724 7744
rect 23020 7828 23072 7880
rect 25044 7871 25096 7880
rect 23388 7803 23440 7812
rect 23388 7769 23397 7803
rect 23397 7769 23431 7803
rect 23431 7769 23440 7803
rect 23388 7760 23440 7769
rect 23572 7803 23624 7812
rect 23572 7769 23581 7803
rect 23581 7769 23615 7803
rect 23615 7769 23624 7803
rect 23572 7760 23624 7769
rect 25044 7837 25053 7871
rect 25053 7837 25087 7871
rect 25087 7837 25096 7871
rect 25044 7828 25096 7837
rect 25320 7828 25372 7880
rect 26424 7828 26476 7880
rect 26884 7871 26936 7880
rect 26884 7837 26893 7871
rect 26893 7837 26927 7871
rect 26927 7837 26936 7871
rect 26884 7828 26936 7837
rect 27804 7896 27856 7948
rect 27068 7871 27120 7880
rect 27068 7837 27082 7871
rect 27082 7837 27116 7871
rect 27116 7837 27120 7871
rect 27068 7828 27120 7837
rect 27252 7871 27304 7880
rect 27252 7837 27261 7871
rect 27261 7837 27295 7871
rect 27295 7837 27304 7871
rect 27252 7828 27304 7837
rect 27896 7828 27948 7880
rect 37280 7828 37332 7880
rect 46296 7871 46348 7880
rect 46296 7837 46305 7871
rect 46305 7837 46339 7871
rect 46339 7837 46348 7871
rect 46296 7828 46348 7837
rect 26240 7760 26292 7812
rect 27160 7760 27212 7812
rect 35900 7760 35952 7812
rect 46756 7760 46808 7812
rect 48136 7803 48188 7812
rect 48136 7769 48145 7803
rect 48145 7769 48179 7803
rect 48179 7769 48188 7803
rect 48136 7760 48188 7769
rect 22008 7692 22060 7744
rect 24400 7735 24452 7744
rect 24400 7701 24409 7735
rect 24409 7701 24443 7735
rect 24443 7701 24452 7735
rect 24400 7692 24452 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 18880 7531 18932 7540
rect 18880 7497 18889 7531
rect 18889 7497 18923 7531
rect 18923 7497 18932 7531
rect 18880 7488 18932 7497
rect 19432 7531 19484 7540
rect 19432 7497 19441 7531
rect 19441 7497 19475 7531
rect 19475 7497 19484 7531
rect 19432 7488 19484 7497
rect 18604 7352 18656 7404
rect 20444 7488 20496 7540
rect 21824 7488 21876 7540
rect 23572 7488 23624 7540
rect 31208 7488 31260 7540
rect 46756 7531 46808 7540
rect 21916 7420 21968 7472
rect 24400 7420 24452 7472
rect 19984 7352 20036 7404
rect 22008 7352 22060 7404
rect 37280 7395 37332 7404
rect 22192 7284 22244 7336
rect 37280 7361 37289 7395
rect 37289 7361 37323 7395
rect 37323 7361 37332 7395
rect 37280 7352 37332 7361
rect 46756 7497 46765 7531
rect 46765 7497 46799 7531
rect 46799 7497 46808 7531
rect 46756 7488 46808 7497
rect 46296 7420 46348 7472
rect 45652 7352 45704 7404
rect 38016 7327 38068 7336
rect 38016 7293 38025 7327
rect 38025 7293 38059 7327
rect 38059 7293 38068 7327
rect 38016 7284 38068 7293
rect 37372 7216 37424 7268
rect 2044 7191 2096 7200
rect 2044 7157 2053 7191
rect 2053 7157 2087 7191
rect 2087 7157 2096 7191
rect 2044 7148 2096 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 2044 6808 2096 6860
rect 2780 6851 2832 6860
rect 2780 6817 2789 6851
rect 2789 6817 2823 6851
rect 2823 6817 2832 6851
rect 2780 6808 2832 6817
rect 2228 6672 2280 6724
rect 18972 6672 19024 6724
rect 22744 6740 22796 6792
rect 23204 6876 23256 6928
rect 23296 6783 23348 6792
rect 23296 6749 23305 6783
rect 23305 6749 23339 6783
rect 23339 6749 23348 6783
rect 23296 6740 23348 6749
rect 23848 6672 23900 6724
rect 46020 6715 46072 6724
rect 46020 6681 46029 6715
rect 46029 6681 46063 6715
rect 46063 6681 46072 6715
rect 46020 6672 46072 6681
rect 47676 6715 47728 6724
rect 47676 6681 47685 6715
rect 47685 6681 47719 6715
rect 47719 6681 47728 6715
rect 47676 6672 47728 6681
rect 23112 6604 23164 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 2228 6443 2280 6452
rect 2228 6409 2237 6443
rect 2237 6409 2271 6443
rect 2271 6409 2280 6443
rect 2228 6400 2280 6409
rect 46020 6400 46072 6452
rect 1492 6264 1544 6316
rect 45836 6307 45888 6316
rect 45836 6273 45845 6307
rect 45845 6273 45879 6307
rect 45879 6273 45888 6307
rect 45836 6264 45888 6273
rect 9128 6128 9180 6180
rect 26056 6128 26108 6180
rect 46296 6060 46348 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 24676 5899 24728 5908
rect 24676 5865 24685 5899
rect 24685 5865 24719 5899
rect 24719 5865 24728 5899
rect 24676 5856 24728 5865
rect 25504 5899 25556 5908
rect 25504 5865 25513 5899
rect 25513 5865 25547 5899
rect 25547 5865 25556 5899
rect 25504 5856 25556 5865
rect 46296 5763 46348 5772
rect 46296 5729 46305 5763
rect 46305 5729 46339 5763
rect 46339 5729 46348 5763
rect 46296 5720 46348 5729
rect 1768 5695 1820 5704
rect 1768 5661 1777 5695
rect 1777 5661 1811 5695
rect 1811 5661 1820 5695
rect 1768 5652 1820 5661
rect 2320 5652 2372 5704
rect 20168 5652 20220 5704
rect 25228 5695 25280 5704
rect 25228 5661 25237 5695
rect 25237 5661 25271 5695
rect 25271 5661 25280 5695
rect 25228 5652 25280 5661
rect 25872 5652 25924 5704
rect 34520 5584 34572 5636
rect 46940 5584 46992 5636
rect 48136 5627 48188 5636
rect 48136 5593 48145 5627
rect 48145 5593 48179 5627
rect 48179 5593 48188 5627
rect 48136 5584 48188 5593
rect 1584 5516 1636 5568
rect 3056 5559 3108 5568
rect 3056 5525 3065 5559
rect 3065 5525 3099 5559
rect 3099 5525 3108 5559
rect 3056 5516 3108 5525
rect 39120 5516 39172 5568
rect 47032 5516 47084 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 46940 5355 46992 5364
rect 46940 5321 46949 5355
rect 46949 5321 46983 5355
rect 46983 5321 46992 5355
rect 46940 5312 46992 5321
rect 3056 5244 3108 5296
rect 47952 5287 48004 5296
rect 47952 5253 47961 5287
rect 47961 5253 47995 5287
rect 47995 5253 48004 5287
rect 47952 5244 48004 5253
rect 1768 5176 1820 5228
rect 17868 5176 17920 5228
rect 30748 5176 30800 5228
rect 46664 5176 46716 5228
rect 47216 5176 47268 5228
rect 2780 5151 2832 5160
rect 2780 5117 2789 5151
rect 2789 5117 2823 5151
rect 2823 5117 2832 5151
rect 2780 5108 2832 5117
rect 32588 5108 32640 5160
rect 46756 5108 46808 5160
rect 25228 5040 25280 5092
rect 1400 4972 1452 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 2688 4768 2740 4820
rect 17132 4768 17184 4820
rect 18512 4768 18564 4820
rect 32220 4768 32272 4820
rect 32956 4768 33008 4820
rect 46848 4768 46900 4820
rect 1400 4675 1452 4684
rect 1400 4641 1409 4675
rect 1409 4641 1443 4675
rect 1443 4641 1452 4675
rect 1400 4632 1452 4641
rect 1584 4675 1636 4684
rect 1584 4641 1593 4675
rect 1593 4641 1627 4675
rect 1627 4641 1636 4675
rect 1584 4632 1636 4641
rect 2780 4675 2832 4684
rect 2780 4641 2789 4675
rect 2789 4641 2823 4675
rect 2823 4641 2832 4675
rect 2780 4632 2832 4641
rect 45008 4564 45060 4616
rect 46940 4496 46992 4548
rect 48320 4496 48372 4548
rect 3700 4428 3752 4480
rect 8024 4428 8076 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 2044 4131 2096 4140
rect 2044 4097 2053 4131
rect 2053 4097 2087 4131
rect 2087 4097 2096 4131
rect 2044 4088 2096 4097
rect 3792 4088 3844 4140
rect 6736 4131 6788 4140
rect 6736 4097 6745 4131
rect 6745 4097 6779 4131
rect 6779 4097 6788 4131
rect 6736 4088 6788 4097
rect 7380 4088 7432 4140
rect 20076 4156 20128 4208
rect 23572 4156 23624 4208
rect 9956 4088 10008 4140
rect 10324 4088 10376 4140
rect 11336 4088 11388 4140
rect 7748 4020 7800 4072
rect 18420 4088 18472 4140
rect 20628 4088 20680 4140
rect 30748 4131 30800 4140
rect 30748 4097 30757 4131
rect 30757 4097 30791 4131
rect 30791 4097 30800 4131
rect 30748 4088 30800 4097
rect 20536 4020 20588 4072
rect 28816 4020 28868 4072
rect 28908 4020 28960 4072
rect 37924 4088 37976 4140
rect 41696 4131 41748 4140
rect 35440 4020 35492 4072
rect 37372 4020 37424 4072
rect 37464 4020 37516 4072
rect 41696 4097 41705 4131
rect 41705 4097 41739 4131
rect 41739 4097 41748 4131
rect 41696 4088 41748 4097
rect 45836 4131 45888 4140
rect 45836 4097 45845 4131
rect 45845 4097 45879 4131
rect 45879 4097 45888 4131
rect 45836 4088 45888 4097
rect 45928 4088 45980 4140
rect 46940 4131 46992 4140
rect 46940 4097 46949 4131
rect 46949 4097 46983 4131
rect 46983 4097 46992 4131
rect 46940 4088 46992 4097
rect 38752 4063 38804 4072
rect 38752 4029 38761 4063
rect 38761 4029 38795 4063
rect 38795 4029 38804 4063
rect 38752 4020 38804 4029
rect 39764 4063 39816 4072
rect 1584 3927 1636 3936
rect 1584 3893 1593 3927
rect 1593 3893 1627 3927
rect 1627 3893 1636 3927
rect 1584 3884 1636 3893
rect 1676 3884 1728 3936
rect 2872 3884 2924 3936
rect 3516 3927 3568 3936
rect 3516 3893 3525 3927
rect 3525 3893 3559 3927
rect 3559 3893 3568 3927
rect 3516 3884 3568 3893
rect 4620 3884 4672 3936
rect 4988 3927 5040 3936
rect 4988 3893 4997 3927
rect 4997 3893 5031 3927
rect 5031 3893 5040 3927
rect 4988 3884 5040 3893
rect 6552 3884 6604 3936
rect 7564 3927 7616 3936
rect 7564 3893 7573 3927
rect 7573 3893 7607 3927
rect 7607 3893 7616 3927
rect 7564 3884 7616 3893
rect 17500 3952 17552 4004
rect 32036 3952 32088 4004
rect 32128 3952 32180 4004
rect 36176 3952 36228 4004
rect 11704 3884 11756 3936
rect 12164 3884 12216 3936
rect 14188 3884 14240 3936
rect 19340 3884 19392 3936
rect 19984 3884 20036 3936
rect 29552 3927 29604 3936
rect 29552 3893 29561 3927
rect 29561 3893 29595 3927
rect 29595 3893 29604 3927
rect 29552 3884 29604 3893
rect 29736 3884 29788 3936
rect 31300 3884 31352 3936
rect 32312 3884 32364 3936
rect 36544 3884 36596 3936
rect 39764 4029 39773 4063
rect 39773 4029 39807 4063
rect 39807 4029 39816 4063
rect 39764 4020 39816 4029
rect 42432 4063 42484 4072
rect 42432 4029 42441 4063
rect 42441 4029 42475 4063
rect 42475 4029 42484 4063
rect 42432 4020 42484 4029
rect 41512 3884 41564 3936
rect 42708 4020 42760 4072
rect 46756 4020 46808 4072
rect 47584 3952 47636 4004
rect 45376 3927 45428 3936
rect 45376 3893 45385 3927
rect 45385 3893 45419 3927
rect 45419 3893 45428 3927
rect 45376 3884 45428 3893
rect 46204 3884 46256 3936
rect 48044 3927 48096 3936
rect 48044 3893 48053 3927
rect 48053 3893 48087 3927
rect 48087 3893 48096 3927
rect 48044 3884 48096 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 1952 3680 2004 3732
rect 6276 3680 6328 3732
rect 6736 3680 6788 3732
rect 10508 3680 10560 3732
rect 20352 3680 20404 3732
rect 20812 3680 20864 3732
rect 3516 3612 3568 3664
rect 3884 3612 3936 3664
rect 13084 3612 13136 3664
rect 1676 3544 1728 3596
rect 1860 3587 1912 3596
rect 1860 3553 1869 3587
rect 1869 3553 1903 3587
rect 1903 3553 1912 3587
rect 1860 3544 1912 3553
rect 4620 3544 4672 3596
rect 5172 3587 5224 3596
rect 5172 3553 5181 3587
rect 5181 3553 5215 3587
rect 5215 3553 5224 3587
rect 5172 3544 5224 3553
rect 7380 3544 7432 3596
rect 9956 3544 10008 3596
rect 11612 3544 11664 3596
rect 13360 3544 13412 3596
rect 3792 3519 3844 3528
rect 3792 3485 3801 3519
rect 3801 3485 3835 3519
rect 3835 3485 3844 3519
rect 3792 3476 3844 3485
rect 6644 3476 6696 3528
rect 11796 3519 11848 3528
rect 11796 3485 11805 3519
rect 11805 3485 11839 3519
rect 11839 3485 11848 3519
rect 11796 3476 11848 3485
rect 11980 3476 12032 3528
rect 12624 3476 12676 3528
rect 19432 3612 19484 3664
rect 27988 3612 28040 3664
rect 36176 3612 36228 3664
rect 38752 3680 38804 3732
rect 41696 3680 41748 3732
rect 47124 3680 47176 3732
rect 38844 3612 38896 3664
rect 17040 3544 17092 3596
rect 19984 3587 20036 3596
rect 19984 3553 19993 3587
rect 19993 3553 20027 3587
rect 20027 3553 20036 3587
rect 19984 3544 20036 3553
rect 20628 3587 20680 3596
rect 20628 3553 20637 3587
rect 20637 3553 20671 3587
rect 20671 3553 20680 3587
rect 20628 3544 20680 3553
rect 14280 3476 14332 3528
rect 17132 3476 17184 3528
rect 17408 3476 17460 3528
rect 18328 3476 18380 3528
rect 19892 3476 19944 3528
rect 23204 3476 23256 3528
rect 23572 3519 23624 3528
rect 23572 3485 23581 3519
rect 23581 3485 23615 3519
rect 23615 3485 23624 3519
rect 23572 3476 23624 3485
rect 27712 3544 27764 3596
rect 31300 3587 31352 3596
rect 31300 3553 31309 3587
rect 31309 3553 31343 3587
rect 31343 3553 31352 3587
rect 31300 3544 31352 3553
rect 31576 3587 31628 3596
rect 31576 3553 31585 3587
rect 31585 3553 31619 3587
rect 31619 3553 31628 3587
rect 31576 3544 31628 3553
rect 36544 3587 36596 3596
rect 36544 3553 36553 3587
rect 36553 3553 36587 3587
rect 36587 3553 36596 3587
rect 36544 3544 36596 3553
rect 36728 3544 36780 3596
rect 38108 3544 38160 3596
rect 39028 3544 39080 3596
rect 41512 3587 41564 3596
rect 25964 3519 26016 3528
rect 25964 3485 25973 3519
rect 25973 3485 26007 3519
rect 26007 3485 26016 3519
rect 25964 3476 26016 3485
rect 27436 3476 27488 3528
rect 27988 3476 28040 3528
rect 28816 3476 28868 3528
rect 36360 3519 36412 3528
rect 36360 3485 36369 3519
rect 36369 3485 36403 3519
rect 36403 3485 36412 3519
rect 36360 3476 36412 3485
rect 38844 3476 38896 3528
rect 39856 3519 39908 3528
rect 39856 3485 39865 3519
rect 39865 3485 39899 3519
rect 39899 3485 39908 3519
rect 39856 3476 39908 3485
rect 41512 3553 41521 3587
rect 41521 3553 41555 3587
rect 41555 3553 41564 3587
rect 41512 3544 41564 3553
rect 41880 3544 41932 3596
rect 45652 3612 45704 3664
rect 45376 3544 45428 3596
rect 46204 3587 46256 3596
rect 46204 3553 46213 3587
rect 46213 3553 46247 3587
rect 46247 3553 46256 3587
rect 46204 3544 46256 3553
rect 46388 3544 46440 3596
rect 2044 3408 2096 3460
rect 3516 3340 3568 3392
rect 4988 3408 5040 3460
rect 7104 3408 7156 3460
rect 11888 3340 11940 3392
rect 14464 3340 14516 3392
rect 17500 3340 17552 3392
rect 20352 3408 20404 3460
rect 26240 3408 26292 3460
rect 23020 3340 23072 3392
rect 23388 3340 23440 3392
rect 26424 3340 26476 3392
rect 27436 3340 27488 3392
rect 29644 3340 29696 3392
rect 29920 3340 29972 3392
rect 40132 3340 40184 3392
rect 45928 3476 45980 3528
rect 44180 3340 44232 3392
rect 45192 3340 45244 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 1952 3179 2004 3188
rect 1952 3145 1961 3179
rect 1961 3145 1995 3179
rect 1995 3145 2004 3179
rect 1952 3136 2004 3145
rect 2596 3136 2648 3188
rect 20352 3179 20404 3188
rect 2780 3068 2832 3120
rect 3516 3111 3568 3120
rect 3516 3077 3525 3111
rect 3525 3077 3559 3111
rect 3559 3077 3568 3111
rect 3516 3068 3568 3077
rect 7564 3068 7616 3120
rect 12164 3111 12216 3120
rect 12164 3077 12173 3111
rect 12173 3077 12207 3111
rect 12207 3077 12216 3111
rect 12164 3068 12216 3077
rect 12256 3068 12308 3120
rect 14188 3068 14240 3120
rect 14464 3111 14516 3120
rect 14464 3077 14473 3111
rect 14473 3077 14507 3111
rect 14507 3077 14516 3111
rect 14464 3068 14516 3077
rect 17500 3111 17552 3120
rect 17500 3077 17509 3111
rect 17509 3077 17543 3111
rect 17543 3077 17552 3111
rect 17500 3068 17552 3077
rect 20352 3145 20361 3179
rect 20361 3145 20395 3179
rect 20395 3145 20404 3179
rect 20352 3136 20404 3145
rect 20444 3136 20496 3188
rect 23388 3111 23440 3120
rect 1952 3000 2004 3052
rect 6644 3043 6696 3052
rect 6644 3009 6653 3043
rect 6653 3009 6687 3043
rect 6687 3009 6696 3043
rect 6644 3000 6696 3009
rect 8392 3000 8444 3052
rect 11980 3043 12032 3052
rect 3332 2975 3384 2984
rect 3332 2941 3341 2975
rect 3341 2941 3375 2975
rect 3375 2941 3384 2975
rect 3332 2932 3384 2941
rect 664 2864 716 2916
rect 2688 2839 2740 2848
rect 2688 2805 2697 2839
rect 2697 2805 2731 2839
rect 2731 2805 2740 2839
rect 2688 2796 2740 2805
rect 3240 2864 3292 2916
rect 6460 2932 6512 2984
rect 11980 3009 11989 3043
rect 11989 3009 12023 3043
rect 12023 3009 12032 3043
rect 11980 3000 12032 3009
rect 14280 3043 14332 3052
rect 14280 3009 14289 3043
rect 14289 3009 14323 3043
rect 14323 3009 14332 3043
rect 14280 3000 14332 3009
rect 17040 3000 17092 3052
rect 20536 3000 20588 3052
rect 10968 2932 11020 2984
rect 12256 2932 12308 2984
rect 12716 2932 12768 2984
rect 12900 2975 12952 2984
rect 12900 2941 12909 2975
rect 12909 2941 12943 2975
rect 12943 2941 12952 2975
rect 12900 2932 12952 2941
rect 15476 2975 15528 2984
rect 15476 2941 15485 2975
rect 15485 2941 15519 2975
rect 15519 2941 15528 2975
rect 15476 2932 15528 2941
rect 18052 2975 18104 2984
rect 18052 2941 18061 2975
rect 18061 2941 18095 2975
rect 18095 2941 18104 2975
rect 18052 2932 18104 2941
rect 12440 2864 12492 2916
rect 23388 3077 23397 3111
rect 23397 3077 23431 3111
rect 23431 3077 23440 3111
rect 23388 3068 23440 3077
rect 23204 3043 23256 3052
rect 23204 3009 23213 3043
rect 23213 3009 23247 3043
rect 23247 3009 23256 3043
rect 23204 3000 23256 3009
rect 25964 3000 26016 3052
rect 23848 2975 23900 2984
rect 23848 2941 23857 2975
rect 23857 2941 23891 2975
rect 23891 2941 23900 2975
rect 23848 2932 23900 2941
rect 28172 2932 28224 2984
rect 28724 3136 28776 3188
rect 48044 3136 48096 3188
rect 29920 3111 29972 3120
rect 29920 3077 29929 3111
rect 29929 3077 29963 3111
rect 29963 3077 29972 3111
rect 29920 3068 29972 3077
rect 32312 3111 32364 3120
rect 32312 3077 32321 3111
rect 32321 3077 32355 3111
rect 32355 3077 32364 3111
rect 32312 3068 32364 3077
rect 40132 3111 40184 3120
rect 40132 3077 40141 3111
rect 40141 3077 40175 3111
rect 40175 3077 40184 3111
rect 40132 3068 40184 3077
rect 44180 3111 44232 3120
rect 44180 3077 44189 3111
rect 44189 3077 44223 3111
rect 44223 3077 44232 3111
rect 44180 3068 44232 3077
rect 44364 3068 44416 3120
rect 46664 3068 46716 3120
rect 29736 3043 29788 3052
rect 29736 3009 29745 3043
rect 29745 3009 29779 3043
rect 29779 3009 29788 3043
rect 29736 3000 29788 3009
rect 32128 3043 32180 3052
rect 32128 3009 32137 3043
rect 32137 3009 32171 3043
rect 32171 3009 32180 3043
rect 32128 3000 32180 3009
rect 36360 3000 36412 3052
rect 42432 3000 42484 3052
rect 45744 3000 45796 3052
rect 46572 3043 46624 3052
rect 46572 3009 46581 3043
rect 46581 3009 46615 3043
rect 46615 3009 46624 3043
rect 46572 3000 46624 3009
rect 49608 3000 49660 3052
rect 30288 2975 30340 2984
rect 30288 2941 30297 2975
rect 30297 2941 30331 2975
rect 30331 2941 30340 2975
rect 30288 2932 30340 2941
rect 33508 2975 33560 2984
rect 33508 2941 33517 2975
rect 33517 2941 33551 2975
rect 33551 2941 33560 2975
rect 33508 2932 33560 2941
rect 39948 2975 40000 2984
rect 39948 2941 39957 2975
rect 39957 2941 39991 2975
rect 39991 2941 40000 2975
rect 39948 2932 40000 2941
rect 41144 2975 41196 2984
rect 41144 2941 41153 2975
rect 41153 2941 41187 2975
rect 41187 2941 41196 2975
rect 41144 2932 41196 2941
rect 44272 2932 44324 2984
rect 44456 2975 44508 2984
rect 44456 2941 44465 2975
rect 44465 2941 44499 2975
rect 44499 2941 44508 2975
rect 44456 2932 44508 2941
rect 5816 2839 5868 2848
rect 5816 2805 5825 2839
rect 5825 2805 5859 2839
rect 5859 2805 5868 2839
rect 5816 2796 5868 2805
rect 9128 2839 9180 2848
rect 9128 2805 9137 2839
rect 9137 2805 9171 2839
rect 9171 2805 9180 2839
rect 9128 2796 9180 2805
rect 9956 2796 10008 2848
rect 12624 2796 12676 2848
rect 12716 2796 12768 2848
rect 20444 2796 20496 2848
rect 28908 2796 28960 2848
rect 29644 2796 29696 2848
rect 29828 2796 29880 2848
rect 32036 2864 32088 2916
rect 33048 2796 33100 2848
rect 37924 2796 37976 2848
rect 44364 2796 44416 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 3332 2592 3384 2644
rect 18236 2592 18288 2644
rect 21364 2592 21416 2644
rect 46848 2592 46900 2644
rect 1308 2524 1360 2576
rect 1584 2456 1636 2508
rect 6184 2524 6236 2576
rect 17776 2567 17828 2576
rect 5816 2456 5868 2508
rect 6552 2499 6604 2508
rect 6552 2465 6561 2499
rect 6561 2465 6595 2499
rect 6595 2465 6604 2499
rect 6552 2456 6604 2465
rect 11796 2456 11848 2508
rect 12256 2499 12308 2508
rect 12256 2465 12265 2499
rect 12265 2465 12299 2499
rect 12299 2465 12308 2499
rect 12256 2456 12308 2465
rect 14740 2499 14792 2508
rect 14740 2465 14749 2499
rect 14749 2465 14783 2499
rect 14783 2465 14792 2499
rect 14740 2456 14792 2465
rect 17776 2533 17785 2567
rect 17785 2533 17819 2567
rect 17819 2533 17828 2567
rect 17776 2524 17828 2533
rect 23664 2524 23716 2576
rect 25872 2567 25924 2576
rect 25872 2533 25881 2567
rect 25881 2533 25915 2567
rect 25915 2533 25924 2567
rect 25872 2524 25924 2533
rect 22744 2456 22796 2508
rect 23756 2456 23808 2508
rect 4528 2388 4580 2440
rect 7748 2388 7800 2440
rect 19984 2388 20036 2440
rect 22560 2388 22612 2440
rect 23204 2388 23256 2440
rect 24492 2388 24544 2440
rect 24676 2388 24728 2440
rect 25136 2388 25188 2440
rect 2872 2320 2924 2372
rect 3424 2320 3476 2372
rect 8668 2320 8720 2372
rect 9680 2320 9732 2372
rect 11704 2363 11756 2372
rect 11704 2329 11713 2363
rect 11713 2329 11747 2363
rect 11747 2329 11756 2363
rect 11704 2320 11756 2329
rect 14188 2320 14240 2372
rect 17408 2320 17460 2372
rect 27068 2431 27120 2440
rect 27068 2397 27077 2431
rect 27077 2397 27111 2431
rect 27111 2397 27120 2431
rect 27068 2388 27120 2397
rect 27344 2456 27396 2508
rect 29552 2499 29604 2508
rect 29552 2465 29561 2499
rect 29561 2465 29595 2499
rect 29595 2465 29604 2499
rect 29552 2456 29604 2465
rect 29736 2499 29788 2508
rect 29736 2465 29745 2499
rect 29745 2465 29779 2499
rect 29779 2465 29788 2499
rect 29736 2456 29788 2465
rect 30932 2499 30984 2508
rect 30932 2465 30941 2499
rect 30941 2465 30975 2499
rect 30975 2465 30984 2499
rect 30932 2456 30984 2465
rect 33876 2456 33928 2508
rect 35900 2456 35952 2508
rect 39948 2499 40000 2508
rect 39948 2465 39957 2499
rect 39957 2465 39991 2499
rect 39991 2465 40000 2499
rect 39948 2456 40000 2465
rect 44272 2499 44324 2508
rect 44272 2465 44281 2499
rect 44281 2465 44315 2499
rect 44315 2465 44324 2499
rect 44272 2456 44324 2465
rect 45008 2499 45060 2508
rect 45008 2465 45017 2499
rect 45017 2465 45051 2499
rect 45051 2465 45060 2499
rect 45008 2456 45060 2465
rect 45192 2499 45244 2508
rect 45192 2465 45201 2499
rect 45201 2465 45235 2499
rect 45235 2465 45244 2499
rect 45192 2456 45244 2465
rect 45376 2456 45428 2508
rect 4804 2295 4856 2304
rect 4804 2261 4813 2295
rect 4813 2261 4847 2295
rect 4847 2261 4856 2295
rect 4804 2252 4856 2261
rect 26516 2320 26568 2372
rect 27160 2320 27212 2372
rect 22836 2295 22888 2304
rect 22836 2261 22845 2295
rect 22845 2261 22879 2295
rect 22879 2261 22888 2295
rect 22836 2252 22888 2261
rect 24032 2252 24084 2304
rect 24676 2252 24728 2304
rect 25320 2252 25372 2304
rect 27712 2388 27764 2440
rect 32864 2388 32916 2440
rect 34796 2388 34848 2440
rect 36084 2388 36136 2440
rect 38660 2388 38712 2440
rect 27528 2320 27580 2372
rect 31392 2252 31444 2304
rect 34152 2320 34204 2372
rect 43168 2320 43220 2372
rect 47768 2363 47820 2372
rect 47768 2329 47777 2363
rect 47777 2329 47811 2363
rect 47811 2329 47820 2363
rect 47768 2320 47820 2329
rect 34060 2295 34112 2304
rect 34060 2261 34069 2295
rect 34069 2261 34103 2295
rect 34103 2261 34112 2295
rect 34060 2252 34112 2261
rect 34520 2252 34572 2304
rect 43444 2295 43496 2304
rect 43444 2261 43453 2295
rect 43453 2261 43487 2295
rect 43487 2261 43496 2295
rect 43444 2252 43496 2261
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 23940 2048 23992 2100
rect 34060 2048 34112 2100
rect 22836 1980 22888 2032
rect 30656 1980 30708 2032
rect 24308 1912 24360 1964
rect 43444 1912 43496 1964
<< metal2 >>
rect 18 51200 74 52000
rect 662 51200 718 52000
rect 1306 51200 1362 52000
rect 1950 51200 2006 52000
rect 2594 51200 2650 52000
rect 3238 51354 3294 52000
rect 3790 51776 3846 51785
rect 3790 51711 3846 51720
rect 3238 51326 3648 51354
rect 3238 51200 3294 51326
rect 32 48278 60 51200
rect 676 49230 704 51200
rect 664 49224 716 49230
rect 664 49166 716 49172
rect 20 48272 72 48278
rect 20 48214 72 48220
rect 1320 47802 1348 51200
rect 1768 49088 1820 49094
rect 1768 49030 1820 49036
rect 1676 48748 1728 48754
rect 1676 48690 1728 48696
rect 1308 47796 1360 47802
rect 1308 47738 1360 47744
rect 1398 47696 1454 47705
rect 1398 47631 1454 47640
rect 1412 47054 1440 47631
rect 1400 47048 1452 47054
rect 1400 46990 1452 46996
rect 1400 45960 1452 45966
rect 1400 45902 1452 45908
rect 1412 45665 1440 45902
rect 1398 45656 1454 45665
rect 1398 45591 1454 45600
rect 1400 45280 1452 45286
rect 1400 45222 1452 45228
rect 1412 44946 1440 45222
rect 1400 44940 1452 44946
rect 1400 44882 1452 44888
rect 1400 42016 1452 42022
rect 1400 41958 1452 41964
rect 1412 41682 1440 41958
rect 1400 41676 1452 41682
rect 1400 41618 1452 41624
rect 1584 41540 1636 41546
rect 1584 41482 1636 41488
rect 1596 41274 1624 41482
rect 1584 41268 1636 41274
rect 1584 41210 1636 41216
rect 1492 41064 1544 41070
rect 1492 41006 1544 41012
rect 1400 40520 1452 40526
rect 1400 40462 1452 40468
rect 1412 40225 1440 40462
rect 1398 40216 1454 40225
rect 1398 40151 1454 40160
rect 1504 37942 1532 41006
rect 1584 40384 1636 40390
rect 1584 40326 1636 40332
rect 1492 37936 1544 37942
rect 1492 37878 1544 37884
rect 1400 37324 1452 37330
rect 1400 37266 1452 37272
rect 1412 36825 1440 37266
rect 1398 36816 1454 36825
rect 1398 36751 1454 36760
rect 1400 34400 1452 34406
rect 1400 34342 1452 34348
rect 1412 34066 1440 34342
rect 1400 34060 1452 34066
rect 1400 34002 1452 34008
rect 1400 27464 1452 27470
rect 1400 27406 1452 27412
rect 1412 27062 1440 27406
rect 1400 27056 1452 27062
rect 1400 26998 1452 27004
rect 1400 26784 1452 26790
rect 1400 26726 1452 26732
rect 1412 26450 1440 26726
rect 1400 26444 1452 26450
rect 1400 26386 1452 26392
rect 1400 24200 1452 24206
rect 1400 24142 1452 24148
rect 1412 23905 1440 24142
rect 1398 23896 1454 23905
rect 1398 23831 1454 23840
rect 1400 22636 1452 22642
rect 1400 22578 1452 22584
rect 1412 22545 1440 22578
rect 1398 22536 1454 22545
rect 1398 22471 1454 22480
rect 1400 19168 1452 19174
rect 1400 19110 1452 19116
rect 1412 18834 1440 19110
rect 1400 18828 1452 18834
rect 1400 18770 1452 18776
rect 20 15972 72 15978
rect 20 15914 72 15920
rect 32 800 60 15914
rect 1400 12776 1452 12782
rect 1400 12718 1452 12724
rect 1412 12345 1440 12718
rect 1398 12336 1454 12345
rect 1398 12271 1454 12280
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1412 7585 1440 7822
rect 1398 7576 1454 7585
rect 1398 7511 1454 7520
rect 1504 6322 1532 37878
rect 1596 31482 1624 40326
rect 1688 37806 1716 48690
rect 1676 37800 1728 37806
rect 1676 37742 1728 37748
rect 1676 37256 1728 37262
rect 1676 37198 1728 37204
rect 1688 36854 1716 37198
rect 1676 36848 1728 36854
rect 1676 36790 1728 36796
rect 1780 36802 1808 49030
rect 1964 48822 1992 51200
rect 2870 50416 2926 50425
rect 2870 50351 2926 50360
rect 2780 49156 2832 49162
rect 2780 49098 2832 49104
rect 1952 48816 2004 48822
rect 1952 48758 2004 48764
rect 2228 48680 2280 48686
rect 2228 48622 2280 48628
rect 2136 48544 2188 48550
rect 2136 48486 2188 48492
rect 1952 48000 2004 48006
rect 1952 47942 2004 47948
rect 1964 47666 1992 47942
rect 2148 47734 2176 48486
rect 2136 47728 2188 47734
rect 2136 47670 2188 47676
rect 1952 47660 2004 47666
rect 1952 47602 2004 47608
rect 2240 47258 2268 48622
rect 2792 48278 2820 49098
rect 2884 48686 2912 50351
rect 3620 49230 3648 51326
rect 3608 49224 3660 49230
rect 3608 49166 3660 49172
rect 2964 49156 3016 49162
rect 2964 49098 3016 49104
rect 2872 48680 2924 48686
rect 2872 48622 2924 48628
rect 2780 48272 2832 48278
rect 2780 48214 2832 48220
rect 2228 47252 2280 47258
rect 2228 47194 2280 47200
rect 2412 47048 2464 47054
rect 2412 46990 2464 46996
rect 2780 47048 2832 47054
rect 2780 46990 2832 46996
rect 2044 45280 2096 45286
rect 2044 45222 2096 45228
rect 2056 44470 2084 45222
rect 2044 44464 2096 44470
rect 2044 44406 2096 44412
rect 1858 44296 1914 44305
rect 1858 44231 1914 44240
rect 1872 43790 1900 44231
rect 1860 43784 1912 43790
rect 1860 43726 1912 43732
rect 2136 43784 2188 43790
rect 2136 43726 2188 43732
rect 1952 43648 2004 43654
rect 1858 43616 1914 43625
rect 1952 43590 2004 43596
rect 1858 43551 1914 43560
rect 1872 43382 1900 43551
rect 1860 43376 1912 43382
rect 1860 43318 1912 43324
rect 1860 41676 1912 41682
rect 1860 41618 1912 41624
rect 1872 41585 1900 41618
rect 1858 41576 1914 41585
rect 1858 41511 1914 41520
rect 1860 41132 1912 41138
rect 1860 41074 1912 41080
rect 1872 40905 1900 41074
rect 1858 40896 1914 40905
rect 1858 40831 1914 40840
rect 1860 37868 1912 37874
rect 1860 37810 1912 37816
rect 1872 37505 1900 37810
rect 1858 37496 1914 37505
rect 1858 37431 1914 37440
rect 1780 36774 1900 36802
rect 1676 36712 1728 36718
rect 1676 36654 1728 36660
rect 1584 31476 1636 31482
rect 1584 31418 1636 31424
rect 1584 26308 1636 26314
rect 1584 26250 1636 26256
rect 1596 26042 1624 26250
rect 1584 26036 1636 26042
rect 1584 25978 1636 25984
rect 1582 25936 1638 25945
rect 1582 25871 1584 25880
rect 1636 25871 1638 25880
rect 1584 25842 1636 25848
rect 1584 24608 1636 24614
rect 1584 24550 1636 24556
rect 1596 24410 1624 24550
rect 1584 24404 1636 24410
rect 1584 24346 1636 24352
rect 1584 23248 1636 23254
rect 1584 23190 1636 23196
rect 1596 22778 1624 23190
rect 1584 22772 1636 22778
rect 1584 22714 1636 22720
rect 1688 17338 1716 36654
rect 1872 35894 1900 36774
rect 1964 36718 1992 43590
rect 2044 39432 2096 39438
rect 2044 39374 2096 39380
rect 2056 38962 2084 39374
rect 2044 38956 2096 38962
rect 2044 38898 2096 38904
rect 1952 36712 2004 36718
rect 1952 36654 2004 36660
rect 2148 36530 2176 43726
rect 2228 43104 2280 43110
rect 2228 43046 2280 43052
rect 1780 35866 1900 35894
rect 1964 36502 2176 36530
rect 1780 24410 1808 35866
rect 1964 35578 1992 36502
rect 2136 36236 2188 36242
rect 2136 36178 2188 36184
rect 2148 35894 2176 36178
rect 2056 35866 2176 35894
rect 2056 35698 2084 35866
rect 2044 35692 2096 35698
rect 2044 35634 2096 35640
rect 1964 35550 2084 35578
rect 1952 35488 2004 35494
rect 1952 35430 2004 35436
rect 1964 35290 1992 35430
rect 1952 35284 2004 35290
rect 1952 35226 2004 35232
rect 1860 35012 1912 35018
rect 1860 34954 1912 34960
rect 1872 34785 1900 34954
rect 1858 34776 1914 34785
rect 1858 34711 1914 34720
rect 2056 34610 2084 35550
rect 2044 34604 2096 34610
rect 2044 34546 2096 34552
rect 1860 34536 1912 34542
rect 1860 34478 1912 34484
rect 1872 33522 1900 34478
rect 2136 34400 2188 34406
rect 2136 34342 2188 34348
rect 2148 34066 2176 34342
rect 2136 34060 2188 34066
rect 2136 34002 2188 34008
rect 1860 33516 1912 33522
rect 1860 33458 1912 33464
rect 2044 32904 2096 32910
rect 2044 32846 2096 32852
rect 2056 32434 2084 32846
rect 2044 32428 2096 32434
rect 2044 32370 2096 32376
rect 1860 31816 1912 31822
rect 1860 31758 1912 31764
rect 2044 31816 2096 31822
rect 2044 31758 2096 31764
rect 1872 31385 1900 31758
rect 1858 31376 1914 31385
rect 1858 31311 1914 31320
rect 1952 31272 2004 31278
rect 1952 31214 2004 31220
rect 1964 30938 1992 31214
rect 1952 30932 2004 30938
rect 1952 30874 2004 30880
rect 1952 30184 2004 30190
rect 1952 30126 2004 30132
rect 1964 29850 1992 30126
rect 1952 29844 2004 29850
rect 1952 29786 2004 29792
rect 2056 29050 2084 31758
rect 1964 29022 2084 29050
rect 1860 27532 1912 27538
rect 1860 27474 1912 27480
rect 1872 27305 1900 27474
rect 1858 27296 1914 27305
rect 1858 27231 1914 27240
rect 1964 26246 1992 29022
rect 2044 28960 2096 28966
rect 2044 28902 2096 28908
rect 2056 28626 2084 28902
rect 2044 28620 2096 28626
rect 2044 28562 2096 28568
rect 2136 28484 2188 28490
rect 2136 28426 2188 28432
rect 2148 28218 2176 28426
rect 2136 28212 2188 28218
rect 2136 28154 2188 28160
rect 2044 28076 2096 28082
rect 2044 28018 2096 28024
rect 2056 27674 2084 28018
rect 2044 27668 2096 27674
rect 2044 27610 2096 27616
rect 2136 27396 2188 27402
rect 2136 27338 2188 27344
rect 2148 27130 2176 27338
rect 2136 27124 2188 27130
rect 2136 27066 2188 27072
rect 1952 26240 2004 26246
rect 1952 26182 2004 26188
rect 2240 24750 2268 43046
rect 2320 40996 2372 41002
rect 2320 40938 2372 40944
rect 2332 26858 2360 40938
rect 2320 26852 2372 26858
rect 2320 26794 2372 26800
rect 2228 24744 2280 24750
rect 2228 24686 2280 24692
rect 1768 24404 1820 24410
rect 1768 24346 1820 24352
rect 2044 23520 2096 23526
rect 2044 23462 2096 23468
rect 2056 23186 2084 23462
rect 2044 23180 2096 23186
rect 2044 23122 2096 23128
rect 2320 23044 2372 23050
rect 2320 22986 2372 22992
rect 2332 22778 2360 22986
rect 2320 22772 2372 22778
rect 2320 22714 2372 22720
rect 2136 22636 2188 22642
rect 2136 22578 2188 22584
rect 2148 22166 2176 22578
rect 2136 22160 2188 22166
rect 2136 22102 2188 22108
rect 1952 18216 2004 18222
rect 1952 18158 2004 18164
rect 1964 17882 1992 18158
rect 1952 17876 2004 17882
rect 1952 17818 2004 17824
rect 1768 17672 1820 17678
rect 1768 17614 1820 17620
rect 2044 17672 2096 17678
rect 2044 17614 2096 17620
rect 1676 17332 1728 17338
rect 1676 17274 1728 17280
rect 1780 17202 1808 17614
rect 1952 17536 2004 17542
rect 1952 17478 2004 17484
rect 1964 17270 1992 17478
rect 1952 17264 2004 17270
rect 1952 17206 2004 17212
rect 1768 17196 1820 17202
rect 1768 17138 1820 17144
rect 1858 17096 1914 17105
rect 1858 17031 1914 17040
rect 1872 16590 1900 17031
rect 1860 16584 1912 16590
rect 1860 16526 1912 16532
rect 2056 13938 2084 17614
rect 2044 13932 2096 13938
rect 2044 13874 2096 13880
rect 1584 13728 1636 13734
rect 1584 13670 1636 13676
rect 1596 13394 1624 13670
rect 1584 13388 1636 13394
rect 1584 13330 1636 13336
rect 1860 11076 1912 11082
rect 1860 11018 1912 11024
rect 1872 10985 1900 11018
rect 1858 10976 1914 10985
rect 1858 10911 1914 10920
rect 1584 10600 1636 10606
rect 1584 10542 1636 10548
rect 1596 10266 1624 10542
rect 1584 10260 1636 10266
rect 1584 10202 1636 10208
rect 1952 10056 2004 10062
rect 1952 9998 2004 10004
rect 1964 9586 1992 9998
rect 1952 9580 2004 9586
rect 1952 9522 2004 9528
rect 2056 9466 2084 13874
rect 1964 9438 2084 9466
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 1872 8265 1900 8434
rect 1858 8256 1914 8265
rect 1858 8191 1914 8200
rect 1492 6316 1544 6322
rect 1492 6258 1544 6264
rect 1768 5704 1820 5710
rect 1768 5646 1820 5652
rect 1584 5568 1636 5574
rect 1584 5510 1636 5516
rect 1400 5024 1452 5030
rect 1400 4966 1452 4972
rect 1412 4690 1440 4966
rect 1596 4690 1624 5510
rect 1780 5234 1808 5646
rect 1768 5228 1820 5234
rect 1768 5170 1820 5176
rect 1400 4684 1452 4690
rect 1400 4626 1452 4632
rect 1584 4684 1636 4690
rect 1584 4626 1636 4632
rect 1964 4570 1992 9438
rect 2148 8022 2176 22102
rect 2320 19508 2372 19514
rect 2320 19450 2372 19456
rect 2228 19168 2280 19174
rect 2228 19110 2280 19116
rect 2240 18834 2268 19110
rect 2228 18828 2280 18834
rect 2228 18770 2280 18776
rect 2136 8016 2188 8022
rect 2136 7958 2188 7964
rect 2044 7200 2096 7206
rect 2044 7142 2096 7148
rect 2056 6866 2084 7142
rect 2044 6860 2096 6866
rect 2044 6802 2096 6808
rect 2228 6724 2280 6730
rect 2228 6666 2280 6672
rect 2240 6458 2268 6666
rect 2228 6452 2280 6458
rect 2228 6394 2280 6400
rect 2332 5710 2360 19450
rect 2424 15638 2452 46990
rect 2792 46646 2820 46990
rect 2780 46640 2832 46646
rect 2780 46582 2832 46588
rect 2504 46504 2556 46510
rect 2504 46446 2556 46452
rect 2516 46170 2544 46446
rect 2778 46336 2834 46345
rect 2778 46271 2834 46280
rect 2504 46164 2556 46170
rect 2504 46106 2556 46112
rect 2504 45960 2556 45966
rect 2504 45902 2556 45908
rect 2516 45626 2544 45902
rect 2504 45620 2556 45626
rect 2504 45562 2556 45568
rect 2792 44946 2820 46271
rect 2870 44976 2926 44985
rect 2780 44940 2832 44946
rect 2870 44911 2926 44920
rect 2780 44882 2832 44888
rect 2780 44804 2832 44810
rect 2780 44746 2832 44752
rect 2792 43994 2820 44746
rect 2884 44334 2912 44911
rect 2872 44328 2924 44334
rect 2872 44270 2924 44276
rect 2780 43988 2832 43994
rect 2780 43930 2832 43936
rect 2976 39030 3004 49098
rect 3054 49056 3110 49065
rect 3054 48991 3110 49000
rect 3068 47598 3096 48991
rect 3422 48376 3478 48385
rect 3422 48311 3424 48320
rect 3476 48311 3478 48320
rect 3424 48282 3476 48288
rect 3608 48136 3660 48142
rect 3608 48078 3660 48084
rect 3148 48068 3200 48074
rect 3148 48010 3200 48016
rect 3240 48068 3292 48074
rect 3240 48010 3292 48016
rect 3056 47592 3108 47598
rect 3056 47534 3108 47540
rect 3160 47258 3188 48010
rect 3252 47802 3280 48010
rect 3240 47796 3292 47802
rect 3240 47738 3292 47744
rect 3148 47252 3200 47258
rect 3148 47194 3200 47200
rect 3240 45960 3292 45966
rect 3240 45902 3292 45908
rect 3252 45558 3280 45902
rect 3240 45552 3292 45558
rect 3240 45494 3292 45500
rect 3054 39536 3110 39545
rect 3054 39471 3110 39480
rect 2964 39024 3016 39030
rect 2964 38966 3016 38972
rect 3068 38894 3096 39471
rect 2964 38888 3016 38894
rect 2964 38830 3016 38836
rect 3056 38888 3108 38894
rect 3056 38830 3108 38836
rect 2976 38554 3004 38830
rect 2964 38548 3016 38554
rect 2964 38490 3016 38496
rect 3620 37126 3648 48078
rect 3804 46646 3832 51711
rect 3882 51200 3938 52000
rect 4526 51354 4582 52000
rect 4526 51326 4936 51354
rect 4526 51200 4582 51326
rect 4066 51096 4122 51105
rect 4066 51031 4122 51040
rect 4080 48210 4108 51031
rect 4214 49532 4522 49552
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49456 4522 49476
rect 4908 49230 4936 51326
rect 5170 51200 5226 52000
rect 5814 51200 5870 52000
rect 6458 51200 6514 52000
rect 7102 51200 7158 52000
rect 7746 51200 7802 52000
rect 8390 51200 8446 52000
rect 9034 51200 9090 52000
rect 9678 51200 9734 52000
rect 10322 51354 10378 52000
rect 10322 51326 10732 51354
rect 10322 51200 10378 51326
rect 4896 49224 4948 49230
rect 4896 49166 4948 49172
rect 4712 49156 4764 49162
rect 4712 49098 4764 49104
rect 4620 48544 4672 48550
rect 4620 48486 4672 48492
rect 4214 48444 4522 48464
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48368 4522 48388
rect 4068 48204 4120 48210
rect 4068 48146 4120 48152
rect 4436 48136 4488 48142
rect 4436 48078 4488 48084
rect 4448 47666 4476 48078
rect 4436 47660 4488 47666
rect 4436 47602 4488 47608
rect 4214 47356 4522 47376
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47280 4522 47300
rect 4066 47016 4122 47025
rect 4066 46951 4122 46960
rect 3792 46640 3844 46646
rect 3792 46582 3844 46588
rect 3976 45960 4028 45966
rect 3976 45902 4028 45908
rect 3884 45416 3936 45422
rect 3884 45358 3936 45364
rect 3896 45082 3924 45358
rect 3884 45076 3936 45082
rect 3884 45018 3936 45024
rect 3792 44872 3844 44878
rect 3792 44814 3844 44820
rect 3608 37120 3660 37126
rect 3608 37062 3660 37068
rect 2504 36576 2556 36582
rect 2504 36518 2556 36524
rect 2516 36242 2544 36518
rect 2504 36236 2556 36242
rect 2504 36178 2556 36184
rect 3804 36174 3832 44814
rect 3988 44538 4016 45902
rect 4080 45422 4108 46951
rect 4214 46268 4522 46288
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46192 4522 46212
rect 4068 45416 4120 45422
rect 4068 45358 4120 45364
rect 4214 45180 4522 45200
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45104 4522 45124
rect 3976 44532 4028 44538
rect 3976 44474 4028 44480
rect 4214 44092 4522 44112
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44016 4522 44036
rect 4214 43004 4522 43024
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42928 4522 42948
rect 4214 41916 4522 41936
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41840 4522 41860
rect 4214 40828 4522 40848
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40752 4522 40772
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 4066 38176 4122 38185
rect 4066 38111 4122 38120
rect 4080 37398 4108 38111
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4068 37392 4120 37398
rect 4068 37334 4120 37340
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 3700 36168 3752 36174
rect 2778 36136 2834 36145
rect 3700 36110 3752 36116
rect 3792 36168 3844 36174
rect 3792 36110 3844 36116
rect 2778 36071 2834 36080
rect 2792 35630 2820 36071
rect 3056 36032 3108 36038
rect 3056 35974 3108 35980
rect 3068 35766 3096 35974
rect 3712 35766 3740 36110
rect 3056 35760 3108 35766
rect 3056 35702 3108 35708
rect 3700 35760 3752 35766
rect 3700 35702 3752 35708
rect 2780 35624 2832 35630
rect 2780 35566 2832 35572
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 2504 34604 2556 34610
rect 2504 34546 2556 34552
rect 2516 26926 2544 34546
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 2778 34096 2834 34105
rect 2778 34031 2780 34040
rect 2832 34031 2834 34040
rect 2780 34002 2832 34008
rect 2780 33448 2832 33454
rect 2778 33416 2780 33425
rect 2832 33416 2834 33425
rect 2778 33351 2834 33360
rect 2780 33312 2832 33318
rect 2780 33254 2832 33260
rect 2792 33114 2820 33254
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 2780 33108 2832 33114
rect 2780 33050 2832 33056
rect 2688 32904 2740 32910
rect 2688 32846 2740 32852
rect 2596 27668 2648 27674
rect 2596 27610 2648 27616
rect 2504 26920 2556 26926
rect 2504 26862 2556 26868
rect 2504 25900 2556 25906
rect 2504 25842 2556 25848
rect 2412 15632 2464 15638
rect 2412 15574 2464 15580
rect 2516 11150 2544 25842
rect 2608 17678 2636 27610
rect 2596 17672 2648 17678
rect 2596 17614 2648 17620
rect 2700 16726 2728 32846
rect 2870 32736 2926 32745
rect 2870 32671 2926 32680
rect 2884 32366 2912 32671
rect 2780 32360 2832 32366
rect 2780 32302 2832 32308
rect 2872 32360 2924 32366
rect 2872 32302 2924 32308
rect 2792 32026 2820 32302
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 3054 32056 3110 32065
rect 2780 32020 2832 32026
rect 4214 32048 4522 32068
rect 3054 31991 3110 32000
rect 2780 31962 2832 31968
rect 3068 31278 3096 31991
rect 2872 31272 2924 31278
rect 2872 31214 2924 31220
rect 3056 31272 3108 31278
rect 3056 31214 3108 31220
rect 2884 30938 2912 31214
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 2872 30932 2924 30938
rect 2872 30874 2924 30880
rect 2780 30184 2832 30190
rect 2780 30126 2832 30132
rect 2872 30184 2924 30190
rect 2872 30126 2924 30132
rect 2792 29850 2820 30126
rect 2884 30025 2912 30126
rect 2870 30016 2926 30025
rect 2870 29951 2926 29960
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 2780 29844 2832 29850
rect 2780 29786 2832 29792
rect 2872 29640 2924 29646
rect 2872 29582 2924 29588
rect 2778 28656 2834 28665
rect 2778 28591 2780 28600
rect 2832 28591 2834 28600
rect 2780 28562 2832 28568
rect 2778 26616 2834 26625
rect 2778 26551 2834 26560
rect 2792 26450 2820 26551
rect 2780 26444 2832 26450
rect 2780 26386 2832 26392
rect 2778 23216 2834 23225
rect 2778 23151 2780 23160
rect 2832 23151 2834 23160
rect 2780 23122 2832 23128
rect 2778 19136 2834 19145
rect 2778 19071 2834 19080
rect 2792 18834 2820 19071
rect 2780 18828 2832 18834
rect 2780 18770 2832 18776
rect 2780 18216 2832 18222
rect 2780 18158 2832 18164
rect 2792 17785 2820 18158
rect 2778 17776 2834 17785
rect 2778 17711 2834 17720
rect 2780 17128 2832 17134
rect 2780 17070 2832 17076
rect 2688 16720 2740 16726
rect 2688 16662 2740 16668
rect 2792 16425 2820 17070
rect 2778 16416 2834 16425
rect 2778 16351 2834 16360
rect 2884 14958 2912 29582
rect 4066 29336 4122 29345
rect 4066 29271 4122 29280
rect 4080 24138 4108 29271
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4068 24132 4120 24138
rect 4068 24074 4120 24080
rect 3056 24064 3108 24070
rect 3056 24006 3108 24012
rect 2872 14952 2924 14958
rect 2872 14894 2924 14900
rect 2872 13728 2924 13734
rect 2778 13696 2834 13705
rect 2872 13670 2924 13676
rect 2778 13631 2834 13640
rect 2792 13394 2820 13631
rect 2884 13462 2912 13670
rect 2872 13456 2924 13462
rect 2872 13398 2924 13404
rect 2780 13388 2832 13394
rect 2780 13330 2832 13336
rect 2504 11144 2556 11150
rect 2504 11086 2556 11092
rect 2596 11008 2648 11014
rect 2596 10950 2648 10956
rect 2608 10742 2636 10950
rect 2596 10736 2648 10742
rect 2596 10678 2648 10684
rect 2964 10600 3016 10606
rect 2964 10542 3016 10548
rect 2870 10296 2926 10305
rect 2870 10231 2926 10240
rect 2780 9920 2832 9926
rect 2780 9862 2832 9868
rect 2792 9654 2820 9862
rect 2780 9648 2832 9654
rect 2780 9590 2832 9596
rect 2884 9518 2912 10231
rect 2976 9625 3004 10542
rect 3068 10062 3096 24006
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4632 22982 4660 48486
rect 4724 23866 4752 49098
rect 5184 47734 5212 51200
rect 6472 49230 6500 51200
rect 7116 49994 7144 51200
rect 7116 49966 7236 49994
rect 6460 49224 6512 49230
rect 6460 49166 6512 49172
rect 7104 49224 7156 49230
rect 7104 49166 7156 49172
rect 5264 49088 5316 49094
rect 5264 49030 5316 49036
rect 6460 49088 6512 49094
rect 6460 49030 6512 49036
rect 5172 47728 5224 47734
rect 5172 47670 5224 47676
rect 5276 38010 5304 49030
rect 5356 48068 5408 48074
rect 5356 48010 5408 48016
rect 5368 47802 5396 48010
rect 5356 47796 5408 47802
rect 5356 47738 5408 47744
rect 5264 38004 5316 38010
rect 5264 37946 5316 37952
rect 6368 28212 6420 28218
rect 6368 28154 6420 28160
rect 6184 26580 6236 26586
rect 6184 26522 6236 26528
rect 5724 26240 5776 26246
rect 5724 26182 5776 26188
rect 5736 25974 5764 26182
rect 5724 25968 5776 25974
rect 5724 25910 5776 25916
rect 6196 25770 6224 26522
rect 6276 26444 6328 26450
rect 6276 26386 6328 26392
rect 6184 25764 6236 25770
rect 6184 25706 6236 25712
rect 4712 23860 4764 23866
rect 4712 23802 4764 23808
rect 4620 22976 4672 22982
rect 4620 22918 4672 22924
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 4068 21888 4120 21894
rect 3974 21856 4030 21865
rect 4068 21830 4120 21836
rect 3974 21791 4030 21800
rect 3988 21418 4016 21791
rect 3976 21412 4028 21418
rect 3976 21354 4028 21360
rect 4080 21185 4108 21830
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4066 21176 4122 21185
rect 4214 21168 4522 21188
rect 4066 21111 4122 21120
rect 5632 20936 5684 20942
rect 5632 20878 5684 20884
rect 5644 20466 5672 20878
rect 5632 20460 5684 20466
rect 5632 20402 5684 20408
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 4066 19816 4122 19825
rect 3976 19780 4028 19786
rect 4066 19751 4122 19760
rect 3976 19722 4028 19728
rect 3988 19514 4016 19722
rect 4080 19514 4108 19751
rect 3976 19508 4028 19514
rect 3976 19450 4028 19456
rect 4068 19508 4120 19514
rect 4068 19450 4120 19456
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 4066 18456 4122 18465
rect 4066 18391 4122 18400
rect 4080 18154 4108 18391
rect 4068 18148 4120 18154
rect 4068 18090 4120 18096
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4068 13456 4120 13462
rect 4068 13398 4120 13404
rect 4080 13025 4108 13398
rect 4066 13016 4122 13025
rect 4066 12951 4122 12960
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 4068 9648 4120 9654
rect 2962 9616 3018 9625
rect 4068 9590 4120 9596
rect 2962 9551 3018 9560
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 4080 8945 4108 9590
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4066 8936 4122 8945
rect 4066 8871 4122 8880
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 2778 6896 2834 6905
rect 2778 6831 2780 6840
rect 2832 6831 2834 6840
rect 2780 6802 2832 6808
rect 3620 6225 3648 8570
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 3606 6216 3662 6225
rect 3606 6151 3662 6160
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 2320 5704 2372 5710
rect 2320 5646 2372 5652
rect 3056 5568 3108 5574
rect 2778 5536 2834 5545
rect 3056 5510 3108 5516
rect 2778 5471 2834 5480
rect 2792 5166 2820 5471
rect 3068 5302 3096 5510
rect 3056 5296 3108 5302
rect 3056 5238 3108 5244
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 2778 4856 2834 4865
rect 2688 4820 2740 4826
rect 4214 4848 4522 4868
rect 2778 4791 2834 4800
rect 2688 4762 2740 4768
rect 1964 4542 2084 4570
rect 2056 4146 2084 4542
rect 2044 4140 2096 4146
rect 2044 4082 2096 4088
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 1676 3936 1728 3942
rect 1676 3878 1728 3884
rect 664 2916 716 2922
rect 664 2858 716 2864
rect 676 800 704 2858
rect 1308 2576 1360 2582
rect 1308 2518 1360 2524
rect 1320 800 1348 2518
rect 1596 2514 1624 3878
rect 1688 3602 1716 3878
rect 1952 3732 2004 3738
rect 1952 3674 2004 3680
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 1860 3596 1912 3602
rect 1860 3538 1912 3544
rect 1872 3505 1900 3538
rect 1858 3496 1914 3505
rect 1858 3431 1914 3440
rect 1964 3194 1992 3674
rect 2056 3466 2084 4082
rect 2044 3460 2096 3466
rect 2044 3402 2096 3408
rect 1952 3188 2004 3194
rect 1952 3130 2004 3136
rect 2596 3188 2648 3194
rect 2596 3130 2648 3136
rect 1952 3052 2004 3058
rect 1952 2994 2004 3000
rect 1584 2508 1636 2514
rect 1584 2450 1636 2456
rect 1964 800 1992 2994
rect 2608 800 2636 3130
rect 2700 2854 2728 4762
rect 2792 4690 2820 4791
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 3700 4480 3752 4486
rect 3700 4422 3752 4428
rect 3712 4185 3740 4422
rect 3698 4176 3754 4185
rect 3698 4111 3754 4120
rect 3792 4140 3844 4146
rect 3792 4082 3844 4088
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 3516 3936 3568 3942
rect 3516 3878 3568 3884
rect 2780 3120 2832 3126
rect 2780 3062 2832 3068
rect 2688 2848 2740 2854
rect 2688 2790 2740 2796
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 1950 0 2006 800
rect 2594 0 2650 800
rect 2792 785 2820 3062
rect 2884 2378 2912 3878
rect 3528 3670 3556 3878
rect 3516 3664 3568 3670
rect 3516 3606 3568 3612
rect 3804 3534 3832 4082
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 3884 3664 3936 3670
rect 3884 3606 3936 3612
rect 3792 3528 3844 3534
rect 3792 3470 3844 3476
rect 3516 3392 3568 3398
rect 3516 3334 3568 3340
rect 3528 3126 3556 3334
rect 3516 3120 3568 3126
rect 3516 3062 3568 3068
rect 3332 2984 3384 2990
rect 3332 2926 3384 2932
rect 3240 2916 3292 2922
rect 3240 2858 3292 2864
rect 2872 2372 2924 2378
rect 2872 2314 2924 2320
rect 3252 800 3280 2858
rect 3344 2650 3372 2926
rect 3332 2644 3384 2650
rect 3332 2586 3384 2592
rect 3424 2372 3476 2378
rect 3424 2314 3476 2320
rect 3436 2145 3464 2314
rect 3422 2136 3478 2145
rect 3422 2071 3478 2080
rect 3896 800 3924 3606
rect 4632 3602 4660 3878
rect 4620 3596 4672 3602
rect 4620 3538 4672 3544
rect 5000 3466 5028 3878
rect 6288 3738 6316 26386
rect 6380 26314 6408 28154
rect 6472 26382 6500 49030
rect 6552 48680 6604 48686
rect 6552 48622 6604 48628
rect 6564 47802 6592 48622
rect 6552 47796 6604 47802
rect 6552 47738 6604 47744
rect 7116 47666 7144 49166
rect 7208 48686 7236 49966
rect 7196 48680 7248 48686
rect 7196 48622 7248 48628
rect 7564 48612 7616 48618
rect 7564 48554 7616 48560
rect 7576 48278 7604 48554
rect 7564 48272 7616 48278
rect 7564 48214 7616 48220
rect 6920 47660 6972 47666
rect 6920 47602 6972 47608
rect 7104 47660 7156 47666
rect 7104 47602 7156 47608
rect 6932 47190 6960 47602
rect 7760 47598 7788 51200
rect 7656 47592 7708 47598
rect 7656 47534 7708 47540
rect 7748 47592 7800 47598
rect 7748 47534 7800 47540
rect 7668 47258 7696 47534
rect 7656 47252 7708 47258
rect 7656 47194 7708 47200
rect 6920 47184 6972 47190
rect 6920 47126 6972 47132
rect 7932 47048 7984 47054
rect 7932 46990 7984 46996
rect 7944 43314 7972 46990
rect 7932 43308 7984 43314
rect 7932 43250 7984 43256
rect 6920 38276 6972 38282
rect 6920 38218 6972 38224
rect 6460 26376 6512 26382
rect 6460 26318 6512 26324
rect 6368 26308 6420 26314
rect 6368 26250 6420 26256
rect 6932 25294 6960 38218
rect 7656 32768 7708 32774
rect 7656 32710 7708 32716
rect 7668 31822 7696 32710
rect 7656 31816 7708 31822
rect 7656 31758 7708 31764
rect 7656 30728 7708 30734
rect 7656 30670 7708 30676
rect 7012 29164 7064 29170
rect 7012 29106 7064 29112
rect 7024 28626 7052 29106
rect 7012 28620 7064 28626
rect 7012 28562 7064 28568
rect 7564 26784 7616 26790
rect 7564 26726 7616 26732
rect 7576 26450 7604 26726
rect 7564 26444 7616 26450
rect 7564 26386 7616 26392
rect 7012 25832 7064 25838
rect 7012 25774 7064 25780
rect 7024 25498 7052 25774
rect 7012 25492 7064 25498
rect 7012 25434 7064 25440
rect 6644 25288 6696 25294
rect 6644 25230 6696 25236
rect 6920 25288 6972 25294
rect 6920 25230 6972 25236
rect 6656 21554 6684 25230
rect 7668 24818 7696 30670
rect 7656 24812 7708 24818
rect 7656 24754 7708 24760
rect 6736 21956 6788 21962
rect 6736 21898 6788 21904
rect 6748 21690 6776 21898
rect 6736 21684 6788 21690
rect 6736 21626 6788 21632
rect 6644 21548 6696 21554
rect 6644 21490 6696 21496
rect 6656 20942 6684 21490
rect 6644 20936 6696 20942
rect 6644 20878 6696 20884
rect 6644 20800 6696 20806
rect 6644 20742 6696 20748
rect 6656 19922 6684 20742
rect 6644 19916 6696 19922
rect 6644 19858 6696 19864
rect 6920 19916 6972 19922
rect 6920 19858 6972 19864
rect 6932 13462 6960 19858
rect 7564 17536 7616 17542
rect 7564 17478 7616 17484
rect 7576 17338 7604 17478
rect 7564 17332 7616 17338
rect 7564 17274 7616 17280
rect 7668 15570 7696 24754
rect 7656 15564 7708 15570
rect 7656 15506 7708 15512
rect 6920 13456 6972 13462
rect 6920 13398 6972 13404
rect 7944 12782 7972 43250
rect 8404 41414 8432 51200
rect 8944 49088 8996 49094
rect 8944 49030 8996 49036
rect 8956 48754 8984 49030
rect 8944 48748 8996 48754
rect 8944 48690 8996 48696
rect 9692 48686 9720 51200
rect 10324 49224 10376 49230
rect 10324 49166 10376 49172
rect 9128 48680 9180 48686
rect 9128 48622 9180 48628
rect 9680 48680 9732 48686
rect 9680 48622 9732 48628
rect 9036 48544 9088 48550
rect 9036 48486 9088 48492
rect 9048 48346 9076 48486
rect 9140 48346 9168 48622
rect 9036 48340 9088 48346
rect 9036 48282 9088 48288
rect 9128 48340 9180 48346
rect 9128 48282 9180 48288
rect 10336 48210 10364 49166
rect 10704 48210 10732 51326
rect 10966 51200 11022 52000
rect 11610 51200 11666 52000
rect 12254 51354 12310 52000
rect 12254 51326 12388 51354
rect 12254 51200 12310 51326
rect 10324 48204 10376 48210
rect 10324 48146 10376 48152
rect 10692 48204 10744 48210
rect 10692 48146 10744 48152
rect 10980 48006 11008 51200
rect 11624 49230 11652 51200
rect 11520 49224 11572 49230
rect 11520 49166 11572 49172
rect 11612 49224 11664 49230
rect 11612 49166 11664 49172
rect 11532 48754 11560 49166
rect 11888 49088 11940 49094
rect 11888 49030 11940 49036
rect 11520 48748 11572 48754
rect 11520 48690 11572 48696
rect 11704 48680 11756 48686
rect 11704 48622 11756 48628
rect 11612 48068 11664 48074
rect 11612 48010 11664 48016
rect 10968 48000 11020 48006
rect 10968 47942 11020 47948
rect 11624 47802 11652 48010
rect 11716 47802 11744 48622
rect 11612 47796 11664 47802
rect 11612 47738 11664 47744
rect 11704 47796 11756 47802
rect 11704 47738 11756 47744
rect 11520 47660 11572 47666
rect 11520 47602 11572 47608
rect 8404 41386 8524 41414
rect 8300 36780 8352 36786
rect 8300 36722 8352 36728
rect 8312 34134 8340 36722
rect 8496 34406 8524 41386
rect 8944 38344 8996 38350
rect 8944 38286 8996 38292
rect 8956 37874 8984 38286
rect 8944 37868 8996 37874
rect 8944 37810 8996 37816
rect 8956 37466 8984 37810
rect 9128 37664 9180 37670
rect 9128 37606 9180 37612
rect 8944 37460 8996 37466
rect 8944 37402 8996 37408
rect 9140 37330 9168 37606
rect 9128 37324 9180 37330
rect 9128 37266 9180 37272
rect 8944 37256 8996 37262
rect 8944 37198 8996 37204
rect 8956 36922 8984 37198
rect 8944 36916 8996 36922
rect 8944 36858 8996 36864
rect 9036 36780 9088 36786
rect 9036 36722 9088 36728
rect 9048 35834 9076 36722
rect 9036 35828 9088 35834
rect 9036 35770 9088 35776
rect 9404 35692 9456 35698
rect 9404 35634 9456 35640
rect 8484 34400 8536 34406
rect 8484 34342 8536 34348
rect 8300 34128 8352 34134
rect 8300 34070 8352 34076
rect 8312 33522 8340 34070
rect 9220 33992 9272 33998
rect 9220 33934 9272 33940
rect 8300 33516 8352 33522
rect 8300 33458 8352 33464
rect 8300 32224 8352 32230
rect 8300 32166 8352 32172
rect 8208 31272 8260 31278
rect 8208 31214 8260 31220
rect 8220 29714 8248 31214
rect 8312 31210 8340 32166
rect 8300 31204 8352 31210
rect 8300 31146 8352 31152
rect 8944 30048 8996 30054
rect 8944 29990 8996 29996
rect 8956 29782 8984 29990
rect 8944 29776 8996 29782
rect 8944 29718 8996 29724
rect 8208 29708 8260 29714
rect 8208 29650 8260 29656
rect 8220 29238 8248 29650
rect 8956 29578 8984 29718
rect 8300 29572 8352 29578
rect 8300 29514 8352 29520
rect 8944 29572 8996 29578
rect 8944 29514 8996 29520
rect 8208 29232 8260 29238
rect 8208 29174 8260 29180
rect 8312 28506 8340 29514
rect 8484 29504 8536 29510
rect 8484 29446 8536 29452
rect 8496 29034 8524 29446
rect 8484 29028 8536 29034
rect 8484 28970 8536 28976
rect 8312 28478 8432 28506
rect 8404 28422 8432 28478
rect 8392 28416 8444 28422
rect 8392 28358 8444 28364
rect 8404 25770 8432 28358
rect 8392 25764 8444 25770
rect 8392 25706 8444 25712
rect 8496 24886 8524 28970
rect 9232 28558 9260 33934
rect 9416 31754 9444 35634
rect 11532 35154 11560 47602
rect 11704 36712 11756 36718
rect 11704 36654 11756 36660
rect 11716 36378 11744 36654
rect 11704 36372 11756 36378
rect 11704 36314 11756 36320
rect 11520 35148 11572 35154
rect 11520 35090 11572 35096
rect 10232 34060 10284 34066
rect 10232 34002 10284 34008
rect 10244 33590 10272 34002
rect 10876 33992 10928 33998
rect 10876 33934 10928 33940
rect 10324 33924 10376 33930
rect 10324 33866 10376 33872
rect 10336 33658 10364 33866
rect 10784 33856 10836 33862
rect 10784 33798 10836 33804
rect 10324 33652 10376 33658
rect 10324 33594 10376 33600
rect 10232 33584 10284 33590
rect 10232 33526 10284 33532
rect 9772 33312 9824 33318
rect 9772 33254 9824 33260
rect 9680 31816 9732 31822
rect 9680 31758 9732 31764
rect 9416 31726 9628 31754
rect 9312 29708 9364 29714
rect 9312 29650 9364 29656
rect 9220 28552 9272 28558
rect 9324 28540 9352 29650
rect 9496 29504 9548 29510
rect 9496 29446 9548 29452
rect 9402 29200 9458 29209
rect 9508 29170 9536 29446
rect 9402 29135 9404 29144
rect 9456 29135 9458 29144
rect 9496 29164 9548 29170
rect 9404 29106 9456 29112
rect 9496 29106 9548 29112
rect 9416 28762 9444 29106
rect 9404 28756 9456 28762
rect 9404 28698 9456 28704
rect 9404 28552 9456 28558
rect 9324 28512 9404 28540
rect 9220 28494 9272 28500
rect 9404 28494 9456 28500
rect 9036 27464 9088 27470
rect 9036 27406 9088 27412
rect 8666 27024 8722 27033
rect 9048 26994 9076 27406
rect 9232 27334 9260 28494
rect 9494 27976 9550 27985
rect 9494 27911 9550 27920
rect 9312 27532 9364 27538
rect 9312 27474 9364 27480
rect 9220 27328 9272 27334
rect 9220 27270 9272 27276
rect 8666 26959 8668 26968
rect 8720 26959 8722 26968
rect 8852 26988 8904 26994
rect 8668 26930 8720 26936
rect 8852 26930 8904 26936
rect 9036 26988 9088 26994
rect 9036 26930 9088 26936
rect 8864 26625 8892 26930
rect 9128 26920 9180 26926
rect 9128 26862 9180 26868
rect 8850 26616 8906 26625
rect 8850 26551 8906 26560
rect 8668 25832 8720 25838
rect 8668 25774 8720 25780
rect 8484 24880 8536 24886
rect 8484 24822 8536 24828
rect 8208 24268 8260 24274
rect 8208 24210 8260 24216
rect 8220 23526 8248 24210
rect 8300 23792 8352 23798
rect 8300 23734 8352 23740
rect 8208 23520 8260 23526
rect 8208 23462 8260 23468
rect 8220 23118 8248 23462
rect 8208 23112 8260 23118
rect 8208 23054 8260 23060
rect 8024 23044 8076 23050
rect 8024 22986 8076 22992
rect 8036 22778 8064 22986
rect 8024 22772 8076 22778
rect 8024 22714 8076 22720
rect 8036 20942 8064 22714
rect 8312 22710 8340 23734
rect 8390 23080 8446 23089
rect 8390 23015 8392 23024
rect 8444 23015 8446 23024
rect 8392 22986 8444 22992
rect 8300 22704 8352 22710
rect 8300 22646 8352 22652
rect 8208 22432 8260 22438
rect 8208 22374 8260 22380
rect 8220 22098 8248 22374
rect 8208 22092 8260 22098
rect 8208 22034 8260 22040
rect 8484 21684 8536 21690
rect 8484 21626 8536 21632
rect 8024 20936 8076 20942
rect 8024 20878 8076 20884
rect 8208 20868 8260 20874
rect 8208 20810 8260 20816
rect 8024 20392 8076 20398
rect 8024 20334 8076 20340
rect 7932 12776 7984 12782
rect 7932 12718 7984 12724
rect 7748 8016 7800 8022
rect 7748 7958 7800 7964
rect 6736 4140 6788 4146
rect 6736 4082 6788 4088
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 6552 3936 6604 3942
rect 6552 3878 6604 3884
rect 6276 3732 6328 3738
rect 6276 3674 6328 3680
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 4988 3460 5040 3466
rect 4988 3402 5040 3408
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 4802 2408 4858 2417
rect 4540 800 4568 2382
rect 4802 2343 4858 2352
rect 4816 2310 4844 2343
rect 4804 2304 4856 2310
rect 4804 2246 4856 2252
rect 5184 800 5212 3538
rect 6460 2984 6512 2990
rect 6460 2926 6512 2932
rect 5816 2848 5868 2854
rect 5816 2790 5868 2796
rect 5828 2514 5856 2790
rect 6184 2576 6236 2582
rect 6184 2518 6236 2524
rect 5816 2508 5868 2514
rect 5816 2450 5868 2456
rect 5828 870 5948 898
rect 5828 800 5856 870
rect 2778 776 2834 785
rect 2778 711 2834 720
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 5920 762 5948 870
rect 6196 762 6224 2518
rect 6472 800 6500 2926
rect 6564 2514 6592 3878
rect 6748 3738 6776 4082
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 7392 3602 7420 4082
rect 7760 4078 7788 7958
rect 8036 4486 8064 20334
rect 8220 20262 8248 20810
rect 8208 20256 8260 20262
rect 8208 20198 8260 20204
rect 8220 19990 8248 20198
rect 8208 19984 8260 19990
rect 8208 19926 8260 19932
rect 8300 18148 8352 18154
rect 8300 18090 8352 18096
rect 8312 17814 8340 18090
rect 8300 17808 8352 17814
rect 8300 17750 8352 17756
rect 8496 12850 8524 21626
rect 8484 12844 8536 12850
rect 8484 12786 8536 12792
rect 8024 4480 8076 4486
rect 8024 4422 8076 4428
rect 7748 4072 7800 4078
rect 7748 4014 7800 4020
rect 7564 3936 7616 3942
rect 7564 3878 7616 3884
rect 7380 3596 7432 3602
rect 7380 3538 7432 3544
rect 6644 3528 6696 3534
rect 6644 3470 6696 3476
rect 6656 3058 6684 3470
rect 7104 3460 7156 3466
rect 7104 3402 7156 3408
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 6552 2508 6604 2514
rect 6552 2450 6604 2456
rect 7116 800 7144 3402
rect 7576 3126 7604 3878
rect 7564 3120 7616 3126
rect 7564 3062 7616 3068
rect 8392 3052 8444 3058
rect 8392 2994 8444 3000
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 7760 800 7788 2382
rect 8404 800 8432 2994
rect 8680 2378 8708 25774
rect 9140 24857 9168 26862
rect 9324 26518 9352 27474
rect 9508 27130 9536 27911
rect 9496 27124 9548 27130
rect 9496 27066 9548 27072
rect 9312 26512 9364 26518
rect 9218 26480 9274 26489
rect 9312 26454 9364 26460
rect 9218 26415 9220 26424
rect 9272 26415 9274 26424
rect 9220 26386 9272 26392
rect 9220 26308 9272 26314
rect 9220 26250 9272 26256
rect 9126 24848 9182 24857
rect 9126 24783 9182 24792
rect 8760 24744 8812 24750
rect 8760 24686 8812 24692
rect 8772 12434 8800 24686
rect 8852 24200 8904 24206
rect 8852 24142 8904 24148
rect 8864 23118 8892 24142
rect 8944 23724 8996 23730
rect 8944 23666 8996 23672
rect 8956 23254 8984 23666
rect 8944 23248 8996 23254
rect 8944 23190 8996 23196
rect 8852 23112 8904 23118
rect 8852 23054 8904 23060
rect 8944 22704 8996 22710
rect 8944 22646 8996 22652
rect 8852 22636 8904 22642
rect 8852 22578 8904 22584
rect 8864 22098 8892 22578
rect 8956 22114 8984 22646
rect 9036 22160 9088 22166
rect 8956 22108 9036 22114
rect 8956 22102 9088 22108
rect 8852 22092 8904 22098
rect 8852 22034 8904 22040
rect 8956 22086 9076 22102
rect 8956 20942 8984 22086
rect 9140 22012 9168 24783
rect 9232 22030 9260 26250
rect 9324 25498 9352 26454
rect 9600 25702 9628 31726
rect 9692 30326 9720 31758
rect 9680 30320 9732 30326
rect 9680 30262 9732 30268
rect 9680 29164 9732 29170
rect 9680 29106 9732 29112
rect 9692 28558 9720 29106
rect 9784 29102 9812 33254
rect 10244 33114 10272 33526
rect 10796 33522 10824 33798
rect 10508 33516 10560 33522
rect 10508 33458 10560 33464
rect 10692 33516 10744 33522
rect 10692 33458 10744 33464
rect 10784 33516 10836 33522
rect 10784 33458 10836 33464
rect 10232 33108 10284 33114
rect 10232 33050 10284 33056
rect 10324 32428 10376 32434
rect 10520 32416 10548 33458
rect 10704 32502 10732 33458
rect 10888 33318 10916 33934
rect 11244 33584 11296 33590
rect 11244 33526 11296 33532
rect 10968 33516 11020 33522
rect 10968 33458 11020 33464
rect 10876 33312 10928 33318
rect 10876 33254 10928 33260
rect 10888 32858 10916 33254
rect 10796 32842 10916 32858
rect 10784 32836 10916 32842
rect 10836 32830 10916 32836
rect 10784 32778 10836 32784
rect 10692 32496 10744 32502
rect 10692 32438 10744 32444
rect 10376 32388 10548 32416
rect 10324 32370 10376 32376
rect 10232 32224 10284 32230
rect 10232 32166 10284 32172
rect 10244 31822 10272 32166
rect 10520 31958 10548 32388
rect 10600 32428 10652 32434
rect 10600 32370 10652 32376
rect 10612 32026 10640 32370
rect 10600 32020 10652 32026
rect 10600 31962 10652 31968
rect 10508 31952 10560 31958
rect 10508 31894 10560 31900
rect 10232 31816 10284 31822
rect 10232 31758 10284 31764
rect 10704 31686 10732 32438
rect 10980 32434 11008 33458
rect 11256 33114 11284 33526
rect 11244 33108 11296 33114
rect 11244 33050 11296 33056
rect 11060 32972 11112 32978
rect 11060 32914 11112 32920
rect 10968 32428 11020 32434
rect 10968 32370 11020 32376
rect 10980 31822 11008 32370
rect 11072 32230 11100 32914
rect 11796 32428 11848 32434
rect 11796 32370 11848 32376
rect 11612 32292 11664 32298
rect 11612 32234 11664 32240
rect 11060 32224 11112 32230
rect 11060 32166 11112 32172
rect 10876 31816 10928 31822
rect 10876 31758 10928 31764
rect 10968 31816 11020 31822
rect 10968 31758 11020 31764
rect 10324 31680 10376 31686
rect 10324 31622 10376 31628
rect 10692 31680 10744 31686
rect 10692 31622 10744 31628
rect 10336 31414 10364 31622
rect 10888 31414 10916 31758
rect 10324 31408 10376 31414
rect 10324 31350 10376 31356
rect 10876 31408 10928 31414
rect 10876 31350 10928 31356
rect 10968 31340 11020 31346
rect 10968 31282 11020 31288
rect 10416 31204 10468 31210
rect 10416 31146 10468 31152
rect 10140 31136 10192 31142
rect 10140 31078 10192 31084
rect 9772 29096 9824 29102
rect 9772 29038 9824 29044
rect 10152 28558 10180 31078
rect 10428 30938 10456 31146
rect 10784 31136 10836 31142
rect 10784 31078 10836 31084
rect 10416 30932 10468 30938
rect 10416 30874 10468 30880
rect 10508 30932 10560 30938
rect 10508 30874 10560 30880
rect 10520 30258 10548 30874
rect 10796 30734 10824 31078
rect 10980 30938 11008 31282
rect 10968 30932 11020 30938
rect 10968 30874 11020 30880
rect 11072 30870 11100 32166
rect 11520 31952 11572 31958
rect 11520 31894 11572 31900
rect 11532 31278 11560 31894
rect 11624 31754 11652 32234
rect 11704 31952 11756 31958
rect 11704 31894 11756 31900
rect 11716 31822 11744 31894
rect 11808 31822 11836 32370
rect 11704 31816 11756 31822
rect 11704 31758 11756 31764
rect 11796 31816 11848 31822
rect 11796 31758 11848 31764
rect 11612 31748 11664 31754
rect 11612 31690 11664 31696
rect 11520 31272 11572 31278
rect 11520 31214 11572 31220
rect 11060 30864 11112 30870
rect 11060 30806 11112 30812
rect 10784 30728 10836 30734
rect 10784 30670 10836 30676
rect 10508 30252 10560 30258
rect 10508 30194 10560 30200
rect 10232 30184 10284 30190
rect 10232 30126 10284 30132
rect 9680 28552 9732 28558
rect 9680 28494 9732 28500
rect 10140 28552 10192 28558
rect 10140 28494 10192 28500
rect 9772 28076 9824 28082
rect 9956 28076 10008 28082
rect 9824 28036 9904 28064
rect 9772 28018 9824 28024
rect 9772 27872 9824 27878
rect 9678 27840 9734 27849
rect 9772 27814 9824 27820
rect 9678 27775 9734 27784
rect 9692 27606 9720 27775
rect 9680 27600 9732 27606
rect 9680 27542 9732 27548
rect 9678 26888 9734 26897
rect 9678 26823 9680 26832
rect 9732 26823 9734 26832
rect 9680 26794 9732 26800
rect 9784 26586 9812 27814
rect 9876 26790 9904 28036
rect 9956 28018 10008 28024
rect 9968 27985 9996 28018
rect 9954 27976 10010 27985
rect 9954 27911 10010 27920
rect 9956 27872 10008 27878
rect 9954 27840 9956 27849
rect 10008 27840 10010 27849
rect 9954 27775 10010 27784
rect 10046 26888 10102 26897
rect 10046 26823 10048 26832
rect 10100 26823 10102 26832
rect 10048 26794 10100 26800
rect 9864 26784 9916 26790
rect 9864 26726 9916 26732
rect 9772 26580 9824 26586
rect 9772 26522 9824 26528
rect 10152 26314 10180 28494
rect 10244 28422 10272 30126
rect 10324 29096 10376 29102
rect 10324 29038 10376 29044
rect 10232 28416 10284 28422
rect 10232 28358 10284 28364
rect 10244 27402 10272 28358
rect 10336 28082 10364 29038
rect 10324 28076 10376 28082
rect 10324 28018 10376 28024
rect 10324 27464 10376 27470
rect 10324 27406 10376 27412
rect 10232 27396 10284 27402
rect 10232 27338 10284 27344
rect 10336 27130 10364 27406
rect 10508 27396 10560 27402
rect 10508 27338 10560 27344
rect 10324 27124 10376 27130
rect 10324 27066 10376 27072
rect 10336 26382 10364 27066
rect 10416 27056 10468 27062
rect 10414 27024 10416 27033
rect 10468 27024 10470 27033
rect 10414 26959 10470 26968
rect 10520 26790 10548 27338
rect 10692 26988 10744 26994
rect 10692 26930 10744 26936
rect 10600 26920 10652 26926
rect 10600 26862 10652 26868
rect 10508 26784 10560 26790
rect 10508 26726 10560 26732
rect 10612 26625 10640 26862
rect 10598 26616 10654 26625
rect 10598 26551 10654 26560
rect 10612 26518 10640 26551
rect 10600 26512 10652 26518
rect 10600 26454 10652 26460
rect 10324 26376 10376 26382
rect 10324 26318 10376 26324
rect 10140 26308 10192 26314
rect 10140 26250 10192 26256
rect 10336 25906 10364 26318
rect 10704 26314 10732 26930
rect 10692 26308 10744 26314
rect 10692 26250 10744 26256
rect 10324 25900 10376 25906
rect 10324 25842 10376 25848
rect 10140 25832 10192 25838
rect 10140 25774 10192 25780
rect 9588 25696 9640 25702
rect 9588 25638 9640 25644
rect 9954 25528 10010 25537
rect 9312 25492 9364 25498
rect 10152 25498 10180 25774
rect 9954 25463 9956 25472
rect 9312 25434 9364 25440
rect 10008 25463 10010 25472
rect 10140 25492 10192 25498
rect 9956 25434 10008 25440
rect 10140 25434 10192 25440
rect 9312 25356 9364 25362
rect 9312 25298 9364 25304
rect 9324 25226 9352 25298
rect 9312 25220 9364 25226
rect 9312 25162 9364 25168
rect 9496 25220 9548 25226
rect 9496 25162 9548 25168
rect 9312 23248 9364 23254
rect 9312 23190 9364 23196
rect 9048 21984 9168 22012
rect 9220 22024 9272 22030
rect 8944 20936 8996 20942
rect 8944 20878 8996 20884
rect 8944 20460 8996 20466
rect 8944 20402 8996 20408
rect 8956 20058 8984 20402
rect 8944 20052 8996 20058
rect 8944 19994 8996 20000
rect 9048 19854 9076 21984
rect 9220 21966 9272 21972
rect 9324 21894 9352 23190
rect 9404 22432 9456 22438
rect 9404 22374 9456 22380
rect 9416 21894 9444 22374
rect 9312 21888 9364 21894
rect 9312 21830 9364 21836
rect 9404 21888 9456 21894
rect 9404 21830 9456 21836
rect 9324 21622 9352 21830
rect 9312 21616 9364 21622
rect 9312 21558 9364 21564
rect 9220 21344 9272 21350
rect 9220 21286 9272 21292
rect 9232 20942 9260 21286
rect 9220 20936 9272 20942
rect 9220 20878 9272 20884
rect 9128 20868 9180 20874
rect 9128 20810 9180 20816
rect 9140 20534 9168 20810
rect 9128 20528 9180 20534
rect 9128 20470 9180 20476
rect 9036 19848 9088 19854
rect 9036 19790 9088 19796
rect 9140 19310 9168 20470
rect 9324 19854 9352 21558
rect 9404 21548 9456 21554
rect 9508 21536 9536 25162
rect 9968 24206 9996 25434
rect 10692 25356 10744 25362
rect 10692 25298 10744 25304
rect 10048 25288 10100 25294
rect 10048 25230 10100 25236
rect 10060 24886 10088 25230
rect 10048 24880 10100 24886
rect 10048 24822 10100 24828
rect 10704 24410 10732 25298
rect 10796 25294 10824 30670
rect 11624 30666 11652 31690
rect 11808 31346 11836 31758
rect 11796 31340 11848 31346
rect 11796 31282 11848 31288
rect 11704 31136 11756 31142
rect 11704 31078 11756 31084
rect 11612 30660 11664 30666
rect 11612 30602 11664 30608
rect 11716 30326 11744 31078
rect 11796 30660 11848 30666
rect 11796 30602 11848 30608
rect 11808 30394 11836 30602
rect 11796 30388 11848 30394
rect 11796 30330 11848 30336
rect 11704 30320 11756 30326
rect 11704 30262 11756 30268
rect 11152 28008 11204 28014
rect 11152 27950 11204 27956
rect 11164 27606 11192 27950
rect 11900 27614 11928 49030
rect 12360 48668 12388 51326
rect 12898 51200 12954 52000
rect 13542 51354 13598 52000
rect 13280 51326 13598 51354
rect 12440 48680 12492 48686
rect 12360 48640 12440 48668
rect 12440 48622 12492 48628
rect 12912 48142 12940 51200
rect 13280 49230 13308 51326
rect 13542 51200 13598 51326
rect 14186 51200 14242 52000
rect 14830 51354 14886 52000
rect 15474 51354 15530 52000
rect 14830 51326 15148 51354
rect 14830 51200 14886 51326
rect 14200 49298 14228 51200
rect 14188 49292 14240 49298
rect 14188 49234 14240 49240
rect 13268 49224 13320 49230
rect 13268 49166 13320 49172
rect 13452 49088 13504 49094
rect 13452 49030 13504 49036
rect 12900 48136 12952 48142
rect 12900 48078 12952 48084
rect 13360 48000 13412 48006
rect 13360 47942 13412 47948
rect 12072 47660 12124 47666
rect 12072 47602 12124 47608
rect 12084 35766 12112 47602
rect 13268 47456 13320 47462
rect 13268 47398 13320 47404
rect 13280 45966 13308 47398
rect 13268 45960 13320 45966
rect 13268 45902 13320 45908
rect 13084 45824 13136 45830
rect 13084 45766 13136 45772
rect 13096 45558 13124 45766
rect 13084 45552 13136 45558
rect 13084 45494 13136 45500
rect 13176 45416 13228 45422
rect 13176 45358 13228 45364
rect 13188 45082 13216 45358
rect 13176 45076 13228 45082
rect 13176 45018 13228 45024
rect 13372 36854 13400 47942
rect 13360 36848 13412 36854
rect 13360 36790 13412 36796
rect 12716 36576 12768 36582
rect 13464 36530 13492 49030
rect 14188 48680 14240 48686
rect 14188 48622 14240 48628
rect 14372 48680 14424 48686
rect 15120 48668 15148 51326
rect 15304 51326 15530 51354
rect 15200 48680 15252 48686
rect 15120 48640 15200 48668
rect 14372 48622 14424 48628
rect 15200 48622 15252 48628
rect 13728 48068 13780 48074
rect 13728 48010 13780 48016
rect 13740 38826 13768 48010
rect 14200 47666 14228 48622
rect 14384 48346 14412 48622
rect 15108 48544 15160 48550
rect 15108 48486 15160 48492
rect 14372 48340 14424 48346
rect 14372 48282 14424 48288
rect 14464 48136 14516 48142
rect 14464 48078 14516 48084
rect 14188 47660 14240 47666
rect 14188 47602 14240 47608
rect 14476 47122 14504 48078
rect 15120 47530 15148 48486
rect 15108 47524 15160 47530
rect 15108 47466 15160 47472
rect 14464 47116 14516 47122
rect 14464 47058 14516 47064
rect 13820 45416 13872 45422
rect 13820 45358 13872 45364
rect 13728 38820 13780 38826
rect 13728 38762 13780 38768
rect 13832 36582 13860 45358
rect 14004 37732 14056 37738
rect 14004 37674 14056 37680
rect 14096 37732 14148 37738
rect 14096 37674 14148 37680
rect 14016 37398 14044 37674
rect 14004 37392 14056 37398
rect 14004 37334 14056 37340
rect 14108 36650 14136 37674
rect 15304 37330 15332 51326
rect 15474 51200 15530 51326
rect 16118 51354 16174 52000
rect 16118 51326 16528 51354
rect 16118 51200 16174 51326
rect 16500 49314 16528 51326
rect 16762 51200 16818 52000
rect 17406 51200 17462 52000
rect 18050 51200 18106 52000
rect 18694 51200 18750 52000
rect 19338 51354 19394 52000
rect 19982 51354 20038 52000
rect 19338 51326 19472 51354
rect 19338 51200 19394 51326
rect 16500 49286 16712 49314
rect 16684 49230 16712 49286
rect 16580 49224 16632 49230
rect 16580 49166 16632 49172
rect 16672 49224 16724 49230
rect 16672 49166 16724 49172
rect 16212 48340 16264 48346
rect 16212 48282 16264 48288
rect 16028 48068 16080 48074
rect 16028 48010 16080 48016
rect 16040 47802 16068 48010
rect 16028 47796 16080 47802
rect 16028 47738 16080 47744
rect 15568 47660 15620 47666
rect 15568 47602 15620 47608
rect 15580 38282 15608 47602
rect 16120 38344 16172 38350
rect 16120 38286 16172 38292
rect 15568 38276 15620 38282
rect 15568 38218 15620 38224
rect 15580 37806 15608 38218
rect 15568 37800 15620 37806
rect 15568 37742 15620 37748
rect 15292 37324 15344 37330
rect 15292 37266 15344 37272
rect 15108 37256 15160 37262
rect 15108 37198 15160 37204
rect 15120 36922 15148 37198
rect 15292 37188 15344 37194
rect 15292 37130 15344 37136
rect 15108 36916 15160 36922
rect 15108 36858 15160 36864
rect 14464 36780 14516 36786
rect 14384 36740 14464 36768
rect 14096 36644 14148 36650
rect 14096 36586 14148 36592
rect 12716 36518 12768 36524
rect 12072 35760 12124 35766
rect 12072 35702 12124 35708
rect 12164 35080 12216 35086
rect 12164 35022 12216 35028
rect 12176 34202 12204 35022
rect 12256 35012 12308 35018
rect 12256 34954 12308 34960
rect 12268 34746 12296 34954
rect 12256 34740 12308 34746
rect 12256 34682 12308 34688
rect 12532 34740 12584 34746
rect 12532 34682 12584 34688
rect 12440 34468 12492 34474
rect 12440 34410 12492 34416
rect 12164 34196 12216 34202
rect 12164 34138 12216 34144
rect 12176 33590 12204 34138
rect 12164 33584 12216 33590
rect 12164 33526 12216 33532
rect 11980 33516 12032 33522
rect 12348 33516 12400 33522
rect 12032 33476 12112 33504
rect 11980 33458 12032 33464
rect 11980 31340 12032 31346
rect 11980 31282 12032 31288
rect 11992 30598 12020 31282
rect 12084 30954 12112 33476
rect 12348 33458 12400 33464
rect 12256 33448 12308 33454
rect 12256 33390 12308 33396
rect 12164 33108 12216 33114
rect 12164 33050 12216 33056
rect 12176 32502 12204 33050
rect 12268 32842 12296 33390
rect 12360 33046 12388 33458
rect 12348 33040 12400 33046
rect 12348 32982 12400 32988
rect 12452 32978 12480 34410
rect 12544 33114 12572 34682
rect 12532 33108 12584 33114
rect 12532 33050 12584 33056
rect 12440 32972 12492 32978
rect 12492 32932 12572 32960
rect 12440 32914 12492 32920
rect 12256 32836 12308 32842
rect 12256 32778 12308 32784
rect 12164 32496 12216 32502
rect 12164 32438 12216 32444
rect 12176 31754 12204 32438
rect 12256 32428 12308 32434
rect 12256 32370 12308 32376
rect 12164 31748 12216 31754
rect 12164 31690 12216 31696
rect 12268 31686 12296 32370
rect 12544 32026 12572 32932
rect 12532 32020 12584 32026
rect 12532 31962 12584 31968
rect 12440 31884 12492 31890
rect 12440 31826 12492 31832
rect 12256 31680 12308 31686
rect 12256 31622 12308 31628
rect 12084 30926 12204 30954
rect 12072 30864 12124 30870
rect 12072 30806 12124 30812
rect 11980 30592 12032 30598
rect 11980 30534 12032 30540
rect 11992 29034 12020 30534
rect 12084 30326 12112 30806
rect 12176 30734 12204 30926
rect 12164 30728 12216 30734
rect 12164 30670 12216 30676
rect 12268 30394 12296 31622
rect 12348 30592 12400 30598
rect 12348 30534 12400 30540
rect 12256 30388 12308 30394
rect 12256 30330 12308 30336
rect 12072 30320 12124 30326
rect 12072 30262 12124 30268
rect 12256 30184 12308 30190
rect 12256 30126 12308 30132
rect 12164 29640 12216 29646
rect 12164 29582 12216 29588
rect 12176 29238 12204 29582
rect 12268 29510 12296 30126
rect 12360 29578 12388 30534
rect 12348 29572 12400 29578
rect 12348 29514 12400 29520
rect 12256 29504 12308 29510
rect 12256 29446 12308 29452
rect 12164 29232 12216 29238
rect 12164 29174 12216 29180
rect 11980 29028 12032 29034
rect 11980 28970 12032 28976
rect 11152 27600 11204 27606
rect 11152 27542 11204 27548
rect 11808 27586 11928 27614
rect 10876 27328 10928 27334
rect 10876 27270 10928 27276
rect 10888 26994 10916 27270
rect 10876 26988 10928 26994
rect 10876 26930 10928 26936
rect 10888 26382 10916 26930
rect 10876 26376 10928 26382
rect 10876 26318 10928 26324
rect 11060 25832 11112 25838
rect 11060 25774 11112 25780
rect 10876 25696 10928 25702
rect 10876 25638 10928 25644
rect 10888 25362 10916 25638
rect 11072 25498 11100 25774
rect 11060 25492 11112 25498
rect 11060 25434 11112 25440
rect 10876 25356 10928 25362
rect 10876 25298 10928 25304
rect 10784 25288 10836 25294
rect 10784 25230 10836 25236
rect 11520 24948 11572 24954
rect 11520 24890 11572 24896
rect 11532 24750 11560 24890
rect 11520 24744 11572 24750
rect 11520 24686 11572 24692
rect 10692 24404 10744 24410
rect 10692 24346 10744 24352
rect 9956 24200 10008 24206
rect 9956 24142 10008 24148
rect 11532 23594 11560 24686
rect 11520 23588 11572 23594
rect 11520 23530 11572 23536
rect 11808 23118 11836 27586
rect 12176 27538 12204 29174
rect 12164 27532 12216 27538
rect 12164 27474 12216 27480
rect 12268 27418 12296 29446
rect 12452 27470 12480 31826
rect 12544 31822 12572 31962
rect 12532 31816 12584 31822
rect 12532 31758 12584 31764
rect 12728 31754 12756 36518
rect 13280 36502 13492 36530
rect 13820 36576 13872 36582
rect 13820 36518 13872 36524
rect 12992 34604 13044 34610
rect 12992 34546 13044 34552
rect 12900 34536 12952 34542
rect 12900 34478 12952 34484
rect 12912 33658 12940 34478
rect 13004 34066 13032 34546
rect 12992 34060 13044 34066
rect 12992 34002 13044 34008
rect 12808 33652 12860 33658
rect 12808 33594 12860 33600
rect 12900 33652 12952 33658
rect 12900 33594 12952 33600
rect 12820 33318 12848 33594
rect 13004 33538 13032 34002
rect 12912 33510 13032 33538
rect 13084 33516 13136 33522
rect 12808 33312 12860 33318
rect 12808 33254 12860 33260
rect 12808 32224 12860 32230
rect 12808 32166 12860 32172
rect 12636 31726 12756 31754
rect 12532 30252 12584 30258
rect 12532 30194 12584 30200
rect 12544 29782 12572 30194
rect 12532 29776 12584 29782
rect 12532 29718 12584 29724
rect 12544 29170 12572 29718
rect 12532 29164 12584 29170
rect 12532 29106 12584 29112
rect 12176 27390 12296 27418
rect 12440 27464 12492 27470
rect 12440 27406 12492 27412
rect 12072 26512 12124 26518
rect 12072 26454 12124 26460
rect 12084 25702 12112 26454
rect 12176 26314 12204 27390
rect 12348 26376 12400 26382
rect 12348 26318 12400 26324
rect 12164 26308 12216 26314
rect 12164 26250 12216 26256
rect 12072 25696 12124 25702
rect 12072 25638 12124 25644
rect 12176 25226 12204 26250
rect 12256 26240 12308 26246
rect 12256 26182 12308 26188
rect 12268 25498 12296 26182
rect 12256 25492 12308 25498
rect 12256 25434 12308 25440
rect 12164 25220 12216 25226
rect 12164 25162 12216 25168
rect 12268 24614 12296 25434
rect 12360 25226 12388 26318
rect 12532 25900 12584 25906
rect 12532 25842 12584 25848
rect 12544 25498 12572 25842
rect 12532 25492 12584 25498
rect 12532 25434 12584 25440
rect 12348 25220 12400 25226
rect 12348 25162 12400 25168
rect 12256 24608 12308 24614
rect 12256 24550 12308 24556
rect 12268 24274 12296 24550
rect 12360 24410 12388 25162
rect 12348 24404 12400 24410
rect 12348 24346 12400 24352
rect 12256 24268 12308 24274
rect 12256 24210 12308 24216
rect 12254 24168 12310 24177
rect 12254 24103 12256 24112
rect 12308 24103 12310 24112
rect 12256 24074 12308 24080
rect 12072 23248 12124 23254
rect 12072 23190 12124 23196
rect 12084 23118 12112 23190
rect 9772 23112 9824 23118
rect 11796 23112 11848 23118
rect 9772 23054 9824 23060
rect 9862 23080 9918 23089
rect 9784 22030 9812 23054
rect 11796 23054 11848 23060
rect 11980 23112 12032 23118
rect 11980 23054 12032 23060
rect 12072 23112 12124 23118
rect 12072 23054 12124 23060
rect 12348 23112 12400 23118
rect 12348 23054 12400 23060
rect 9862 23015 9864 23024
rect 9916 23015 9918 23024
rect 9864 22986 9916 22992
rect 11612 22976 11664 22982
rect 11612 22918 11664 22924
rect 11624 22710 11652 22918
rect 11992 22778 12020 23054
rect 11980 22772 12032 22778
rect 11980 22714 12032 22720
rect 11612 22704 11664 22710
rect 11612 22646 11664 22652
rect 11520 22636 11572 22642
rect 11520 22578 11572 22584
rect 10784 22568 10836 22574
rect 10784 22510 10836 22516
rect 9772 22024 9824 22030
rect 9772 21966 9824 21972
rect 9456 21508 9536 21536
rect 9784 21536 9812 21966
rect 10140 21888 10192 21894
rect 10140 21830 10192 21836
rect 10152 21622 10180 21830
rect 10140 21616 10192 21622
rect 10140 21558 10192 21564
rect 9864 21548 9916 21554
rect 9784 21508 9864 21536
rect 9404 21490 9456 21496
rect 9404 20800 9456 20806
rect 9404 20742 9456 20748
rect 9416 19854 9444 20742
rect 9784 19854 9812 21508
rect 9864 21490 9916 21496
rect 10796 20942 10824 22510
rect 11532 22166 11560 22578
rect 11520 22160 11572 22166
rect 11520 22102 11572 22108
rect 11612 21956 11664 21962
rect 11612 21898 11664 21904
rect 11624 21690 11652 21898
rect 11992 21690 12020 22714
rect 12360 22681 12388 23054
rect 12346 22672 12402 22681
rect 12346 22607 12402 22616
rect 11612 21684 11664 21690
rect 11612 21626 11664 21632
rect 11980 21684 12032 21690
rect 11980 21626 12032 21632
rect 12360 21554 12388 22607
rect 12636 22094 12664 31726
rect 12716 31136 12768 31142
rect 12716 31078 12768 31084
rect 12728 30666 12756 31078
rect 12820 30734 12848 32166
rect 12912 31958 12940 33510
rect 13084 33458 13136 33464
rect 12992 33448 13044 33454
rect 12992 33390 13044 33396
rect 13004 32570 13032 33390
rect 13096 32842 13124 33458
rect 13176 32904 13228 32910
rect 13176 32846 13228 32852
rect 13084 32836 13136 32842
rect 13084 32778 13136 32784
rect 12992 32564 13044 32570
rect 12992 32506 13044 32512
rect 13096 32434 13124 32778
rect 13084 32428 13136 32434
rect 13084 32370 13136 32376
rect 12992 32292 13044 32298
rect 12992 32234 13044 32240
rect 13004 31958 13032 32234
rect 12900 31952 12952 31958
rect 12900 31894 12952 31900
rect 12992 31952 13044 31958
rect 12992 31894 13044 31900
rect 12912 31822 12940 31894
rect 12900 31816 12952 31822
rect 12900 31758 12952 31764
rect 12992 31476 13044 31482
rect 12992 31418 13044 31424
rect 12808 30728 12860 30734
rect 12808 30670 12860 30676
rect 12716 30660 12768 30666
rect 12716 30602 12768 30608
rect 13004 29578 13032 31418
rect 13096 31346 13124 32370
rect 13188 32230 13216 32846
rect 13176 32224 13228 32230
rect 13176 32166 13228 32172
rect 13084 31340 13136 31346
rect 13084 31282 13136 31288
rect 13084 30728 13136 30734
rect 13188 30716 13216 32166
rect 13280 31482 13308 36502
rect 14188 34944 14240 34950
rect 14188 34886 14240 34892
rect 13636 34604 13688 34610
rect 13636 34546 13688 34552
rect 13820 34604 13872 34610
rect 13820 34546 13872 34552
rect 13648 33318 13676 34546
rect 13832 33998 13860 34546
rect 14200 34542 14228 34886
rect 13912 34536 13964 34542
rect 13912 34478 13964 34484
rect 14188 34536 14240 34542
rect 14188 34478 14240 34484
rect 13820 33992 13872 33998
rect 13820 33934 13872 33940
rect 13832 33454 13860 33934
rect 13820 33448 13872 33454
rect 13820 33390 13872 33396
rect 13636 33312 13688 33318
rect 13636 33254 13688 33260
rect 13544 32904 13596 32910
rect 13544 32846 13596 32852
rect 13556 32502 13584 32846
rect 13544 32496 13596 32502
rect 13544 32438 13596 32444
rect 13648 32366 13676 33254
rect 13728 33040 13780 33046
rect 13728 32982 13780 32988
rect 13740 32774 13768 32982
rect 13728 32768 13780 32774
rect 13728 32710 13780 32716
rect 13544 32360 13596 32366
rect 13544 32302 13596 32308
rect 13636 32360 13688 32366
rect 13636 32302 13688 32308
rect 13556 31822 13584 32302
rect 13544 31816 13596 31822
rect 13544 31758 13596 31764
rect 13648 31482 13676 32302
rect 13268 31476 13320 31482
rect 13268 31418 13320 31424
rect 13636 31476 13688 31482
rect 13636 31418 13688 31424
rect 13360 31340 13412 31346
rect 13360 31282 13412 31288
rect 13268 31272 13320 31278
rect 13268 31214 13320 31220
rect 13136 30688 13216 30716
rect 13084 30670 13136 30676
rect 12992 29572 13044 29578
rect 12992 29514 13044 29520
rect 12992 28960 13044 28966
rect 12992 28902 13044 28908
rect 13004 28082 13032 28902
rect 13096 28218 13124 30670
rect 13176 30592 13228 30598
rect 13176 30534 13228 30540
rect 13084 28212 13136 28218
rect 13084 28154 13136 28160
rect 12992 28076 13044 28082
rect 12992 28018 13044 28024
rect 12900 27940 12952 27946
rect 12900 27882 12952 27888
rect 12912 26042 12940 27882
rect 12900 26036 12952 26042
rect 12900 25978 12952 25984
rect 13084 25152 13136 25158
rect 13084 25094 13136 25100
rect 13096 24750 13124 25094
rect 13084 24744 13136 24750
rect 13084 24686 13136 24692
rect 12900 24200 12952 24206
rect 12900 24142 12952 24148
rect 12912 23050 12940 24142
rect 12992 24132 13044 24138
rect 12992 24074 13044 24080
rect 13004 23730 13032 24074
rect 12992 23724 13044 23730
rect 12992 23666 13044 23672
rect 12900 23044 12952 23050
rect 12900 22986 12952 22992
rect 12912 22438 12940 22986
rect 12716 22432 12768 22438
rect 12716 22374 12768 22380
rect 12900 22432 12952 22438
rect 12900 22374 12952 22380
rect 12452 22066 12664 22094
rect 12348 21548 12400 21554
rect 12348 21490 12400 21496
rect 11152 21480 11204 21486
rect 11152 21422 11204 21428
rect 11164 21146 11192 21422
rect 11152 21140 11204 21146
rect 11152 21082 11204 21088
rect 10784 20936 10836 20942
rect 10784 20878 10836 20884
rect 10324 20800 10376 20806
rect 10324 20742 10376 20748
rect 10336 20602 10364 20742
rect 10324 20596 10376 20602
rect 10324 20538 10376 20544
rect 10796 20534 10824 20878
rect 10784 20528 10836 20534
rect 10784 20470 10836 20476
rect 10692 20460 10744 20466
rect 10692 20402 10744 20408
rect 10140 20256 10192 20262
rect 10140 20198 10192 20204
rect 9312 19848 9364 19854
rect 9312 19790 9364 19796
rect 9404 19848 9456 19854
rect 9404 19790 9456 19796
rect 9772 19848 9824 19854
rect 9772 19790 9824 19796
rect 9128 19304 9180 19310
rect 9128 19246 9180 19252
rect 9140 17746 9168 19246
rect 9324 18834 9352 19790
rect 9404 19372 9456 19378
rect 9404 19314 9456 19320
rect 9864 19372 9916 19378
rect 9864 19314 9916 19320
rect 9416 18970 9444 19314
rect 9772 19168 9824 19174
rect 9772 19110 9824 19116
rect 9404 18964 9456 18970
rect 9404 18906 9456 18912
rect 9312 18828 9364 18834
rect 9312 18770 9364 18776
rect 9784 18766 9812 19110
rect 9772 18760 9824 18766
rect 9772 18702 9824 18708
rect 9128 17740 9180 17746
rect 9128 17682 9180 17688
rect 9876 17678 9904 19314
rect 10152 18766 10180 20198
rect 10232 19848 10284 19854
rect 10232 19790 10284 19796
rect 10244 18766 10272 19790
rect 10704 19378 10732 20402
rect 10692 19372 10744 19378
rect 10692 19314 10744 19320
rect 10140 18760 10192 18766
rect 10140 18702 10192 18708
rect 10232 18760 10284 18766
rect 10232 18702 10284 18708
rect 11244 18760 11296 18766
rect 11244 18702 11296 18708
rect 11256 17746 11284 18702
rect 11244 17740 11296 17746
rect 11244 17682 11296 17688
rect 11336 17740 11388 17746
rect 11336 17682 11388 17688
rect 9864 17672 9916 17678
rect 9864 17614 9916 17620
rect 8852 17604 8904 17610
rect 8852 17546 8904 17552
rect 10048 17604 10100 17610
rect 10048 17546 10100 17552
rect 8864 17338 8892 17546
rect 10060 17338 10088 17546
rect 10416 17536 10468 17542
rect 10416 17478 10468 17484
rect 10508 17536 10560 17542
rect 10508 17478 10560 17484
rect 10428 17377 10456 17478
rect 10414 17368 10470 17377
rect 8852 17332 8904 17338
rect 8852 17274 8904 17280
rect 10048 17332 10100 17338
rect 10414 17303 10470 17312
rect 10048 17274 10100 17280
rect 10520 17202 10548 17478
rect 9772 17196 9824 17202
rect 9772 17138 9824 17144
rect 9956 17196 10008 17202
rect 9956 17138 10008 17144
rect 10508 17196 10560 17202
rect 10508 17138 10560 17144
rect 9784 12850 9812 17138
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 8772 12406 9076 12434
rect 8668 2372 8720 2378
rect 8668 2314 8720 2320
rect 9048 800 9076 12406
rect 9128 6180 9180 6186
rect 9128 6122 9180 6128
rect 9140 2854 9168 6122
rect 9968 4146 9996 17138
rect 11256 16658 11284 17682
rect 11244 16652 11296 16658
rect 11244 16594 11296 16600
rect 10508 12776 10560 12782
rect 10508 12718 10560 12724
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 10324 4140 10376 4146
rect 10324 4082 10376 4088
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 9968 2854 9996 3538
rect 9128 2848 9180 2854
rect 9128 2790 9180 2796
rect 9956 2848 10008 2854
rect 9956 2790 10008 2796
rect 9680 2372 9732 2378
rect 9680 2314 9732 2320
rect 9692 800 9720 2314
rect 10336 800 10364 4082
rect 10520 3738 10548 12718
rect 11348 4146 11376 17682
rect 11980 17672 12032 17678
rect 11980 17614 12032 17620
rect 11992 17202 12020 17614
rect 11520 17196 11572 17202
rect 11520 17138 11572 17144
rect 11980 17196 12032 17202
rect 11980 17138 12032 17144
rect 11532 16250 11560 17138
rect 11888 17060 11940 17066
rect 11888 17002 11940 17008
rect 11704 16992 11756 16998
rect 11704 16934 11756 16940
rect 11716 16590 11744 16934
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11900 16522 11928 17002
rect 11888 16516 11940 16522
rect 11888 16458 11940 16464
rect 11704 16448 11756 16454
rect 11704 16390 11756 16396
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 11520 16244 11572 16250
rect 11520 16186 11572 16192
rect 11532 16114 11560 16186
rect 11716 16182 11744 16390
rect 11808 16250 11836 16390
rect 11796 16244 11848 16250
rect 11796 16186 11848 16192
rect 11704 16176 11756 16182
rect 11704 16118 11756 16124
rect 11520 16108 11572 16114
rect 11520 16050 11572 16056
rect 11612 12844 11664 12850
rect 11612 12786 11664 12792
rect 11624 12238 11652 12786
rect 11612 12232 11664 12238
rect 11612 12174 11664 12180
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 11716 11218 11744 12038
rect 11704 11212 11756 11218
rect 11704 11154 11756 11160
rect 12452 7562 12480 22066
rect 12532 20256 12584 20262
rect 12532 20198 12584 20204
rect 12544 19446 12572 20198
rect 12532 19440 12584 19446
rect 12532 19382 12584 19388
rect 12624 19304 12676 19310
rect 12624 19246 12676 19252
rect 12636 18970 12664 19246
rect 12624 18964 12676 18970
rect 12624 18906 12676 18912
rect 12636 18766 12664 18906
rect 12624 18760 12676 18766
rect 12624 18702 12676 18708
rect 12728 17202 12756 22374
rect 12808 21888 12860 21894
rect 12808 21830 12860 21836
rect 12820 21350 12848 21830
rect 12808 21344 12860 21350
rect 12808 21286 12860 21292
rect 12820 17746 12848 21286
rect 12808 17740 12860 17746
rect 12808 17682 12860 17688
rect 12912 17270 12940 22374
rect 13004 22234 13032 23666
rect 12992 22228 13044 22234
rect 12992 22170 13044 22176
rect 12992 20936 13044 20942
rect 12992 20878 13044 20884
rect 13004 18834 13032 20878
rect 12992 18828 13044 18834
rect 12992 18770 13044 18776
rect 13004 18358 13032 18770
rect 12992 18352 13044 18358
rect 12992 18294 13044 18300
rect 12900 17264 12952 17270
rect 12900 17206 12952 17212
rect 12716 17196 12768 17202
rect 12716 17138 12768 17144
rect 12532 13388 12584 13394
rect 12532 13330 12584 13336
rect 12544 9654 12572 13330
rect 12728 11898 12756 17138
rect 13188 15910 13216 30534
rect 13280 30326 13308 31214
rect 13372 30734 13400 31282
rect 13648 30938 13676 31418
rect 13636 30932 13688 30938
rect 13636 30874 13688 30880
rect 13360 30728 13412 30734
rect 13360 30670 13412 30676
rect 13268 30320 13320 30326
rect 13268 30262 13320 30268
rect 13280 29714 13308 30262
rect 13268 29708 13320 29714
rect 13268 29650 13320 29656
rect 13280 29170 13308 29650
rect 13268 29164 13320 29170
rect 13268 29106 13320 29112
rect 13268 26036 13320 26042
rect 13268 25978 13320 25984
rect 13280 25702 13308 25978
rect 13544 25900 13596 25906
rect 13544 25842 13596 25848
rect 13268 25696 13320 25702
rect 13268 25638 13320 25644
rect 13268 24812 13320 24818
rect 13556 24800 13584 25842
rect 13636 25832 13688 25838
rect 13740 25820 13768 32710
rect 13924 32450 13952 34478
rect 14200 34066 14228 34478
rect 14188 34060 14240 34066
rect 14188 34002 14240 34008
rect 14200 32910 14228 34002
rect 14280 33312 14332 33318
rect 14280 33254 14332 33260
rect 14188 32904 14240 32910
rect 14188 32846 14240 32852
rect 13832 32434 13952 32450
rect 13820 32428 13952 32434
rect 13872 32422 13952 32428
rect 13820 32370 13872 32376
rect 14292 32298 14320 33254
rect 14280 32292 14332 32298
rect 14280 32234 14332 32240
rect 14280 31816 14332 31822
rect 14280 31758 14332 31764
rect 14292 31142 14320 31758
rect 14280 31136 14332 31142
rect 14280 31078 14332 31084
rect 14384 30870 14412 36740
rect 14464 36722 14516 36728
rect 15200 36576 15252 36582
rect 15200 36518 15252 36524
rect 15212 36174 15240 36518
rect 15200 36168 15252 36174
rect 15200 36110 15252 36116
rect 15016 36032 15068 36038
rect 15016 35974 15068 35980
rect 14832 35692 14884 35698
rect 14832 35634 14884 35640
rect 14464 34604 14516 34610
rect 14464 34546 14516 34552
rect 14648 34604 14700 34610
rect 14648 34546 14700 34552
rect 14476 31482 14504 34546
rect 14660 34202 14688 34546
rect 14648 34196 14700 34202
rect 14648 34138 14700 34144
rect 14556 33516 14608 33522
rect 14556 33458 14608 33464
rect 14568 32570 14596 33458
rect 14740 32904 14792 32910
rect 14740 32846 14792 32852
rect 14556 32564 14608 32570
rect 14556 32506 14608 32512
rect 14752 32434 14780 32846
rect 14740 32428 14792 32434
rect 14740 32370 14792 32376
rect 14844 31754 14872 35634
rect 14752 31726 14872 31754
rect 14924 31748 14976 31754
rect 14464 31476 14516 31482
rect 14464 31418 14516 31424
rect 14464 31340 14516 31346
rect 14464 31282 14516 31288
rect 14476 31210 14504 31282
rect 14464 31204 14516 31210
rect 14464 31146 14516 31152
rect 14372 30864 14424 30870
rect 14372 30806 14424 30812
rect 14372 30728 14424 30734
rect 14372 30670 14424 30676
rect 14384 30394 14412 30670
rect 14372 30388 14424 30394
rect 14372 30330 14424 30336
rect 14372 30252 14424 30258
rect 14372 30194 14424 30200
rect 14188 30184 14240 30190
rect 14188 30126 14240 30132
rect 14200 29850 14228 30126
rect 14188 29844 14240 29850
rect 14188 29786 14240 29792
rect 14280 29640 14332 29646
rect 14280 29582 14332 29588
rect 14096 29164 14148 29170
rect 14096 29106 14148 29112
rect 14108 28762 14136 29106
rect 14096 28756 14148 28762
rect 14096 28698 14148 28704
rect 14188 27328 14240 27334
rect 14188 27270 14240 27276
rect 14200 27062 14228 27270
rect 14188 27056 14240 27062
rect 14188 26998 14240 27004
rect 14096 26784 14148 26790
rect 14096 26726 14148 26732
rect 14108 26382 14136 26726
rect 14096 26376 14148 26382
rect 14096 26318 14148 26324
rect 13688 25792 13768 25820
rect 13636 25774 13688 25780
rect 14200 25226 14228 26998
rect 14292 26790 14320 29582
rect 14384 28914 14412 30194
rect 14476 28966 14504 28997
rect 14464 28960 14516 28966
rect 14384 28908 14464 28914
rect 14384 28902 14516 28908
rect 14384 28886 14504 28902
rect 14476 28626 14504 28886
rect 14464 28620 14516 28626
rect 14464 28562 14516 28568
rect 14556 27056 14608 27062
rect 14556 26998 14608 27004
rect 14280 26784 14332 26790
rect 14280 26726 14332 26732
rect 14372 26376 14424 26382
rect 14372 26318 14424 26324
rect 14280 26240 14332 26246
rect 14280 26182 14332 26188
rect 14292 25498 14320 26182
rect 14280 25492 14332 25498
rect 14280 25434 14332 25440
rect 14188 25220 14240 25226
rect 14188 25162 14240 25168
rect 13728 24812 13780 24818
rect 13556 24772 13728 24800
rect 13268 24754 13320 24760
rect 13728 24754 13780 24760
rect 13280 24410 13308 24754
rect 13360 24744 13412 24750
rect 13360 24686 13412 24692
rect 13268 24404 13320 24410
rect 13268 24346 13320 24352
rect 13176 15904 13228 15910
rect 13176 15846 13228 15852
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 13084 11212 13136 11218
rect 13084 11154 13136 11160
rect 12532 9648 12584 9654
rect 12532 9590 12584 9596
rect 12452 7534 13032 7562
rect 11336 4140 11388 4146
rect 11336 4082 11388 4088
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 12164 3936 12216 3942
rect 12164 3878 12216 3884
rect 10508 3732 10560 3738
rect 10508 3674 10560 3680
rect 11612 3596 11664 3602
rect 11612 3538 11664 3544
rect 10968 2984 11020 2990
rect 10968 2926 11020 2932
rect 10980 800 11008 2926
rect 11624 800 11652 3538
rect 11716 2378 11744 3878
rect 11796 3528 11848 3534
rect 11796 3470 11848 3476
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 11808 2514 11836 3470
rect 11888 3392 11940 3398
rect 11888 3334 11940 3340
rect 11900 2938 11928 3334
rect 11992 3058 12020 3470
rect 12176 3126 12204 3878
rect 12624 3528 12676 3534
rect 12624 3470 12676 3476
rect 12164 3120 12216 3126
rect 12164 3062 12216 3068
rect 12256 3120 12308 3126
rect 12256 3062 12308 3068
rect 11980 3052 12032 3058
rect 11980 2994 12032 3000
rect 12268 2990 12296 3062
rect 12256 2984 12308 2990
rect 11900 2910 12020 2938
rect 12256 2926 12308 2932
rect 11992 2666 12020 2910
rect 12440 2916 12492 2922
rect 12440 2858 12492 2864
rect 12452 2666 12480 2858
rect 12636 2854 12664 3470
rect 12716 2984 12768 2990
rect 12716 2926 12768 2932
rect 12900 2984 12952 2990
rect 12900 2926 12952 2932
rect 12728 2854 12756 2926
rect 12624 2848 12676 2854
rect 12624 2790 12676 2796
rect 12716 2848 12768 2854
rect 12716 2790 12768 2796
rect 11992 2638 12480 2666
rect 11796 2508 11848 2514
rect 11796 2450 11848 2456
rect 12256 2508 12308 2514
rect 12256 2450 12308 2456
rect 11704 2372 11756 2378
rect 11704 2314 11756 2320
rect 12268 800 12296 2450
rect 12912 800 12940 2926
rect 13004 2774 13032 7534
rect 13096 3670 13124 11154
rect 13084 3664 13136 3670
rect 13084 3606 13136 3612
rect 13372 3602 13400 24686
rect 13452 24608 13504 24614
rect 13452 24550 13504 24556
rect 13544 24608 13596 24614
rect 13544 24550 13596 24556
rect 13464 24410 13492 24550
rect 13452 24404 13504 24410
rect 13452 24346 13504 24352
rect 13556 23526 13584 24550
rect 13740 24410 13768 24754
rect 14188 24744 14240 24750
rect 14188 24686 14240 24692
rect 13728 24404 13780 24410
rect 13728 24346 13780 24352
rect 13740 23526 13768 24346
rect 13912 24268 13964 24274
rect 13912 24210 13964 24216
rect 13924 23730 13952 24210
rect 14200 24206 14228 24686
rect 14188 24200 14240 24206
rect 14188 24142 14240 24148
rect 14292 24070 14320 25434
rect 14384 25226 14412 26318
rect 14568 25906 14596 26998
rect 14556 25900 14608 25906
rect 14556 25842 14608 25848
rect 14752 25786 14780 31726
rect 14924 31690 14976 31696
rect 14832 31680 14884 31686
rect 14832 31622 14884 31628
rect 14844 31346 14872 31622
rect 14832 31340 14884 31346
rect 14832 31282 14884 31288
rect 14844 29646 14872 31282
rect 14936 31210 14964 31690
rect 15028 31686 15056 35974
rect 15304 35834 15332 37130
rect 15844 36100 15896 36106
rect 15844 36042 15896 36048
rect 16028 36100 16080 36106
rect 16028 36042 16080 36048
rect 15292 35828 15344 35834
rect 15292 35770 15344 35776
rect 15856 35290 15884 36042
rect 16040 35630 16068 36042
rect 16028 35624 16080 35630
rect 16028 35566 16080 35572
rect 15844 35284 15896 35290
rect 15844 35226 15896 35232
rect 15108 35012 15160 35018
rect 15108 34954 15160 34960
rect 15120 34066 15148 34954
rect 16040 34542 16068 35566
rect 16028 34536 16080 34542
rect 16028 34478 16080 34484
rect 15660 34400 15712 34406
rect 15660 34342 15712 34348
rect 15108 34060 15160 34066
rect 15108 34002 15160 34008
rect 15120 32434 15148 34002
rect 15384 33992 15436 33998
rect 15384 33934 15436 33940
rect 15396 33318 15424 33934
rect 15384 33312 15436 33318
rect 15384 33254 15436 33260
rect 15396 32910 15424 33254
rect 15384 32904 15436 32910
rect 15384 32846 15436 32852
rect 15108 32428 15160 32434
rect 15108 32370 15160 32376
rect 15108 32224 15160 32230
rect 15108 32166 15160 32172
rect 15016 31680 15068 31686
rect 15016 31622 15068 31628
rect 15016 31340 15068 31346
rect 15120 31328 15148 32166
rect 15292 31952 15344 31958
rect 15292 31894 15344 31900
rect 15068 31300 15148 31328
rect 15200 31340 15252 31346
rect 15016 31282 15068 31288
rect 15200 31282 15252 31288
rect 14924 31204 14976 31210
rect 14924 31146 14976 31152
rect 14924 30864 14976 30870
rect 14924 30806 14976 30812
rect 14832 29640 14884 29646
rect 14832 29582 14884 29588
rect 14832 26512 14884 26518
rect 14832 26454 14884 26460
rect 14844 25906 14872 26454
rect 14832 25900 14884 25906
rect 14832 25842 14884 25848
rect 14752 25758 14872 25786
rect 14464 25696 14516 25702
rect 14464 25638 14516 25644
rect 14476 25498 14504 25638
rect 14554 25528 14610 25537
rect 14464 25492 14516 25498
rect 14554 25463 14556 25472
rect 14464 25434 14516 25440
rect 14608 25463 14610 25472
rect 14556 25434 14608 25440
rect 14372 25220 14424 25226
rect 14372 25162 14424 25168
rect 14384 24954 14412 25162
rect 14844 25158 14872 25758
rect 14832 25152 14884 25158
rect 14832 25094 14884 25100
rect 14372 24948 14424 24954
rect 14372 24890 14424 24896
rect 14648 24404 14700 24410
rect 14648 24346 14700 24352
rect 14280 24064 14332 24070
rect 14280 24006 14332 24012
rect 14660 23730 14688 24346
rect 13912 23724 13964 23730
rect 13912 23666 13964 23672
rect 14648 23724 14700 23730
rect 14648 23666 14700 23672
rect 13544 23520 13596 23526
rect 13544 23462 13596 23468
rect 13728 23520 13780 23526
rect 13728 23462 13780 23468
rect 14740 23520 14792 23526
rect 14740 23462 14792 23468
rect 13452 23112 13504 23118
rect 13452 23054 13504 23060
rect 13464 22642 13492 23054
rect 13452 22636 13504 22642
rect 13452 22578 13504 22584
rect 13464 21962 13492 22578
rect 13452 21956 13504 21962
rect 13452 21898 13504 21904
rect 13464 21622 13492 21898
rect 13452 21616 13504 21622
rect 13452 21558 13504 21564
rect 13556 21554 13584 23462
rect 13740 22710 13768 23462
rect 14188 23044 14240 23050
rect 14188 22986 14240 22992
rect 14200 22778 14228 22986
rect 14188 22772 14240 22778
rect 14188 22714 14240 22720
rect 14464 22772 14516 22778
rect 14464 22714 14516 22720
rect 13728 22704 13780 22710
rect 13728 22646 13780 22652
rect 14280 22704 14332 22710
rect 14280 22646 14332 22652
rect 13544 21548 13596 21554
rect 13544 21490 13596 21496
rect 13556 18766 13584 21490
rect 13636 19848 13688 19854
rect 13636 19790 13688 19796
rect 13544 18760 13596 18766
rect 13544 18702 13596 18708
rect 13648 17864 13676 19790
rect 13740 19378 13768 22646
rect 13820 21480 13872 21486
rect 13820 21422 13872 21428
rect 13832 19854 13860 21422
rect 13912 20868 13964 20874
rect 13912 20810 13964 20816
rect 13924 20602 13952 20810
rect 13912 20596 13964 20602
rect 13912 20538 13964 20544
rect 14188 20460 14240 20466
rect 14188 20402 14240 20408
rect 13820 19848 13872 19854
rect 13820 19790 13872 19796
rect 13728 19372 13780 19378
rect 13728 19314 13780 19320
rect 13832 18426 13860 19790
rect 13820 18420 13872 18426
rect 13820 18362 13872 18368
rect 13728 17876 13780 17882
rect 13648 17836 13728 17864
rect 13728 17818 13780 17824
rect 13740 17134 13768 17818
rect 13728 17128 13780 17134
rect 13728 17070 13780 17076
rect 14004 13252 14056 13258
rect 14004 13194 14056 13200
rect 14016 12986 14044 13194
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 14200 11150 14228 20402
rect 14292 20330 14320 22646
rect 14476 22642 14504 22714
rect 14554 22672 14610 22681
rect 14464 22636 14516 22642
rect 14554 22607 14610 22616
rect 14464 22578 14516 22584
rect 14568 20466 14596 22607
rect 14752 21622 14780 23462
rect 14740 21616 14792 21622
rect 14740 21558 14792 21564
rect 14844 20602 14872 25094
rect 14936 22094 14964 30806
rect 15028 29646 15056 31282
rect 15212 30938 15240 31282
rect 15200 30932 15252 30938
rect 15200 30874 15252 30880
rect 15304 30870 15332 31894
rect 15292 30864 15344 30870
rect 15292 30806 15344 30812
rect 15200 30048 15252 30054
rect 15200 29990 15252 29996
rect 15108 29844 15160 29850
rect 15108 29786 15160 29792
rect 15120 29714 15148 29786
rect 15108 29708 15160 29714
rect 15108 29650 15160 29656
rect 15016 29640 15068 29646
rect 15016 29582 15068 29588
rect 15120 29152 15148 29650
rect 15028 29124 15148 29152
rect 15028 28966 15056 29124
rect 15108 29028 15160 29034
rect 15108 28970 15160 28976
rect 15016 28960 15068 28966
rect 15016 28902 15068 28908
rect 15028 28558 15056 28902
rect 15016 28552 15068 28558
rect 15016 28494 15068 28500
rect 15120 27402 15148 28970
rect 15212 28490 15240 29990
rect 15304 29238 15332 30806
rect 15292 29232 15344 29238
rect 15292 29174 15344 29180
rect 15200 28484 15252 28490
rect 15200 28426 15252 28432
rect 15200 28008 15252 28014
rect 15200 27950 15252 27956
rect 15108 27396 15160 27402
rect 15108 27338 15160 27344
rect 15212 27334 15240 27950
rect 15200 27328 15252 27334
rect 15200 27270 15252 27276
rect 15016 26920 15068 26926
rect 15016 26862 15068 26868
rect 15028 26314 15056 26862
rect 15108 26784 15160 26790
rect 15108 26726 15160 26732
rect 15016 26308 15068 26314
rect 15016 26250 15068 26256
rect 15120 26234 15148 26726
rect 15212 26382 15240 27270
rect 15396 27130 15424 32846
rect 15568 29640 15620 29646
rect 15568 29582 15620 29588
rect 15476 29504 15528 29510
rect 15476 29446 15528 29452
rect 15488 29238 15516 29446
rect 15476 29232 15528 29238
rect 15476 29174 15528 29180
rect 15580 29102 15608 29582
rect 15568 29096 15620 29102
rect 15568 29038 15620 29044
rect 15580 28082 15608 29038
rect 15672 28762 15700 34342
rect 16040 34066 16068 34478
rect 16028 34060 16080 34066
rect 16028 34002 16080 34008
rect 16040 33590 16068 34002
rect 16028 33584 16080 33590
rect 16028 33526 16080 33532
rect 16040 32434 16068 33526
rect 16028 32428 16080 32434
rect 16028 32370 16080 32376
rect 16028 31340 16080 31346
rect 16028 31282 16080 31288
rect 16040 30258 16068 31282
rect 16028 30252 16080 30258
rect 16028 30194 16080 30200
rect 15936 29844 15988 29850
rect 15936 29786 15988 29792
rect 15948 29170 15976 29786
rect 16040 29646 16068 30194
rect 16028 29640 16080 29646
rect 16028 29582 16080 29588
rect 15752 29164 15804 29170
rect 15936 29164 15988 29170
rect 15804 29124 15884 29152
rect 15752 29106 15804 29112
rect 15660 28756 15712 28762
rect 15660 28698 15712 28704
rect 15856 28558 15884 29124
rect 15936 29106 15988 29112
rect 15844 28552 15896 28558
rect 15844 28494 15896 28500
rect 16028 28552 16080 28558
rect 16028 28494 16080 28500
rect 15568 28076 15620 28082
rect 15568 28018 15620 28024
rect 15384 27124 15436 27130
rect 15384 27066 15436 27072
rect 15200 26376 15252 26382
rect 15200 26318 15252 26324
rect 15292 26376 15344 26382
rect 15292 26318 15344 26324
rect 15304 26234 15332 26318
rect 15396 26314 15424 27066
rect 15384 26308 15436 26314
rect 15384 26250 15436 26256
rect 15120 26206 15332 26234
rect 15120 24614 15148 26206
rect 15108 24608 15160 24614
rect 15108 24550 15160 24556
rect 15108 23656 15160 23662
rect 15108 23598 15160 23604
rect 15120 23254 15148 23598
rect 15108 23248 15160 23254
rect 15108 23190 15160 23196
rect 15568 23044 15620 23050
rect 15568 22986 15620 22992
rect 15580 22778 15608 22986
rect 15568 22772 15620 22778
rect 15568 22714 15620 22720
rect 15752 22772 15804 22778
rect 15752 22714 15804 22720
rect 15014 22672 15070 22681
rect 15764 22642 15792 22714
rect 15014 22607 15016 22616
rect 15068 22607 15070 22616
rect 15752 22636 15804 22642
rect 15016 22578 15068 22584
rect 15752 22578 15804 22584
rect 14936 22066 15056 22094
rect 14832 20596 14884 20602
rect 14832 20538 14884 20544
rect 14556 20460 14608 20466
rect 14556 20402 14608 20408
rect 14280 20324 14332 20330
rect 14280 20266 14332 20272
rect 14372 19780 14424 19786
rect 14372 19722 14424 19728
rect 14384 18902 14412 19722
rect 14464 19304 14516 19310
rect 14464 19246 14516 19252
rect 14372 18896 14424 18902
rect 14372 18838 14424 18844
rect 14384 18358 14412 18838
rect 14476 18766 14504 19246
rect 14648 19168 14700 19174
rect 14648 19110 14700 19116
rect 14464 18760 14516 18766
rect 14464 18702 14516 18708
rect 14372 18352 14424 18358
rect 14372 18294 14424 18300
rect 14384 17762 14412 18294
rect 14476 18222 14504 18702
rect 14660 18290 14688 19110
rect 14648 18284 14700 18290
rect 14648 18226 14700 18232
rect 14924 18284 14976 18290
rect 14924 18226 14976 18232
rect 14464 18216 14516 18222
rect 14936 18193 14964 18226
rect 14464 18158 14516 18164
rect 14922 18184 14978 18193
rect 14292 17734 14412 17762
rect 14476 17746 14504 18158
rect 14922 18119 14978 18128
rect 14924 18080 14976 18086
rect 14924 18022 14976 18028
rect 14646 17912 14702 17921
rect 14646 17847 14702 17856
rect 14660 17814 14688 17847
rect 14648 17808 14700 17814
rect 14648 17750 14700 17756
rect 14464 17740 14516 17746
rect 14292 16998 14320 17734
rect 14464 17682 14516 17688
rect 14372 17672 14424 17678
rect 14372 17614 14424 17620
rect 14280 16992 14332 16998
rect 14280 16934 14332 16940
rect 14292 16182 14320 16934
rect 14384 16658 14412 17614
rect 14476 17270 14504 17682
rect 14936 17610 14964 18022
rect 15028 17610 15056 22066
rect 15568 21140 15620 21146
rect 15568 21082 15620 21088
rect 15580 20806 15608 21082
rect 15568 20800 15620 20806
rect 15568 20742 15620 20748
rect 15108 19712 15160 19718
rect 15108 19654 15160 19660
rect 15120 19378 15148 19654
rect 15108 19372 15160 19378
rect 15108 19314 15160 19320
rect 15292 19372 15344 19378
rect 15292 19314 15344 19320
rect 15304 18766 15332 19314
rect 15580 19242 15608 20742
rect 15568 19236 15620 19242
rect 15568 19178 15620 19184
rect 15292 18760 15344 18766
rect 15292 18702 15344 18708
rect 15304 18290 15332 18702
rect 15856 18290 15884 28494
rect 16040 28218 16068 28494
rect 16028 28212 16080 28218
rect 16028 28154 16080 28160
rect 15936 22636 15988 22642
rect 15936 22578 15988 22584
rect 15948 22234 15976 22578
rect 15936 22228 15988 22234
rect 15936 22170 15988 22176
rect 16132 22094 16160 38286
rect 16224 22778 16252 48282
rect 16592 48210 16620 49166
rect 16776 48770 16804 51200
rect 16776 48742 17264 48770
rect 17236 48686 17264 48742
rect 16948 48680 17000 48686
rect 16948 48622 17000 48628
rect 17224 48680 17276 48686
rect 17224 48622 17276 48628
rect 16960 48278 16988 48622
rect 16948 48272 17000 48278
rect 16948 48214 17000 48220
rect 17420 48210 17448 51200
rect 18064 49298 18092 51200
rect 18052 49292 18104 49298
rect 18052 49234 18104 49240
rect 19444 49230 19472 51326
rect 19982 51326 20116 51354
rect 19982 51200 20038 51326
rect 20088 49230 20116 51326
rect 20626 51200 20682 52000
rect 21270 51200 21326 52000
rect 21914 51354 21970 52000
rect 21914 51326 22048 51354
rect 21914 51200 21970 51326
rect 20444 49428 20496 49434
rect 20444 49370 20496 49376
rect 19432 49224 19484 49230
rect 19432 49166 19484 49172
rect 20076 49224 20128 49230
rect 20076 49166 20128 49172
rect 19574 48988 19882 49008
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48912 19882 48932
rect 19432 48680 19484 48686
rect 19432 48622 19484 48628
rect 19340 48612 19392 48618
rect 19340 48554 19392 48560
rect 17960 48544 18012 48550
rect 17960 48486 18012 48492
rect 16580 48204 16632 48210
rect 16580 48146 16632 48152
rect 17408 48204 17460 48210
rect 17408 48146 17460 48152
rect 17972 47802 18000 48486
rect 19352 48278 19380 48554
rect 19340 48272 19392 48278
rect 19340 48214 19392 48220
rect 19444 47802 19472 48622
rect 20076 48136 20128 48142
rect 20076 48078 20128 48084
rect 19574 47900 19882 47920
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47824 19882 47844
rect 17960 47796 18012 47802
rect 17960 47738 18012 47744
rect 19432 47796 19484 47802
rect 19432 47738 19484 47744
rect 18420 47728 18472 47734
rect 18420 47670 18472 47676
rect 20088 47682 20116 48078
rect 20168 48068 20220 48074
rect 20168 48010 20220 48016
rect 20180 47802 20208 48010
rect 20260 48000 20312 48006
rect 20260 47942 20312 47948
rect 20352 48000 20404 48006
rect 20352 47942 20404 47948
rect 20272 47802 20300 47942
rect 20168 47796 20220 47802
rect 20168 47738 20220 47744
rect 20260 47796 20312 47802
rect 20260 47738 20312 47744
rect 20364 47682 20392 47942
rect 16948 47592 17000 47598
rect 16948 47534 17000 47540
rect 16960 47258 16988 47534
rect 16948 47252 17000 47258
rect 16948 47194 17000 47200
rect 18052 47252 18104 47258
rect 18052 47194 18104 47200
rect 17868 47184 17920 47190
rect 17868 47126 17920 47132
rect 17224 39296 17276 39302
rect 17224 39238 17276 39244
rect 17236 38962 17264 39238
rect 17224 38956 17276 38962
rect 17224 38898 17276 38904
rect 17236 37874 17264 38898
rect 17408 38276 17460 38282
rect 17408 38218 17460 38224
rect 17224 37868 17276 37874
rect 17224 37810 17276 37816
rect 17236 37262 17264 37810
rect 17420 37806 17448 38218
rect 17408 37800 17460 37806
rect 17408 37742 17460 37748
rect 17420 37398 17448 37742
rect 17408 37392 17460 37398
rect 17460 37352 17540 37380
rect 17408 37334 17460 37340
rect 17224 37256 17276 37262
rect 17224 37198 17276 37204
rect 16488 36848 16540 36854
rect 16488 36790 16540 36796
rect 16500 36378 16528 36790
rect 17236 36786 17264 37198
rect 17224 36780 17276 36786
rect 17224 36722 17276 36728
rect 16856 36712 16908 36718
rect 16856 36654 16908 36660
rect 16488 36372 16540 36378
rect 16488 36314 16540 36320
rect 16500 35766 16528 36314
rect 16488 35760 16540 35766
rect 16488 35702 16540 35708
rect 16764 35692 16816 35698
rect 16764 35634 16816 35640
rect 16304 35488 16356 35494
rect 16304 35430 16356 35436
rect 16316 35086 16344 35430
rect 16776 35086 16804 35634
rect 16304 35080 16356 35086
rect 16304 35022 16356 35028
rect 16764 35080 16816 35086
rect 16764 35022 16816 35028
rect 16776 33522 16804 35022
rect 16764 33516 16816 33522
rect 16764 33458 16816 33464
rect 16580 31748 16632 31754
rect 16580 31690 16632 31696
rect 16672 31748 16724 31754
rect 16672 31690 16724 31696
rect 16592 30870 16620 31690
rect 16684 31414 16712 31690
rect 16776 31414 16804 33458
rect 16672 31408 16724 31414
rect 16672 31350 16724 31356
rect 16764 31408 16816 31414
rect 16764 31350 16816 31356
rect 16776 30938 16804 31350
rect 16764 30932 16816 30938
rect 16764 30874 16816 30880
rect 16580 30864 16632 30870
rect 16580 30806 16632 30812
rect 16776 30734 16804 30874
rect 16672 30728 16724 30734
rect 16672 30670 16724 30676
rect 16764 30728 16816 30734
rect 16764 30670 16816 30676
rect 16684 30190 16712 30670
rect 16672 30184 16724 30190
rect 16672 30126 16724 30132
rect 16580 29844 16632 29850
rect 16580 29786 16632 29792
rect 16488 29708 16540 29714
rect 16488 29650 16540 29656
rect 16500 29102 16528 29650
rect 16592 29306 16620 29786
rect 16684 29306 16712 30126
rect 16764 30048 16816 30054
rect 16764 29990 16816 29996
rect 16580 29300 16632 29306
rect 16580 29242 16632 29248
rect 16672 29300 16724 29306
rect 16672 29242 16724 29248
rect 16488 29096 16540 29102
rect 16488 29038 16540 29044
rect 16488 28960 16540 28966
rect 16488 28902 16540 28908
rect 16500 28558 16528 28902
rect 16488 28552 16540 28558
rect 16488 28494 16540 28500
rect 16500 27470 16528 28494
rect 16488 27464 16540 27470
rect 16488 27406 16540 27412
rect 16672 25832 16724 25838
rect 16672 25774 16724 25780
rect 16684 25294 16712 25774
rect 16580 25288 16632 25294
rect 16580 25230 16632 25236
rect 16672 25288 16724 25294
rect 16672 25230 16724 25236
rect 16592 24954 16620 25230
rect 16580 24948 16632 24954
rect 16580 24890 16632 24896
rect 16212 22772 16264 22778
rect 16212 22714 16264 22720
rect 16210 22672 16266 22681
rect 16210 22607 16212 22616
rect 16264 22607 16266 22616
rect 16212 22578 16264 22584
rect 16224 22234 16252 22578
rect 16212 22228 16264 22234
rect 16212 22170 16264 22176
rect 16040 22066 16160 22094
rect 15936 20936 15988 20942
rect 15936 20878 15988 20884
rect 15948 19514 15976 20878
rect 15936 19508 15988 19514
rect 15936 19450 15988 19456
rect 16040 18358 16068 22066
rect 16776 20482 16804 29990
rect 16868 24177 16896 36654
rect 17408 36168 17460 36174
rect 17408 36110 17460 36116
rect 17040 36100 17092 36106
rect 17040 36042 17092 36048
rect 16948 36032 17000 36038
rect 16948 35974 17000 35980
rect 16960 35766 16988 35974
rect 16948 35760 17000 35766
rect 16948 35702 17000 35708
rect 17052 34950 17080 36042
rect 17420 35290 17448 36110
rect 17408 35284 17460 35290
rect 17408 35226 17460 35232
rect 17040 34944 17092 34950
rect 17040 34886 17092 34892
rect 17052 34610 17080 34886
rect 17040 34604 17092 34610
rect 17040 34546 17092 34552
rect 17224 34604 17276 34610
rect 17224 34546 17276 34552
rect 17052 31686 17080 34546
rect 17236 33658 17264 34546
rect 17316 34400 17368 34406
rect 17316 34342 17368 34348
rect 17328 34066 17356 34342
rect 17316 34060 17368 34066
rect 17316 34002 17368 34008
rect 17224 33652 17276 33658
rect 17224 33594 17276 33600
rect 17224 32428 17276 32434
rect 17224 32370 17276 32376
rect 17236 32026 17264 32370
rect 17224 32020 17276 32026
rect 17224 31962 17276 31968
rect 17316 32020 17368 32026
rect 17316 31962 17368 31968
rect 17328 31906 17356 31962
rect 17236 31878 17356 31906
rect 17236 31754 17264 31878
rect 17512 31754 17540 37352
rect 17880 36718 17908 47126
rect 17868 36712 17920 36718
rect 17868 36654 17920 36660
rect 17592 36168 17644 36174
rect 17592 36110 17644 36116
rect 17604 35018 17632 36110
rect 17960 35828 18012 35834
rect 17960 35770 18012 35776
rect 17972 35086 18000 35770
rect 17960 35080 18012 35086
rect 17960 35022 18012 35028
rect 17592 35012 17644 35018
rect 17592 34954 17644 34960
rect 17604 34542 17632 34954
rect 17960 34604 18012 34610
rect 17960 34546 18012 34552
rect 17592 34536 17644 34542
rect 17592 34478 17644 34484
rect 17972 32570 18000 34546
rect 17960 32564 18012 32570
rect 17960 32506 18012 32512
rect 17144 31726 17264 31754
rect 17316 31748 17368 31754
rect 17040 31680 17092 31686
rect 17040 31622 17092 31628
rect 17052 31346 17080 31622
rect 17040 31340 17092 31346
rect 17040 31282 17092 31288
rect 17052 30258 17080 31282
rect 17040 30252 17092 30258
rect 17040 30194 17092 30200
rect 17144 30054 17172 31726
rect 17316 31690 17368 31696
rect 17420 31726 17540 31754
rect 17224 31340 17276 31346
rect 17328 31328 17356 31690
rect 17276 31300 17356 31328
rect 17224 31282 17276 31288
rect 17236 30598 17264 31282
rect 17224 30592 17276 30598
rect 17224 30534 17276 30540
rect 17132 30048 17184 30054
rect 17132 29990 17184 29996
rect 17236 29850 17264 30534
rect 17224 29844 17276 29850
rect 17224 29786 17276 29792
rect 17420 29730 17448 31726
rect 17684 31204 17736 31210
rect 17684 31146 17736 31152
rect 17500 30184 17552 30190
rect 17500 30126 17552 30132
rect 17052 29702 17448 29730
rect 17052 27674 17080 29702
rect 17132 29640 17184 29646
rect 17132 29582 17184 29588
rect 17144 29170 17172 29582
rect 17224 29504 17276 29510
rect 17408 29504 17460 29510
rect 17276 29464 17356 29492
rect 17224 29446 17276 29452
rect 17328 29306 17356 29464
rect 17512 29492 17540 30126
rect 17696 29646 17724 31146
rect 17972 30734 18000 32506
rect 17960 30728 18012 30734
rect 17960 30670 18012 30676
rect 17776 29776 17828 29782
rect 17776 29718 17828 29724
rect 17592 29640 17644 29646
rect 17592 29582 17644 29588
rect 17684 29640 17736 29646
rect 17684 29582 17736 29588
rect 17460 29464 17540 29492
rect 17408 29446 17460 29452
rect 17224 29300 17276 29306
rect 17224 29242 17276 29248
rect 17316 29300 17368 29306
rect 17316 29242 17368 29248
rect 17132 29164 17184 29170
rect 17132 29106 17184 29112
rect 17236 28490 17264 29242
rect 17224 28484 17276 28490
rect 17224 28426 17276 28432
rect 17040 27668 17092 27674
rect 17040 27610 17092 27616
rect 17420 27470 17448 29446
rect 17500 29232 17552 29238
rect 17500 29174 17552 29180
rect 17512 29102 17540 29174
rect 17500 29096 17552 29102
rect 17500 29038 17552 29044
rect 17512 28218 17540 29038
rect 17604 29034 17632 29582
rect 17788 29209 17816 29718
rect 17868 29504 17920 29510
rect 17868 29446 17920 29452
rect 17960 29504 18012 29510
rect 17960 29446 18012 29452
rect 17880 29238 17908 29446
rect 17868 29232 17920 29238
rect 17774 29200 17830 29209
rect 17684 29164 17736 29170
rect 17868 29174 17920 29180
rect 17774 29135 17776 29144
rect 17684 29106 17736 29112
rect 17828 29135 17830 29144
rect 17776 29106 17828 29112
rect 17592 29028 17644 29034
rect 17592 28970 17644 28976
rect 17604 28422 17632 28970
rect 17592 28416 17644 28422
rect 17592 28358 17644 28364
rect 17500 28212 17552 28218
rect 17500 28154 17552 28160
rect 17604 27878 17632 28358
rect 17696 28014 17724 29106
rect 17684 28008 17736 28014
rect 17684 27950 17736 27956
rect 17592 27872 17644 27878
rect 17592 27814 17644 27820
rect 17408 27464 17460 27470
rect 17408 27406 17460 27412
rect 17696 27334 17724 27950
rect 17788 27606 17816 29106
rect 17972 29102 18000 29446
rect 17960 29096 18012 29102
rect 17960 29038 18012 29044
rect 17776 27600 17828 27606
rect 17776 27542 17828 27548
rect 17684 27328 17736 27334
rect 17684 27270 17736 27276
rect 17590 26480 17646 26489
rect 17590 26415 17646 26424
rect 17604 26382 17632 26415
rect 17592 26376 17644 26382
rect 17592 26318 17644 26324
rect 17682 26344 17738 26353
rect 17682 26279 17738 26288
rect 16948 26240 17000 26246
rect 16948 26182 17000 26188
rect 16960 25906 16988 26182
rect 16948 25900 17000 25906
rect 16948 25842 17000 25848
rect 17040 25696 17092 25702
rect 17040 25638 17092 25644
rect 17052 25362 17080 25638
rect 17040 25356 17092 25362
rect 17040 25298 17092 25304
rect 17406 24848 17462 24857
rect 17696 24818 17724 26279
rect 18064 26042 18092 47194
rect 18236 47184 18288 47190
rect 18236 47126 18288 47132
rect 18248 46646 18276 47126
rect 18236 46640 18288 46646
rect 18236 46582 18288 46588
rect 18248 45966 18276 46582
rect 18432 45966 18460 47670
rect 19064 47660 19116 47666
rect 19064 47602 19116 47608
rect 19340 47660 19392 47666
rect 20088 47654 20392 47682
rect 19340 47602 19392 47608
rect 19076 47462 19104 47602
rect 19064 47456 19116 47462
rect 19064 47398 19116 47404
rect 18236 45960 18288 45966
rect 18236 45902 18288 45908
rect 18420 45960 18472 45966
rect 18420 45902 18472 45908
rect 18880 39908 18932 39914
rect 18880 39850 18932 39856
rect 18236 39432 18288 39438
rect 18236 39374 18288 39380
rect 18328 39432 18380 39438
rect 18328 39374 18380 39380
rect 18144 37188 18196 37194
rect 18144 37130 18196 37136
rect 18156 36310 18184 37130
rect 18144 36304 18196 36310
rect 18144 36246 18196 36252
rect 18144 36168 18196 36174
rect 18144 36110 18196 36116
rect 18156 31754 18184 36110
rect 18248 36106 18276 39374
rect 18340 38758 18368 39374
rect 18604 38956 18656 38962
rect 18604 38898 18656 38904
rect 18328 38752 18380 38758
rect 18328 38694 18380 38700
rect 18340 38214 18368 38694
rect 18328 38208 18380 38214
rect 18328 38150 18380 38156
rect 18236 36100 18288 36106
rect 18236 36042 18288 36048
rect 18340 32842 18368 38150
rect 18616 37874 18644 38898
rect 18892 38894 18920 39850
rect 18880 38888 18932 38894
rect 18880 38830 18932 38836
rect 18604 37868 18656 37874
rect 18604 37810 18656 37816
rect 18616 37262 18644 37810
rect 18604 37256 18656 37262
rect 18604 37198 18656 37204
rect 18616 36786 18644 37198
rect 18788 36848 18840 36854
rect 18788 36790 18840 36796
rect 18604 36780 18656 36786
rect 18604 36722 18656 36728
rect 18616 36378 18644 36722
rect 18604 36372 18656 36378
rect 18604 36314 18656 36320
rect 18420 35080 18472 35086
rect 18420 35022 18472 35028
rect 18328 32836 18380 32842
rect 18328 32778 18380 32784
rect 18328 31952 18380 31958
rect 18328 31894 18380 31900
rect 18156 31726 18276 31754
rect 18144 26512 18196 26518
rect 18144 26454 18196 26460
rect 18156 26353 18184 26454
rect 18142 26344 18198 26353
rect 18142 26279 18198 26288
rect 18144 26240 18196 26246
rect 18144 26182 18196 26188
rect 17960 26036 18012 26042
rect 17960 25978 18012 25984
rect 18052 26036 18104 26042
rect 18052 25978 18104 25984
rect 17972 25906 18000 25978
rect 17960 25900 18012 25906
rect 17960 25842 18012 25848
rect 18156 25838 18184 26182
rect 18144 25832 18196 25838
rect 18144 25774 18196 25780
rect 18052 25696 18104 25702
rect 18052 25638 18104 25644
rect 17958 25256 18014 25265
rect 17958 25191 18014 25200
rect 17972 25158 18000 25191
rect 17960 25152 18012 25158
rect 17960 25094 18012 25100
rect 17406 24783 17408 24792
rect 17460 24783 17462 24792
rect 17684 24812 17736 24818
rect 17408 24754 17460 24760
rect 17684 24754 17736 24760
rect 17420 24682 17448 24754
rect 18064 24682 18092 25638
rect 17408 24676 17460 24682
rect 17408 24618 17460 24624
rect 18052 24676 18104 24682
rect 18052 24618 18104 24624
rect 18156 24274 18184 25774
rect 18248 25362 18276 31726
rect 18340 31414 18368 31894
rect 18432 31754 18460 35022
rect 18604 33856 18656 33862
rect 18604 33798 18656 33804
rect 18616 33522 18644 33798
rect 18604 33516 18656 33522
rect 18604 33458 18656 33464
rect 18432 31726 18552 31754
rect 18328 31408 18380 31414
rect 18328 31350 18380 31356
rect 18420 30796 18472 30802
rect 18420 30738 18472 30744
rect 18328 29640 18380 29646
rect 18328 29582 18380 29588
rect 18340 28694 18368 29582
rect 18328 28688 18380 28694
rect 18328 28630 18380 28636
rect 18432 28150 18460 30738
rect 18420 28144 18472 28150
rect 18420 28086 18472 28092
rect 18524 26874 18552 31726
rect 18340 26846 18552 26874
rect 18236 25356 18288 25362
rect 18236 25298 18288 25304
rect 18236 25152 18288 25158
rect 18236 25094 18288 25100
rect 18248 24886 18276 25094
rect 18236 24880 18288 24886
rect 18236 24822 18288 24828
rect 18144 24268 18196 24274
rect 18144 24210 18196 24216
rect 16948 24200 17000 24206
rect 16854 24168 16910 24177
rect 16948 24142 17000 24148
rect 17868 24200 17920 24206
rect 17868 24142 17920 24148
rect 16854 24103 16910 24112
rect 16868 23526 16896 24103
rect 16856 23520 16908 23526
rect 16856 23462 16908 23468
rect 16960 23254 16988 24142
rect 17592 24064 17644 24070
rect 17592 24006 17644 24012
rect 17604 23798 17632 24006
rect 17592 23792 17644 23798
rect 17592 23734 17644 23740
rect 17604 23662 17632 23734
rect 17592 23656 17644 23662
rect 17592 23598 17644 23604
rect 16948 23248 17000 23254
rect 16948 23190 17000 23196
rect 16960 21962 16988 23190
rect 17040 23112 17092 23118
rect 17040 23054 17092 23060
rect 17052 22642 17080 23054
rect 17040 22636 17092 22642
rect 17040 22578 17092 22584
rect 16948 21956 17000 21962
rect 16948 21898 17000 21904
rect 16856 20868 16908 20874
rect 16856 20810 16908 20816
rect 16868 20602 16896 20810
rect 16856 20596 16908 20602
rect 16856 20538 16908 20544
rect 16580 20460 16632 20466
rect 16776 20454 16896 20482
rect 16580 20402 16632 20408
rect 16592 19310 16620 20402
rect 16764 19440 16816 19446
rect 16764 19382 16816 19388
rect 16672 19372 16724 19378
rect 16672 19314 16724 19320
rect 16580 19304 16632 19310
rect 16580 19246 16632 19252
rect 16592 18358 16620 19246
rect 16684 18834 16712 19314
rect 16672 18828 16724 18834
rect 16672 18770 16724 18776
rect 16672 18692 16724 18698
rect 16672 18634 16724 18640
rect 16684 18426 16712 18634
rect 16672 18420 16724 18426
rect 16672 18362 16724 18368
rect 16028 18352 16080 18358
rect 16028 18294 16080 18300
rect 16580 18352 16632 18358
rect 16580 18294 16632 18300
rect 15292 18284 15344 18290
rect 15292 18226 15344 18232
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 14924 17604 14976 17610
rect 14924 17546 14976 17552
rect 15016 17604 15068 17610
rect 15016 17546 15068 17552
rect 15304 17338 15332 18226
rect 16040 17882 16068 18294
rect 16028 17876 16080 17882
rect 16028 17818 16080 17824
rect 16120 17876 16172 17882
rect 16120 17818 16172 17824
rect 15382 17640 15438 17649
rect 16132 17610 16160 17818
rect 16776 17814 16804 19382
rect 16764 17808 16816 17814
rect 16764 17750 16816 17756
rect 15382 17575 15438 17584
rect 16120 17604 16172 17610
rect 15292 17332 15344 17338
rect 15292 17274 15344 17280
rect 14464 17264 14516 17270
rect 14464 17206 14516 17212
rect 15396 17202 15424 17575
rect 16120 17546 16172 17552
rect 16580 17604 16632 17610
rect 16580 17546 16632 17552
rect 16026 17368 16082 17377
rect 15936 17332 15988 17338
rect 16026 17303 16082 17312
rect 15936 17274 15988 17280
rect 15948 17202 15976 17274
rect 16040 17270 16068 17303
rect 16028 17264 16080 17270
rect 16028 17206 16080 17212
rect 15384 17196 15436 17202
rect 15384 17138 15436 17144
rect 15936 17196 15988 17202
rect 15936 17138 15988 17144
rect 15384 17060 15436 17066
rect 15384 17002 15436 17008
rect 15844 17060 15896 17066
rect 15844 17002 15896 17008
rect 15200 16992 15252 16998
rect 15200 16934 15252 16940
rect 14372 16652 14424 16658
rect 14372 16594 14424 16600
rect 15212 16590 15240 16934
rect 15200 16584 15252 16590
rect 15200 16526 15252 16532
rect 15396 16182 15424 17002
rect 15476 16992 15528 16998
rect 15476 16934 15528 16940
rect 14280 16176 14332 16182
rect 14280 16118 14332 16124
rect 15384 16176 15436 16182
rect 15384 16118 15436 16124
rect 15488 12850 15516 16934
rect 15856 16250 15884 17002
rect 16592 16794 16620 17546
rect 16580 16788 16632 16794
rect 16580 16730 16632 16736
rect 16672 16448 16724 16454
rect 16672 16390 16724 16396
rect 15844 16244 15896 16250
rect 15844 16186 15896 16192
rect 16684 16114 16712 16390
rect 16672 16108 16724 16114
rect 16672 16050 16724 16056
rect 16868 15994 16896 20454
rect 16960 17649 16988 21898
rect 17052 21010 17080 22578
rect 17604 22030 17632 23598
rect 17684 23520 17736 23526
rect 17684 23462 17736 23468
rect 17592 22024 17644 22030
rect 17592 21966 17644 21972
rect 17500 21888 17552 21894
rect 17500 21830 17552 21836
rect 17040 21004 17092 21010
rect 17040 20946 17092 20952
rect 17052 19514 17080 20946
rect 17132 20460 17184 20466
rect 17132 20402 17184 20408
rect 17040 19508 17092 19514
rect 17040 19450 17092 19456
rect 17040 17740 17092 17746
rect 17040 17682 17092 17688
rect 16946 17640 17002 17649
rect 16946 17575 17002 17584
rect 16684 15966 16896 15994
rect 15476 12844 15528 12850
rect 15476 12786 15528 12792
rect 14188 11144 14240 11150
rect 14188 11086 14240 11092
rect 16684 7750 16712 15966
rect 17052 11558 17080 17682
rect 17040 11552 17092 11558
rect 17040 11494 17092 11500
rect 16672 7744 16724 7750
rect 16672 7686 16724 7692
rect 17144 4826 17172 20402
rect 17316 19848 17368 19854
rect 17316 19790 17368 19796
rect 17328 18766 17356 19790
rect 17512 19700 17540 21830
rect 17592 20256 17644 20262
rect 17592 20198 17644 20204
rect 17604 19854 17632 20198
rect 17592 19848 17644 19854
rect 17592 19790 17644 19796
rect 17512 19672 17632 19700
rect 17316 18760 17368 18766
rect 17316 18702 17368 18708
rect 17224 18692 17276 18698
rect 17224 18634 17276 18640
rect 17236 18290 17264 18634
rect 17224 18284 17276 18290
rect 17224 18226 17276 18232
rect 17224 18148 17276 18154
rect 17224 18090 17276 18096
rect 17236 14260 17264 18090
rect 17328 17678 17356 18702
rect 17408 18216 17460 18222
rect 17406 18184 17408 18193
rect 17460 18184 17462 18193
rect 17406 18119 17462 18128
rect 17500 18080 17552 18086
rect 17500 18022 17552 18028
rect 17512 17678 17540 18022
rect 17316 17672 17368 17678
rect 17500 17672 17552 17678
rect 17368 17632 17448 17660
rect 17316 17614 17368 17620
rect 17420 17134 17448 17632
rect 17500 17614 17552 17620
rect 17408 17128 17460 17134
rect 17408 17070 17460 17076
rect 17420 16726 17448 17070
rect 17408 16720 17460 16726
rect 17408 16662 17460 16668
rect 17604 14278 17632 19672
rect 17696 17218 17724 23462
rect 17776 22976 17828 22982
rect 17776 22918 17828 22924
rect 17788 22642 17816 22918
rect 17776 22636 17828 22642
rect 17776 22578 17828 22584
rect 17880 22438 17908 24142
rect 17960 23588 18012 23594
rect 17960 23530 18012 23536
rect 17972 23050 18000 23530
rect 18236 23112 18288 23118
rect 18236 23054 18288 23060
rect 17960 23044 18012 23050
rect 17960 22986 18012 22992
rect 17868 22432 17920 22438
rect 17868 22374 17920 22380
rect 18248 22234 18276 23054
rect 18236 22228 18288 22234
rect 18236 22170 18288 22176
rect 18052 21956 18104 21962
rect 18052 21898 18104 21904
rect 18064 21622 18092 21898
rect 18052 21616 18104 21622
rect 18052 21558 18104 21564
rect 18144 21344 18196 21350
rect 18144 21286 18196 21292
rect 18156 20534 18184 21286
rect 18144 20528 18196 20534
rect 18144 20470 18196 20476
rect 18236 20460 18288 20466
rect 18236 20402 18288 20408
rect 17868 19848 17920 19854
rect 17868 19790 17920 19796
rect 17880 19514 17908 19790
rect 17868 19508 17920 19514
rect 17868 19450 17920 19456
rect 17776 18624 17828 18630
rect 17776 18566 17828 18572
rect 17788 18426 17816 18566
rect 17776 18420 17828 18426
rect 17776 18362 17828 18368
rect 17696 17190 17816 17218
rect 17684 16788 17736 16794
rect 17684 16730 17736 16736
rect 17696 15094 17724 16730
rect 17684 15088 17736 15094
rect 17684 15030 17736 15036
rect 17316 14272 17368 14278
rect 17236 14232 17316 14260
rect 17316 14214 17368 14220
rect 17408 14272 17460 14278
rect 17408 14214 17460 14220
rect 17592 14272 17644 14278
rect 17592 14214 17644 14220
rect 17224 13728 17276 13734
rect 17224 13670 17276 13676
rect 17236 13258 17264 13670
rect 17224 13252 17276 13258
rect 17224 13194 17276 13200
rect 17328 13190 17356 14214
rect 17420 13938 17448 14214
rect 17408 13932 17460 13938
rect 17408 13874 17460 13880
rect 17500 13932 17552 13938
rect 17500 13874 17552 13880
rect 17316 13184 17368 13190
rect 17316 13126 17368 13132
rect 17132 4820 17184 4826
rect 17132 4762 17184 4768
rect 17512 4010 17540 13874
rect 17788 9330 17816 17190
rect 17868 16516 17920 16522
rect 17868 16458 17920 16464
rect 17880 14890 17908 16458
rect 17868 14884 17920 14890
rect 17868 14826 17920 14832
rect 17880 12238 17908 14826
rect 17960 14476 18012 14482
rect 17960 14418 18012 14424
rect 17972 13938 18000 14418
rect 17960 13932 18012 13938
rect 17960 13874 18012 13880
rect 18144 13864 18196 13870
rect 18144 13806 18196 13812
rect 18052 13184 18104 13190
rect 18052 13126 18104 13132
rect 18064 12918 18092 13126
rect 18156 12986 18184 13806
rect 18144 12980 18196 12986
rect 18144 12922 18196 12928
rect 18052 12912 18104 12918
rect 18052 12854 18104 12860
rect 17868 12232 17920 12238
rect 17868 12174 17920 12180
rect 18052 11348 18104 11354
rect 18052 11290 18104 11296
rect 17960 11144 18012 11150
rect 17960 11086 18012 11092
rect 17972 9654 18000 11086
rect 18064 10742 18092 11290
rect 18052 10736 18104 10742
rect 18052 10678 18104 10684
rect 17960 9648 18012 9654
rect 17960 9590 18012 9596
rect 17960 9376 18012 9382
rect 17788 9302 17908 9330
rect 17960 9318 18012 9324
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 17500 4004 17552 4010
rect 17500 3946 17552 3952
rect 14188 3936 14240 3942
rect 14188 3878 14240 3884
rect 13360 3596 13412 3602
rect 13360 3538 13412 3544
rect 14200 3126 14228 3878
rect 17040 3596 17092 3602
rect 17040 3538 17092 3544
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 14188 3120 14240 3126
rect 14188 3062 14240 3068
rect 14292 3058 14320 3470
rect 14464 3392 14516 3398
rect 14464 3334 14516 3340
rect 14476 3126 14504 3334
rect 14464 3120 14516 3126
rect 14464 3062 14516 3068
rect 17052 3058 17080 3538
rect 17132 3528 17184 3534
rect 17408 3528 17460 3534
rect 17184 3488 17408 3516
rect 17132 3470 17184 3476
rect 17408 3470 17460 3476
rect 17500 3392 17552 3398
rect 17500 3334 17552 3340
rect 17512 3126 17540 3334
rect 17500 3120 17552 3126
rect 17500 3062 17552 3068
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 15476 2984 15528 2990
rect 15476 2926 15528 2932
rect 13004 2746 13216 2774
rect 5920 734 6224 762
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13188 762 13216 2746
rect 14738 2544 14794 2553
rect 14738 2479 14740 2488
rect 14792 2479 14794 2488
rect 14740 2450 14792 2456
rect 14188 2372 14240 2378
rect 14188 2314 14240 2320
rect 13464 870 13584 898
rect 13464 762 13492 870
rect 13556 800 13584 870
rect 14200 800 14228 2314
rect 15488 800 15516 2926
rect 17788 2582 17816 9114
rect 17880 5234 17908 9302
rect 17972 8498 18000 9318
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 18144 8424 18196 8430
rect 18144 8366 18196 8372
rect 18156 8090 18184 8366
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 17868 5228 17920 5234
rect 17868 5170 17920 5176
rect 18052 2984 18104 2990
rect 18052 2926 18104 2932
rect 17776 2576 17828 2582
rect 17776 2518 17828 2524
rect 17408 2372 17460 2378
rect 17408 2314 17460 2320
rect 17420 800 17448 2314
rect 18064 800 18092 2926
rect 18248 2650 18276 20402
rect 18340 17202 18368 26846
rect 18616 26738 18644 33458
rect 18696 32224 18748 32230
rect 18696 32166 18748 32172
rect 18708 31278 18736 32166
rect 18696 31272 18748 31278
rect 18696 31214 18748 31220
rect 18708 30666 18736 31214
rect 18696 30660 18748 30666
rect 18696 30602 18748 30608
rect 18432 26710 18644 26738
rect 18432 24750 18460 26710
rect 18800 26500 18828 36790
rect 18892 33318 18920 38830
rect 18972 34672 19024 34678
rect 18972 34614 19024 34620
rect 18984 33590 19012 34614
rect 18972 33584 19024 33590
rect 18972 33526 19024 33532
rect 19076 33402 19104 47398
rect 19248 47048 19300 47054
rect 19248 46990 19300 46996
rect 19260 46578 19288 46990
rect 19248 46572 19300 46578
rect 19248 46514 19300 46520
rect 19260 46170 19288 46514
rect 19248 46164 19300 46170
rect 19248 46106 19300 46112
rect 19260 45966 19288 46106
rect 19248 45960 19300 45966
rect 19248 45902 19300 45908
rect 19156 45892 19208 45898
rect 19156 45834 19208 45840
rect 19168 36174 19196 45834
rect 19260 45490 19288 45902
rect 19248 45484 19300 45490
rect 19248 45426 19300 45432
rect 19248 38344 19300 38350
rect 19248 38286 19300 38292
rect 19156 36168 19208 36174
rect 19156 36110 19208 36116
rect 19156 36032 19208 36038
rect 19156 35974 19208 35980
rect 19168 35086 19196 35974
rect 19260 35834 19288 38286
rect 19248 35828 19300 35834
rect 19248 35770 19300 35776
rect 19248 35692 19300 35698
rect 19248 35634 19300 35640
rect 19156 35080 19208 35086
rect 19156 35022 19208 35028
rect 19260 34950 19288 35634
rect 19248 34944 19300 34950
rect 19248 34886 19300 34892
rect 18984 33374 19104 33402
rect 18880 33312 18932 33318
rect 18880 33254 18932 33260
rect 18880 32768 18932 32774
rect 18880 32710 18932 32716
rect 18892 31414 18920 32710
rect 18880 31408 18932 31414
rect 18880 31350 18932 31356
rect 18524 26472 18828 26500
rect 18420 24744 18472 24750
rect 18420 24686 18472 24692
rect 18420 21548 18472 21554
rect 18420 21490 18472 21496
rect 18432 21078 18460 21490
rect 18420 21072 18472 21078
rect 18420 21014 18472 21020
rect 18524 18442 18552 26472
rect 18984 26364 19012 33374
rect 19064 33312 19116 33318
rect 19064 33254 19116 33260
rect 18616 26336 19012 26364
rect 18616 20058 18644 26336
rect 19076 26228 19104 33254
rect 19352 30394 19380 47602
rect 20076 47456 20128 47462
rect 20076 47398 20128 47404
rect 20088 46986 20116 47398
rect 20076 46980 20128 46986
rect 20076 46922 20128 46928
rect 19574 46812 19882 46832
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46736 19882 46756
rect 20076 46504 20128 46510
rect 20076 46446 20128 46452
rect 19984 45892 20036 45898
rect 19984 45834 20036 45840
rect 19574 45724 19882 45744
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45648 19882 45668
rect 19574 44636 19882 44656
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44560 19882 44580
rect 19574 43548 19882 43568
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43472 19882 43492
rect 19574 42460 19882 42480
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42384 19882 42404
rect 19574 41372 19882 41392
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41296 19882 41316
rect 19574 40284 19882 40304
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40208 19882 40228
rect 19432 39296 19484 39302
rect 19432 39238 19484 39244
rect 19444 38418 19472 39238
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 19996 38842 20024 45834
rect 20088 45626 20116 46446
rect 20076 45620 20128 45626
rect 20076 45562 20128 45568
rect 20088 38978 20116 45562
rect 20088 38950 20208 38978
rect 19996 38814 20116 38842
rect 19984 38752 20036 38758
rect 19984 38694 20036 38700
rect 19432 38412 19484 38418
rect 19432 38354 19484 38360
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 19708 37936 19760 37942
rect 19706 37904 19708 37913
rect 19760 37904 19762 37913
rect 19706 37839 19762 37848
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 19996 36242 20024 38694
rect 19984 36236 20036 36242
rect 19984 36178 20036 36184
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19984 35148 20036 35154
rect 19984 35090 20036 35096
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 19708 34536 19760 34542
rect 19708 34478 19760 34484
rect 19720 33998 19748 34478
rect 19708 33992 19760 33998
rect 19708 33934 19760 33940
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 19996 33522 20024 35090
rect 19984 33516 20036 33522
rect 19984 33458 20036 33464
rect 19996 33046 20024 33458
rect 19984 33040 20036 33046
rect 19984 32982 20036 32988
rect 20088 32858 20116 38814
rect 19996 32830 20116 32858
rect 19432 32768 19484 32774
rect 19432 32710 19484 32716
rect 19444 31890 19472 32710
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 19432 31884 19484 31890
rect 19432 31826 19484 31832
rect 19996 31754 20024 32830
rect 20180 32756 20208 38950
rect 20272 35766 20300 47654
rect 20456 42090 20484 49370
rect 20536 49088 20588 49094
rect 20536 49030 20588 49036
rect 20548 46934 20576 49030
rect 20640 48210 20668 51200
rect 21364 49292 21416 49298
rect 21364 49234 21416 49240
rect 20996 49224 21048 49230
rect 20996 49166 21048 49172
rect 21008 48278 21036 49166
rect 21088 49156 21140 49162
rect 21088 49098 21140 49104
rect 20996 48272 21048 48278
rect 20996 48214 21048 48220
rect 20628 48204 20680 48210
rect 20628 48146 20680 48152
rect 20548 46906 20668 46934
rect 20640 42242 20668 46906
rect 20548 42214 20668 42242
rect 20444 42084 20496 42090
rect 20444 42026 20496 42032
rect 20444 39976 20496 39982
rect 20444 39918 20496 39924
rect 20456 39506 20484 39918
rect 20444 39500 20496 39506
rect 20444 39442 20496 39448
rect 20456 37262 20484 39442
rect 20444 37256 20496 37262
rect 20444 37198 20496 37204
rect 20352 37188 20404 37194
rect 20352 37130 20404 37136
rect 20364 37097 20392 37130
rect 20350 37088 20406 37097
rect 20350 37023 20406 37032
rect 20456 36854 20484 37198
rect 20444 36848 20496 36854
rect 20444 36790 20496 36796
rect 20352 36712 20404 36718
rect 20352 36654 20404 36660
rect 20260 35760 20312 35766
rect 20260 35702 20312 35708
rect 19444 31726 20024 31754
rect 20088 32728 20208 32756
rect 19340 30388 19392 30394
rect 19340 30330 19392 30336
rect 19340 29640 19392 29646
rect 19340 29582 19392 29588
rect 19352 28966 19380 29582
rect 19340 28960 19392 28966
rect 19340 28902 19392 28908
rect 19352 28082 19380 28902
rect 19340 28076 19392 28082
rect 19340 28018 19392 28024
rect 19444 26874 19472 31726
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19524 30320 19576 30326
rect 19524 30262 19576 30268
rect 19536 29850 19564 30262
rect 19708 30252 19760 30258
rect 19708 30194 19760 30200
rect 19720 30161 19748 30194
rect 19984 30184 20036 30190
rect 19706 30152 19762 30161
rect 19984 30126 20036 30132
rect 19706 30087 19762 30096
rect 19996 29850 20024 30126
rect 19524 29844 19576 29850
rect 19524 29786 19576 29792
rect 19984 29844 20036 29850
rect 19984 29786 20036 29792
rect 19982 29744 20038 29753
rect 19982 29679 20038 29688
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19892 29164 19944 29170
rect 19892 29106 19944 29112
rect 19616 28960 19668 28966
rect 19616 28902 19668 28908
rect 19628 28490 19656 28902
rect 19904 28558 19932 29106
rect 19892 28552 19944 28558
rect 19892 28494 19944 28500
rect 19616 28484 19668 28490
rect 19616 28426 19668 28432
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 19996 28257 20024 29679
rect 19982 28248 20038 28257
rect 19982 28183 20038 28192
rect 19984 28076 20036 28082
rect 19984 28018 20036 28024
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 19524 26988 19576 26994
rect 19524 26930 19576 26936
rect 19352 26846 19472 26874
rect 19156 26308 19208 26314
rect 19156 26250 19208 26256
rect 18892 26200 19104 26228
rect 18892 25906 18920 26200
rect 19064 26036 19116 26042
rect 19064 25978 19116 25984
rect 19076 25906 19104 25978
rect 18880 25900 18932 25906
rect 18880 25842 18932 25848
rect 19064 25900 19116 25906
rect 19064 25842 19116 25848
rect 18788 25696 18840 25702
rect 18788 25638 18840 25644
rect 18800 25226 18828 25638
rect 19168 25226 19196 26250
rect 19248 25900 19300 25906
rect 19248 25842 19300 25848
rect 18788 25220 18840 25226
rect 18788 25162 18840 25168
rect 19156 25220 19208 25226
rect 19156 25162 19208 25168
rect 19168 24818 19196 25162
rect 19260 24954 19288 25842
rect 19248 24948 19300 24954
rect 19248 24890 19300 24896
rect 19156 24812 19208 24818
rect 19156 24754 19208 24760
rect 18788 24744 18840 24750
rect 18788 24686 18840 24692
rect 18696 23112 18748 23118
rect 18696 23054 18748 23060
rect 18708 22166 18736 23054
rect 18696 22160 18748 22166
rect 18696 22102 18748 22108
rect 18708 20466 18736 22102
rect 18696 20460 18748 20466
rect 18696 20402 18748 20408
rect 18604 20052 18656 20058
rect 18604 19994 18656 20000
rect 18432 18414 18552 18442
rect 18432 17921 18460 18414
rect 18512 18284 18564 18290
rect 18512 18226 18564 18232
rect 18604 18284 18656 18290
rect 18604 18226 18656 18232
rect 18418 17912 18474 17921
rect 18418 17847 18474 17856
rect 18524 17338 18552 18226
rect 18512 17332 18564 17338
rect 18512 17274 18564 17280
rect 18328 17196 18380 17202
rect 18328 17138 18380 17144
rect 18616 16998 18644 18226
rect 18696 18080 18748 18086
rect 18696 18022 18748 18028
rect 18604 16992 18656 16998
rect 18604 16934 18656 16940
rect 18328 16108 18380 16114
rect 18328 16050 18380 16056
rect 18340 15502 18368 16050
rect 18512 16040 18564 16046
rect 18512 15982 18564 15988
rect 18420 15564 18472 15570
rect 18420 15506 18472 15512
rect 18328 15496 18380 15502
rect 18328 15438 18380 15444
rect 18340 15026 18368 15438
rect 18328 15020 18380 15026
rect 18328 14962 18380 14968
rect 18328 11008 18380 11014
rect 18328 10950 18380 10956
rect 18340 3534 18368 10950
rect 18432 4146 18460 15506
rect 18524 4826 18552 15982
rect 18708 15638 18736 18022
rect 18696 15632 18748 15638
rect 18696 15574 18748 15580
rect 18696 13184 18748 13190
rect 18696 13126 18748 13132
rect 18604 12640 18656 12646
rect 18604 12582 18656 12588
rect 18616 9722 18644 12582
rect 18604 9716 18656 9722
rect 18604 9658 18656 9664
rect 18616 7886 18644 9658
rect 18708 9586 18736 13126
rect 18800 12434 18828 24686
rect 19168 24206 19196 24754
rect 19156 24200 19208 24206
rect 19156 24142 19208 24148
rect 19168 23866 19196 24142
rect 19156 23860 19208 23866
rect 19156 23802 19208 23808
rect 19248 23724 19300 23730
rect 19248 23666 19300 23672
rect 19156 23180 19208 23186
rect 19156 23122 19208 23128
rect 18880 22432 18932 22438
rect 18880 22374 18932 22380
rect 18892 21962 18920 22374
rect 18880 21956 18932 21962
rect 18880 21898 18932 21904
rect 18892 21554 18920 21898
rect 19168 21894 19196 23122
rect 19260 22982 19288 23666
rect 19248 22976 19300 22982
rect 19248 22918 19300 22924
rect 19156 21888 19208 21894
rect 19156 21830 19208 21836
rect 19064 21616 19116 21622
rect 19064 21558 19116 21564
rect 18880 21548 18932 21554
rect 18880 21490 18932 21496
rect 18972 21480 19024 21486
rect 18972 21422 19024 21428
rect 18984 21146 19012 21422
rect 18972 21140 19024 21146
rect 18972 21082 19024 21088
rect 19076 20466 19104 21558
rect 19168 20602 19196 21830
rect 19260 21622 19288 22918
rect 19248 21616 19300 21622
rect 19248 21558 19300 21564
rect 19156 20596 19208 20602
rect 19156 20538 19208 20544
rect 19064 20460 19116 20466
rect 19064 20402 19116 20408
rect 19248 20460 19300 20466
rect 19248 20402 19300 20408
rect 19156 20392 19208 20398
rect 19156 20334 19208 20340
rect 18972 16992 19024 16998
rect 18972 16934 19024 16940
rect 18984 16522 19012 16934
rect 18972 16516 19024 16522
rect 18972 16458 19024 16464
rect 18984 16114 19012 16458
rect 18972 16108 19024 16114
rect 18972 16050 19024 16056
rect 19168 15094 19196 20334
rect 19260 20058 19288 20402
rect 19248 20052 19300 20058
rect 19248 19994 19300 20000
rect 19156 15088 19208 15094
rect 19156 15030 19208 15036
rect 19168 14958 19196 15030
rect 19156 14952 19208 14958
rect 19156 14894 19208 14900
rect 18800 12406 18920 12434
rect 18788 11076 18840 11082
rect 18788 11018 18840 11024
rect 18800 10810 18828 11018
rect 18788 10804 18840 10810
rect 18788 10746 18840 10752
rect 18892 10554 18920 12406
rect 19064 11688 19116 11694
rect 19064 11630 19116 11636
rect 18972 11552 19024 11558
rect 18972 11494 19024 11500
rect 18984 11218 19012 11494
rect 18972 11212 19024 11218
rect 18972 11154 19024 11160
rect 19076 10690 19104 11630
rect 19168 11014 19196 14894
rect 19248 14272 19300 14278
rect 19248 14214 19300 14220
rect 19260 14006 19288 14214
rect 19248 14000 19300 14006
rect 19248 13942 19300 13948
rect 19248 13728 19300 13734
rect 19248 13670 19300 13676
rect 19260 13326 19288 13670
rect 19248 13320 19300 13326
rect 19248 13262 19300 13268
rect 19260 12374 19288 13262
rect 19248 12368 19300 12374
rect 19248 12310 19300 12316
rect 19260 11082 19288 12310
rect 19352 12209 19380 26846
rect 19536 26586 19564 26930
rect 19524 26580 19576 26586
rect 19524 26522 19576 26528
rect 19536 26382 19564 26522
rect 19524 26376 19576 26382
rect 19996 26364 20024 28018
rect 20088 26500 20116 32728
rect 20168 32428 20220 32434
rect 20168 32370 20220 32376
rect 20180 31414 20208 32370
rect 20168 31408 20220 31414
rect 20168 31350 20220 31356
rect 20180 30734 20208 31350
rect 20168 30728 20220 30734
rect 20168 30670 20220 30676
rect 20168 30252 20220 30258
rect 20168 30194 20220 30200
rect 20180 29306 20208 30194
rect 20168 29300 20220 29306
rect 20168 29242 20220 29248
rect 20168 28688 20220 28694
rect 20168 28630 20220 28636
rect 20180 28150 20208 28630
rect 20168 28144 20220 28150
rect 20168 28086 20220 28092
rect 20272 26874 20300 35702
rect 20364 34066 20392 36654
rect 20456 35290 20484 36790
rect 20444 35284 20496 35290
rect 20444 35226 20496 35232
rect 20352 34060 20404 34066
rect 20352 34002 20404 34008
rect 20364 32434 20392 34002
rect 20444 33516 20496 33522
rect 20444 33458 20496 33464
rect 20456 33114 20484 33458
rect 20444 33108 20496 33114
rect 20444 33050 20496 33056
rect 20352 32428 20404 32434
rect 20352 32370 20404 32376
rect 20352 32224 20404 32230
rect 20352 32166 20404 32172
rect 20364 30297 20392 32166
rect 20548 31362 20576 42214
rect 20628 42084 20680 42090
rect 20628 42026 20680 42032
rect 20640 35698 20668 42026
rect 21100 41614 21128 49098
rect 21088 41608 21140 41614
rect 21088 41550 21140 41556
rect 20996 40044 21048 40050
rect 20996 39986 21048 39992
rect 21272 40044 21324 40050
rect 21272 39986 21324 39992
rect 20904 39840 20956 39846
rect 20904 39782 20956 39788
rect 20720 39364 20772 39370
rect 20720 39306 20772 39312
rect 20732 39098 20760 39306
rect 20720 39092 20772 39098
rect 20720 39034 20772 39040
rect 20916 38962 20944 39782
rect 20904 38956 20956 38962
rect 20904 38898 20956 38904
rect 21008 38418 21036 39986
rect 21284 39302 21312 39986
rect 21272 39296 21324 39302
rect 21272 39238 21324 39244
rect 21088 38956 21140 38962
rect 21088 38898 21140 38904
rect 21100 38826 21128 38898
rect 21088 38820 21140 38826
rect 21088 38762 21140 38768
rect 20996 38412 21048 38418
rect 20996 38354 21048 38360
rect 20720 37800 20772 37806
rect 20720 37742 20772 37748
rect 20732 37466 20760 37742
rect 20720 37460 20772 37466
rect 20720 37402 20772 37408
rect 21100 36786 21128 38762
rect 21088 36780 21140 36786
rect 21088 36722 21140 36728
rect 21272 36032 21324 36038
rect 21272 35974 21324 35980
rect 21088 35828 21140 35834
rect 21088 35770 21140 35776
rect 20994 35728 21050 35737
rect 20628 35692 20680 35698
rect 20628 35634 20680 35640
rect 20916 35672 20994 35680
rect 20916 35652 20996 35672
rect 20720 35624 20772 35630
rect 20720 35566 20772 35572
rect 20628 35488 20680 35494
rect 20628 35430 20680 35436
rect 20640 35086 20668 35430
rect 20628 35080 20680 35086
rect 20628 35022 20680 35028
rect 20732 34932 20760 35566
rect 20640 34904 20760 34932
rect 20812 34944 20864 34950
rect 20640 33998 20668 34904
rect 20812 34886 20864 34892
rect 20824 34610 20852 34886
rect 20812 34604 20864 34610
rect 20812 34546 20864 34552
rect 20628 33992 20680 33998
rect 20628 33934 20680 33940
rect 20640 33046 20668 33934
rect 20628 33040 20680 33046
rect 20628 32982 20680 32988
rect 20809 32904 20861 32910
rect 20916 32892 20944 35652
rect 21048 35663 21050 35672
rect 20996 35634 21048 35640
rect 21100 34542 21128 35770
rect 21180 34604 21232 34610
rect 21180 34546 21232 34552
rect 21088 34536 21140 34542
rect 21088 34478 21140 34484
rect 20996 33312 21048 33318
rect 20996 33254 21048 33260
rect 21008 32978 21036 33254
rect 20996 32972 21048 32978
rect 20996 32914 21048 32920
rect 20861 32864 20944 32892
rect 20809 32846 20861 32852
rect 20548 31334 20668 31362
rect 20536 31272 20588 31278
rect 20536 31214 20588 31220
rect 20548 30433 20576 31214
rect 20534 30424 20590 30433
rect 20444 30388 20496 30394
rect 20534 30359 20590 30368
rect 20444 30330 20496 30336
rect 20350 30288 20406 30297
rect 20350 30223 20406 30232
rect 20456 30138 20484 30330
rect 20364 30110 20484 30138
rect 20364 29594 20392 30110
rect 20444 30048 20496 30054
rect 20444 29990 20496 29996
rect 20536 30048 20588 30054
rect 20536 29990 20588 29996
rect 20456 29714 20484 29990
rect 20444 29708 20496 29714
rect 20444 29650 20496 29656
rect 20548 29646 20576 29990
rect 20536 29640 20588 29646
rect 20364 29566 20484 29594
rect 20536 29582 20588 29588
rect 20350 29336 20406 29345
rect 20350 29271 20406 29280
rect 20364 27033 20392 29271
rect 20350 27024 20406 27033
rect 20350 26959 20406 26968
rect 20272 26846 20392 26874
rect 20088 26472 20208 26500
rect 20076 26376 20128 26382
rect 19996 26336 20076 26364
rect 19524 26318 19576 26324
rect 20076 26318 20128 26324
rect 19432 26240 19484 26246
rect 19432 26182 19484 26188
rect 19444 25906 19472 26182
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19892 25968 19944 25974
rect 19892 25910 19944 25916
rect 19432 25900 19484 25906
rect 19432 25842 19484 25848
rect 19444 24818 19472 25842
rect 19904 25702 19932 25910
rect 19984 25764 20036 25770
rect 19984 25706 20036 25712
rect 19892 25696 19944 25702
rect 19892 25638 19944 25644
rect 19996 25537 20024 25706
rect 19982 25528 20038 25537
rect 19524 25492 19576 25498
rect 19982 25463 20038 25472
rect 19524 25434 19576 25440
rect 19536 25226 19564 25434
rect 20088 25294 20116 26318
rect 20180 25344 20208 26472
rect 20260 26308 20312 26314
rect 20260 26250 20312 26256
rect 20272 26042 20300 26250
rect 20260 26036 20312 26042
rect 20260 25978 20312 25984
rect 20260 25900 20312 25906
rect 20260 25842 20312 25848
rect 20272 25673 20300 25842
rect 20258 25664 20314 25673
rect 20258 25599 20314 25608
rect 20180 25316 20300 25344
rect 20076 25288 20128 25294
rect 20076 25230 20128 25236
rect 19524 25220 19576 25226
rect 19524 25162 19576 25168
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19892 24880 19944 24886
rect 19890 24848 19892 24857
rect 19944 24848 19946 24857
rect 19432 24812 19484 24818
rect 19890 24783 19946 24792
rect 19432 24754 19484 24760
rect 19444 23662 19472 24754
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 20088 23848 20116 25230
rect 20168 25220 20220 25226
rect 20168 25162 20220 25168
rect 20180 24954 20208 25162
rect 20168 24948 20220 24954
rect 20168 24890 20220 24896
rect 20168 24064 20220 24070
rect 20168 24006 20220 24012
rect 19904 23820 20116 23848
rect 19432 23656 19484 23662
rect 19432 23598 19484 23604
rect 19904 23186 19932 23820
rect 20180 23594 20208 24006
rect 20168 23588 20220 23594
rect 20168 23530 20220 23536
rect 20272 23254 20300 25316
rect 19984 23248 20036 23254
rect 19984 23190 20036 23196
rect 20260 23248 20312 23254
rect 20260 23190 20312 23196
rect 19892 23180 19944 23186
rect 19892 23122 19944 23128
rect 19432 23112 19484 23118
rect 19432 23054 19484 23060
rect 19444 22760 19472 23054
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19444 22732 19555 22760
rect 19527 22692 19555 22732
rect 19527 22681 19564 22692
rect 19522 22672 19578 22681
rect 19432 22636 19484 22642
rect 19522 22607 19578 22616
rect 19432 22578 19484 22584
rect 19444 22098 19472 22578
rect 19432 22092 19484 22098
rect 19432 22034 19484 22040
rect 19536 21978 19564 22607
rect 19798 22264 19854 22273
rect 19798 22199 19800 22208
rect 19852 22199 19854 22208
rect 19800 22170 19852 22176
rect 19892 22160 19944 22166
rect 19892 22102 19944 22108
rect 19904 22030 19932 22102
rect 19444 21950 19564 21978
rect 19892 22024 19944 22030
rect 19892 21966 19944 21972
rect 19444 15473 19472 21950
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19890 19408 19946 19417
rect 19890 19343 19946 19352
rect 19904 18737 19932 19343
rect 19890 18728 19946 18737
rect 19890 18663 19946 18672
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19524 16040 19576 16046
rect 19524 15982 19576 15988
rect 19536 15706 19564 15982
rect 19524 15700 19576 15706
rect 19524 15642 19576 15648
rect 19430 15464 19486 15473
rect 19430 15399 19486 15408
rect 19432 15360 19484 15366
rect 19432 15302 19484 15308
rect 19444 14906 19472 15302
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19614 15056 19670 15065
rect 19614 14991 19670 15000
rect 19444 14878 19564 14906
rect 19432 14816 19484 14822
rect 19432 14758 19484 14764
rect 19444 14414 19472 14758
rect 19432 14408 19484 14414
rect 19432 14350 19484 14356
rect 19536 14260 19564 14878
rect 19628 14385 19656 14991
rect 19614 14376 19670 14385
rect 19614 14311 19616 14320
rect 19668 14311 19670 14320
rect 19616 14282 19668 14288
rect 19444 14232 19564 14260
rect 19444 12646 19472 14232
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 19616 12912 19668 12918
rect 19616 12854 19668 12860
rect 19432 12640 19484 12646
rect 19432 12582 19484 12588
rect 19338 12200 19394 12209
rect 19628 12170 19656 12854
rect 19338 12135 19394 12144
rect 19616 12164 19668 12170
rect 19616 12106 19668 12112
rect 19340 12096 19392 12102
rect 19340 12038 19392 12044
rect 19248 11076 19300 11082
rect 19248 11018 19300 11024
rect 19156 11008 19208 11014
rect 19156 10950 19208 10956
rect 19260 10810 19288 11018
rect 19248 10804 19300 10810
rect 19248 10746 19300 10752
rect 18984 10674 19104 10690
rect 18972 10668 19104 10674
rect 19024 10662 19104 10668
rect 18972 10610 19024 10616
rect 18892 10526 19012 10554
rect 18696 9580 18748 9586
rect 18696 9522 18748 9528
rect 18696 8016 18748 8022
rect 18696 7958 18748 7964
rect 18604 7880 18656 7886
rect 18604 7822 18656 7828
rect 18616 7410 18644 7822
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 18512 4820 18564 4826
rect 18512 4762 18564 4768
rect 18420 4140 18472 4146
rect 18420 4082 18472 4088
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 18236 2644 18288 2650
rect 18236 2586 18288 2592
rect 18708 800 18736 7958
rect 18880 7812 18932 7818
rect 18880 7754 18932 7760
rect 18892 7546 18920 7754
rect 18880 7540 18932 7546
rect 18880 7482 18932 7488
rect 18984 6730 19012 10526
rect 19076 10282 19104 10662
rect 19076 10254 19196 10282
rect 19168 9994 19196 10254
rect 19156 9988 19208 9994
rect 19156 9930 19208 9936
rect 19168 8974 19196 9930
rect 19260 9042 19288 10746
rect 19352 10606 19380 12038
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19890 11792 19946 11801
rect 19890 11727 19892 11736
rect 19944 11727 19946 11736
rect 19892 11698 19944 11704
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19444 10674 19472 11086
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19432 10668 19484 10674
rect 19432 10610 19484 10616
rect 19800 10668 19852 10674
rect 19800 10610 19852 10616
rect 19340 10600 19392 10606
rect 19340 10542 19392 10548
rect 19352 10198 19380 10542
rect 19340 10192 19392 10198
rect 19340 10134 19392 10140
rect 19432 9988 19484 9994
rect 19432 9930 19484 9936
rect 19340 9920 19392 9926
rect 19340 9862 19392 9868
rect 19352 9625 19380 9862
rect 19338 9616 19394 9625
rect 19338 9551 19394 9560
rect 19444 9382 19472 9930
rect 19812 9908 19840 10610
rect 19996 10146 20024 23190
rect 20168 23112 20220 23118
rect 20168 23054 20220 23060
rect 20258 23080 20314 23089
rect 20076 22976 20128 22982
rect 20076 22918 20128 22924
rect 20088 20602 20116 22918
rect 20076 20596 20128 20602
rect 20076 20538 20128 20544
rect 20076 20460 20128 20466
rect 20076 20402 20128 20408
rect 20088 19174 20116 20402
rect 20076 19168 20128 19174
rect 20076 19110 20128 19116
rect 20088 18766 20116 19110
rect 20076 18760 20128 18766
rect 20076 18702 20128 18708
rect 20076 17740 20128 17746
rect 20076 17682 20128 17688
rect 20088 16794 20116 17682
rect 20180 16998 20208 23054
rect 20258 23015 20314 23024
rect 20168 16992 20220 16998
rect 20168 16934 20220 16940
rect 20076 16788 20128 16794
rect 20076 16730 20128 16736
rect 20076 16040 20128 16046
rect 20076 15982 20128 15988
rect 20088 12918 20116 15982
rect 20168 15972 20220 15978
rect 20168 15914 20220 15920
rect 20180 14482 20208 15914
rect 20168 14476 20220 14482
rect 20168 14418 20220 14424
rect 20166 14376 20222 14385
rect 20166 14311 20222 14320
rect 20076 12912 20128 12918
rect 20076 12854 20128 12860
rect 20074 12744 20130 12753
rect 20074 12679 20130 12688
rect 20088 12374 20116 12679
rect 20076 12368 20128 12374
rect 20076 12310 20128 12316
rect 20076 12164 20128 12170
rect 20076 12106 20128 12112
rect 20088 10742 20116 12106
rect 20180 11098 20208 14311
rect 20272 11218 20300 23015
rect 20364 22094 20392 26846
rect 20456 22982 20484 29566
rect 20640 29322 20668 31334
rect 20916 30394 20944 32864
rect 21100 31906 21128 34478
rect 21008 31878 21128 31906
rect 20904 30388 20956 30394
rect 20904 30330 20956 30336
rect 20916 30190 20944 30330
rect 20904 30184 20956 30190
rect 20904 30126 20956 30132
rect 21008 29753 21036 31878
rect 21088 31816 21140 31822
rect 21088 31758 21140 31764
rect 20994 29744 21050 29753
rect 20994 29679 21050 29688
rect 20640 29294 20852 29322
rect 20628 29232 20680 29238
rect 20628 29174 20680 29180
rect 20536 28484 20588 28490
rect 20536 28426 20588 28432
rect 20548 26330 20576 28426
rect 20640 27878 20668 29174
rect 20720 28552 20772 28558
rect 20720 28494 20772 28500
rect 20628 27872 20680 27878
rect 20628 27814 20680 27820
rect 20640 27470 20668 27814
rect 20732 27606 20760 28494
rect 20720 27600 20772 27606
rect 20720 27542 20772 27548
rect 20628 27464 20680 27470
rect 20628 27406 20680 27412
rect 20548 26302 20668 26330
rect 20536 26240 20588 26246
rect 20536 26182 20588 26188
rect 20548 25906 20576 26182
rect 20536 25900 20588 25906
rect 20536 25842 20588 25848
rect 20536 25152 20588 25158
rect 20536 25094 20588 25100
rect 20548 24818 20576 25094
rect 20536 24812 20588 24818
rect 20536 24754 20588 24760
rect 20444 22976 20496 22982
rect 20444 22918 20496 22924
rect 20364 22066 20484 22094
rect 20352 21956 20404 21962
rect 20352 21898 20404 21904
rect 20364 21690 20392 21898
rect 20352 21684 20404 21690
rect 20352 21626 20404 21632
rect 20352 20256 20404 20262
rect 20352 20198 20404 20204
rect 20364 19854 20392 20198
rect 20352 19848 20404 19854
rect 20352 19790 20404 19796
rect 20350 19680 20406 19689
rect 20350 19615 20406 19624
rect 20364 18358 20392 19615
rect 20352 18352 20404 18358
rect 20352 18294 20404 18300
rect 20364 17377 20392 18294
rect 20350 17368 20406 17377
rect 20350 17303 20406 17312
rect 20456 17218 20484 22066
rect 20536 20460 20588 20466
rect 20536 20402 20588 20408
rect 20548 19990 20576 20402
rect 20536 19984 20588 19990
rect 20536 19926 20588 19932
rect 20548 18834 20576 19926
rect 20640 19825 20668 26302
rect 20824 26246 20852 29294
rect 20904 29164 20956 29170
rect 20904 29106 20956 29112
rect 20916 27674 20944 29106
rect 20904 27668 20956 27674
rect 20904 27610 20956 27616
rect 20812 26240 20864 26246
rect 20812 26182 20864 26188
rect 20720 25900 20772 25906
rect 20720 25842 20772 25848
rect 20732 24818 20760 25842
rect 20812 25832 20864 25838
rect 20812 25774 20864 25780
rect 20720 24812 20772 24818
rect 20720 24754 20772 24760
rect 20824 24750 20852 25774
rect 20812 24744 20864 24750
rect 20812 24686 20864 24692
rect 20916 23118 20944 27610
rect 20996 26920 21048 26926
rect 20996 26862 21048 26868
rect 20904 23112 20956 23118
rect 20904 23054 20956 23060
rect 20720 22432 20772 22438
rect 20720 22374 20772 22380
rect 20732 21418 20760 22374
rect 20904 22024 20956 22030
rect 21008 22012 21036 26862
rect 21100 26790 21128 31758
rect 21192 28558 21220 34546
rect 21284 34202 21312 35974
rect 21272 34196 21324 34202
rect 21272 34138 21324 34144
rect 21376 32230 21404 49234
rect 22020 48822 22048 51326
rect 22558 51200 22614 52000
rect 23202 51354 23258 52000
rect 23846 51354 23902 52000
rect 24490 51354 24546 52000
rect 23202 51326 23428 51354
rect 23202 51200 23258 51326
rect 22572 49298 22600 51200
rect 22376 49292 22428 49298
rect 22376 49234 22428 49240
rect 22560 49292 22612 49298
rect 22560 49234 22612 49240
rect 22192 49156 22244 49162
rect 22192 49098 22244 49104
rect 22008 48816 22060 48822
rect 22008 48758 22060 48764
rect 22100 48544 22152 48550
rect 22100 48486 22152 48492
rect 21732 47660 21784 47666
rect 21732 47602 21784 47608
rect 21548 45416 21600 45422
rect 21548 45358 21600 45364
rect 21456 37460 21508 37466
rect 21456 37402 21508 37408
rect 21364 32224 21416 32230
rect 21364 32166 21416 32172
rect 21180 28552 21232 28558
rect 21180 28494 21232 28500
rect 21088 26784 21140 26790
rect 21088 26726 21140 26732
rect 21180 25424 21232 25430
rect 21180 25366 21232 25372
rect 21192 25265 21220 25366
rect 21272 25288 21324 25294
rect 21178 25256 21234 25265
rect 21272 25230 21324 25236
rect 21178 25191 21234 25200
rect 21180 22160 21232 22166
rect 21180 22102 21232 22108
rect 20956 21984 21036 22012
rect 20904 21966 20956 21972
rect 20720 21412 20772 21418
rect 20720 21354 20772 21360
rect 20626 19816 20682 19825
rect 20626 19751 20682 19760
rect 20628 19712 20680 19718
rect 20628 19654 20680 19660
rect 20640 19378 20668 19654
rect 20628 19372 20680 19378
rect 20628 19314 20680 19320
rect 20536 18828 20588 18834
rect 20536 18770 20588 18776
rect 20732 18290 20760 21354
rect 21192 21026 21220 22102
rect 20824 20998 21220 21026
rect 20824 18902 20852 20998
rect 20996 20936 21048 20942
rect 20996 20878 21048 20884
rect 21088 20936 21140 20942
rect 21088 20878 21140 20884
rect 21008 20466 21036 20878
rect 20996 20460 21048 20466
rect 20996 20402 21048 20408
rect 20996 20256 21048 20262
rect 21100 20244 21128 20878
rect 21284 20482 21312 25230
rect 21364 24132 21416 24138
rect 21364 24074 21416 24080
rect 21048 20216 21128 20244
rect 21192 20454 21312 20482
rect 20996 20198 21048 20204
rect 20904 19780 20956 19786
rect 20904 19722 20956 19728
rect 20916 19310 20944 19722
rect 20904 19304 20956 19310
rect 20904 19246 20956 19252
rect 21008 18970 21036 20198
rect 21192 19990 21220 20454
rect 21272 20392 21324 20398
rect 21272 20334 21324 20340
rect 21180 19984 21232 19990
rect 21180 19926 21232 19932
rect 21088 19236 21140 19242
rect 21088 19178 21140 19184
rect 20996 18964 21048 18970
rect 20996 18906 21048 18912
rect 20812 18896 20864 18902
rect 20812 18838 20864 18844
rect 20996 18352 21048 18358
rect 20996 18294 21048 18300
rect 20720 18284 20772 18290
rect 20720 18226 20772 18232
rect 20904 18284 20956 18290
rect 20904 18226 20956 18232
rect 20720 18080 20772 18086
rect 20720 18022 20772 18028
rect 20628 17604 20680 17610
rect 20628 17546 20680 17552
rect 20364 17190 20484 17218
rect 20536 17196 20588 17202
rect 20260 11212 20312 11218
rect 20260 11154 20312 11160
rect 20180 11070 20300 11098
rect 20076 10736 20128 10742
rect 20076 10678 20128 10684
rect 20168 10668 20220 10674
rect 20168 10610 20220 10616
rect 20180 10266 20208 10610
rect 20168 10260 20220 10266
rect 20168 10202 20220 10208
rect 19996 10118 20208 10146
rect 20074 10024 20130 10033
rect 20074 9959 20130 9968
rect 19812 9880 20024 9908
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19996 9722 20024 9880
rect 19984 9716 20036 9722
rect 19984 9658 20036 9664
rect 19614 9616 19670 9625
rect 19996 9586 20024 9658
rect 19614 9551 19616 9560
rect 19668 9551 19670 9560
rect 19984 9580 20036 9586
rect 19616 9522 19668 9528
rect 19984 9522 20036 9528
rect 19432 9376 19484 9382
rect 19432 9318 19484 9324
rect 19248 9036 19300 9042
rect 19248 8978 19300 8984
rect 19156 8968 19208 8974
rect 19156 8910 19208 8916
rect 19996 8906 20024 9522
rect 19984 8900 20036 8906
rect 19984 8842 20036 8848
rect 19432 8832 19484 8838
rect 19432 8774 19484 8780
rect 19340 8424 19392 8430
rect 19340 8366 19392 8372
rect 18972 6724 19024 6730
rect 18972 6666 19024 6672
rect 19352 3942 19380 8366
rect 19444 7546 19472 8774
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19432 7540 19484 7546
rect 19432 7482 19484 7488
rect 19430 7440 19486 7449
rect 19996 7410 20024 8842
rect 19430 7375 19486 7384
rect 19984 7404 20036 7410
rect 19340 3936 19392 3942
rect 19340 3878 19392 3884
rect 19444 3670 19472 7375
rect 19984 7346 20036 7352
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 20088 4214 20116 9959
rect 20180 5710 20208 10118
rect 20272 9586 20300 11070
rect 20364 10441 20392 17190
rect 20536 17138 20588 17144
rect 20444 16992 20496 16998
rect 20444 16934 20496 16940
rect 20350 10432 20406 10441
rect 20350 10367 20406 10376
rect 20456 10282 20484 16934
rect 20548 16794 20576 17138
rect 20640 17066 20668 17546
rect 20628 17060 20680 17066
rect 20628 17002 20680 17008
rect 20626 16960 20682 16969
rect 20626 16895 20682 16904
rect 20536 16788 20588 16794
rect 20536 16730 20588 16736
rect 20640 15978 20668 16895
rect 20732 16590 20760 18022
rect 20916 17542 20944 18226
rect 20904 17536 20956 17542
rect 20904 17478 20956 17484
rect 21008 17338 21036 18294
rect 21100 17785 21128 19178
rect 21086 17776 21142 17785
rect 21086 17711 21142 17720
rect 20812 17332 20864 17338
rect 20812 17274 20864 17280
rect 20996 17332 21048 17338
rect 20996 17274 21048 17280
rect 20824 16998 20852 17274
rect 20904 17128 20956 17134
rect 20904 17070 20956 17076
rect 20812 16992 20864 16998
rect 20812 16934 20864 16940
rect 20720 16584 20772 16590
rect 20720 16526 20772 16532
rect 20812 16516 20864 16522
rect 20812 16458 20864 16464
rect 20720 16108 20772 16114
rect 20720 16050 20772 16056
rect 20628 15972 20680 15978
rect 20628 15914 20680 15920
rect 20732 15586 20760 16050
rect 20640 15558 20760 15586
rect 20536 15360 20588 15366
rect 20536 15302 20588 15308
rect 20548 15162 20576 15302
rect 20536 15156 20588 15162
rect 20536 15098 20588 15104
rect 20640 15008 20668 15558
rect 20720 15496 20772 15502
rect 20720 15438 20772 15444
rect 20732 15162 20760 15438
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 20548 14980 20668 15008
rect 20548 14550 20576 14980
rect 20720 14952 20772 14958
rect 20720 14894 20772 14900
rect 20628 14816 20680 14822
rect 20628 14758 20680 14764
rect 20536 14544 20588 14550
rect 20536 14486 20588 14492
rect 20640 14006 20668 14758
rect 20732 14346 20760 14894
rect 20824 14414 20852 16458
rect 20916 16114 20944 17070
rect 21008 16590 21036 17274
rect 20996 16584 21048 16590
rect 20996 16526 21048 16532
rect 20996 16448 21048 16454
rect 20996 16390 21048 16396
rect 20904 16108 20956 16114
rect 20904 16050 20956 16056
rect 20904 15496 20956 15502
rect 20904 15438 20956 15444
rect 20916 14618 20944 15438
rect 20904 14612 20956 14618
rect 20904 14554 20956 14560
rect 20812 14408 20864 14414
rect 20812 14350 20864 14356
rect 20720 14340 20772 14346
rect 20720 14282 20772 14288
rect 20628 14000 20680 14006
rect 20628 13942 20680 13948
rect 20536 13932 20588 13938
rect 20536 13874 20588 13880
rect 20548 13530 20576 13874
rect 20628 13864 20680 13870
rect 20628 13806 20680 13812
rect 20536 13524 20588 13530
rect 20536 13466 20588 13472
rect 20640 13190 20668 13806
rect 20732 13394 20760 14282
rect 20904 14272 20956 14278
rect 20904 14214 20956 14220
rect 21008 14226 21036 16390
rect 21192 15706 21220 19926
rect 21284 17338 21312 20334
rect 21272 17332 21324 17338
rect 21272 17274 21324 17280
rect 21180 15700 21232 15706
rect 21180 15642 21232 15648
rect 21088 15496 21140 15502
rect 21088 15438 21140 15444
rect 21100 14346 21128 15438
rect 21180 15020 21232 15026
rect 21180 14962 21232 14968
rect 21192 14618 21220 14962
rect 21180 14612 21232 14618
rect 21180 14554 21232 14560
rect 21272 14544 21324 14550
rect 21272 14486 21324 14492
rect 21180 14408 21232 14414
rect 21180 14350 21232 14356
rect 21088 14340 21140 14346
rect 21088 14282 21140 14288
rect 20916 13938 20944 14214
rect 21008 14198 21128 14226
rect 20904 13932 20956 13938
rect 20904 13874 20956 13880
rect 20996 13728 21048 13734
rect 20996 13670 21048 13676
rect 20720 13388 20772 13394
rect 20720 13330 20772 13336
rect 21008 13326 21036 13670
rect 20996 13320 21048 13326
rect 20996 13262 21048 13268
rect 20628 13184 20680 13190
rect 20628 13126 20680 13132
rect 21100 12306 21128 14198
rect 21192 12986 21220 14350
rect 21284 14074 21312 14486
rect 21272 14068 21324 14074
rect 21272 14010 21324 14016
rect 21180 12980 21232 12986
rect 21180 12922 21232 12928
rect 21088 12300 21140 12306
rect 21088 12242 21140 12248
rect 20536 11756 20588 11762
rect 20536 11698 20588 11704
rect 20548 11665 20576 11698
rect 20534 11656 20590 11665
rect 20534 11591 20590 11600
rect 21270 11656 21326 11665
rect 21270 11591 21326 11600
rect 20536 11552 20588 11558
rect 20536 11494 20588 11500
rect 20364 10254 20484 10282
rect 20260 9580 20312 9586
rect 20260 9522 20312 9528
rect 20364 8378 20392 10254
rect 20548 10198 20576 11494
rect 20720 11212 20772 11218
rect 20720 11154 20772 11160
rect 20444 10192 20496 10198
rect 20444 10134 20496 10140
rect 20536 10192 20588 10198
rect 20536 10134 20588 10140
rect 20456 9518 20484 10134
rect 20444 9512 20496 9518
rect 20444 9454 20496 9460
rect 20456 8566 20484 9454
rect 20732 9330 20760 11154
rect 21284 10810 21312 11591
rect 21272 10804 21324 10810
rect 21272 10746 21324 10752
rect 20904 10736 20956 10742
rect 20904 10678 20956 10684
rect 20548 9302 20760 9330
rect 20444 8560 20496 8566
rect 20444 8502 20496 8508
rect 20272 8362 20392 8378
rect 20260 8356 20392 8362
rect 20312 8350 20392 8356
rect 20260 8298 20312 8304
rect 20352 8288 20404 8294
rect 20352 8230 20404 8236
rect 20364 8090 20392 8230
rect 20352 8084 20404 8090
rect 20352 8026 20404 8032
rect 20456 7546 20484 8502
rect 20444 7540 20496 7546
rect 20444 7482 20496 7488
rect 20168 5704 20220 5710
rect 20168 5646 20220 5652
rect 20076 4208 20128 4214
rect 20076 4150 20128 4156
rect 20548 4078 20576 9302
rect 20916 8922 20944 10678
rect 20996 10056 21048 10062
rect 20996 9998 21048 10004
rect 21008 9722 21036 9998
rect 20996 9716 21048 9722
rect 20996 9658 21048 9664
rect 20732 8894 20944 8922
rect 20996 8900 21048 8906
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 20640 8294 20668 8774
rect 20628 8288 20680 8294
rect 20628 8230 20680 8236
rect 20640 7954 20668 8230
rect 20628 7948 20680 7954
rect 20628 7890 20680 7896
rect 20732 7834 20760 8894
rect 20996 8842 21048 8848
rect 21180 8900 21232 8906
rect 21180 8842 21232 8848
rect 20812 8832 20864 8838
rect 20812 8774 20864 8780
rect 20824 8498 20852 8774
rect 21008 8498 21036 8842
rect 21192 8498 21220 8842
rect 20812 8492 20864 8498
rect 20812 8434 20864 8440
rect 20996 8492 21048 8498
rect 20996 8434 21048 8440
rect 21180 8492 21232 8498
rect 21180 8434 21232 8440
rect 20640 7806 20760 7834
rect 20640 4146 20668 7806
rect 20628 4140 20680 4146
rect 20628 4082 20680 4088
rect 20536 4072 20588 4078
rect 20536 4014 20588 4020
rect 19984 3936 20036 3942
rect 19984 3878 20036 3884
rect 19432 3664 19484 3670
rect 19432 3606 19484 3612
rect 19996 3602 20024 3878
rect 20352 3732 20404 3738
rect 20352 3674 20404 3680
rect 20364 3641 20392 3674
rect 20350 3632 20406 3641
rect 19984 3596 20036 3602
rect 20350 3567 20406 3576
rect 19984 3538 20036 3544
rect 19892 3528 19944 3534
rect 19890 3496 19892 3505
rect 19944 3496 19946 3505
rect 19890 3431 19946 3440
rect 20352 3460 20404 3466
rect 20352 3402 20404 3408
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 20364 3194 20392 3402
rect 20352 3188 20404 3194
rect 20352 3130 20404 3136
rect 20444 3188 20496 3194
rect 20444 3130 20496 3136
rect 20456 2854 20484 3130
rect 20548 3058 20576 4014
rect 20640 3720 20668 4082
rect 20812 3732 20864 3738
rect 20640 3692 20812 3720
rect 20812 3674 20864 3680
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 20536 3052 20588 3058
rect 20536 2994 20588 3000
rect 20444 2848 20496 2854
rect 20444 2790 20496 2796
rect 19984 2440 20036 2446
rect 19984 2382 20036 2388
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 19996 800 20024 2382
rect 20640 800 20668 3538
rect 21376 2650 21404 24074
rect 21468 22094 21496 37402
rect 21560 35698 21588 45358
rect 21640 38412 21692 38418
rect 21640 38354 21692 38360
rect 21548 35692 21600 35698
rect 21548 35634 21600 35640
rect 21652 34610 21680 38354
rect 21744 36922 21772 47602
rect 21824 40588 21876 40594
rect 21824 40530 21876 40536
rect 21836 39030 21864 40530
rect 22008 39296 22060 39302
rect 22008 39238 22060 39244
rect 21824 39024 21876 39030
rect 21824 38966 21876 38972
rect 21836 38554 21864 38966
rect 21824 38548 21876 38554
rect 21824 38490 21876 38496
rect 21836 37942 21864 38490
rect 21824 37936 21876 37942
rect 21824 37878 21876 37884
rect 21824 37664 21876 37670
rect 21824 37606 21876 37612
rect 21836 37262 21864 37606
rect 21824 37256 21876 37262
rect 21824 37198 21876 37204
rect 21916 37256 21968 37262
rect 21916 37198 21968 37204
rect 21732 36916 21784 36922
rect 21732 36858 21784 36864
rect 21928 36786 21956 37198
rect 21916 36780 21968 36786
rect 21916 36722 21968 36728
rect 21732 36100 21784 36106
rect 21732 36042 21784 36048
rect 21916 36100 21968 36106
rect 21916 36042 21968 36048
rect 21744 35834 21772 36042
rect 21732 35828 21784 35834
rect 21732 35770 21784 35776
rect 21732 35624 21784 35630
rect 21732 35566 21784 35572
rect 21744 34746 21772 35566
rect 21732 34740 21784 34746
rect 21732 34682 21784 34688
rect 21640 34604 21692 34610
rect 21640 34546 21692 34552
rect 21652 33522 21680 34546
rect 21824 34196 21876 34202
rect 21824 34138 21876 34144
rect 21640 33516 21692 33522
rect 21640 33458 21692 33464
rect 21652 31142 21680 33458
rect 21732 32768 21784 32774
rect 21732 32710 21784 32716
rect 21640 31136 21692 31142
rect 21640 31078 21692 31084
rect 21548 29844 21600 29850
rect 21548 29786 21600 29792
rect 21560 29510 21588 29786
rect 21652 29714 21680 31078
rect 21640 29708 21692 29714
rect 21640 29650 21692 29656
rect 21548 29504 21600 29510
rect 21548 29446 21600 29452
rect 21548 24608 21600 24614
rect 21548 24550 21600 24556
rect 21560 24138 21588 24550
rect 21548 24132 21600 24138
rect 21548 24074 21600 24080
rect 21468 22066 21680 22094
rect 21548 21888 21600 21894
rect 21548 21830 21600 21836
rect 21560 21146 21588 21830
rect 21548 21140 21600 21146
rect 21548 21082 21600 21088
rect 21548 21004 21600 21010
rect 21548 20946 21600 20952
rect 21560 20806 21588 20946
rect 21548 20800 21600 20806
rect 21548 20742 21600 20748
rect 21548 20460 21600 20466
rect 21548 20402 21600 20408
rect 21456 20052 21508 20058
rect 21456 19994 21508 20000
rect 21468 19718 21496 19994
rect 21456 19712 21508 19718
rect 21456 19654 21508 19660
rect 21456 18896 21508 18902
rect 21456 18838 21508 18844
rect 21468 16590 21496 18838
rect 21560 18834 21588 20402
rect 21652 20398 21680 22066
rect 21640 20392 21692 20398
rect 21640 20334 21692 20340
rect 21640 19916 21692 19922
rect 21640 19858 21692 19864
rect 21652 18902 21680 19858
rect 21640 18896 21692 18902
rect 21640 18838 21692 18844
rect 21548 18828 21600 18834
rect 21548 18770 21600 18776
rect 21640 18760 21692 18766
rect 21640 18702 21692 18708
rect 21548 18624 21600 18630
rect 21548 18566 21600 18572
rect 21560 18222 21588 18566
rect 21652 18426 21680 18702
rect 21640 18420 21692 18426
rect 21640 18362 21692 18368
rect 21548 18216 21600 18222
rect 21548 18158 21600 18164
rect 21640 17672 21692 17678
rect 21640 17614 21692 17620
rect 21652 17134 21680 17614
rect 21640 17128 21692 17134
rect 21640 17070 21692 17076
rect 21456 16584 21508 16590
rect 21456 16526 21508 16532
rect 21468 14890 21496 16526
rect 21640 15088 21692 15094
rect 21640 15030 21692 15036
rect 21456 14884 21508 14890
rect 21456 14826 21508 14832
rect 21456 14612 21508 14618
rect 21456 14554 21508 14560
rect 21468 13326 21496 14554
rect 21652 14278 21680 15030
rect 21640 14272 21692 14278
rect 21640 14214 21692 14220
rect 21652 13802 21680 14214
rect 21640 13796 21692 13802
rect 21640 13738 21692 13744
rect 21548 13728 21600 13734
rect 21548 13670 21600 13676
rect 21560 13394 21588 13670
rect 21652 13394 21680 13738
rect 21548 13388 21600 13394
rect 21548 13330 21600 13336
rect 21640 13388 21692 13394
rect 21640 13330 21692 13336
rect 21456 13320 21508 13326
rect 21456 13262 21508 13268
rect 21468 12782 21496 13262
rect 21560 12850 21588 13330
rect 21548 12844 21600 12850
rect 21548 12786 21600 12792
rect 21456 12776 21508 12782
rect 21456 12718 21508 12724
rect 21548 12232 21600 12238
rect 21548 12174 21600 12180
rect 21560 11898 21588 12174
rect 21548 11892 21600 11898
rect 21548 11834 21600 11840
rect 21744 10742 21772 32710
rect 21836 30122 21864 34138
rect 21928 31754 21956 36042
rect 22020 34202 22048 39238
rect 22008 34196 22060 34202
rect 22008 34138 22060 34144
rect 22008 32904 22060 32910
rect 22008 32846 22060 32852
rect 22020 32434 22048 32846
rect 22112 32774 22140 48486
rect 22204 47734 22232 49098
rect 22192 47728 22244 47734
rect 22192 47670 22244 47676
rect 22388 47666 22416 49234
rect 23400 49076 23428 51326
rect 23846 51326 24164 51354
rect 23846 51200 23902 51326
rect 23400 49048 23520 49076
rect 23492 48686 23520 49048
rect 22652 48680 22704 48686
rect 22652 48622 22704 48628
rect 22836 48680 22888 48686
rect 22836 48622 22888 48628
rect 23480 48680 23532 48686
rect 23480 48622 23532 48628
rect 22664 48142 22692 48622
rect 22848 48278 22876 48622
rect 22836 48272 22888 48278
rect 22836 48214 22888 48220
rect 22652 48136 22704 48142
rect 22652 48078 22704 48084
rect 22928 48068 22980 48074
rect 22928 48010 22980 48016
rect 22376 47660 22428 47666
rect 22376 47602 22428 47608
rect 22940 46646 22968 48010
rect 24136 47666 24164 51326
rect 24490 51326 24808 51354
rect 24490 51200 24546 51326
rect 24216 49360 24268 49366
rect 24216 49302 24268 49308
rect 24124 47660 24176 47666
rect 24124 47602 24176 47608
rect 23940 47456 23992 47462
rect 23940 47398 23992 47404
rect 22928 46640 22980 46646
rect 22928 46582 22980 46588
rect 22836 45824 22888 45830
rect 22836 45766 22888 45772
rect 22652 42560 22704 42566
rect 22652 42502 22704 42508
rect 22664 40526 22692 42502
rect 22652 40520 22704 40526
rect 22652 40462 22704 40468
rect 22468 40452 22520 40458
rect 22468 40394 22520 40400
rect 22376 40384 22428 40390
rect 22376 40326 22428 40332
rect 22388 40118 22416 40326
rect 22376 40112 22428 40118
rect 22376 40054 22428 40060
rect 22480 38554 22508 40394
rect 22652 40180 22704 40186
rect 22652 40122 22704 40128
rect 22664 39098 22692 40122
rect 22652 39092 22704 39098
rect 22652 39034 22704 39040
rect 22560 38956 22612 38962
rect 22560 38898 22612 38904
rect 22468 38548 22520 38554
rect 22468 38490 22520 38496
rect 22376 38276 22428 38282
rect 22376 38218 22428 38224
rect 22284 37868 22336 37874
rect 22284 37810 22336 37816
rect 22296 36922 22324 37810
rect 22388 37398 22416 38218
rect 22468 37868 22520 37874
rect 22468 37810 22520 37816
rect 22376 37392 22428 37398
rect 22376 37334 22428 37340
rect 22480 37262 22508 37810
rect 22572 37806 22600 38898
rect 22664 38570 22692 39034
rect 22664 38542 22784 38570
rect 22652 38412 22704 38418
rect 22652 38354 22704 38360
rect 22664 38214 22692 38354
rect 22756 38350 22784 38542
rect 22744 38344 22796 38350
rect 22744 38286 22796 38292
rect 22756 38214 22784 38286
rect 22652 38208 22704 38214
rect 22652 38150 22704 38156
rect 22744 38208 22796 38214
rect 22744 38150 22796 38156
rect 22560 37800 22612 37806
rect 22560 37742 22612 37748
rect 22468 37256 22520 37262
rect 22468 37198 22520 37204
rect 22376 37188 22428 37194
rect 22376 37130 22428 37136
rect 22388 36922 22416 37130
rect 22468 37120 22520 37126
rect 22468 37062 22520 37068
rect 22284 36916 22336 36922
rect 22284 36858 22336 36864
rect 22376 36916 22428 36922
rect 22376 36858 22428 36864
rect 22480 36786 22508 37062
rect 22468 36780 22520 36786
rect 22468 36722 22520 36728
rect 22572 36666 22600 37742
rect 22756 36802 22784 38150
rect 22664 36774 22784 36802
rect 22664 36718 22692 36774
rect 22388 36650 22600 36666
rect 22652 36712 22704 36718
rect 22652 36654 22704 36660
rect 22376 36644 22600 36650
rect 22428 36638 22600 36644
rect 22376 36586 22428 36592
rect 22192 36168 22244 36174
rect 22192 36110 22244 36116
rect 22204 34610 22232 36110
rect 22284 35760 22336 35766
rect 22284 35702 22336 35708
rect 22296 35562 22324 35702
rect 22284 35556 22336 35562
rect 22284 35498 22336 35504
rect 22284 34944 22336 34950
rect 22284 34886 22336 34892
rect 22296 34610 22324 34886
rect 22192 34604 22244 34610
rect 22192 34546 22244 34552
rect 22284 34604 22336 34610
rect 22284 34546 22336 34552
rect 22204 33590 22232 34546
rect 22192 33584 22244 33590
rect 22192 33526 22244 33532
rect 22284 32836 22336 32842
rect 22284 32778 22336 32784
rect 22100 32768 22152 32774
rect 22100 32710 22152 32716
rect 22008 32428 22060 32434
rect 22008 32370 22060 32376
rect 22296 32026 22324 32778
rect 22284 32020 22336 32026
rect 22284 31962 22336 31968
rect 21928 31726 22048 31754
rect 21916 30728 21968 30734
rect 21916 30670 21968 30676
rect 21928 30258 21956 30670
rect 21916 30252 21968 30258
rect 21916 30194 21968 30200
rect 21824 30116 21876 30122
rect 21824 30058 21876 30064
rect 21824 29572 21876 29578
rect 21824 29514 21876 29520
rect 21836 29170 21864 29514
rect 21824 29164 21876 29170
rect 21824 29106 21876 29112
rect 21928 25294 21956 30194
rect 21916 25288 21968 25294
rect 21916 25230 21968 25236
rect 21824 24812 21876 24818
rect 21824 24754 21876 24760
rect 21836 24721 21864 24754
rect 21822 24712 21878 24721
rect 21822 24647 21878 24656
rect 21916 24676 21968 24682
rect 21916 24618 21968 24624
rect 21824 24608 21876 24614
rect 21824 24550 21876 24556
rect 21836 23118 21864 24550
rect 21928 24177 21956 24618
rect 21914 24168 21970 24177
rect 21914 24103 21970 24112
rect 21824 23112 21876 23118
rect 21824 23054 21876 23060
rect 21916 22704 21968 22710
rect 21916 22646 21968 22652
rect 21928 22234 21956 22646
rect 21916 22228 21968 22234
rect 21916 22170 21968 22176
rect 21824 21412 21876 21418
rect 21824 21354 21876 21360
rect 21836 19174 21864 21354
rect 21916 19304 21968 19310
rect 21916 19246 21968 19252
rect 21824 19168 21876 19174
rect 21824 19110 21876 19116
rect 21824 18896 21876 18902
rect 21824 18838 21876 18844
rect 21836 18426 21864 18838
rect 21824 18420 21876 18426
rect 21824 18362 21876 18368
rect 21836 18290 21864 18362
rect 21928 18358 21956 19246
rect 21916 18352 21968 18358
rect 21916 18294 21968 18300
rect 21824 18284 21876 18290
rect 21824 18226 21876 18232
rect 21824 17332 21876 17338
rect 21824 17274 21876 17280
rect 21836 13433 21864 17274
rect 22020 15178 22048 31726
rect 22100 31748 22152 31754
rect 22100 31690 22152 31696
rect 22112 31278 22140 31690
rect 22100 31272 22152 31278
rect 22100 31214 22152 31220
rect 22388 30054 22416 36586
rect 22664 36242 22692 36654
rect 22652 36236 22704 36242
rect 22652 36178 22704 36184
rect 22560 35148 22612 35154
rect 22560 35090 22612 35096
rect 22468 33856 22520 33862
rect 22468 33798 22520 33804
rect 22480 31822 22508 33798
rect 22468 31816 22520 31822
rect 22468 31758 22520 31764
rect 22468 30728 22520 30734
rect 22468 30670 22520 30676
rect 22480 30190 22508 30670
rect 22468 30184 22520 30190
rect 22468 30126 22520 30132
rect 22376 30048 22428 30054
rect 22376 29990 22428 29996
rect 22376 29640 22428 29646
rect 22376 29582 22428 29588
rect 22388 29238 22416 29582
rect 22376 29232 22428 29238
rect 22376 29174 22428 29180
rect 22480 29102 22508 30126
rect 22468 29096 22520 29102
rect 22468 29038 22520 29044
rect 22468 25152 22520 25158
rect 22468 25094 22520 25100
rect 22192 24200 22244 24206
rect 22192 24142 22244 24148
rect 22204 23254 22232 24142
rect 22192 23248 22244 23254
rect 22192 23190 22244 23196
rect 22192 22432 22244 22438
rect 22192 22374 22244 22380
rect 22204 21962 22232 22374
rect 22192 21956 22244 21962
rect 22192 21898 22244 21904
rect 22376 21548 22428 21554
rect 22376 21490 22428 21496
rect 22100 21344 22152 21350
rect 22098 21312 22100 21321
rect 22284 21344 22336 21350
rect 22152 21312 22154 21321
rect 22284 21286 22336 21292
rect 22098 21247 22154 21256
rect 22112 19417 22140 21247
rect 22192 21004 22244 21010
rect 22192 20946 22244 20952
rect 22204 19990 22232 20946
rect 22296 20924 22324 21286
rect 22388 21146 22416 21490
rect 22376 21140 22428 21146
rect 22376 21082 22428 21088
rect 22376 20936 22428 20942
rect 22296 20896 22376 20924
rect 22296 20534 22324 20896
rect 22376 20878 22428 20884
rect 22284 20528 22336 20534
rect 22284 20470 22336 20476
rect 22284 20256 22336 20262
rect 22284 20198 22336 20204
rect 22192 19984 22244 19990
rect 22192 19926 22244 19932
rect 22296 19922 22324 20198
rect 22284 19916 22336 19922
rect 22284 19858 22336 19864
rect 22284 19712 22336 19718
rect 22284 19654 22336 19660
rect 22296 19514 22324 19654
rect 22284 19508 22336 19514
rect 22284 19450 22336 19456
rect 22098 19408 22154 19417
rect 22098 19343 22154 19352
rect 22376 19168 22428 19174
rect 22376 19110 22428 19116
rect 22100 18624 22152 18630
rect 22100 18566 22152 18572
rect 22112 18290 22140 18566
rect 22100 18284 22152 18290
rect 22100 18226 22152 18232
rect 22284 18216 22336 18222
rect 22284 18158 22336 18164
rect 22192 18080 22244 18086
rect 22192 18022 22244 18028
rect 22100 17672 22152 17678
rect 22100 17614 22152 17620
rect 22112 17338 22140 17614
rect 22100 17332 22152 17338
rect 22100 17274 22152 17280
rect 22204 17202 22232 18022
rect 22296 17882 22324 18158
rect 22284 17876 22336 17882
rect 22284 17818 22336 17824
rect 22282 17776 22338 17785
rect 22282 17711 22338 17720
rect 22296 17542 22324 17711
rect 22388 17678 22416 19110
rect 22376 17672 22428 17678
rect 22376 17614 22428 17620
rect 22284 17536 22336 17542
rect 22284 17478 22336 17484
rect 22192 17196 22244 17202
rect 22192 17138 22244 17144
rect 22192 15360 22244 15366
rect 22192 15302 22244 15308
rect 21928 15150 22048 15178
rect 22204 15162 22232 15302
rect 22192 15156 22244 15162
rect 21822 13424 21878 13433
rect 21822 13359 21878 13368
rect 21824 13252 21876 13258
rect 21824 13194 21876 13200
rect 21836 12306 21864 13194
rect 21824 12300 21876 12306
rect 21824 12242 21876 12248
rect 21836 11830 21864 12242
rect 21824 11824 21876 11830
rect 21824 11766 21876 11772
rect 21836 11354 21864 11766
rect 21824 11348 21876 11354
rect 21824 11290 21876 11296
rect 21732 10736 21784 10742
rect 21732 10678 21784 10684
rect 21548 8560 21600 8566
rect 21548 8502 21600 8508
rect 21560 8294 21588 8502
rect 21928 8480 21956 15150
rect 22192 15098 22244 15104
rect 22100 15088 22152 15094
rect 22100 15030 22152 15036
rect 22008 14340 22060 14346
rect 22008 14282 22060 14288
rect 22020 14090 22048 14282
rect 22112 14260 22140 15030
rect 22204 14958 22232 15098
rect 22192 14952 22244 14958
rect 22192 14894 22244 14900
rect 22296 14890 22324 17478
rect 22480 17218 22508 25094
rect 22388 17190 22508 17218
rect 22284 14884 22336 14890
rect 22284 14826 22336 14832
rect 22192 14272 22244 14278
rect 22112 14232 22192 14260
rect 22192 14214 22244 14220
rect 22020 14062 22140 14090
rect 22008 14000 22060 14006
rect 22008 13942 22060 13948
rect 22020 11150 22048 13942
rect 22008 11144 22060 11150
rect 22008 11086 22060 11092
rect 21652 8452 21956 8480
rect 22020 8514 22048 11086
rect 22112 9926 22140 14062
rect 22204 12646 22232 14214
rect 22284 13864 22336 13870
rect 22284 13806 22336 13812
rect 22296 13530 22324 13806
rect 22284 13524 22336 13530
rect 22284 13466 22336 13472
rect 22192 12640 22244 12646
rect 22192 12582 22244 12588
rect 22192 12232 22244 12238
rect 22192 12174 22244 12180
rect 22204 11762 22232 12174
rect 22284 12096 22336 12102
rect 22284 12038 22336 12044
rect 22192 11756 22244 11762
rect 22192 11698 22244 11704
rect 22204 10538 22232 11698
rect 22296 11082 22324 12038
rect 22284 11076 22336 11082
rect 22284 11018 22336 11024
rect 22192 10532 22244 10538
rect 22192 10474 22244 10480
rect 22100 9920 22152 9926
rect 22100 9862 22152 9868
rect 22388 9178 22416 17190
rect 22572 17066 22600 35090
rect 22652 33516 22704 33522
rect 22652 33458 22704 33464
rect 22664 24410 22692 33458
rect 22744 31204 22796 31210
rect 22744 31146 22796 31152
rect 22756 29850 22784 31146
rect 22744 29844 22796 29850
rect 22744 29786 22796 29792
rect 22756 29170 22784 29786
rect 22744 29164 22796 29170
rect 22744 29106 22796 29112
rect 22848 28694 22876 45766
rect 22940 38418 22968 46582
rect 23388 40588 23440 40594
rect 23388 40530 23440 40536
rect 23112 40044 23164 40050
rect 23112 39986 23164 39992
rect 23124 39642 23152 39986
rect 23112 39636 23164 39642
rect 23112 39578 23164 39584
rect 23400 39574 23428 40530
rect 23848 40520 23900 40526
rect 23848 40462 23900 40468
rect 23664 39976 23716 39982
rect 23664 39918 23716 39924
rect 23388 39568 23440 39574
rect 23388 39510 23440 39516
rect 23676 39506 23704 39918
rect 23756 39568 23808 39574
rect 23756 39510 23808 39516
rect 23664 39500 23716 39506
rect 23664 39442 23716 39448
rect 23572 39432 23624 39438
rect 23216 39392 23572 39420
rect 23020 39296 23072 39302
rect 23020 39238 23072 39244
rect 23032 38962 23060 39238
rect 23020 38956 23072 38962
rect 23020 38898 23072 38904
rect 23216 38894 23244 39392
rect 23572 39374 23624 39380
rect 23664 39364 23716 39370
rect 23664 39306 23716 39312
rect 23478 39128 23534 39137
rect 23296 39092 23348 39098
rect 23478 39063 23480 39072
rect 23296 39034 23348 39040
rect 23532 39063 23534 39072
rect 23480 39034 23532 39040
rect 23308 38978 23336 39034
rect 23676 38978 23704 39306
rect 23308 38950 23704 38978
rect 23768 38894 23796 39510
rect 23860 39438 23888 40462
rect 23952 39642 23980 47398
rect 24124 41608 24176 41614
rect 24124 41550 24176 41556
rect 24032 40180 24084 40186
rect 24032 40122 24084 40128
rect 23940 39636 23992 39642
rect 23940 39578 23992 39584
rect 23848 39432 23900 39438
rect 23848 39374 23900 39380
rect 23204 38888 23256 38894
rect 23204 38830 23256 38836
rect 23756 38888 23808 38894
rect 23756 38830 23808 38836
rect 23860 38826 23888 39374
rect 23940 39024 23992 39030
rect 23940 38966 23992 38972
rect 23848 38820 23900 38826
rect 23848 38762 23900 38768
rect 23952 38486 23980 38966
rect 23940 38480 23992 38486
rect 23940 38422 23992 38428
rect 24044 38418 24072 40122
rect 22928 38412 22980 38418
rect 22928 38354 22980 38360
rect 24032 38412 24084 38418
rect 24032 38354 24084 38360
rect 23480 38344 23532 38350
rect 23400 38304 23480 38332
rect 23020 37868 23072 37874
rect 23020 37810 23072 37816
rect 23204 37868 23256 37874
rect 23204 37810 23256 37816
rect 23032 37466 23060 37810
rect 23020 37460 23072 37466
rect 23020 37402 23072 37408
rect 23020 36780 23072 36786
rect 23020 36722 23072 36728
rect 23032 35834 23060 36722
rect 23020 35828 23072 35834
rect 23020 35770 23072 35776
rect 23216 34950 23244 37810
rect 23400 37806 23428 38304
rect 23480 38286 23532 38292
rect 23388 37800 23440 37806
rect 23388 37742 23440 37748
rect 23388 37664 23440 37670
rect 23388 37606 23440 37612
rect 23296 36168 23348 36174
rect 23296 36110 23348 36116
rect 23308 35698 23336 36110
rect 23400 35698 23428 37606
rect 23572 37324 23624 37330
rect 23572 37266 23624 37272
rect 23584 37194 23612 37266
rect 23572 37188 23624 37194
rect 23572 37130 23624 37136
rect 23296 35692 23348 35698
rect 23296 35634 23348 35640
rect 23388 35692 23440 35698
rect 23388 35634 23440 35640
rect 23584 35494 23612 37130
rect 24044 35698 24072 38354
rect 24032 35692 24084 35698
rect 24032 35634 24084 35640
rect 23756 35624 23808 35630
rect 23756 35566 23808 35572
rect 23572 35488 23624 35494
rect 23572 35430 23624 35436
rect 23296 35080 23348 35086
rect 23296 35022 23348 35028
rect 22928 34944 22980 34950
rect 22928 34886 22980 34892
rect 23204 34944 23256 34950
rect 23204 34886 23256 34892
rect 22940 33930 22968 34886
rect 23020 34400 23072 34406
rect 23020 34342 23072 34348
rect 23032 33998 23060 34342
rect 23020 33992 23072 33998
rect 23020 33934 23072 33940
rect 22928 33924 22980 33930
rect 22928 33866 22980 33872
rect 23112 32428 23164 32434
rect 23112 32370 23164 32376
rect 23124 32026 23152 32370
rect 23112 32020 23164 32026
rect 23112 31962 23164 31968
rect 22928 31884 22980 31890
rect 22928 31826 22980 31832
rect 22940 30802 22968 31826
rect 23308 31210 23336 35022
rect 23572 34604 23624 34610
rect 23572 34546 23624 34552
rect 23480 34536 23532 34542
rect 23480 34478 23532 34484
rect 23492 34202 23520 34478
rect 23480 34196 23532 34202
rect 23480 34138 23532 34144
rect 23584 32774 23612 34546
rect 23572 32768 23624 32774
rect 23572 32710 23624 32716
rect 23388 32224 23440 32230
rect 23388 32166 23440 32172
rect 23480 32224 23532 32230
rect 23480 32166 23532 32172
rect 23400 31822 23428 32166
rect 23388 31816 23440 31822
rect 23388 31758 23440 31764
rect 23492 31346 23520 32166
rect 23572 31816 23624 31822
rect 23572 31758 23624 31764
rect 23584 31482 23612 31758
rect 23572 31476 23624 31482
rect 23572 31418 23624 31424
rect 23388 31340 23440 31346
rect 23388 31282 23440 31288
rect 23480 31340 23532 31346
rect 23480 31282 23532 31288
rect 23400 31226 23428 31282
rect 23296 31204 23348 31210
rect 23400 31198 23520 31226
rect 23296 31146 23348 31152
rect 23388 31136 23440 31142
rect 23388 31078 23440 31084
rect 22928 30796 22980 30802
rect 22928 30738 22980 30744
rect 22940 30394 22968 30738
rect 23400 30734 23428 31078
rect 23388 30728 23440 30734
rect 23388 30670 23440 30676
rect 23492 30666 23520 31198
rect 23480 30660 23532 30666
rect 23480 30602 23532 30608
rect 22928 30388 22980 30394
rect 22928 30330 22980 30336
rect 23492 30258 23520 30602
rect 23204 30252 23256 30258
rect 23204 30194 23256 30200
rect 23480 30252 23532 30258
rect 23480 30194 23532 30200
rect 23112 30048 23164 30054
rect 23112 29990 23164 29996
rect 23124 29646 23152 29990
rect 23112 29640 23164 29646
rect 23112 29582 23164 29588
rect 23216 29306 23244 30194
rect 23768 30054 23796 35566
rect 23940 35012 23992 35018
rect 23940 34954 23992 34960
rect 23848 34672 23900 34678
rect 23848 34614 23900 34620
rect 23860 34134 23888 34614
rect 23848 34128 23900 34134
rect 23848 34070 23900 34076
rect 23848 33380 23900 33386
rect 23848 33322 23900 33328
rect 23860 32502 23888 33322
rect 23848 32496 23900 32502
rect 23848 32438 23900 32444
rect 23664 30048 23716 30054
rect 23664 29990 23716 29996
rect 23756 30048 23808 30054
rect 23756 29990 23808 29996
rect 23676 29578 23704 29990
rect 23768 29646 23796 29990
rect 23756 29640 23808 29646
rect 23756 29582 23808 29588
rect 23664 29572 23716 29578
rect 23664 29514 23716 29520
rect 23388 29504 23440 29510
rect 23386 29472 23388 29481
rect 23756 29504 23808 29510
rect 23440 29472 23442 29481
rect 23756 29446 23808 29452
rect 23386 29407 23442 29416
rect 23204 29300 23256 29306
rect 23204 29242 23256 29248
rect 23768 29170 23796 29446
rect 23756 29164 23808 29170
rect 23756 29106 23808 29112
rect 23480 28756 23532 28762
rect 23480 28698 23532 28704
rect 22836 28688 22888 28694
rect 22836 28630 22888 28636
rect 23204 28416 23256 28422
rect 23204 28358 23256 28364
rect 23216 28150 23244 28358
rect 23204 28144 23256 28150
rect 23204 28086 23256 28092
rect 23492 28014 23520 28698
rect 23480 28008 23532 28014
rect 23480 27950 23532 27956
rect 22928 27396 22980 27402
rect 22928 27338 22980 27344
rect 22940 27130 22968 27338
rect 23204 27328 23256 27334
rect 23204 27270 23256 27276
rect 22928 27124 22980 27130
rect 22928 27066 22980 27072
rect 23216 26994 23244 27270
rect 23204 26988 23256 26994
rect 23204 26930 23256 26936
rect 23572 26444 23624 26450
rect 23572 26386 23624 26392
rect 22928 25968 22980 25974
rect 22928 25910 22980 25916
rect 22940 25158 22968 25910
rect 23112 25832 23164 25838
rect 23112 25774 23164 25780
rect 22928 25152 22980 25158
rect 22928 25094 22980 25100
rect 23124 24993 23152 25774
rect 23584 25498 23612 26386
rect 23952 26042 23980 34954
rect 24044 32366 24072 35634
rect 24032 32360 24084 32366
rect 24032 32302 24084 32308
rect 24136 31754 24164 41550
rect 24228 38350 24256 49302
rect 24780 49298 24808 51326
rect 25134 51200 25190 52000
rect 25778 51354 25834 52000
rect 25778 51326 26004 51354
rect 25778 51200 25834 51326
rect 24768 49292 24820 49298
rect 24768 49234 24820 49240
rect 24584 49156 24636 49162
rect 24584 49098 24636 49104
rect 24596 48278 24624 49098
rect 25228 49088 25280 49094
rect 25228 49030 25280 49036
rect 25320 49088 25372 49094
rect 25320 49030 25372 49036
rect 24952 48544 25004 48550
rect 24952 48486 25004 48492
rect 24584 48272 24636 48278
rect 24584 48214 24636 48220
rect 24400 48136 24452 48142
rect 24400 48078 24452 48084
rect 24412 48006 24440 48078
rect 24400 48000 24452 48006
rect 24400 47942 24452 47948
rect 24412 39846 24440 47942
rect 24400 39840 24452 39846
rect 24400 39782 24452 39788
rect 24216 38344 24268 38350
rect 24216 38286 24268 38292
rect 24860 37868 24912 37874
rect 24860 37810 24912 37816
rect 24872 37262 24900 37810
rect 24860 37256 24912 37262
rect 24860 37198 24912 37204
rect 24676 37188 24728 37194
rect 24676 37130 24728 37136
rect 24688 36922 24716 37130
rect 24860 37120 24912 37126
rect 24860 37062 24912 37068
rect 24676 36916 24728 36922
rect 24676 36858 24728 36864
rect 24308 36712 24360 36718
rect 24308 36654 24360 36660
rect 24320 35698 24348 36654
rect 24872 36582 24900 37062
rect 24860 36576 24912 36582
rect 24860 36518 24912 36524
rect 24860 36304 24912 36310
rect 24860 36246 24912 36252
rect 24872 35834 24900 36246
rect 24860 35828 24912 35834
rect 24860 35770 24912 35776
rect 24308 35692 24360 35698
rect 24308 35634 24360 35640
rect 24492 35488 24544 35494
rect 24492 35430 24544 35436
rect 24584 35488 24636 35494
rect 24584 35430 24636 35436
rect 24400 34944 24452 34950
rect 24400 34886 24452 34892
rect 24216 34604 24268 34610
rect 24216 34546 24268 34552
rect 24228 33454 24256 34546
rect 24412 34474 24440 34886
rect 24400 34468 24452 34474
rect 24400 34410 24452 34416
rect 24504 34406 24532 35430
rect 24596 35154 24624 35430
rect 24584 35148 24636 35154
rect 24584 35090 24636 35096
rect 24584 34604 24636 34610
rect 24584 34546 24636 34552
rect 24308 34400 24360 34406
rect 24308 34342 24360 34348
rect 24492 34400 24544 34406
rect 24492 34342 24544 34348
rect 24216 33448 24268 33454
rect 24216 33390 24268 33396
rect 24228 32348 24256 33390
rect 24320 32502 24348 34342
rect 24596 34202 24624 34546
rect 24860 34536 24912 34542
rect 24860 34478 24912 34484
rect 24872 34202 24900 34478
rect 24584 34196 24636 34202
rect 24584 34138 24636 34144
rect 24860 34196 24912 34202
rect 24860 34138 24912 34144
rect 24768 33992 24820 33998
rect 24766 33960 24768 33969
rect 24820 33960 24822 33969
rect 24688 33918 24766 33946
rect 24308 32496 24360 32502
rect 24308 32438 24360 32444
rect 24228 32320 24440 32348
rect 24032 31748 24084 31754
rect 24136 31726 24256 31754
rect 24032 31690 24084 31696
rect 24044 30802 24072 31690
rect 24032 30796 24084 30802
rect 24032 30738 24084 30744
rect 24044 30394 24072 30738
rect 24032 30388 24084 30394
rect 24032 30330 24084 30336
rect 24124 30252 24176 30258
rect 24124 30194 24176 30200
rect 24136 29850 24164 30194
rect 24124 29844 24176 29850
rect 24124 29786 24176 29792
rect 24032 29776 24084 29782
rect 24032 29718 24084 29724
rect 24044 29510 24072 29718
rect 24032 29504 24084 29510
rect 24032 29446 24084 29452
rect 23940 26036 23992 26042
rect 23940 25978 23992 25984
rect 23848 25900 23900 25906
rect 23848 25842 23900 25848
rect 24032 25900 24084 25906
rect 24032 25842 24084 25848
rect 23754 25528 23810 25537
rect 23572 25492 23624 25498
rect 23754 25463 23756 25472
rect 23572 25434 23624 25440
rect 23808 25463 23810 25472
rect 23756 25434 23808 25440
rect 23584 25242 23612 25434
rect 23400 25226 23520 25242
rect 23388 25220 23520 25226
rect 23440 25214 23520 25220
rect 23584 25214 23796 25242
rect 23388 25162 23440 25168
rect 23110 24984 23166 24993
rect 23110 24919 23166 24928
rect 22744 24744 22796 24750
rect 22744 24686 22796 24692
rect 22652 24404 22704 24410
rect 22652 24346 22704 24352
rect 22560 17060 22612 17066
rect 22560 17002 22612 17008
rect 22560 15700 22612 15706
rect 22560 15642 22612 15648
rect 22572 15162 22600 15642
rect 22560 15156 22612 15162
rect 22560 15098 22612 15104
rect 22468 14340 22520 14346
rect 22468 14282 22520 14288
rect 22480 14074 22508 14282
rect 22468 14068 22520 14074
rect 22468 14010 22520 14016
rect 22480 13326 22508 14010
rect 22468 13320 22520 13326
rect 22468 13262 22520 13268
rect 22664 12918 22692 24346
rect 22756 24206 22784 24686
rect 23492 24614 23520 25214
rect 23572 25152 23624 25158
rect 23572 25094 23624 25100
rect 23584 24954 23612 25094
rect 23572 24948 23624 24954
rect 23572 24890 23624 24896
rect 23480 24608 23532 24614
rect 23480 24550 23532 24556
rect 23296 24336 23348 24342
rect 23296 24278 23348 24284
rect 22744 24200 22796 24206
rect 22744 24142 22796 24148
rect 23112 23588 23164 23594
rect 23112 23530 23164 23536
rect 23124 23322 23152 23530
rect 23308 23508 23336 24278
rect 23492 23798 23520 24550
rect 23664 24200 23716 24206
rect 23664 24142 23716 24148
rect 23480 23792 23532 23798
rect 23480 23734 23532 23740
rect 23676 23730 23704 24142
rect 23664 23724 23716 23730
rect 23664 23666 23716 23672
rect 23388 23520 23440 23526
rect 23308 23488 23388 23508
rect 23480 23520 23532 23526
rect 23440 23488 23442 23497
rect 23308 23480 23386 23488
rect 23480 23462 23532 23468
rect 23386 23423 23442 23432
rect 23020 23316 23072 23322
rect 23020 23258 23072 23264
rect 23112 23316 23164 23322
rect 23112 23258 23164 23264
rect 23032 22234 23060 23258
rect 23204 23248 23256 23254
rect 23204 23190 23256 23196
rect 23020 22228 23072 22234
rect 23020 22170 23072 22176
rect 22744 21956 22796 21962
rect 22744 21898 22796 21904
rect 22756 21622 22784 21898
rect 22744 21616 22796 21622
rect 22744 21558 22796 21564
rect 23112 21616 23164 21622
rect 23112 21558 23164 21564
rect 22756 19378 22784 21558
rect 23124 21418 23152 21558
rect 23112 21412 23164 21418
rect 23112 21354 23164 21360
rect 23112 20936 23164 20942
rect 23112 20878 23164 20884
rect 23020 19848 23072 19854
rect 23020 19790 23072 19796
rect 22744 19372 22796 19378
rect 22744 19314 22796 19320
rect 23032 19242 23060 19790
rect 23020 19236 23072 19242
rect 23020 19178 23072 19184
rect 23124 18902 23152 20878
rect 23112 18896 23164 18902
rect 23112 18838 23164 18844
rect 23020 18352 23072 18358
rect 23020 18294 23072 18300
rect 23032 17814 23060 18294
rect 23112 18080 23164 18086
rect 23112 18022 23164 18028
rect 23124 17814 23152 18022
rect 23020 17808 23072 17814
rect 23020 17750 23072 17756
rect 23112 17808 23164 17814
rect 23112 17750 23164 17756
rect 22928 17672 22980 17678
rect 22928 17614 22980 17620
rect 22940 17270 22968 17614
rect 23112 17604 23164 17610
rect 23112 17546 23164 17552
rect 22928 17264 22980 17270
rect 22928 17206 22980 17212
rect 23020 17264 23072 17270
rect 23020 17206 23072 17212
rect 23032 16658 23060 17206
rect 23124 17202 23152 17546
rect 23112 17196 23164 17202
rect 23112 17138 23164 17144
rect 23020 16652 23072 16658
rect 23020 16594 23072 16600
rect 23020 15904 23072 15910
rect 23020 15846 23072 15852
rect 22928 14952 22980 14958
rect 22928 14894 22980 14900
rect 22744 14476 22796 14482
rect 22744 14418 22796 14424
rect 22652 12912 22704 12918
rect 22652 12854 22704 12860
rect 22468 12844 22520 12850
rect 22468 12786 22520 12792
rect 22480 11626 22508 12786
rect 22560 12708 22612 12714
rect 22560 12650 22612 12656
rect 22572 12374 22600 12650
rect 22560 12368 22612 12374
rect 22560 12310 22612 12316
rect 22652 12096 22704 12102
rect 22652 12038 22704 12044
rect 22468 11620 22520 11626
rect 22468 11562 22520 11568
rect 22664 11558 22692 12038
rect 22756 11694 22784 14418
rect 22836 14272 22888 14278
rect 22836 14214 22888 14220
rect 22848 13462 22876 14214
rect 22836 13456 22888 13462
rect 22836 13398 22888 13404
rect 22940 12850 22968 14894
rect 22928 12844 22980 12850
rect 22928 12786 22980 12792
rect 23032 12306 23060 15846
rect 23112 14612 23164 14618
rect 23112 14554 23164 14560
rect 23124 14414 23152 14554
rect 23112 14408 23164 14414
rect 23112 14350 23164 14356
rect 23020 12300 23072 12306
rect 23020 12242 23072 12248
rect 22744 11688 22796 11694
rect 22744 11630 22796 11636
rect 22756 11558 22784 11630
rect 22652 11552 22704 11558
rect 22652 11494 22704 11500
rect 22744 11552 22796 11558
rect 22744 11494 22796 11500
rect 23032 10470 23060 12242
rect 23216 12238 23244 23190
rect 23492 23118 23520 23462
rect 23572 23316 23624 23322
rect 23572 23258 23624 23264
rect 23480 23112 23532 23118
rect 23480 23054 23532 23060
rect 23584 22794 23612 23258
rect 23492 22766 23612 22794
rect 23492 22642 23520 22766
rect 23480 22636 23532 22642
rect 23480 22578 23532 22584
rect 23296 22092 23348 22098
rect 23296 22034 23348 22040
rect 23308 21350 23336 22034
rect 23388 21888 23440 21894
rect 23388 21830 23440 21836
rect 23296 21344 23348 21350
rect 23296 21286 23348 21292
rect 23308 21146 23336 21286
rect 23296 21140 23348 21146
rect 23296 21082 23348 21088
rect 23308 20602 23336 21082
rect 23296 20596 23348 20602
rect 23296 20538 23348 20544
rect 23308 19378 23336 20538
rect 23296 19372 23348 19378
rect 23296 19314 23348 19320
rect 23400 19310 23428 21830
rect 23492 21010 23520 22578
rect 23572 22500 23624 22506
rect 23572 22442 23624 22448
rect 23480 21004 23532 21010
rect 23480 20946 23532 20952
rect 23480 20800 23532 20806
rect 23480 20742 23532 20748
rect 23492 19854 23520 20742
rect 23480 19848 23532 19854
rect 23480 19790 23532 19796
rect 23492 19446 23520 19790
rect 23480 19440 23532 19446
rect 23480 19382 23532 19388
rect 23388 19304 23440 19310
rect 23388 19246 23440 19252
rect 23492 18766 23520 19382
rect 23388 18760 23440 18766
rect 23388 18702 23440 18708
rect 23480 18760 23532 18766
rect 23480 18702 23532 18708
rect 23296 18148 23348 18154
rect 23296 18090 23348 18096
rect 23308 17134 23336 18090
rect 23400 18086 23428 18702
rect 23584 18170 23612 22442
rect 23768 20913 23796 25214
rect 23860 24993 23888 25842
rect 23940 25696 23992 25702
rect 23940 25638 23992 25644
rect 23952 25430 23980 25638
rect 23940 25424 23992 25430
rect 23940 25366 23992 25372
rect 23846 24984 23902 24993
rect 23846 24919 23902 24928
rect 23940 24812 23992 24818
rect 23940 24754 23992 24760
rect 23952 24342 23980 24754
rect 23940 24336 23992 24342
rect 23940 24278 23992 24284
rect 23848 24132 23900 24138
rect 23848 24074 23900 24080
rect 23754 20904 23810 20913
rect 23754 20839 23810 20848
rect 23664 20800 23716 20806
rect 23664 20742 23716 20748
rect 23756 20800 23808 20806
rect 23756 20742 23808 20748
rect 23676 20466 23704 20742
rect 23664 20460 23716 20466
rect 23664 20402 23716 20408
rect 23662 20360 23718 20369
rect 23662 20295 23718 20304
rect 23676 18426 23704 20295
rect 23768 19922 23796 20742
rect 23756 19916 23808 19922
rect 23756 19858 23808 19864
rect 23664 18420 23716 18426
rect 23664 18362 23716 18368
rect 23584 18142 23796 18170
rect 23388 18080 23440 18086
rect 23388 18022 23440 18028
rect 23572 18080 23624 18086
rect 23572 18022 23624 18028
rect 23480 17876 23532 17882
rect 23480 17818 23532 17824
rect 23296 17128 23348 17134
rect 23296 17070 23348 17076
rect 23492 16998 23520 17818
rect 23584 17202 23612 18022
rect 23572 17196 23624 17202
rect 23572 17138 23624 17144
rect 23480 16992 23532 16998
rect 23480 16934 23532 16940
rect 23664 16992 23716 16998
rect 23664 16934 23716 16940
rect 23388 15088 23440 15094
rect 23388 15030 23440 15036
rect 23296 14340 23348 14346
rect 23296 14282 23348 14288
rect 23308 14006 23336 14282
rect 23400 14074 23428 15030
rect 23492 14906 23520 16934
rect 23676 16590 23704 16934
rect 23664 16584 23716 16590
rect 23664 16526 23716 16532
rect 23572 15360 23624 15366
rect 23572 15302 23624 15308
rect 23664 15360 23716 15366
rect 23664 15302 23716 15308
rect 23584 15026 23612 15302
rect 23572 15020 23624 15026
rect 23572 14962 23624 14968
rect 23492 14878 23612 14906
rect 23480 14816 23532 14822
rect 23480 14758 23532 14764
rect 23388 14068 23440 14074
rect 23388 14010 23440 14016
rect 23296 14000 23348 14006
rect 23296 13942 23348 13948
rect 23492 13938 23520 14758
rect 23480 13932 23532 13938
rect 23480 13874 23532 13880
rect 23584 13530 23612 14878
rect 23676 14550 23704 15302
rect 23664 14544 23716 14550
rect 23664 14486 23716 14492
rect 23664 14000 23716 14006
rect 23664 13942 23716 13948
rect 23572 13524 23624 13530
rect 23572 13466 23624 13472
rect 23676 13410 23704 13942
rect 23584 13382 23704 13410
rect 23296 13252 23348 13258
rect 23296 13194 23348 13200
rect 23308 12986 23336 13194
rect 23296 12980 23348 12986
rect 23296 12922 23348 12928
rect 23388 12436 23440 12442
rect 23388 12378 23440 12384
rect 23204 12232 23256 12238
rect 23204 12174 23256 12180
rect 23400 10674 23428 12378
rect 23480 12164 23532 12170
rect 23480 12106 23532 12112
rect 23492 11354 23520 12106
rect 23480 11348 23532 11354
rect 23480 11290 23532 11296
rect 23388 10668 23440 10674
rect 23388 10610 23440 10616
rect 23492 10606 23520 11290
rect 23480 10600 23532 10606
rect 23480 10542 23532 10548
rect 23020 10464 23072 10470
rect 23020 10406 23072 10412
rect 23388 9512 23440 9518
rect 23388 9454 23440 9460
rect 22376 9172 22428 9178
rect 22376 9114 22428 9120
rect 22928 8968 22980 8974
rect 22928 8910 22980 8916
rect 23296 8968 23348 8974
rect 23296 8910 23348 8916
rect 22192 8900 22244 8906
rect 22192 8842 22244 8848
rect 22100 8560 22152 8566
rect 22020 8508 22100 8514
rect 22020 8502 22152 8508
rect 22020 8486 22140 8502
rect 21548 8288 21600 8294
rect 21548 8230 21600 8236
rect 21364 2644 21416 2650
rect 21364 2586 21416 2592
rect 21284 870 21404 898
rect 21284 800 21312 870
rect 13188 734 13492 762
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 21376 762 21404 870
rect 21652 762 21680 8452
rect 21824 8356 21876 8362
rect 21824 8298 21876 8304
rect 21916 8356 21968 8362
rect 21916 8298 21968 8304
rect 21836 7546 21864 8298
rect 21824 7540 21876 7546
rect 21824 7482 21876 7488
rect 21928 7478 21956 8298
rect 22020 7750 22048 8486
rect 22204 8242 22232 8842
rect 22284 8288 22336 8294
rect 22204 8236 22284 8242
rect 22204 8230 22336 8236
rect 22204 8214 22324 8230
rect 22008 7744 22060 7750
rect 22008 7686 22060 7692
rect 21916 7472 21968 7478
rect 21916 7414 21968 7420
rect 22020 7410 22048 7686
rect 22008 7404 22060 7410
rect 22008 7346 22060 7352
rect 22204 7342 22232 8214
rect 22940 8090 22968 8910
rect 23204 8832 23256 8838
rect 23204 8774 23256 8780
rect 23112 8560 23164 8566
rect 23112 8502 23164 8508
rect 22928 8084 22980 8090
rect 22928 8026 22980 8032
rect 23020 7880 23072 7886
rect 23020 7822 23072 7828
rect 22192 7336 22244 7342
rect 22192 7278 22244 7284
rect 22744 6792 22796 6798
rect 22744 6734 22796 6740
rect 22756 2514 22784 6734
rect 23032 3398 23060 7822
rect 23124 6662 23152 8502
rect 23216 6934 23244 8774
rect 23308 7857 23336 8910
rect 23400 8906 23428 9454
rect 23388 8900 23440 8906
rect 23388 8842 23440 8848
rect 23400 7993 23428 8842
rect 23386 7984 23442 7993
rect 23386 7919 23442 7928
rect 23294 7848 23350 7857
rect 23400 7818 23428 7919
rect 23584 7818 23612 13382
rect 23664 13320 23716 13326
rect 23664 13262 23716 13268
rect 23676 12782 23704 13262
rect 23664 12776 23716 12782
rect 23664 12718 23716 12724
rect 23676 9654 23704 12718
rect 23664 9648 23716 9654
rect 23664 9590 23716 9596
rect 23664 8968 23716 8974
rect 23664 8910 23716 8916
rect 23294 7783 23350 7792
rect 23388 7812 23440 7818
rect 23204 6928 23256 6934
rect 23204 6870 23256 6876
rect 23308 6798 23336 7783
rect 23388 7754 23440 7760
rect 23572 7812 23624 7818
rect 23572 7754 23624 7760
rect 23584 7546 23612 7754
rect 23572 7540 23624 7546
rect 23572 7482 23624 7488
rect 23296 6792 23348 6798
rect 23296 6734 23348 6740
rect 23112 6656 23164 6662
rect 23112 6598 23164 6604
rect 23572 4208 23624 4214
rect 23572 4150 23624 4156
rect 23584 3534 23612 4150
rect 23204 3528 23256 3534
rect 23204 3470 23256 3476
rect 23572 3528 23624 3534
rect 23572 3470 23624 3476
rect 23020 3392 23072 3398
rect 23020 3334 23072 3340
rect 23216 3058 23244 3470
rect 23388 3392 23440 3398
rect 23388 3334 23440 3340
rect 23400 3126 23428 3334
rect 23388 3120 23440 3126
rect 23388 3062 23440 3068
rect 23204 3052 23256 3058
rect 23204 2994 23256 3000
rect 23676 2582 23704 8910
rect 23664 2576 23716 2582
rect 23664 2518 23716 2524
rect 23768 2514 23796 18142
rect 23860 17066 23888 24074
rect 24044 24018 24072 25842
rect 24122 25800 24178 25809
rect 24122 25735 24178 25744
rect 24136 25702 24164 25735
rect 24124 25696 24176 25702
rect 24124 25638 24176 25644
rect 24124 25288 24176 25294
rect 24124 25230 24176 25236
rect 23952 23990 24072 24018
rect 23848 17060 23900 17066
rect 23848 17002 23900 17008
rect 23848 14544 23900 14550
rect 23848 14486 23900 14492
rect 23860 13190 23888 14486
rect 23848 13184 23900 13190
rect 23848 13126 23900 13132
rect 23860 12918 23888 13126
rect 23848 12912 23900 12918
rect 23848 12854 23900 12860
rect 23848 12640 23900 12646
rect 23848 12582 23900 12588
rect 23860 12306 23888 12582
rect 23952 12434 23980 23990
rect 24136 23882 24164 25230
rect 24044 23854 24164 23882
rect 24044 18358 24072 23854
rect 24124 22636 24176 22642
rect 24124 22578 24176 22584
rect 24136 22409 24164 22578
rect 24228 22438 24256 31726
rect 24412 31482 24440 32320
rect 24492 32224 24544 32230
rect 24492 32166 24544 32172
rect 24504 31822 24532 32166
rect 24492 31816 24544 31822
rect 24492 31758 24544 31764
rect 24584 31748 24636 31754
rect 24584 31690 24636 31696
rect 24400 31476 24452 31482
rect 24400 31418 24452 31424
rect 24400 31136 24452 31142
rect 24400 31078 24452 31084
rect 24412 30734 24440 31078
rect 24400 30728 24452 30734
rect 24400 30670 24452 30676
rect 24596 30666 24624 31690
rect 24688 31346 24716 33918
rect 24766 33895 24822 33904
rect 24872 32570 24900 34138
rect 24860 32564 24912 32570
rect 24860 32506 24912 32512
rect 24768 32292 24820 32298
rect 24768 32234 24820 32240
rect 24676 31340 24728 31346
rect 24676 31282 24728 31288
rect 24688 30938 24716 31282
rect 24780 31278 24808 32234
rect 24768 31272 24820 31278
rect 24768 31214 24820 31220
rect 24676 30932 24728 30938
rect 24676 30874 24728 30880
rect 24584 30660 24636 30666
rect 24584 30602 24636 30608
rect 24596 30433 24624 30602
rect 24582 30424 24638 30433
rect 24308 30388 24360 30394
rect 24582 30359 24638 30368
rect 24308 30330 24360 30336
rect 24320 30258 24348 30330
rect 24308 30252 24360 30258
rect 24308 30194 24360 30200
rect 24780 29288 24808 31214
rect 24860 30660 24912 30666
rect 24860 30602 24912 30608
rect 24872 30394 24900 30602
rect 24860 30388 24912 30394
rect 24860 30330 24912 30336
rect 24860 29504 24912 29510
rect 24858 29472 24860 29481
rect 24912 29472 24914 29481
rect 24858 29407 24914 29416
rect 24504 29260 24900 29288
rect 24308 28688 24360 28694
rect 24308 28630 24360 28636
rect 24320 25906 24348 28630
rect 24400 26036 24452 26042
rect 24400 25978 24452 25984
rect 24308 25900 24360 25906
rect 24308 25842 24360 25848
rect 24412 25294 24440 25978
rect 24400 25288 24452 25294
rect 24400 25230 24452 25236
rect 24400 25152 24452 25158
rect 24504 25106 24532 29260
rect 24872 29170 24900 29260
rect 24768 29164 24820 29170
rect 24768 29106 24820 29112
rect 24860 29164 24912 29170
rect 24860 29106 24912 29112
rect 24584 27532 24636 27538
rect 24584 27474 24636 27480
rect 24452 25100 24532 25106
rect 24400 25094 24532 25100
rect 24412 25078 24532 25094
rect 24216 22432 24268 22438
rect 24122 22400 24178 22409
rect 24216 22374 24268 22380
rect 24122 22335 24178 22344
rect 24412 22094 24440 25078
rect 24596 24834 24624 27474
rect 24780 27470 24808 29106
rect 24860 27600 24912 27606
rect 24860 27542 24912 27548
rect 24768 27464 24820 27470
rect 24768 27406 24820 27412
rect 24676 27328 24728 27334
rect 24676 27270 24728 27276
rect 24688 27062 24716 27270
rect 24780 27062 24808 27406
rect 24872 27130 24900 27542
rect 24860 27124 24912 27130
rect 24860 27066 24912 27072
rect 24676 27056 24728 27062
rect 24676 26998 24728 27004
rect 24768 27056 24820 27062
rect 24768 26998 24820 27004
rect 24768 26376 24820 26382
rect 24768 26318 24820 26324
rect 24676 26036 24728 26042
rect 24676 25978 24728 25984
rect 24688 25226 24716 25978
rect 24780 25702 24808 26318
rect 24768 25696 24820 25702
rect 24768 25638 24820 25644
rect 24860 25696 24912 25702
rect 24860 25638 24912 25644
rect 24872 25514 24900 25638
rect 24780 25486 24900 25514
rect 24676 25220 24728 25226
rect 24676 25162 24728 25168
rect 24676 24948 24728 24954
rect 24676 24890 24728 24896
rect 24320 22066 24440 22094
rect 24504 24806 24624 24834
rect 24124 21956 24176 21962
rect 24124 21898 24176 21904
rect 24136 20777 24164 21898
rect 24216 21480 24268 21486
rect 24216 21422 24268 21428
rect 24122 20768 24178 20777
rect 24122 20703 24178 20712
rect 24124 20596 24176 20602
rect 24124 20538 24176 20544
rect 24032 18352 24084 18358
rect 24032 18294 24084 18300
rect 24136 18290 24164 20538
rect 24228 20534 24256 21422
rect 24216 20528 24268 20534
rect 24216 20470 24268 20476
rect 24228 19446 24256 20470
rect 24216 19440 24268 19446
rect 24216 19382 24268 19388
rect 24216 18420 24268 18426
rect 24216 18362 24268 18368
rect 24124 18284 24176 18290
rect 24124 18226 24176 18232
rect 24228 18222 24256 18362
rect 24216 18216 24268 18222
rect 24136 18164 24216 18170
rect 24136 18158 24268 18164
rect 24136 18142 24256 18158
rect 24032 18080 24084 18086
rect 24032 18022 24084 18028
rect 24044 17610 24072 18022
rect 24136 17746 24164 18142
rect 24228 18093 24256 18142
rect 24124 17740 24176 17746
rect 24124 17682 24176 17688
rect 24136 17649 24164 17682
rect 24216 17672 24268 17678
rect 24122 17640 24178 17649
rect 24032 17604 24084 17610
rect 24320 17660 24348 22066
rect 24400 21004 24452 21010
rect 24400 20946 24452 20952
rect 24268 17632 24348 17660
rect 24216 17614 24268 17620
rect 24122 17575 24178 17584
rect 24032 17546 24084 17552
rect 24122 17232 24178 17241
rect 24412 17218 24440 20946
rect 24504 20602 24532 24806
rect 24584 24676 24636 24682
rect 24584 24618 24636 24624
rect 24596 24206 24624 24618
rect 24688 24206 24716 24890
rect 24584 24200 24636 24206
rect 24584 24142 24636 24148
rect 24676 24200 24728 24206
rect 24676 24142 24728 24148
rect 24780 23746 24808 25486
rect 24964 25362 24992 48486
rect 25240 48278 25268 49030
rect 25332 48890 25360 49030
rect 25320 48884 25372 48890
rect 25320 48826 25372 48832
rect 25976 48822 26004 51326
rect 26422 51200 26478 52000
rect 27066 51200 27122 52000
rect 27710 51200 27766 52000
rect 28354 51200 28410 52000
rect 28998 51200 29054 52000
rect 29642 51200 29698 52000
rect 30930 51200 30986 52000
rect 31574 51200 31630 52000
rect 32218 51200 32274 52000
rect 32862 51354 32918 52000
rect 32862 51326 33088 51354
rect 32862 51200 32918 51326
rect 26436 49230 26464 51200
rect 26424 49224 26476 49230
rect 26424 49166 26476 49172
rect 26608 49088 26660 49094
rect 26608 49030 26660 49036
rect 25964 48816 26016 48822
rect 25964 48758 26016 48764
rect 25228 48272 25280 48278
rect 25228 48214 25280 48220
rect 26620 41414 26648 49030
rect 27080 48210 27108 51200
rect 27344 49156 27396 49162
rect 27344 49098 27396 49104
rect 27356 48754 27384 49098
rect 27528 49088 27580 49094
rect 27528 49030 27580 49036
rect 27540 48822 27568 49030
rect 27528 48816 27580 48822
rect 27528 48758 27580 48764
rect 27344 48748 27396 48754
rect 27344 48690 27396 48696
rect 27724 48618 27752 51200
rect 27988 49224 28040 49230
rect 27988 49166 28040 49172
rect 27620 48612 27672 48618
rect 27620 48554 27672 48560
rect 27712 48612 27764 48618
rect 27712 48554 27764 48560
rect 27068 48204 27120 48210
rect 27068 48146 27120 48152
rect 27068 48068 27120 48074
rect 27068 48010 27120 48016
rect 27080 47802 27108 48010
rect 27068 47796 27120 47802
rect 27068 47738 27120 47744
rect 27632 47666 27660 48554
rect 27620 47660 27672 47666
rect 27620 47602 27672 47608
rect 26976 47524 27028 47530
rect 26976 47466 27028 47472
rect 26988 47190 27016 47466
rect 26976 47184 27028 47190
rect 26976 47126 27028 47132
rect 26528 41386 26648 41414
rect 28000 41414 28028 49166
rect 28368 47598 28396 51200
rect 29012 49230 29040 51200
rect 29656 49722 29684 51200
rect 29656 49694 30052 49722
rect 29092 49360 29144 49366
rect 29092 49302 29144 49308
rect 29000 49224 29052 49230
rect 29000 49166 29052 49172
rect 28724 48680 28776 48686
rect 28724 48622 28776 48628
rect 28736 48278 28764 48622
rect 28724 48272 28776 48278
rect 28724 48214 28776 48220
rect 28172 47592 28224 47598
rect 28172 47534 28224 47540
rect 28356 47592 28408 47598
rect 28356 47534 28408 47540
rect 28184 47054 28212 47534
rect 28080 47048 28132 47054
rect 28080 46990 28132 46996
rect 28172 47048 28224 47054
rect 28172 46990 28224 46996
rect 28092 45626 28120 46990
rect 28080 45620 28132 45626
rect 28080 45562 28132 45568
rect 28816 45620 28868 45626
rect 28816 45562 28868 45568
rect 28828 45422 28856 45562
rect 28816 45416 28868 45422
rect 28816 45358 28868 45364
rect 28000 41386 28120 41414
rect 25044 39840 25096 39846
rect 25044 39782 25096 39788
rect 25056 39302 25084 39782
rect 25044 39296 25096 39302
rect 25044 39238 25096 39244
rect 25780 39296 25832 39302
rect 25780 39238 25832 39244
rect 25056 35630 25084 39238
rect 25136 38956 25188 38962
rect 25136 38898 25188 38904
rect 25148 38486 25176 38898
rect 25136 38480 25188 38486
rect 25136 38422 25188 38428
rect 25792 38418 25820 39238
rect 26068 38950 26280 38978
rect 26068 38654 26096 38950
rect 26252 38894 26280 38950
rect 26240 38888 26292 38894
rect 26240 38830 26292 38836
rect 26148 38820 26200 38826
rect 26148 38762 26200 38768
rect 25884 38626 26096 38654
rect 25780 38412 25832 38418
rect 25780 38354 25832 38360
rect 25228 38344 25280 38350
rect 25228 38286 25280 38292
rect 25240 37466 25268 38286
rect 25412 37868 25464 37874
rect 25412 37810 25464 37816
rect 25228 37460 25280 37466
rect 25228 37402 25280 37408
rect 25228 37256 25280 37262
rect 25228 37198 25280 37204
rect 25044 35624 25096 35630
rect 25044 35566 25096 35572
rect 25044 34604 25096 34610
rect 25044 34546 25096 34552
rect 25056 34202 25084 34546
rect 25044 34196 25096 34202
rect 25044 34138 25096 34144
rect 25044 33992 25096 33998
rect 25044 33934 25096 33940
rect 25056 32774 25084 33934
rect 25044 32768 25096 32774
rect 25044 32710 25096 32716
rect 25044 31408 25096 31414
rect 25044 31350 25096 31356
rect 25056 30326 25084 31350
rect 25044 30320 25096 30326
rect 25044 30262 25096 30268
rect 25044 30184 25096 30190
rect 25044 30126 25096 30132
rect 25056 29889 25084 30126
rect 25042 29880 25098 29889
rect 25042 29815 25098 29824
rect 25240 26874 25268 37198
rect 25424 35834 25452 37810
rect 25688 37324 25740 37330
rect 25688 37266 25740 37272
rect 25504 37120 25556 37126
rect 25504 37062 25556 37068
rect 25516 36174 25544 37062
rect 25700 36718 25728 37266
rect 25688 36712 25740 36718
rect 25688 36654 25740 36660
rect 25700 36242 25728 36654
rect 25688 36236 25740 36242
rect 25688 36178 25740 36184
rect 25504 36168 25556 36174
rect 25504 36110 25556 36116
rect 25412 35828 25464 35834
rect 25412 35770 25464 35776
rect 25596 35692 25648 35698
rect 25596 35634 25648 35640
rect 25608 35018 25636 35634
rect 25700 35630 25728 36178
rect 25792 36174 25820 38354
rect 25884 38282 25912 38626
rect 26160 38350 26188 38762
rect 26424 38752 26476 38758
rect 26424 38694 26476 38700
rect 26436 38350 26464 38694
rect 26148 38344 26200 38350
rect 26148 38286 26200 38292
rect 26424 38344 26476 38350
rect 26424 38286 26476 38292
rect 25872 38276 25924 38282
rect 25872 38218 25924 38224
rect 25884 37330 25912 38218
rect 26056 37800 26108 37806
rect 26056 37742 26108 37748
rect 25872 37324 25924 37330
rect 25924 37284 26004 37312
rect 25872 37266 25924 37272
rect 25872 36780 25924 36786
rect 25872 36722 25924 36728
rect 25884 36378 25912 36722
rect 25976 36666 26004 37284
rect 26068 36786 26096 37742
rect 26160 37398 26188 38286
rect 26332 38004 26384 38010
rect 26332 37946 26384 37952
rect 26344 37913 26372 37946
rect 26330 37904 26386 37913
rect 26330 37839 26386 37848
rect 26148 37392 26200 37398
rect 26148 37334 26200 37340
rect 26056 36780 26108 36786
rect 26056 36722 26108 36728
rect 25976 36638 26096 36666
rect 25964 36576 26016 36582
rect 25964 36518 26016 36524
rect 25872 36372 25924 36378
rect 25872 36314 25924 36320
rect 25780 36168 25832 36174
rect 25780 36110 25832 36116
rect 25688 35624 25740 35630
rect 25688 35566 25740 35572
rect 25596 35012 25648 35018
rect 25596 34954 25648 34960
rect 25700 34950 25728 35566
rect 25688 34944 25740 34950
rect 25688 34886 25740 34892
rect 25504 34400 25556 34406
rect 25504 34342 25556 34348
rect 25516 33998 25544 34342
rect 25504 33992 25556 33998
rect 25504 33934 25556 33940
rect 25792 33930 25820 36110
rect 25976 35986 26004 36518
rect 26068 36106 26096 36638
rect 26160 36310 26188 37334
rect 26240 37256 26292 37262
rect 26240 37198 26292 37204
rect 26252 36922 26280 37198
rect 26240 36916 26292 36922
rect 26240 36858 26292 36864
rect 26332 36780 26384 36786
rect 26332 36722 26384 36728
rect 26344 36378 26372 36722
rect 26436 36650 26464 38286
rect 26424 36644 26476 36650
rect 26424 36586 26476 36592
rect 26332 36372 26384 36378
rect 26332 36314 26384 36320
rect 26148 36304 26200 36310
rect 26148 36246 26200 36252
rect 26240 36168 26292 36174
rect 26240 36110 26292 36116
rect 26056 36100 26108 36106
rect 26056 36042 26108 36048
rect 25976 35958 26188 35986
rect 25964 34604 26016 34610
rect 25964 34546 26016 34552
rect 25872 34468 25924 34474
rect 25872 34410 25924 34416
rect 25884 33998 25912 34410
rect 25872 33992 25924 33998
rect 25872 33934 25924 33940
rect 25780 33924 25832 33930
rect 25780 33866 25832 33872
rect 25596 33856 25648 33862
rect 25596 33798 25648 33804
rect 25412 32564 25464 32570
rect 25412 32506 25464 32512
rect 25424 32026 25452 32506
rect 25412 32020 25464 32026
rect 25412 31962 25464 31968
rect 25320 31748 25372 31754
rect 25320 31690 25372 31696
rect 25332 31482 25360 31690
rect 25320 31476 25372 31482
rect 25320 31418 25372 31424
rect 25412 30728 25464 30734
rect 25412 30670 25464 30676
rect 25504 30728 25556 30734
rect 25504 30670 25556 30676
rect 25320 30592 25372 30598
rect 25320 30534 25372 30540
rect 25332 30258 25360 30534
rect 25320 30252 25372 30258
rect 25320 30194 25372 30200
rect 25424 29646 25452 30670
rect 25516 30258 25544 30670
rect 25504 30252 25556 30258
rect 25504 30194 25556 30200
rect 25504 29708 25556 29714
rect 25504 29650 25556 29656
rect 25412 29640 25464 29646
rect 25412 29582 25464 29588
rect 25516 29238 25544 29650
rect 25504 29232 25556 29238
rect 25504 29174 25556 29180
rect 25608 27606 25636 33798
rect 25976 32434 26004 34546
rect 26160 34406 26188 35958
rect 26148 34400 26200 34406
rect 26148 34342 26200 34348
rect 26054 34096 26110 34105
rect 26054 34031 26056 34040
rect 26108 34031 26110 34040
rect 26056 34002 26108 34008
rect 26056 33380 26108 33386
rect 26056 33322 26108 33328
rect 25964 32428 26016 32434
rect 25964 32370 26016 32376
rect 25780 31680 25832 31686
rect 25780 31622 25832 31628
rect 25792 31346 25820 31622
rect 26068 31414 26096 33322
rect 26160 32366 26188 34342
rect 26252 33318 26280 36110
rect 26332 35692 26384 35698
rect 26332 35634 26384 35640
rect 26344 33590 26372 35634
rect 26436 34610 26464 36586
rect 26424 34604 26476 34610
rect 26424 34546 26476 34552
rect 26424 34400 26476 34406
rect 26424 34342 26476 34348
rect 26436 33998 26464 34342
rect 26424 33992 26476 33998
rect 26424 33934 26476 33940
rect 26528 33810 26556 41386
rect 26700 39432 26752 39438
rect 26700 39374 26752 39380
rect 26712 39030 26740 39374
rect 26976 39364 27028 39370
rect 26976 39306 27028 39312
rect 26790 39128 26846 39137
rect 26988 39098 27016 39306
rect 26790 39063 26846 39072
rect 26976 39092 27028 39098
rect 26804 39030 26832 39063
rect 26976 39034 27028 39040
rect 26700 39024 26752 39030
rect 26700 38966 26752 38972
rect 26792 39024 26844 39030
rect 26792 38966 26844 38972
rect 26712 37262 26740 38966
rect 27528 38956 27580 38962
rect 27528 38898 27580 38904
rect 27540 38842 27568 38898
rect 27540 38814 27660 38842
rect 26792 37664 26844 37670
rect 26792 37606 26844 37612
rect 26700 37256 26752 37262
rect 26700 37198 26752 37204
rect 26712 36718 26740 37198
rect 26700 36712 26752 36718
rect 26700 36654 26752 36660
rect 26712 34950 26740 36654
rect 26804 36174 26832 37606
rect 27436 37460 27488 37466
rect 27436 37402 27488 37408
rect 26792 36168 26844 36174
rect 26792 36110 26844 36116
rect 27448 36106 27476 37402
rect 27160 36100 27212 36106
rect 27160 36042 27212 36048
rect 27436 36100 27488 36106
rect 27436 36042 27488 36048
rect 26792 35080 26844 35086
rect 26792 35022 26844 35028
rect 26700 34944 26752 34950
rect 26700 34886 26752 34892
rect 26608 34196 26660 34202
rect 26608 34138 26660 34144
rect 26436 33782 26556 33810
rect 26332 33584 26384 33590
rect 26332 33526 26384 33532
rect 26240 33312 26292 33318
rect 26240 33254 26292 33260
rect 26148 32360 26200 32366
rect 26148 32302 26200 32308
rect 26056 31408 26108 31414
rect 26056 31350 26108 31356
rect 25780 31340 25832 31346
rect 25780 31282 25832 31288
rect 25964 31340 26016 31346
rect 25964 31282 26016 31288
rect 25976 30734 26004 31282
rect 25964 30728 26016 30734
rect 25964 30670 26016 30676
rect 26054 30424 26110 30433
rect 26054 30359 26110 30368
rect 26068 30326 26096 30359
rect 26056 30320 26108 30326
rect 26056 30262 26108 30268
rect 25780 30184 25832 30190
rect 25780 30126 25832 30132
rect 26332 30184 26384 30190
rect 26332 30126 26384 30132
rect 25688 30048 25740 30054
rect 25688 29990 25740 29996
rect 25700 29850 25728 29990
rect 25688 29844 25740 29850
rect 25688 29786 25740 29792
rect 25596 27600 25648 27606
rect 25596 27542 25648 27548
rect 25240 26846 25452 26874
rect 25228 25696 25280 25702
rect 25228 25638 25280 25644
rect 24952 25356 25004 25362
rect 24952 25298 25004 25304
rect 24964 24970 24992 25298
rect 25136 25152 25188 25158
rect 25136 25094 25188 25100
rect 24872 24942 24992 24970
rect 24872 24886 24900 24942
rect 24860 24880 24912 24886
rect 25148 24857 25176 25094
rect 24860 24822 24912 24828
rect 25134 24848 25190 24857
rect 24952 24812 25004 24818
rect 25134 24783 25190 24792
rect 24952 24754 25004 24760
rect 24596 23718 24808 23746
rect 24964 23730 24992 24754
rect 25240 24750 25268 25638
rect 25320 25288 25372 25294
rect 25320 25230 25372 25236
rect 25228 24744 25280 24750
rect 25228 24686 25280 24692
rect 25136 24200 25188 24206
rect 25136 24142 25188 24148
rect 24952 23724 25004 23730
rect 24492 20596 24544 20602
rect 24492 20538 24544 20544
rect 24492 20256 24544 20262
rect 24492 20198 24544 20204
rect 24122 17167 24178 17176
rect 24228 17190 24440 17218
rect 24136 17134 24164 17167
rect 24124 17128 24176 17134
rect 24124 17070 24176 17076
rect 24032 14408 24084 14414
rect 24032 14350 24084 14356
rect 24044 14006 24072 14350
rect 24032 14000 24084 14006
rect 24032 13942 24084 13948
rect 24228 13326 24256 17190
rect 24308 17128 24360 17134
rect 24308 17070 24360 17076
rect 24216 13320 24268 13326
rect 24216 13262 24268 13268
rect 23952 12406 24072 12434
rect 23848 12300 23900 12306
rect 23848 12242 23900 12248
rect 23848 9376 23900 9382
rect 23848 9318 23900 9324
rect 23860 7954 23888 9318
rect 23848 7948 23900 7954
rect 23848 7890 23900 7896
rect 23860 6730 23888 7890
rect 24044 7562 24072 12406
rect 24124 12368 24176 12374
rect 24124 12310 24176 12316
rect 24136 11898 24164 12310
rect 24124 11892 24176 11898
rect 24124 11834 24176 11840
rect 24216 11688 24268 11694
rect 24216 11630 24268 11636
rect 24228 10674 24256 11630
rect 24216 10668 24268 10674
rect 24216 10610 24268 10616
rect 24216 10532 24268 10538
rect 24216 10474 24268 10480
rect 24122 9752 24178 9761
rect 24122 9687 24178 9696
rect 23952 7534 24072 7562
rect 23848 6724 23900 6730
rect 23848 6666 23900 6672
rect 23848 2984 23900 2990
rect 23848 2926 23900 2932
rect 22744 2508 22796 2514
rect 22744 2450 22796 2456
rect 23756 2508 23808 2514
rect 23756 2450 23808 2456
rect 22560 2440 22612 2446
rect 22560 2382 22612 2388
rect 23204 2440 23256 2446
rect 23204 2382 23256 2388
rect 22572 800 22600 2382
rect 22836 2304 22888 2310
rect 22836 2246 22888 2252
rect 22848 2038 22876 2246
rect 22836 2032 22888 2038
rect 22836 1974 22888 1980
rect 23216 800 23244 2382
rect 23860 800 23888 2926
rect 23952 2106 23980 7534
rect 24136 2774 24164 9687
rect 24228 8362 24256 10474
rect 24216 8356 24268 8362
rect 24216 8298 24268 8304
rect 24044 2746 24164 2774
rect 24044 2310 24072 2746
rect 24032 2304 24084 2310
rect 24032 2246 24084 2252
rect 23940 2100 23992 2106
rect 23940 2042 23992 2048
rect 24320 1970 24348 17070
rect 24400 14272 24452 14278
rect 24400 14214 24452 14220
rect 24412 12918 24440 14214
rect 24400 12912 24452 12918
rect 24400 12854 24452 12860
rect 24412 12170 24440 12854
rect 24400 12164 24452 12170
rect 24400 12106 24452 12112
rect 24400 11756 24452 11762
rect 24400 11698 24452 11704
rect 24412 10674 24440 11698
rect 24400 10668 24452 10674
rect 24400 10610 24452 10616
rect 24412 10538 24440 10610
rect 24400 10532 24452 10538
rect 24400 10474 24452 10480
rect 24504 9042 24532 20198
rect 24596 19922 24624 23718
rect 24952 23666 25004 23672
rect 25148 23662 25176 24142
rect 25136 23656 25188 23662
rect 25136 23598 25188 23604
rect 25240 23594 25268 24686
rect 25332 24614 25360 25230
rect 25320 24608 25372 24614
rect 25320 24550 25372 24556
rect 25228 23588 25280 23594
rect 25228 23530 25280 23536
rect 24676 23520 24728 23526
rect 24674 23488 24676 23497
rect 24860 23520 24912 23526
rect 24728 23488 24730 23497
rect 24860 23462 24912 23468
rect 25044 23520 25096 23526
rect 25044 23462 25096 23468
rect 24674 23423 24730 23432
rect 24688 22506 24716 23423
rect 24768 23248 24820 23254
rect 24768 23190 24820 23196
rect 24676 22500 24728 22506
rect 24676 22442 24728 22448
rect 24676 21888 24728 21894
rect 24676 21830 24728 21836
rect 24688 21350 24716 21830
rect 24676 21344 24728 21350
rect 24676 21286 24728 21292
rect 24676 20936 24728 20942
rect 24676 20878 24728 20884
rect 24584 19916 24636 19922
rect 24584 19858 24636 19864
rect 24596 17746 24624 19858
rect 24688 19514 24716 20878
rect 24780 20262 24808 23190
rect 24872 23118 24900 23462
rect 25056 23322 25084 23462
rect 25044 23316 25096 23322
rect 25044 23258 25096 23264
rect 24860 23112 24912 23118
rect 24860 23054 24912 23060
rect 25044 22636 25096 22642
rect 25044 22578 25096 22584
rect 24860 21888 24912 21894
rect 24860 21830 24912 21836
rect 24872 21554 24900 21830
rect 24860 21548 24912 21554
rect 24860 21490 24912 21496
rect 24952 21412 25004 21418
rect 24952 21354 25004 21360
rect 24860 21344 24912 21350
rect 24860 21286 24912 21292
rect 24872 20890 24900 21286
rect 24964 21010 24992 21354
rect 24952 21004 25004 21010
rect 24952 20946 25004 20952
rect 24872 20874 24992 20890
rect 24872 20868 25004 20874
rect 24872 20862 24952 20868
rect 24768 20256 24820 20262
rect 24768 20198 24820 20204
rect 24676 19508 24728 19514
rect 24676 19450 24728 19456
rect 24768 19440 24820 19446
rect 24768 19382 24820 19388
rect 24676 18624 24728 18630
rect 24676 18566 24728 18572
rect 24688 18222 24716 18566
rect 24676 18216 24728 18222
rect 24676 18158 24728 18164
rect 24780 17882 24808 19382
rect 24872 19378 24900 20862
rect 24952 20810 25004 20816
rect 24950 20768 25006 20777
rect 24950 20703 25006 20712
rect 24860 19372 24912 19378
rect 24860 19314 24912 19320
rect 24860 19236 24912 19242
rect 24860 19178 24912 19184
rect 24768 17876 24820 17882
rect 24768 17818 24820 17824
rect 24584 17740 24636 17746
rect 24584 17682 24636 17688
rect 24768 17536 24820 17542
rect 24768 17478 24820 17484
rect 24780 17241 24808 17478
rect 24872 17270 24900 19178
rect 24964 17746 24992 20703
rect 24952 17740 25004 17746
rect 24952 17682 25004 17688
rect 24860 17264 24912 17270
rect 24766 17232 24822 17241
rect 24860 17206 24912 17212
rect 24766 17167 24822 17176
rect 24768 17060 24820 17066
rect 24768 17002 24820 17008
rect 24584 15020 24636 15026
rect 24584 14962 24636 14968
rect 24596 14618 24624 14962
rect 24584 14612 24636 14618
rect 24584 14554 24636 14560
rect 24676 14612 24728 14618
rect 24676 14554 24728 14560
rect 24688 14278 24716 14554
rect 24676 14272 24728 14278
rect 24676 14214 24728 14220
rect 24676 11076 24728 11082
rect 24676 11018 24728 11024
rect 24688 10810 24716 11018
rect 24676 10804 24728 10810
rect 24676 10746 24728 10752
rect 24780 9058 24808 17002
rect 24872 15502 24900 17206
rect 24860 15496 24912 15502
rect 24860 15438 24912 15444
rect 24964 15366 24992 17682
rect 25056 17338 25084 22578
rect 25320 22432 25372 22438
rect 25320 22374 25372 22380
rect 25332 22166 25360 22374
rect 25320 22160 25372 22166
rect 25320 22102 25372 22108
rect 25136 22024 25188 22030
rect 25136 21966 25188 21972
rect 25148 21078 25176 21966
rect 25228 21548 25280 21554
rect 25228 21490 25280 21496
rect 25240 21146 25268 21490
rect 25228 21140 25280 21146
rect 25228 21082 25280 21088
rect 25136 21072 25188 21078
rect 25136 21014 25188 21020
rect 25320 21004 25372 21010
rect 25320 20946 25372 20952
rect 25136 20936 25188 20942
rect 25136 20878 25188 20884
rect 25148 18426 25176 20878
rect 25332 20262 25360 20946
rect 25320 20256 25372 20262
rect 25320 20198 25372 20204
rect 25320 18692 25372 18698
rect 25320 18634 25372 18640
rect 25136 18420 25188 18426
rect 25136 18362 25188 18368
rect 25332 18290 25360 18634
rect 25320 18284 25372 18290
rect 25320 18226 25372 18232
rect 25332 17882 25360 18226
rect 25136 17876 25188 17882
rect 25136 17818 25188 17824
rect 25320 17876 25372 17882
rect 25320 17818 25372 17824
rect 25148 17338 25176 17818
rect 25044 17332 25096 17338
rect 25044 17274 25096 17280
rect 25136 17332 25188 17338
rect 25136 17274 25188 17280
rect 25424 17218 25452 26846
rect 25686 25664 25742 25673
rect 25686 25599 25742 25608
rect 25596 25288 25648 25294
rect 25596 25230 25648 25236
rect 25504 24948 25556 24954
rect 25504 24890 25556 24896
rect 25516 22681 25544 24890
rect 25608 24206 25636 25230
rect 25700 24954 25728 25599
rect 25688 24948 25740 24954
rect 25688 24890 25740 24896
rect 25596 24200 25648 24206
rect 25596 24142 25648 24148
rect 25688 23044 25740 23050
rect 25688 22986 25740 22992
rect 25502 22672 25558 22681
rect 25502 22607 25558 22616
rect 25504 22568 25556 22574
rect 25504 22510 25556 22516
rect 25136 17196 25188 17202
rect 25136 17138 25188 17144
rect 25240 17190 25452 17218
rect 25148 16454 25176 17138
rect 25136 16448 25188 16454
rect 25136 16390 25188 16396
rect 25148 16114 25176 16390
rect 25136 16108 25188 16114
rect 25136 16050 25188 16056
rect 25044 15904 25096 15910
rect 25044 15846 25096 15852
rect 25056 15706 25084 15846
rect 25044 15700 25096 15706
rect 25044 15642 25096 15648
rect 24952 15360 25004 15366
rect 24952 15302 25004 15308
rect 25148 15026 25176 16050
rect 25136 15020 25188 15026
rect 25136 14962 25188 14968
rect 24952 14884 25004 14890
rect 24952 14826 25004 14832
rect 24860 14816 24912 14822
rect 24860 14758 24912 14764
rect 24872 12434 24900 14758
rect 24964 14482 24992 14826
rect 24952 14476 25004 14482
rect 24952 14418 25004 14424
rect 25042 14376 25098 14385
rect 25042 14311 25044 14320
rect 25096 14311 25098 14320
rect 25044 14282 25096 14288
rect 25056 12782 25084 14282
rect 25136 13524 25188 13530
rect 25136 13466 25188 13472
rect 25148 12850 25176 13466
rect 25136 12844 25188 12850
rect 25136 12786 25188 12792
rect 25044 12776 25096 12782
rect 25044 12718 25096 12724
rect 24872 12406 25084 12434
rect 24952 12232 25004 12238
rect 24952 12174 25004 12180
rect 24964 11898 24992 12174
rect 24952 11892 25004 11898
rect 24952 11834 25004 11840
rect 25056 11694 25084 12406
rect 25148 12238 25176 12786
rect 25136 12232 25188 12238
rect 25136 12174 25188 12180
rect 25044 11688 25096 11694
rect 25044 11630 25096 11636
rect 24952 9376 25004 9382
rect 24952 9318 25004 9324
rect 24964 9110 24992 9318
rect 24492 9036 24544 9042
rect 24492 8978 24544 8984
rect 24688 9030 24808 9058
rect 24952 9104 25004 9110
rect 24952 9046 25004 9052
rect 24400 7744 24452 7750
rect 24400 7686 24452 7692
rect 24412 7478 24440 7686
rect 24400 7472 24452 7478
rect 24400 7414 24452 7420
rect 24688 5914 24716 9030
rect 25044 8968 25096 8974
rect 25044 8910 25096 8916
rect 25136 8968 25188 8974
rect 25136 8910 25188 8916
rect 24952 8832 25004 8838
rect 24952 8774 25004 8780
rect 24964 8498 24992 8774
rect 24952 8492 25004 8498
rect 24952 8434 25004 8440
rect 25056 8090 25084 8910
rect 25044 8084 25096 8090
rect 25044 8026 25096 8032
rect 25044 7880 25096 7886
rect 25042 7848 25044 7857
rect 25148 7868 25176 8910
rect 25096 7848 25176 7868
rect 25098 7840 25176 7848
rect 25042 7783 25098 7792
rect 25240 7562 25268 17190
rect 25320 15904 25372 15910
rect 25320 15846 25372 15852
rect 25332 13734 25360 15846
rect 25320 13728 25372 13734
rect 25320 13670 25372 13676
rect 25320 13320 25372 13326
rect 25320 13262 25372 13268
rect 25332 12918 25360 13262
rect 25320 12912 25372 12918
rect 25320 12854 25372 12860
rect 25332 12646 25360 12854
rect 25320 12640 25372 12646
rect 25320 12582 25372 12588
rect 25332 12442 25360 12582
rect 25320 12436 25372 12442
rect 25320 12378 25372 12384
rect 25320 11008 25372 11014
rect 25320 10950 25372 10956
rect 25332 10810 25360 10950
rect 25320 10804 25372 10810
rect 25320 10746 25372 10752
rect 25332 10130 25360 10746
rect 25320 10124 25372 10130
rect 25320 10066 25372 10072
rect 25318 7984 25374 7993
rect 25318 7919 25374 7928
rect 25332 7886 25360 7919
rect 25320 7880 25372 7886
rect 25320 7822 25372 7828
rect 25240 7534 25360 7562
rect 24676 5908 24728 5914
rect 24676 5850 24728 5856
rect 25228 5704 25280 5710
rect 25228 5646 25280 5652
rect 25240 5098 25268 5646
rect 25228 5092 25280 5098
rect 25228 5034 25280 5040
rect 24492 2440 24544 2446
rect 24492 2382 24544 2388
rect 24676 2440 24728 2446
rect 24676 2382 24728 2388
rect 25136 2440 25188 2446
rect 25136 2382 25188 2388
rect 24308 1964 24360 1970
rect 24308 1906 24360 1912
rect 24504 800 24532 2382
rect 24688 2310 24716 2382
rect 24676 2304 24728 2310
rect 24676 2246 24728 2252
rect 25148 800 25176 2382
rect 25332 2310 25360 7534
rect 25516 5914 25544 22510
rect 25596 21684 25648 21690
rect 25596 21626 25648 21632
rect 25608 21554 25636 21626
rect 25596 21548 25648 21554
rect 25596 21490 25648 21496
rect 25608 20942 25636 21490
rect 25700 21321 25728 22986
rect 25686 21312 25742 21321
rect 25686 21247 25742 21256
rect 25700 21146 25728 21247
rect 25688 21140 25740 21146
rect 25688 21082 25740 21088
rect 25596 20936 25648 20942
rect 25596 20878 25648 20884
rect 25688 20256 25740 20262
rect 25688 20198 25740 20204
rect 25596 19508 25648 19514
rect 25596 19450 25648 19456
rect 25608 18970 25636 19450
rect 25596 18964 25648 18970
rect 25596 18906 25648 18912
rect 25700 18630 25728 20198
rect 25688 18624 25740 18630
rect 25688 18566 25740 18572
rect 25596 18148 25648 18154
rect 25596 18090 25648 18096
rect 25608 13870 25636 18090
rect 25700 16114 25728 18566
rect 25688 16108 25740 16114
rect 25688 16050 25740 16056
rect 25700 14550 25728 16050
rect 25688 14544 25740 14550
rect 25688 14486 25740 14492
rect 25596 13864 25648 13870
rect 25596 13806 25648 13812
rect 25688 12640 25740 12646
rect 25688 12582 25740 12588
rect 25596 12436 25648 12442
rect 25596 12378 25648 12384
rect 25608 11558 25636 12378
rect 25700 12238 25728 12582
rect 25688 12232 25740 12238
rect 25688 12174 25740 12180
rect 25792 11880 25820 30126
rect 25872 29776 25924 29782
rect 25872 29718 25924 29724
rect 25884 29345 25912 29718
rect 25870 29336 25926 29345
rect 25870 29271 25926 29280
rect 26344 28762 26372 30126
rect 26436 29510 26464 33782
rect 26620 33658 26648 34138
rect 26608 33652 26660 33658
rect 26608 33594 26660 33600
rect 26608 33380 26660 33386
rect 26608 33322 26660 33328
rect 26516 33312 26568 33318
rect 26516 33254 26568 33260
rect 26424 29504 26476 29510
rect 26424 29446 26476 29452
rect 26332 28756 26384 28762
rect 26332 28698 26384 28704
rect 26344 28490 26372 28698
rect 26332 28484 26384 28490
rect 26332 28426 26384 28432
rect 26240 28416 26292 28422
rect 26240 28358 26292 28364
rect 26252 28082 26280 28358
rect 26056 28076 26108 28082
rect 26056 28018 26108 28024
rect 26240 28076 26292 28082
rect 26240 28018 26292 28024
rect 25964 25900 26016 25906
rect 25964 25842 26016 25848
rect 25976 25362 26004 25842
rect 25964 25356 26016 25362
rect 25964 25298 26016 25304
rect 25964 23792 26016 23798
rect 25964 23734 26016 23740
rect 25976 21894 26004 23734
rect 25964 21888 26016 21894
rect 25964 21830 26016 21836
rect 25872 20936 25924 20942
rect 25872 20878 25924 20884
rect 25964 20936 26016 20942
rect 25964 20878 26016 20884
rect 25884 20602 25912 20878
rect 25872 20596 25924 20602
rect 25872 20538 25924 20544
rect 25884 19786 25912 20538
rect 25976 20466 26004 20878
rect 25964 20460 26016 20466
rect 25964 20402 26016 20408
rect 25872 19780 25924 19786
rect 25872 19722 25924 19728
rect 25964 19168 26016 19174
rect 25964 19110 26016 19116
rect 25872 18964 25924 18970
rect 25872 18906 25924 18912
rect 25884 15450 25912 18906
rect 25976 18766 26004 19110
rect 25964 18760 26016 18766
rect 25964 18702 26016 18708
rect 25884 15422 26004 15450
rect 25872 15360 25924 15366
rect 25872 15302 25924 15308
rect 25884 12442 25912 15302
rect 25976 15026 26004 15422
rect 25964 15020 26016 15026
rect 25964 14962 26016 14968
rect 25964 12640 26016 12646
rect 25964 12582 26016 12588
rect 25872 12436 25924 12442
rect 25872 12378 25924 12384
rect 25700 11852 25820 11880
rect 25596 11552 25648 11558
rect 25596 11494 25648 11500
rect 25700 8566 25728 11852
rect 25976 11778 26004 12582
rect 25792 11762 26004 11778
rect 25780 11756 26004 11762
rect 25832 11750 26004 11756
rect 25780 11698 25832 11704
rect 25976 11354 26004 11750
rect 25964 11348 26016 11354
rect 25964 11290 26016 11296
rect 25688 8560 25740 8566
rect 25688 8502 25740 8508
rect 26068 6186 26096 28018
rect 26240 27872 26292 27878
rect 26240 27814 26292 27820
rect 26252 27402 26280 27814
rect 26240 27396 26292 27402
rect 26240 27338 26292 27344
rect 26436 26858 26464 29446
rect 26332 26852 26384 26858
rect 26332 26794 26384 26800
rect 26424 26852 26476 26858
rect 26424 26794 26476 26800
rect 26344 26314 26372 26794
rect 26332 26308 26384 26314
rect 26332 26250 26384 26256
rect 26330 24304 26386 24313
rect 26330 24239 26386 24248
rect 26344 24206 26372 24239
rect 26240 24200 26292 24206
rect 26240 24142 26292 24148
rect 26332 24200 26384 24206
rect 26332 24142 26384 24148
rect 26252 23322 26280 24142
rect 26240 23316 26292 23322
rect 26240 23258 26292 23264
rect 26344 23186 26372 24142
rect 26424 23248 26476 23254
rect 26424 23190 26476 23196
rect 26332 23180 26384 23186
rect 26332 23122 26384 23128
rect 26436 22710 26464 23190
rect 26424 22704 26476 22710
rect 26146 22672 26202 22681
rect 26424 22646 26476 22652
rect 26146 22607 26148 22616
rect 26200 22607 26202 22616
rect 26148 22578 26200 22584
rect 26148 21004 26200 21010
rect 26148 20946 26200 20952
rect 26160 18698 26188 20946
rect 26424 20800 26476 20806
rect 26424 20742 26476 20748
rect 26436 19854 26464 20742
rect 26424 19848 26476 19854
rect 26424 19790 26476 19796
rect 26424 19304 26476 19310
rect 26424 19246 26476 19252
rect 26436 18902 26464 19246
rect 26424 18896 26476 18902
rect 26424 18838 26476 18844
rect 26148 18692 26200 18698
rect 26148 18634 26200 18640
rect 26160 18358 26188 18634
rect 26148 18352 26200 18358
rect 26148 18294 26200 18300
rect 26148 18216 26200 18222
rect 26148 18158 26200 18164
rect 26160 17610 26188 18158
rect 26148 17604 26200 17610
rect 26148 17546 26200 17552
rect 26160 15366 26188 17546
rect 26148 15360 26200 15366
rect 26148 15302 26200 15308
rect 26148 14544 26200 14550
rect 26148 14486 26200 14492
rect 26160 12306 26188 14486
rect 26238 13424 26294 13433
rect 26238 13359 26294 13368
rect 26148 12300 26200 12306
rect 26148 12242 26200 12248
rect 26252 12186 26280 13359
rect 26332 12708 26384 12714
rect 26332 12650 26384 12656
rect 26344 12238 26372 12650
rect 26160 12158 26280 12186
rect 26332 12232 26384 12238
rect 26332 12174 26384 12180
rect 26424 12164 26476 12170
rect 26160 11286 26188 12158
rect 26424 12106 26476 12112
rect 26240 12096 26292 12102
rect 26240 12038 26292 12044
rect 26148 11280 26200 11286
rect 26148 11222 26200 11228
rect 26252 11150 26280 12038
rect 26332 11756 26384 11762
rect 26332 11698 26384 11704
rect 26344 11218 26372 11698
rect 26332 11212 26384 11218
rect 26332 11154 26384 11160
rect 26436 11150 26464 12106
rect 26240 11144 26292 11150
rect 26240 11086 26292 11092
rect 26424 11144 26476 11150
rect 26424 11086 26476 11092
rect 26424 9580 26476 9586
rect 26424 9522 26476 9528
rect 26436 8974 26464 9522
rect 26424 8968 26476 8974
rect 26424 8910 26476 8916
rect 26240 8356 26292 8362
rect 26240 8298 26292 8304
rect 26252 7818 26280 8298
rect 26436 7886 26464 8910
rect 26424 7880 26476 7886
rect 26424 7822 26476 7828
rect 26240 7812 26292 7818
rect 26240 7754 26292 7760
rect 26056 6180 26108 6186
rect 26056 6122 26108 6128
rect 25504 5908 25556 5914
rect 25504 5850 25556 5856
rect 25872 5704 25924 5710
rect 25872 5646 25924 5652
rect 25884 2582 25912 5646
rect 26238 3632 26294 3641
rect 26238 3567 26294 3576
rect 25964 3528 26016 3534
rect 25964 3470 26016 3476
rect 25976 3058 26004 3470
rect 26252 3466 26280 3567
rect 26240 3460 26292 3466
rect 26240 3402 26292 3408
rect 26424 3392 26476 3398
rect 26424 3334 26476 3340
rect 25964 3052 26016 3058
rect 25964 2994 26016 3000
rect 25872 2576 25924 2582
rect 25872 2518 25924 2524
rect 25320 2304 25372 2310
rect 25320 2246 25372 2252
rect 26436 800 26464 3334
rect 26528 2378 26556 33254
rect 26620 29714 26648 33322
rect 26712 31822 26740 34886
rect 26804 32910 26832 35022
rect 27068 34128 27120 34134
rect 27066 34096 27068 34105
rect 27120 34096 27122 34105
rect 27066 34031 27122 34040
rect 26884 33992 26936 33998
rect 26884 33934 26936 33940
rect 26896 33590 26924 33934
rect 26884 33584 26936 33590
rect 26884 33526 26936 33532
rect 26792 32904 26844 32910
rect 26792 32846 26844 32852
rect 27172 32842 27200 36042
rect 27632 35222 27660 38814
rect 27896 38276 27948 38282
rect 27896 38218 27948 38224
rect 27908 37942 27936 38218
rect 27896 37936 27948 37942
rect 27896 37878 27948 37884
rect 27804 36780 27856 36786
rect 27804 36722 27856 36728
rect 27710 35728 27766 35737
rect 27710 35663 27712 35672
rect 27764 35663 27766 35672
rect 27712 35634 27764 35640
rect 27620 35216 27672 35222
rect 27620 35158 27672 35164
rect 27252 35012 27304 35018
rect 27252 34954 27304 34960
rect 27344 35012 27396 35018
rect 27344 34954 27396 34960
rect 27264 34746 27292 34954
rect 27252 34740 27304 34746
rect 27252 34682 27304 34688
rect 27252 33652 27304 33658
rect 27252 33594 27304 33600
rect 27160 32836 27212 32842
rect 27160 32778 27212 32784
rect 26700 31816 26752 31822
rect 26700 31758 26752 31764
rect 27172 31142 27200 32778
rect 27160 31136 27212 31142
rect 27160 31078 27212 31084
rect 26700 30592 26752 30598
rect 26700 30534 26752 30540
rect 26608 29708 26660 29714
rect 26608 29650 26660 29656
rect 26712 28014 26740 30534
rect 26792 29708 26844 29714
rect 26792 29650 26844 29656
rect 26804 29578 26832 29650
rect 26976 29640 27028 29646
rect 26976 29582 27028 29588
rect 26792 29572 26844 29578
rect 26792 29514 26844 29520
rect 26988 29034 27016 29582
rect 27068 29300 27120 29306
rect 27068 29242 27120 29248
rect 26976 29028 27028 29034
rect 26976 28970 27028 28976
rect 26988 28014 27016 28970
rect 27080 28626 27108 29242
rect 27068 28620 27120 28626
rect 27068 28562 27120 28568
rect 27264 28558 27292 33594
rect 27356 33454 27384 34954
rect 27436 34060 27488 34066
rect 27436 34002 27488 34008
rect 27344 33448 27396 33454
rect 27344 33390 27396 33396
rect 27448 31958 27476 34002
rect 27528 33856 27580 33862
rect 27528 33798 27580 33804
rect 27540 33590 27568 33798
rect 27528 33584 27580 33590
rect 27528 33526 27580 33532
rect 27528 33448 27580 33454
rect 27528 33390 27580 33396
rect 27540 33046 27568 33390
rect 27528 33040 27580 33046
rect 27528 32982 27580 32988
rect 27540 32434 27568 32982
rect 27528 32428 27580 32434
rect 27528 32370 27580 32376
rect 27436 31952 27488 31958
rect 27436 31894 27488 31900
rect 27724 30802 27752 35634
rect 27816 33658 27844 36722
rect 27896 36032 27948 36038
rect 27896 35974 27948 35980
rect 27908 35018 27936 35974
rect 27896 35012 27948 35018
rect 27896 34954 27948 34960
rect 27804 33652 27856 33658
rect 27804 33594 27856 33600
rect 27908 31346 27936 34954
rect 27988 31680 28040 31686
rect 27988 31622 28040 31628
rect 27896 31340 27948 31346
rect 27896 31282 27948 31288
rect 27712 30796 27764 30802
rect 27712 30738 27764 30744
rect 27908 30734 27936 31282
rect 27896 30728 27948 30734
rect 27896 30670 27948 30676
rect 27528 30592 27580 30598
rect 27528 30534 27580 30540
rect 27540 30190 27568 30534
rect 28000 30394 28028 31622
rect 27988 30388 28040 30394
rect 27988 30330 28040 30336
rect 27620 30252 27672 30258
rect 27620 30194 27672 30200
rect 27528 30184 27580 30190
rect 27342 30152 27398 30161
rect 27528 30126 27580 30132
rect 27342 30087 27398 30096
rect 27356 28626 27384 30087
rect 27436 30048 27488 30054
rect 27436 29990 27488 29996
rect 27448 29170 27476 29990
rect 27528 29572 27580 29578
rect 27528 29514 27580 29520
rect 27540 29238 27568 29514
rect 27528 29232 27580 29238
rect 27528 29174 27580 29180
rect 27436 29164 27488 29170
rect 27436 29106 27488 29112
rect 27632 29102 27660 30194
rect 27804 30116 27856 30122
rect 27804 30058 27856 30064
rect 27816 29850 27844 30058
rect 27986 29880 28042 29889
rect 27712 29844 27764 29850
rect 27712 29786 27764 29792
rect 27804 29844 27856 29850
rect 27986 29815 27988 29824
rect 27804 29786 27856 29792
rect 28040 29815 28042 29824
rect 27988 29786 28040 29792
rect 27620 29096 27672 29102
rect 27620 29038 27672 29044
rect 27344 28620 27396 28626
rect 27344 28562 27396 28568
rect 27724 28558 27752 29786
rect 28092 28778 28120 41386
rect 28908 37868 28960 37874
rect 28908 37810 28960 37816
rect 28920 37738 28948 37810
rect 28356 37732 28408 37738
rect 28356 37674 28408 37680
rect 28908 37732 28960 37738
rect 28908 37674 28960 37680
rect 28368 37398 28396 37674
rect 28356 37392 28408 37398
rect 28356 37334 28408 37340
rect 28368 35834 28396 37334
rect 28816 37188 28868 37194
rect 28816 37130 28868 37136
rect 28356 35828 28408 35834
rect 28356 35770 28408 35776
rect 28724 35692 28776 35698
rect 28724 35634 28776 35640
rect 28356 35624 28408 35630
rect 28356 35566 28408 35572
rect 28368 35086 28396 35566
rect 28356 35080 28408 35086
rect 28356 35022 28408 35028
rect 28736 35018 28764 35634
rect 28828 35630 28856 37130
rect 28920 36666 28948 37674
rect 29000 37664 29052 37670
rect 29000 37606 29052 37612
rect 29012 37262 29040 37606
rect 29000 37256 29052 37262
rect 29000 37198 29052 37204
rect 28920 36638 29040 36666
rect 28908 36576 28960 36582
rect 28908 36518 28960 36524
rect 28920 35766 28948 36518
rect 29012 35834 29040 36638
rect 29000 35828 29052 35834
rect 29000 35770 29052 35776
rect 28908 35760 28960 35766
rect 28908 35702 28960 35708
rect 28816 35624 28868 35630
rect 28816 35566 28868 35572
rect 28828 35222 28856 35566
rect 28816 35216 28868 35222
rect 28816 35158 28868 35164
rect 28920 35018 28948 35702
rect 28724 35012 28776 35018
rect 28724 34954 28776 34960
rect 28908 35012 28960 35018
rect 28908 34954 28960 34960
rect 28920 34610 28948 34954
rect 28908 34604 28960 34610
rect 28908 34546 28960 34552
rect 28448 34468 28500 34474
rect 28448 34410 28500 34416
rect 28460 34066 28488 34410
rect 28448 34060 28500 34066
rect 28448 34002 28500 34008
rect 29000 34060 29052 34066
rect 29000 34002 29052 34008
rect 28354 33960 28410 33969
rect 28354 33895 28356 33904
rect 28408 33895 28410 33904
rect 28356 33866 28408 33872
rect 28448 33516 28500 33522
rect 28448 33458 28500 33464
rect 28264 33380 28316 33386
rect 28264 33322 28316 33328
rect 28172 33312 28224 33318
rect 28172 33254 28224 33260
rect 28184 32910 28212 33254
rect 28276 32910 28304 33322
rect 28460 33114 28488 33458
rect 28448 33108 28500 33114
rect 28448 33050 28500 33056
rect 28632 33040 28684 33046
rect 28632 32982 28684 32988
rect 28172 32904 28224 32910
rect 28172 32846 28224 32852
rect 28264 32904 28316 32910
rect 28264 32846 28316 32852
rect 28184 31890 28212 32846
rect 28540 32224 28592 32230
rect 28540 32166 28592 32172
rect 28552 31890 28580 32166
rect 28172 31884 28224 31890
rect 28172 31826 28224 31832
rect 28540 31884 28592 31890
rect 28540 31826 28592 31832
rect 28644 31822 28672 32982
rect 29012 32366 29040 34002
rect 29000 32360 29052 32366
rect 29000 32302 29052 32308
rect 28632 31816 28684 31822
rect 28632 31758 28684 31764
rect 28264 31680 28316 31686
rect 28264 31622 28316 31628
rect 28172 30592 28224 30598
rect 28172 30534 28224 30540
rect 28184 30258 28212 30534
rect 28172 30252 28224 30258
rect 28172 30194 28224 30200
rect 28000 28750 28120 28778
rect 27252 28552 27304 28558
rect 27252 28494 27304 28500
rect 27712 28552 27764 28558
rect 27764 28512 27844 28540
rect 27712 28494 27764 28500
rect 27344 28484 27396 28490
rect 27344 28426 27396 28432
rect 26700 28008 26752 28014
rect 26700 27950 26752 27956
rect 26976 28008 27028 28014
rect 26976 27950 27028 27956
rect 26988 27470 27016 27950
rect 27356 27674 27384 28426
rect 27436 28416 27488 28422
rect 27436 28358 27488 28364
rect 27712 28416 27764 28422
rect 27712 28358 27764 28364
rect 27448 27674 27476 28358
rect 27724 28150 27752 28358
rect 27816 28150 27844 28512
rect 27712 28144 27764 28150
rect 27712 28086 27764 28092
rect 27804 28144 27856 28150
rect 27804 28086 27856 28092
rect 27712 27872 27764 27878
rect 27712 27814 27764 27820
rect 27344 27668 27396 27674
rect 27344 27610 27396 27616
rect 27436 27668 27488 27674
rect 27436 27610 27488 27616
rect 26792 27464 26844 27470
rect 26792 27406 26844 27412
rect 26976 27464 27028 27470
rect 26976 27406 27028 27412
rect 27068 27464 27120 27470
rect 27068 27406 27120 27412
rect 26700 24676 26752 24682
rect 26700 24618 26752 24624
rect 26608 24268 26660 24274
rect 26712 24256 26740 24618
rect 26804 24274 26832 27406
rect 27080 26994 27108 27406
rect 27068 26988 27120 26994
rect 27068 26930 27120 26936
rect 27252 26920 27304 26926
rect 27252 26862 27304 26868
rect 27264 26586 27292 26862
rect 27252 26580 27304 26586
rect 27252 26522 27304 26528
rect 27448 26382 27476 27610
rect 27724 27402 27752 27814
rect 27712 27396 27764 27402
rect 27712 27338 27764 27344
rect 27436 26376 27488 26382
rect 27436 26318 27488 26324
rect 28000 25974 28028 28750
rect 28184 28082 28212 30194
rect 28172 28076 28224 28082
rect 28172 28018 28224 28024
rect 28080 27940 28132 27946
rect 28080 27882 28132 27888
rect 28092 27674 28120 27882
rect 28080 27668 28132 27674
rect 28080 27610 28132 27616
rect 28080 26920 28132 26926
rect 28080 26862 28132 26868
rect 27988 25968 28040 25974
rect 27988 25910 28040 25916
rect 27160 24812 27212 24818
rect 27160 24754 27212 24760
rect 27436 24812 27488 24818
rect 27436 24754 27488 24760
rect 27620 24812 27672 24818
rect 27620 24754 27672 24760
rect 27068 24608 27120 24614
rect 27068 24550 27120 24556
rect 26660 24228 26740 24256
rect 26608 24210 26660 24216
rect 26712 23730 26740 24228
rect 26792 24268 26844 24274
rect 26792 24210 26844 24216
rect 26804 23730 26832 24210
rect 27080 23730 27108 24550
rect 27172 23866 27200 24754
rect 27160 23860 27212 23866
rect 27160 23802 27212 23808
rect 26700 23724 26752 23730
rect 26700 23666 26752 23672
rect 26792 23724 26844 23730
rect 26792 23666 26844 23672
rect 27068 23724 27120 23730
rect 27068 23666 27120 23672
rect 26976 23044 27028 23050
rect 26976 22986 27028 22992
rect 26988 22642 27016 22986
rect 27448 22778 27476 24754
rect 27632 24313 27660 24754
rect 27618 24304 27674 24313
rect 27618 24239 27674 24248
rect 27988 24064 28040 24070
rect 27988 24006 28040 24012
rect 28000 23866 28028 24006
rect 27988 23860 28040 23866
rect 27988 23802 28040 23808
rect 27988 23656 28040 23662
rect 27988 23598 28040 23604
rect 27896 23520 27948 23526
rect 27816 23480 27896 23508
rect 27712 23316 27764 23322
rect 27712 23258 27764 23264
rect 27436 22772 27488 22778
rect 27436 22714 27488 22720
rect 26976 22636 27028 22642
rect 26976 22578 27028 22584
rect 27724 22234 27752 23258
rect 27816 22642 27844 23480
rect 27896 23462 27948 23468
rect 28000 23254 28028 23598
rect 27988 23248 28040 23254
rect 27988 23190 28040 23196
rect 28092 22930 28120 26862
rect 28172 24064 28224 24070
rect 28172 24006 28224 24012
rect 28184 23118 28212 24006
rect 28276 23322 28304 31622
rect 28644 31482 28672 31758
rect 28632 31476 28684 31482
rect 28632 31418 28684 31424
rect 28816 31340 28868 31346
rect 28816 31282 28868 31288
rect 28828 31142 28856 31282
rect 28816 31136 28868 31142
rect 28816 31078 28868 31084
rect 28540 30184 28592 30190
rect 28540 30126 28592 30132
rect 28552 29714 28580 30126
rect 28540 29708 28592 29714
rect 28540 29650 28592 29656
rect 28828 29646 28856 31078
rect 28816 29640 28868 29646
rect 28816 29582 28868 29588
rect 28356 28552 28408 28558
rect 28356 28494 28408 28500
rect 28368 27674 28396 28494
rect 28356 27668 28408 27674
rect 28356 27610 28408 27616
rect 28632 27464 28684 27470
rect 28632 27406 28684 27412
rect 28644 27334 28672 27406
rect 28632 27328 28684 27334
rect 28632 27270 28684 27276
rect 28908 24812 28960 24818
rect 28908 24754 28960 24760
rect 28630 24712 28686 24721
rect 28630 24647 28686 24656
rect 28448 24132 28500 24138
rect 28448 24074 28500 24080
rect 28460 23730 28488 24074
rect 28540 24064 28592 24070
rect 28540 24006 28592 24012
rect 28448 23724 28500 23730
rect 28448 23666 28500 23672
rect 28264 23316 28316 23322
rect 28264 23258 28316 23264
rect 28172 23112 28224 23118
rect 28224 23072 28304 23100
rect 28172 23054 28224 23060
rect 28092 22902 28212 22930
rect 27804 22636 27856 22642
rect 27804 22578 27856 22584
rect 27712 22228 27764 22234
rect 27712 22170 27764 22176
rect 27620 21616 27672 21622
rect 27620 21558 27672 21564
rect 27632 20942 27660 21558
rect 27620 20936 27672 20942
rect 27620 20878 27672 20884
rect 27712 20868 27764 20874
rect 27712 20810 27764 20816
rect 26700 20256 26752 20262
rect 26700 20198 26752 20204
rect 27528 20256 27580 20262
rect 27528 20198 27580 20204
rect 26712 19854 26740 20198
rect 27436 19916 27488 19922
rect 27540 19904 27568 20198
rect 27724 20058 27752 20810
rect 27816 20466 27844 22578
rect 28080 22432 28132 22438
rect 28080 22374 28132 22380
rect 27804 20460 27856 20466
rect 27804 20402 27856 20408
rect 27988 20392 28040 20398
rect 27988 20334 28040 20340
rect 27804 20324 27856 20330
rect 27804 20266 27856 20272
rect 27712 20052 27764 20058
rect 27712 19994 27764 20000
rect 27488 19876 27568 19904
rect 27436 19858 27488 19864
rect 26700 19848 26752 19854
rect 26700 19790 26752 19796
rect 27620 19848 27672 19854
rect 27620 19790 27672 19796
rect 26712 19446 26740 19790
rect 27528 19712 27580 19718
rect 27528 19654 27580 19660
rect 26700 19440 26752 19446
rect 26700 19382 26752 19388
rect 27344 19372 27396 19378
rect 27344 19314 27396 19320
rect 27356 19174 27384 19314
rect 27344 19168 27396 19174
rect 27344 19110 27396 19116
rect 26700 18964 26752 18970
rect 26700 18906 26752 18912
rect 26792 18964 26844 18970
rect 26792 18906 26844 18912
rect 26712 17882 26740 18906
rect 26804 18834 26832 18906
rect 26792 18828 26844 18834
rect 26792 18770 26844 18776
rect 26700 17876 26752 17882
rect 26700 17818 26752 17824
rect 26608 16040 26660 16046
rect 26608 15982 26660 15988
rect 26620 15502 26648 15982
rect 26712 15706 26740 17818
rect 26804 17678 26832 18770
rect 27356 18766 27384 19110
rect 27540 18970 27568 19654
rect 27528 18964 27580 18970
rect 27528 18906 27580 18912
rect 26884 18760 26936 18766
rect 27068 18760 27120 18766
rect 26936 18720 27016 18748
rect 26884 18702 26936 18708
rect 26988 17678 27016 18720
rect 27068 18702 27120 18708
rect 27344 18760 27396 18766
rect 27344 18702 27396 18708
rect 26792 17672 26844 17678
rect 26792 17614 26844 17620
rect 26976 17672 27028 17678
rect 26976 17614 27028 17620
rect 26804 17338 26832 17614
rect 26792 17332 26844 17338
rect 26792 17274 26844 17280
rect 26700 15700 26752 15706
rect 26700 15642 26752 15648
rect 26608 15496 26660 15502
rect 26608 15438 26660 15444
rect 26712 14482 26740 15642
rect 26884 15496 26936 15502
rect 26884 15438 26936 15444
rect 26896 14618 26924 15438
rect 26884 14612 26936 14618
rect 26884 14554 26936 14560
rect 26700 14476 26752 14482
rect 26700 14418 26752 14424
rect 26712 13530 26740 14418
rect 26988 14385 27016 17614
rect 27080 15978 27108 18702
rect 27356 17678 27384 18702
rect 27540 18358 27568 18906
rect 27528 18352 27580 18358
rect 27528 18294 27580 18300
rect 27632 18170 27660 19790
rect 27816 18850 27844 20266
rect 28000 19310 28028 20334
rect 27988 19304 28040 19310
rect 27988 19246 28040 19252
rect 27540 18142 27660 18170
rect 27724 18822 27844 18850
rect 27344 17672 27396 17678
rect 27344 17614 27396 17620
rect 27160 17196 27212 17202
rect 27160 17138 27212 17144
rect 27344 17196 27396 17202
rect 27344 17138 27396 17144
rect 27172 16658 27200 17138
rect 27252 17060 27304 17066
rect 27252 17002 27304 17008
rect 27160 16652 27212 16658
rect 27160 16594 27212 16600
rect 27158 16280 27214 16289
rect 27158 16215 27160 16224
rect 27212 16215 27214 16224
rect 27160 16186 27212 16192
rect 27068 15972 27120 15978
rect 27068 15914 27120 15920
rect 27080 14618 27108 15914
rect 27160 14816 27212 14822
rect 27160 14758 27212 14764
rect 27068 14612 27120 14618
rect 27068 14554 27120 14560
rect 27172 14414 27200 14758
rect 27160 14408 27212 14414
rect 26974 14376 27030 14385
rect 27160 14350 27212 14356
rect 26974 14311 27030 14320
rect 27160 14272 27212 14278
rect 27160 14214 27212 14220
rect 27172 14074 27200 14214
rect 27160 14068 27212 14074
rect 27160 14010 27212 14016
rect 27160 13932 27212 13938
rect 27160 13874 27212 13880
rect 26700 13524 26752 13530
rect 26700 13466 26752 13472
rect 27172 13258 27200 13874
rect 27160 13252 27212 13258
rect 27160 13194 27212 13200
rect 26976 13184 27028 13190
rect 26976 13126 27028 13132
rect 26700 12844 26752 12850
rect 26700 12786 26752 12792
rect 26608 12436 26660 12442
rect 26608 12378 26660 12384
rect 26620 11801 26648 12378
rect 26606 11792 26662 11801
rect 26712 11762 26740 12786
rect 26988 11830 27016 13126
rect 27068 12368 27120 12374
rect 27068 12310 27120 12316
rect 27080 12102 27108 12310
rect 27160 12232 27212 12238
rect 27160 12174 27212 12180
rect 27068 12096 27120 12102
rect 27068 12038 27120 12044
rect 26792 11824 26844 11830
rect 26792 11766 26844 11772
rect 26976 11824 27028 11830
rect 26976 11766 27028 11772
rect 26606 11727 26662 11736
rect 26700 11756 26752 11762
rect 26700 11698 26752 11704
rect 26804 11150 26832 11766
rect 26976 11552 27028 11558
rect 26976 11494 27028 11500
rect 26988 11150 27016 11494
rect 27172 11354 27200 12174
rect 27160 11348 27212 11354
rect 27160 11290 27212 11296
rect 27160 11212 27212 11218
rect 27160 11154 27212 11160
rect 26608 11144 26660 11150
rect 26608 11086 26660 11092
rect 26792 11144 26844 11150
rect 26792 11086 26844 11092
rect 26976 11144 27028 11150
rect 26976 11086 27028 11092
rect 26620 10606 26648 11086
rect 26608 10600 26660 10606
rect 26608 10542 26660 10548
rect 26608 9920 26660 9926
rect 26608 9862 26660 9868
rect 26620 8906 26648 9862
rect 26608 8900 26660 8906
rect 26608 8842 26660 8848
rect 26620 8294 26648 8842
rect 26804 8362 26832 11086
rect 26976 11008 27028 11014
rect 26976 10950 27028 10956
rect 26988 10062 27016 10950
rect 27172 10266 27200 11154
rect 27160 10260 27212 10266
rect 27160 10202 27212 10208
rect 26976 10056 27028 10062
rect 26976 9998 27028 10004
rect 26976 9512 27028 9518
rect 26976 9454 27028 9460
rect 26988 8498 27016 9454
rect 27068 8832 27120 8838
rect 27068 8774 27120 8780
rect 26976 8492 27028 8498
rect 26976 8434 27028 8440
rect 26792 8356 26844 8362
rect 26792 8298 26844 8304
rect 26608 8288 26660 8294
rect 26608 8230 26660 8236
rect 27080 7886 27108 8774
rect 27264 8650 27292 17002
rect 27356 15910 27384 17138
rect 27436 16584 27488 16590
rect 27436 16526 27488 16532
rect 27448 16250 27476 16526
rect 27436 16244 27488 16250
rect 27436 16186 27488 16192
rect 27344 15904 27396 15910
rect 27344 15846 27396 15852
rect 27448 15706 27476 16186
rect 27436 15700 27488 15706
rect 27436 15642 27488 15648
rect 27540 14958 27568 18142
rect 27620 18080 27672 18086
rect 27620 18022 27672 18028
rect 27632 17882 27660 18022
rect 27620 17876 27672 17882
rect 27620 17818 27672 17824
rect 27618 17640 27674 17649
rect 27618 17575 27674 17584
rect 27528 14952 27580 14958
rect 27528 14894 27580 14900
rect 27436 14612 27488 14618
rect 27436 14554 27488 14560
rect 27448 13938 27476 14554
rect 27540 14414 27568 14894
rect 27632 14822 27660 17575
rect 27620 14816 27672 14822
rect 27620 14758 27672 14764
rect 27528 14408 27580 14414
rect 27528 14350 27580 14356
rect 27620 14272 27672 14278
rect 27620 14214 27672 14220
rect 27632 14074 27660 14214
rect 27620 14068 27672 14074
rect 27620 14010 27672 14016
rect 27436 13932 27488 13938
rect 27436 13874 27488 13880
rect 27344 13388 27396 13394
rect 27344 13330 27396 13336
rect 27356 12986 27384 13330
rect 27632 13326 27660 14010
rect 27620 13320 27672 13326
rect 27620 13262 27672 13268
rect 27344 12980 27396 12986
rect 27344 12922 27396 12928
rect 27356 11762 27384 12922
rect 27632 12782 27660 13262
rect 27724 13190 27752 18822
rect 27804 18760 27856 18766
rect 27804 18702 27856 18708
rect 27816 18426 27844 18702
rect 27804 18420 27856 18426
rect 27804 18362 27856 18368
rect 28092 17270 28120 22374
rect 28080 17264 28132 17270
rect 28080 17206 28132 17212
rect 28092 16590 28120 17206
rect 28080 16584 28132 16590
rect 28080 16526 28132 16532
rect 28080 16108 28132 16114
rect 28080 16050 28132 16056
rect 28092 15570 28120 16050
rect 28080 15564 28132 15570
rect 28080 15506 28132 15512
rect 27988 15020 28040 15026
rect 27988 14962 28040 14968
rect 27896 13728 27948 13734
rect 27896 13670 27948 13676
rect 27908 13394 27936 13670
rect 27896 13388 27948 13394
rect 27896 13330 27948 13336
rect 27712 13184 27764 13190
rect 27712 13126 27764 13132
rect 27804 12912 27856 12918
rect 27804 12854 27856 12860
rect 27712 12844 27764 12850
rect 27712 12786 27764 12792
rect 27620 12776 27672 12782
rect 27620 12718 27672 12724
rect 27528 12708 27580 12714
rect 27528 12650 27580 12656
rect 27540 12186 27568 12650
rect 27724 12238 27752 12786
rect 27816 12288 27844 12854
rect 27908 12782 27936 13330
rect 28000 13258 28028 14962
rect 28080 14272 28132 14278
rect 28080 14214 28132 14220
rect 28092 13938 28120 14214
rect 28080 13932 28132 13938
rect 28080 13874 28132 13880
rect 27988 13252 28040 13258
rect 27988 13194 28040 13200
rect 27896 12776 27948 12782
rect 27896 12718 27948 12724
rect 28000 12306 28028 13194
rect 27896 12300 27948 12306
rect 27816 12260 27896 12288
rect 27896 12242 27948 12248
rect 27988 12300 28040 12306
rect 27988 12242 28040 12248
rect 27448 12158 27568 12186
rect 27712 12232 27764 12238
rect 27712 12174 27764 12180
rect 27908 12186 27936 12242
rect 27908 12158 28028 12186
rect 27448 11898 27476 12158
rect 27528 12096 27580 12102
rect 27528 12038 27580 12044
rect 27436 11892 27488 11898
rect 27436 11834 27488 11840
rect 27344 11756 27396 11762
rect 27344 11698 27396 11704
rect 27540 11082 27568 12038
rect 27894 11928 27950 11937
rect 27894 11863 27950 11872
rect 27908 11830 27936 11863
rect 27896 11824 27948 11830
rect 27896 11766 27948 11772
rect 28000 11558 28028 12158
rect 28080 12096 28132 12102
rect 28080 12038 28132 12044
rect 28092 11937 28120 12038
rect 28078 11928 28134 11937
rect 28078 11863 28134 11872
rect 28080 11824 28132 11830
rect 28080 11766 28132 11772
rect 28092 11665 28120 11766
rect 28078 11656 28134 11665
rect 28078 11591 28134 11600
rect 27896 11552 27948 11558
rect 27896 11494 27948 11500
rect 27988 11552 28040 11558
rect 27988 11494 28040 11500
rect 27908 11218 27936 11494
rect 27896 11212 27948 11218
rect 27896 11154 27948 11160
rect 27528 11076 27580 11082
rect 27528 11018 27580 11024
rect 27540 10742 27568 11018
rect 27528 10736 27580 10742
rect 27528 10678 27580 10684
rect 27804 9580 27856 9586
rect 27804 9522 27856 9528
rect 27816 9382 27844 9522
rect 27908 9518 27936 11154
rect 27988 9580 28040 9586
rect 27988 9522 28040 9528
rect 27896 9512 27948 9518
rect 27896 9454 27948 9460
rect 27712 9376 27764 9382
rect 27712 9318 27764 9324
rect 27804 9376 27856 9382
rect 27804 9318 27856 9324
rect 27724 8974 27752 9318
rect 28000 9178 28028 9522
rect 27988 9172 28040 9178
rect 27988 9114 28040 9120
rect 27804 9036 27856 9042
rect 27804 8978 27856 8984
rect 27712 8968 27764 8974
rect 27712 8910 27764 8916
rect 27264 8622 27384 8650
rect 27252 8492 27304 8498
rect 27252 8434 27304 8440
rect 27264 8090 27292 8434
rect 27252 8084 27304 8090
rect 27252 8026 27304 8032
rect 26884 7880 26936 7886
rect 26884 7822 26936 7828
rect 27068 7880 27120 7886
rect 27252 7880 27304 7886
rect 27068 7822 27120 7828
rect 27250 7848 27252 7857
rect 27304 7848 27306 7857
rect 26896 7562 26924 7822
rect 27160 7812 27212 7818
rect 27250 7783 27306 7792
rect 27160 7754 27212 7760
rect 27172 7562 27200 7754
rect 26896 7534 27200 7562
rect 27356 2514 27384 8622
rect 27816 7954 27844 8978
rect 27896 8968 27948 8974
rect 27896 8910 27948 8916
rect 27804 7948 27856 7954
rect 27804 7890 27856 7896
rect 27908 7886 27936 8910
rect 27896 7880 27948 7886
rect 27896 7822 27948 7828
rect 27988 3664 28040 3670
rect 27908 3624 27988 3652
rect 27712 3596 27764 3602
rect 27908 3584 27936 3624
rect 27988 3606 28040 3612
rect 27764 3556 27936 3584
rect 27712 3538 27764 3544
rect 27436 3528 27488 3534
rect 27988 3528 28040 3534
rect 27436 3470 27488 3476
rect 27986 3496 27988 3505
rect 28040 3496 28042 3505
rect 27448 3398 27476 3470
rect 27986 3431 28042 3440
rect 27436 3392 27488 3398
rect 27436 3334 27488 3340
rect 28184 2990 28212 22902
rect 28276 21894 28304 23072
rect 28460 22642 28488 23666
rect 28448 22636 28500 22642
rect 28448 22578 28500 22584
rect 28552 22094 28580 24006
rect 28644 23594 28672 24647
rect 28632 23588 28684 23594
rect 28632 23530 28684 23536
rect 28632 23112 28684 23118
rect 28816 23112 28868 23118
rect 28684 23072 28764 23100
rect 28632 23054 28684 23060
rect 28460 22066 28580 22094
rect 28264 21888 28316 21894
rect 28264 21830 28316 21836
rect 28276 19378 28304 21830
rect 28356 19508 28408 19514
rect 28356 19450 28408 19456
rect 28264 19372 28316 19378
rect 28264 19314 28316 19320
rect 28276 18970 28304 19314
rect 28264 18964 28316 18970
rect 28264 18906 28316 18912
rect 28368 18834 28396 19450
rect 28356 18828 28408 18834
rect 28356 18770 28408 18776
rect 28264 18760 28316 18766
rect 28264 18702 28316 18708
rect 28276 18358 28304 18702
rect 28368 18358 28396 18770
rect 28264 18352 28316 18358
rect 28264 18294 28316 18300
rect 28356 18352 28408 18358
rect 28356 18294 28408 18300
rect 28276 16250 28304 18294
rect 28356 17740 28408 17746
rect 28356 17682 28408 17688
rect 28368 16794 28396 17682
rect 28356 16788 28408 16794
rect 28356 16730 28408 16736
rect 28264 16244 28316 16250
rect 28264 16186 28316 16192
rect 28276 15484 28304 16186
rect 28356 15496 28408 15502
rect 28276 15456 28356 15484
rect 28276 14890 28304 15456
rect 28356 15438 28408 15444
rect 28460 15026 28488 22066
rect 28632 20936 28684 20942
rect 28632 20878 28684 20884
rect 28644 19378 28672 20878
rect 28736 20516 28764 23072
rect 28920 23100 28948 24754
rect 28998 23896 29054 23905
rect 28998 23831 29054 23840
rect 29012 23798 29040 23831
rect 29000 23792 29052 23798
rect 29000 23734 29052 23740
rect 29104 23662 29132 49302
rect 29920 49156 29972 49162
rect 29920 49098 29972 49104
rect 29644 49088 29696 49094
rect 29644 49030 29696 49036
rect 29276 39296 29328 39302
rect 29276 39238 29328 39244
rect 29184 37800 29236 37806
rect 29184 37742 29236 37748
rect 29196 37466 29224 37742
rect 29184 37460 29236 37466
rect 29184 37402 29236 37408
rect 29184 36100 29236 36106
rect 29184 36042 29236 36048
rect 29196 35494 29224 36042
rect 29288 35494 29316 39238
rect 29656 38729 29684 49030
rect 29828 48680 29880 48686
rect 29828 48622 29880 48628
rect 29736 48136 29788 48142
rect 29736 48078 29788 48084
rect 29642 38720 29698 38729
rect 29642 38655 29698 38664
rect 29460 38344 29512 38350
rect 29460 38286 29512 38292
rect 29368 37868 29420 37874
rect 29368 37810 29420 37816
rect 29380 37670 29408 37810
rect 29472 37806 29500 38286
rect 29460 37800 29512 37806
rect 29460 37742 29512 37748
rect 29368 37664 29420 37670
rect 29368 37606 29420 37612
rect 29184 35488 29236 35494
rect 29184 35430 29236 35436
rect 29276 35488 29328 35494
rect 29276 35430 29328 35436
rect 29288 34746 29316 35430
rect 29276 34740 29328 34746
rect 29276 34682 29328 34688
rect 29288 34406 29316 34682
rect 29276 34400 29328 34406
rect 29276 34342 29328 34348
rect 29184 32496 29236 32502
rect 29184 32438 29236 32444
rect 29196 32298 29224 32438
rect 29184 32292 29236 32298
rect 29184 32234 29236 32240
rect 29380 31958 29408 37606
rect 29748 36106 29776 48078
rect 29840 47802 29868 48622
rect 29932 48278 29960 49098
rect 30024 48686 30052 49694
rect 30944 49298 30972 51200
rect 30656 49292 30708 49298
rect 30656 49234 30708 49240
rect 30932 49292 30984 49298
rect 30932 49234 30984 49240
rect 30012 48680 30064 48686
rect 30012 48622 30064 48628
rect 29920 48272 29972 48278
rect 29920 48214 29972 48220
rect 29828 47796 29880 47802
rect 29828 47738 29880 47744
rect 30012 47660 30064 47666
rect 30012 47602 30064 47608
rect 29828 47592 29880 47598
rect 29828 47534 29880 47540
rect 29840 47190 29868 47534
rect 29828 47184 29880 47190
rect 29828 47126 29880 47132
rect 29736 36100 29788 36106
rect 29736 36042 29788 36048
rect 29840 35986 29868 47126
rect 30024 47122 30052 47602
rect 30668 47190 30696 49234
rect 32128 49088 32180 49094
rect 32128 49030 32180 49036
rect 32140 48754 32168 49030
rect 32128 48748 32180 48754
rect 32128 48690 32180 48696
rect 32232 48210 32260 51200
rect 32312 48680 32364 48686
rect 33060 48668 33088 51326
rect 33506 51200 33562 52000
rect 34150 51354 34206 52000
rect 34794 51354 34850 52000
rect 33888 51326 34206 51354
rect 33324 49224 33376 49230
rect 33324 49166 33376 49172
rect 33140 48680 33192 48686
rect 33060 48640 33140 48668
rect 32312 48622 32364 48628
rect 33140 48622 33192 48628
rect 32220 48204 32272 48210
rect 32220 48146 32272 48152
rect 31024 48136 31076 48142
rect 31024 48078 31076 48084
rect 31036 47666 31064 48078
rect 32324 47802 32352 48622
rect 32496 48136 32548 48142
rect 32496 48078 32548 48084
rect 32312 47796 32364 47802
rect 32312 47738 32364 47744
rect 31852 47728 31904 47734
rect 31852 47670 31904 47676
rect 31024 47660 31076 47666
rect 31024 47602 31076 47608
rect 30748 47524 30800 47530
rect 30748 47466 30800 47472
rect 30760 47190 30788 47466
rect 30656 47184 30708 47190
rect 30656 47126 30708 47132
rect 30748 47184 30800 47190
rect 30748 47126 30800 47132
rect 30012 47116 30064 47122
rect 30012 47058 30064 47064
rect 31024 46980 31076 46986
rect 31024 46922 31076 46928
rect 30196 38956 30248 38962
rect 30196 38898 30248 38904
rect 30932 38956 30984 38962
rect 30932 38898 30984 38904
rect 29920 38208 29972 38214
rect 29918 38176 29920 38185
rect 30012 38208 30064 38214
rect 29972 38176 29974 38185
rect 30012 38150 30064 38156
rect 29918 38111 29974 38120
rect 30024 37670 30052 38150
rect 30012 37664 30064 37670
rect 30012 37606 30064 37612
rect 29920 37256 29972 37262
rect 29920 37198 29972 37204
rect 29656 35958 29868 35986
rect 29368 31952 29420 31958
rect 29368 31894 29420 31900
rect 29552 31952 29604 31958
rect 29552 31894 29604 31900
rect 29564 29714 29592 31894
rect 29552 29708 29604 29714
rect 29552 29650 29604 29656
rect 29552 28688 29604 28694
rect 29552 28630 29604 28636
rect 29564 28082 29592 28630
rect 29656 28234 29684 35958
rect 29736 35080 29788 35086
rect 29736 35022 29788 35028
rect 29748 33538 29776 35022
rect 29828 34944 29880 34950
rect 29828 34886 29880 34892
rect 29840 34678 29868 34886
rect 29828 34672 29880 34678
rect 29828 34614 29880 34620
rect 29932 34542 29960 37198
rect 30208 37126 30236 38898
rect 30288 37800 30340 37806
rect 30288 37742 30340 37748
rect 30300 37330 30328 37742
rect 30564 37664 30616 37670
rect 30564 37606 30616 37612
rect 30288 37324 30340 37330
rect 30288 37266 30340 37272
rect 30012 37120 30064 37126
rect 30012 37062 30064 37068
rect 30196 37120 30248 37126
rect 30196 37062 30248 37068
rect 30024 36718 30052 37062
rect 30300 36718 30328 37266
rect 30576 37194 30604 37606
rect 30564 37188 30616 37194
rect 30564 37130 30616 37136
rect 30944 37126 30972 38898
rect 30932 37120 30984 37126
rect 30932 37062 30984 37068
rect 30944 36786 30972 37062
rect 30932 36780 30984 36786
rect 30932 36722 30984 36728
rect 30012 36712 30064 36718
rect 30012 36654 30064 36660
rect 30288 36712 30340 36718
rect 30288 36654 30340 36660
rect 30024 34746 30052 36654
rect 30300 35562 30328 36654
rect 30288 35556 30340 35562
rect 30288 35498 30340 35504
rect 30300 35222 30328 35498
rect 30288 35216 30340 35222
rect 30288 35158 30340 35164
rect 30748 35080 30800 35086
rect 30748 35022 30800 35028
rect 30196 34944 30248 34950
rect 30196 34886 30248 34892
rect 30012 34740 30064 34746
rect 30012 34682 30064 34688
rect 30104 34604 30156 34610
rect 30104 34546 30156 34552
rect 29920 34536 29972 34542
rect 29840 34484 29920 34490
rect 29840 34478 29972 34484
rect 29840 34462 29960 34478
rect 29840 33998 29868 34462
rect 29828 33992 29880 33998
rect 29828 33934 29880 33940
rect 29840 33658 29868 33934
rect 30012 33924 30064 33930
rect 30012 33866 30064 33872
rect 29828 33652 29880 33658
rect 29828 33594 29880 33600
rect 30024 33538 30052 33866
rect 30116 33658 30144 34546
rect 30104 33652 30156 33658
rect 30104 33594 30156 33600
rect 29748 33510 30052 33538
rect 29736 32768 29788 32774
rect 29736 32710 29788 32716
rect 29748 32502 29776 32710
rect 29736 32496 29788 32502
rect 29736 32438 29788 32444
rect 29840 30326 29868 33510
rect 30116 32910 30144 33594
rect 30208 32910 30236 34886
rect 30288 34060 30340 34066
rect 30288 34002 30340 34008
rect 30300 32978 30328 34002
rect 30760 33998 30788 35022
rect 30944 34678 30972 36722
rect 31036 35222 31064 46922
rect 31116 38752 31168 38758
rect 31116 38694 31168 38700
rect 31128 37874 31156 38694
rect 31666 38448 31722 38457
rect 31300 38412 31352 38418
rect 31666 38383 31722 38392
rect 31300 38354 31352 38360
rect 31116 37868 31168 37874
rect 31116 37810 31168 37816
rect 31208 37800 31260 37806
rect 31312 37788 31340 38354
rect 31680 38350 31708 38383
rect 31484 38344 31536 38350
rect 31484 38286 31536 38292
rect 31668 38344 31720 38350
rect 31668 38286 31720 38292
rect 31392 38276 31444 38282
rect 31392 38218 31444 38224
rect 31260 37760 31340 37788
rect 31208 37742 31260 37748
rect 31312 37398 31340 37760
rect 31300 37392 31352 37398
rect 31300 37334 31352 37340
rect 31208 37188 31260 37194
rect 31208 37130 31260 37136
rect 31220 36650 31248 37130
rect 31208 36644 31260 36650
rect 31208 36586 31260 36592
rect 31312 36310 31340 37334
rect 31404 37330 31432 38218
rect 31496 37806 31524 38286
rect 31484 37800 31536 37806
rect 31484 37742 31536 37748
rect 31392 37324 31444 37330
rect 31392 37266 31444 37272
rect 31496 37262 31524 37742
rect 31576 37732 31628 37738
rect 31576 37674 31628 37680
rect 31484 37256 31536 37262
rect 31484 37198 31536 37204
rect 31300 36304 31352 36310
rect 31300 36246 31352 36252
rect 31116 36168 31168 36174
rect 31168 36128 31432 36156
rect 31116 36110 31168 36116
rect 31024 35216 31076 35222
rect 31024 35158 31076 35164
rect 30932 34672 30984 34678
rect 30932 34614 30984 34620
rect 30840 34400 30892 34406
rect 30840 34342 30892 34348
rect 30748 33992 30800 33998
rect 30748 33934 30800 33940
rect 30564 33856 30616 33862
rect 30564 33798 30616 33804
rect 30576 33590 30604 33798
rect 30564 33584 30616 33590
rect 30564 33526 30616 33532
rect 30380 33312 30432 33318
rect 30380 33254 30432 33260
rect 30288 32972 30340 32978
rect 30288 32914 30340 32920
rect 30104 32904 30156 32910
rect 30104 32846 30156 32852
rect 30196 32904 30248 32910
rect 30196 32846 30248 32852
rect 29920 32428 29972 32434
rect 29920 32370 29972 32376
rect 30012 32428 30064 32434
rect 30012 32370 30064 32376
rect 29932 32026 29960 32370
rect 29920 32020 29972 32026
rect 29920 31962 29972 31968
rect 29828 30320 29880 30326
rect 29828 30262 29880 30268
rect 29932 30122 29960 31962
rect 30024 31822 30052 32370
rect 30208 31890 30236 32846
rect 30300 32366 30328 32914
rect 30392 32910 30420 33254
rect 30576 32978 30604 33526
rect 30656 33516 30708 33522
rect 30656 33458 30708 33464
rect 30668 33114 30696 33458
rect 30656 33108 30708 33114
rect 30656 33050 30708 33056
rect 30564 32972 30616 32978
rect 30564 32914 30616 32920
rect 30380 32904 30432 32910
rect 30380 32846 30432 32852
rect 30656 32428 30708 32434
rect 30656 32370 30708 32376
rect 30288 32360 30340 32366
rect 30288 32302 30340 32308
rect 30668 32298 30696 32370
rect 30656 32292 30708 32298
rect 30656 32234 30708 32240
rect 30472 32224 30524 32230
rect 30472 32166 30524 32172
rect 30196 31884 30248 31890
rect 30196 31826 30248 31832
rect 30012 31816 30064 31822
rect 30012 31758 30064 31764
rect 30484 31346 30512 32166
rect 30668 31346 30696 32234
rect 30760 31414 30788 33934
rect 30852 33522 30880 34342
rect 30840 33516 30892 33522
rect 30840 33458 30892 33464
rect 31024 33516 31076 33522
rect 31024 33458 31076 33464
rect 31036 33114 31064 33458
rect 30932 33108 30984 33114
rect 30932 33050 30984 33056
rect 31024 33108 31076 33114
rect 31024 33050 31076 33056
rect 30748 31408 30800 31414
rect 30748 31350 30800 31356
rect 30472 31340 30524 31346
rect 30472 31282 30524 31288
rect 30656 31340 30708 31346
rect 30656 31282 30708 31288
rect 30472 31204 30524 31210
rect 30472 31146 30524 31152
rect 30484 30938 30512 31146
rect 30472 30932 30524 30938
rect 30472 30874 30524 30880
rect 30484 30734 30512 30874
rect 30472 30728 30524 30734
rect 30472 30670 30524 30676
rect 29920 30116 29972 30122
rect 30104 30116 30156 30122
rect 29972 30076 30052 30104
rect 29920 30058 29972 30064
rect 29920 29504 29972 29510
rect 29920 29446 29972 29452
rect 29932 29306 29960 29446
rect 30024 29306 30052 30076
rect 30104 30058 30156 30064
rect 29920 29300 29972 29306
rect 29920 29242 29972 29248
rect 30012 29300 30064 29306
rect 30012 29242 30064 29248
rect 29656 28206 29868 28234
rect 29552 28076 29604 28082
rect 29552 28018 29604 28024
rect 29736 28076 29788 28082
rect 29736 28018 29788 28024
rect 29644 27872 29696 27878
rect 29644 27814 29696 27820
rect 29656 27470 29684 27814
rect 29748 27674 29776 28018
rect 29736 27668 29788 27674
rect 29736 27610 29788 27616
rect 29644 27464 29696 27470
rect 29644 27406 29696 27412
rect 29840 26382 29868 28206
rect 29932 28014 29960 29242
rect 30116 28694 30144 30058
rect 30196 30048 30248 30054
rect 30196 29990 30248 29996
rect 30208 29714 30236 29990
rect 30196 29708 30248 29714
rect 30196 29650 30248 29656
rect 30380 29572 30432 29578
rect 30380 29514 30432 29520
rect 30104 28688 30156 28694
rect 30104 28630 30156 28636
rect 30392 28558 30420 29514
rect 30380 28552 30432 28558
rect 30380 28494 30432 28500
rect 29920 28008 29972 28014
rect 29920 27950 29972 27956
rect 30564 27600 30616 27606
rect 30564 27542 30616 27548
rect 30576 27130 30604 27542
rect 30564 27124 30616 27130
rect 30564 27066 30616 27072
rect 29920 26920 29972 26926
rect 29920 26862 29972 26868
rect 29932 26586 29960 26862
rect 29920 26580 29972 26586
rect 29920 26522 29972 26528
rect 29828 26376 29880 26382
rect 29828 26318 29880 26324
rect 30748 26376 30800 26382
rect 30748 26318 30800 26324
rect 29840 25974 29868 26318
rect 30196 26240 30248 26246
rect 30196 26182 30248 26188
rect 30380 26240 30432 26246
rect 30380 26182 30432 26188
rect 29828 25968 29880 25974
rect 29828 25910 29880 25916
rect 29840 25158 29868 25910
rect 30104 25832 30156 25838
rect 30104 25774 30156 25780
rect 30116 25498 30144 25774
rect 30208 25498 30236 26182
rect 30392 26042 30420 26182
rect 30380 26036 30432 26042
rect 30380 25978 30432 25984
rect 30104 25492 30156 25498
rect 30104 25434 30156 25440
rect 30196 25492 30248 25498
rect 30196 25434 30248 25440
rect 29828 25152 29880 25158
rect 29828 25094 29880 25100
rect 29276 24880 29328 24886
rect 29196 24840 29276 24868
rect 29196 24342 29224 24840
rect 29276 24822 29328 24828
rect 30392 24818 30420 25978
rect 30760 25906 30788 26318
rect 30748 25900 30800 25906
rect 30748 25842 30800 25848
rect 30760 25294 30788 25842
rect 30748 25288 30800 25294
rect 30748 25230 30800 25236
rect 29368 24812 29420 24818
rect 29368 24754 29420 24760
rect 30196 24812 30248 24818
rect 30196 24754 30248 24760
rect 30380 24812 30432 24818
rect 30380 24754 30432 24760
rect 29276 24676 29328 24682
rect 29276 24618 29328 24624
rect 29184 24336 29236 24342
rect 29184 24278 29236 24284
rect 29288 24290 29316 24618
rect 29380 24449 29408 24754
rect 29552 24744 29604 24750
rect 29552 24686 29604 24692
rect 29366 24440 29422 24449
rect 29366 24375 29422 24384
rect 29564 24290 29592 24686
rect 29828 24608 29880 24614
rect 29828 24550 29880 24556
rect 29288 24262 29592 24290
rect 29092 23656 29144 23662
rect 29092 23598 29144 23604
rect 29000 23112 29052 23118
rect 28920 23080 29000 23100
rect 29052 23080 29054 23089
rect 28920 23072 28998 23080
rect 28816 23054 28868 23060
rect 28828 22778 28856 23054
rect 29472 23050 29500 24262
rect 29840 24206 29868 24550
rect 29552 24200 29604 24206
rect 29552 24142 29604 24148
rect 29828 24200 29880 24206
rect 29828 24142 29880 24148
rect 29564 23882 29592 24142
rect 29564 23854 29776 23882
rect 29552 23724 29604 23730
rect 29552 23666 29604 23672
rect 29564 23322 29592 23666
rect 29748 23662 29776 23854
rect 29736 23656 29788 23662
rect 29736 23598 29788 23604
rect 29644 23520 29696 23526
rect 29644 23462 29696 23468
rect 29552 23316 29604 23322
rect 29552 23258 29604 23264
rect 28998 23015 29054 23024
rect 29460 23044 29512 23050
rect 29460 22986 29512 22992
rect 29656 22982 29684 23462
rect 29748 23322 29776 23598
rect 29736 23316 29788 23322
rect 29736 23258 29788 23264
rect 29368 22976 29420 22982
rect 29368 22918 29420 22924
rect 29644 22976 29696 22982
rect 29644 22918 29696 22924
rect 28816 22772 28868 22778
rect 28816 22714 28868 22720
rect 29380 22642 29408 22918
rect 29748 22710 29776 23258
rect 30208 23118 30236 24754
rect 30472 23860 30524 23866
rect 30472 23802 30524 23808
rect 30196 23112 30248 23118
rect 30194 23080 30196 23089
rect 30248 23080 30250 23089
rect 30194 23015 30250 23024
rect 29736 22704 29788 22710
rect 29736 22646 29788 22652
rect 30380 22704 30432 22710
rect 30380 22646 30432 22652
rect 29368 22636 29420 22642
rect 29368 22578 29420 22584
rect 30392 22234 30420 22646
rect 30380 22228 30432 22234
rect 30380 22170 30432 22176
rect 30378 21992 30434 22001
rect 30378 21927 30380 21936
rect 30432 21927 30434 21936
rect 30380 21898 30432 21904
rect 29000 20800 29052 20806
rect 29000 20742 29052 20748
rect 29012 20534 29040 20742
rect 29000 20528 29052 20534
rect 28736 20488 28856 20516
rect 28724 20324 28776 20330
rect 28724 20266 28776 20272
rect 28736 19854 28764 20266
rect 28724 19848 28776 19854
rect 28724 19790 28776 19796
rect 28632 19372 28684 19378
rect 28632 19314 28684 19320
rect 28644 18748 28672 19314
rect 28724 18760 28776 18766
rect 28644 18720 28724 18748
rect 28540 18284 28592 18290
rect 28540 18226 28592 18232
rect 28552 16658 28580 18226
rect 28644 17746 28672 18720
rect 28724 18702 28776 18708
rect 28724 18080 28776 18086
rect 28724 18022 28776 18028
rect 28632 17740 28684 17746
rect 28632 17682 28684 17688
rect 28540 16652 28592 16658
rect 28540 16594 28592 16600
rect 28632 16652 28684 16658
rect 28632 16594 28684 16600
rect 28644 15994 28672 16594
rect 28736 16046 28764 18022
rect 28552 15978 28672 15994
rect 28724 16040 28776 16046
rect 28724 15982 28776 15988
rect 28540 15972 28672 15978
rect 28592 15966 28672 15972
rect 28540 15914 28592 15920
rect 28448 15020 28500 15026
rect 28448 14962 28500 14968
rect 28264 14884 28316 14890
rect 28264 14826 28316 14832
rect 28448 14544 28500 14550
rect 28448 14486 28500 14492
rect 28356 14408 28408 14414
rect 28354 14376 28356 14385
rect 28408 14376 28410 14385
rect 28354 14311 28410 14320
rect 28460 12238 28488 14486
rect 28552 13394 28580 15914
rect 28736 15366 28764 15982
rect 28724 15360 28776 15366
rect 28724 15302 28776 15308
rect 28632 13932 28684 13938
rect 28632 13874 28684 13880
rect 28540 13388 28592 13394
rect 28540 13330 28592 13336
rect 28540 13184 28592 13190
rect 28540 13126 28592 13132
rect 28552 12374 28580 13126
rect 28644 12850 28672 13874
rect 28632 12844 28684 12850
rect 28632 12786 28684 12792
rect 28828 12434 28856 20488
rect 29000 20470 29052 20476
rect 29012 19786 29040 20470
rect 30484 20466 30512 23802
rect 30656 22160 30708 22166
rect 30654 22128 30656 22137
rect 30708 22128 30710 22137
rect 30654 22063 30710 22072
rect 30745 22024 30797 22030
rect 30745 21966 30797 21972
rect 30760 21486 30788 21966
rect 30748 21480 30800 21486
rect 30748 21422 30800 21428
rect 30760 21010 30788 21422
rect 30748 21004 30800 21010
rect 30748 20946 30800 20952
rect 29184 20460 29236 20466
rect 29184 20402 29236 20408
rect 30472 20460 30524 20466
rect 30472 20402 30524 20408
rect 29092 20256 29144 20262
rect 29092 20198 29144 20204
rect 29000 19780 29052 19786
rect 29000 19722 29052 19728
rect 28908 19372 28960 19378
rect 28908 19314 28960 19320
rect 28920 18970 28948 19314
rect 28908 18964 28960 18970
rect 28908 18906 28960 18912
rect 29012 18222 29040 19722
rect 29000 18216 29052 18222
rect 29000 18158 29052 18164
rect 29104 17338 29132 20198
rect 29196 19446 29224 20402
rect 30380 20392 30432 20398
rect 30380 20334 30432 20340
rect 30392 19854 30420 20334
rect 30380 19848 30432 19854
rect 30380 19790 30432 19796
rect 29184 19440 29236 19446
rect 29184 19382 29236 19388
rect 29644 17604 29696 17610
rect 29644 17546 29696 17552
rect 29092 17332 29144 17338
rect 29092 17274 29144 17280
rect 29460 17264 29512 17270
rect 29460 17206 29512 17212
rect 28908 16788 28960 16794
rect 28908 16730 28960 16736
rect 28920 16250 28948 16730
rect 29472 16590 29500 17206
rect 29552 16992 29604 16998
rect 29552 16934 29604 16940
rect 29460 16584 29512 16590
rect 29460 16526 29512 16532
rect 28908 16244 28960 16250
rect 28908 16186 28960 16192
rect 29000 16108 29052 16114
rect 28920 16068 29000 16096
rect 28920 14550 28948 16068
rect 29000 16050 29052 16056
rect 29184 16040 29236 16046
rect 29184 15982 29236 15988
rect 29092 15972 29144 15978
rect 29092 15914 29144 15920
rect 29104 15638 29132 15914
rect 29196 15910 29224 15982
rect 29564 15910 29592 16934
rect 29656 16250 29684 17546
rect 29828 17536 29880 17542
rect 29828 17478 29880 17484
rect 29840 16590 29868 17478
rect 30288 17196 30340 17202
rect 30288 17138 30340 17144
rect 30196 16992 30248 16998
rect 30196 16934 30248 16940
rect 30208 16590 30236 16934
rect 30300 16794 30328 17138
rect 30288 16788 30340 16794
rect 30288 16730 30340 16736
rect 29828 16584 29880 16590
rect 29828 16526 29880 16532
rect 30196 16584 30248 16590
rect 30196 16526 30248 16532
rect 30380 16516 30432 16522
rect 30380 16458 30432 16464
rect 30392 16289 30420 16458
rect 30378 16280 30434 16289
rect 29644 16244 29696 16250
rect 30378 16215 30434 16224
rect 29644 16186 29696 16192
rect 29184 15904 29236 15910
rect 29184 15846 29236 15852
rect 29552 15904 29604 15910
rect 29552 15846 29604 15852
rect 29092 15632 29144 15638
rect 29092 15574 29144 15580
rect 29196 15502 29224 15846
rect 29564 15502 29592 15846
rect 29184 15496 29236 15502
rect 29184 15438 29236 15444
rect 29552 15496 29604 15502
rect 29552 15438 29604 15444
rect 28908 14544 28960 14550
rect 28908 14486 28960 14492
rect 29564 14006 29592 15438
rect 29552 14000 29604 14006
rect 29552 13942 29604 13948
rect 28908 13728 28960 13734
rect 28908 13670 28960 13676
rect 28920 12986 28948 13670
rect 30484 13326 30512 20402
rect 30760 19990 30788 20946
rect 30748 19984 30800 19990
rect 30748 19926 30800 19932
rect 30748 16448 30800 16454
rect 30748 16390 30800 16396
rect 30760 16114 30788 16390
rect 30840 16176 30892 16182
rect 30840 16118 30892 16124
rect 30748 16108 30800 16114
rect 30748 16050 30800 16056
rect 30852 16046 30880 16118
rect 30840 16040 30892 16046
rect 30840 15982 30892 15988
rect 30852 15026 30880 15982
rect 30840 15020 30892 15026
rect 30840 14962 30892 14968
rect 30748 13728 30800 13734
rect 30748 13670 30800 13676
rect 30760 13326 30788 13670
rect 30472 13320 30524 13326
rect 30472 13262 30524 13268
rect 30748 13320 30800 13326
rect 30748 13262 30800 13268
rect 28908 12980 28960 12986
rect 28908 12922 28960 12928
rect 28736 12406 28856 12434
rect 28540 12368 28592 12374
rect 28540 12310 28592 12316
rect 28552 12238 28580 12310
rect 28264 12232 28316 12238
rect 28264 12174 28316 12180
rect 28448 12232 28500 12238
rect 28448 12174 28500 12180
rect 28540 12232 28592 12238
rect 28540 12174 28592 12180
rect 28276 9382 28304 12174
rect 28356 11756 28408 11762
rect 28356 11698 28408 11704
rect 28368 11014 28396 11698
rect 28356 11008 28408 11014
rect 28356 10950 28408 10956
rect 28264 9376 28316 9382
rect 28264 9318 28316 9324
rect 28736 3194 28764 12406
rect 28920 11150 28948 12922
rect 30484 12442 30512 13262
rect 30564 13184 30616 13190
rect 30564 13126 30616 13132
rect 30472 12436 30524 12442
rect 30472 12378 30524 12384
rect 30380 12368 30432 12374
rect 30380 12310 30432 12316
rect 30392 11796 30420 12310
rect 30380 11790 30432 11796
rect 30380 11732 30432 11738
rect 30472 11756 30524 11762
rect 30472 11698 30524 11704
rect 29644 11688 29696 11694
rect 29644 11630 29696 11636
rect 29552 11212 29604 11218
rect 29552 11154 29604 11160
rect 28908 11144 28960 11150
rect 28908 11086 28960 11092
rect 29564 10606 29592 11154
rect 29656 11082 29684 11630
rect 29736 11620 29788 11626
rect 29736 11562 29788 11568
rect 29644 11076 29696 11082
rect 29644 11018 29696 11024
rect 29552 10600 29604 10606
rect 29552 10542 29604 10548
rect 29748 8498 29776 11562
rect 30012 11552 30064 11558
rect 30012 11494 30064 11500
rect 30104 11552 30156 11558
rect 30104 11494 30156 11500
rect 30024 10742 30052 11494
rect 30116 11286 30144 11494
rect 30484 11354 30512 11698
rect 30576 11694 30604 13126
rect 30840 12844 30892 12850
rect 30840 12786 30892 12792
rect 30852 12374 30880 12786
rect 30840 12368 30892 12374
rect 30840 12310 30892 12316
rect 30656 12164 30708 12170
rect 30656 12106 30708 12112
rect 30668 11762 30696 12106
rect 30748 12096 30800 12102
rect 30748 12038 30800 12044
rect 30656 11756 30708 11762
rect 30656 11698 30708 11704
rect 30564 11688 30616 11694
rect 30564 11630 30616 11636
rect 30472 11348 30524 11354
rect 30472 11290 30524 11296
rect 30104 11280 30156 11286
rect 30104 11222 30156 11228
rect 30760 11150 30788 12038
rect 30748 11144 30800 11150
rect 30748 11086 30800 11092
rect 30380 11076 30432 11082
rect 30380 11018 30432 11024
rect 30012 10736 30064 10742
rect 30012 10678 30064 10684
rect 30392 10470 30420 11018
rect 30380 10464 30432 10470
rect 30380 10406 30432 10412
rect 30012 9376 30064 9382
rect 30012 9318 30064 9324
rect 30024 9042 30052 9318
rect 30012 9036 30064 9042
rect 30012 8978 30064 8984
rect 30288 9036 30340 9042
rect 30288 8978 30340 8984
rect 30300 8634 30328 8978
rect 30392 8906 30420 10406
rect 30656 9376 30708 9382
rect 30656 9318 30708 9324
rect 30380 8900 30432 8906
rect 30380 8842 30432 8848
rect 30288 8628 30340 8634
rect 30288 8570 30340 8576
rect 30668 8566 30696 9318
rect 30656 8560 30708 8566
rect 30656 8502 30708 8508
rect 29736 8492 29788 8498
rect 29736 8434 29788 8440
rect 29828 8356 29880 8362
rect 29828 8298 29880 8304
rect 28816 4072 28868 4078
rect 28816 4014 28868 4020
rect 28908 4072 28960 4078
rect 28908 4014 28960 4020
rect 28828 3534 28856 4014
rect 28816 3528 28868 3534
rect 28816 3470 28868 3476
rect 28724 3188 28776 3194
rect 28724 3130 28776 3136
rect 28172 2984 28224 2990
rect 28172 2926 28224 2932
rect 28920 2854 28948 4014
rect 29552 3936 29604 3942
rect 29552 3878 29604 3884
rect 29736 3936 29788 3942
rect 29736 3878 29788 3884
rect 28908 2848 28960 2854
rect 28908 2790 28960 2796
rect 29564 2514 29592 3878
rect 29644 3392 29696 3398
rect 29644 3334 29696 3340
rect 29656 2938 29684 3334
rect 29748 3058 29776 3878
rect 29736 3052 29788 3058
rect 29736 2994 29788 3000
rect 29656 2910 29776 2938
rect 29644 2848 29696 2854
rect 29644 2790 29696 2796
rect 27344 2508 27396 2514
rect 27344 2450 27396 2456
rect 29552 2508 29604 2514
rect 29552 2450 29604 2456
rect 27068 2440 27120 2446
rect 27712 2440 27764 2446
rect 27068 2382 27120 2388
rect 26516 2372 26568 2378
rect 26516 2314 26568 2320
rect 27080 800 27108 2382
rect 27172 2378 27568 2394
rect 27712 2382 27764 2388
rect 27160 2372 27580 2378
rect 27212 2366 27528 2372
rect 27160 2314 27212 2320
rect 27528 2314 27580 2320
rect 27724 800 27752 2382
rect 29656 800 29684 2790
rect 29748 2514 29776 2910
rect 29840 2854 29868 8298
rect 30748 5228 30800 5234
rect 30748 5170 30800 5176
rect 30760 4146 30788 5170
rect 30748 4140 30800 4146
rect 30748 4082 30800 4088
rect 29920 3392 29972 3398
rect 29920 3334 29972 3340
rect 29932 3126 29960 3334
rect 29920 3120 29972 3126
rect 29920 3062 29972 3068
rect 30288 2984 30340 2990
rect 30288 2926 30340 2932
rect 29828 2848 29880 2854
rect 29828 2790 29880 2796
rect 29736 2508 29788 2514
rect 29736 2450 29788 2456
rect 30300 800 30328 2926
rect 30944 2774 30972 33050
rect 31208 31816 31260 31822
rect 31208 31758 31260 31764
rect 31220 31278 31248 31758
rect 31208 31272 31260 31278
rect 31208 31214 31260 31220
rect 31024 30796 31076 30802
rect 31024 30738 31076 30744
rect 31036 29578 31064 30738
rect 31024 29572 31076 29578
rect 31024 29514 31076 29520
rect 31024 28960 31076 28966
rect 31024 28902 31076 28908
rect 31036 28490 31064 28902
rect 31220 28762 31248 31214
rect 31300 31136 31352 31142
rect 31300 31078 31352 31084
rect 31312 30870 31340 31078
rect 31300 30864 31352 30870
rect 31300 30806 31352 30812
rect 31208 28756 31260 28762
rect 31208 28698 31260 28704
rect 31220 28490 31248 28698
rect 31024 28484 31076 28490
rect 31024 28426 31076 28432
rect 31208 28484 31260 28490
rect 31208 28426 31260 28432
rect 31208 27396 31260 27402
rect 31208 27338 31260 27344
rect 31220 26314 31248 27338
rect 31116 26308 31168 26314
rect 31116 26250 31168 26256
rect 31208 26308 31260 26314
rect 31208 26250 31260 26256
rect 31024 23792 31076 23798
rect 31024 23734 31076 23740
rect 31036 16182 31064 23734
rect 31128 22094 31156 26250
rect 31404 22094 31432 36128
rect 31496 35494 31524 37198
rect 31588 36174 31616 37674
rect 31864 36564 31892 47670
rect 32508 47598 32536 48078
rect 33336 47666 33364 49166
rect 33416 48612 33468 48618
rect 33416 48554 33468 48560
rect 33324 47660 33376 47666
rect 33324 47602 33376 47608
rect 32496 47592 32548 47598
rect 32496 47534 32548 47540
rect 31944 38344 31996 38350
rect 31944 38286 31996 38292
rect 32128 38344 32180 38350
rect 32128 38286 32180 38292
rect 31956 36922 31984 38286
rect 32036 38208 32088 38214
rect 32034 38176 32036 38185
rect 32088 38176 32090 38185
rect 32034 38111 32090 38120
rect 32036 37732 32088 37738
rect 32140 37720 32168 38286
rect 32088 37692 32168 37720
rect 32036 37674 32088 37680
rect 31944 36916 31996 36922
rect 31944 36858 31996 36864
rect 31772 36536 31892 36564
rect 31576 36168 31628 36174
rect 31576 36110 31628 36116
rect 31484 35488 31536 35494
rect 31484 35430 31536 35436
rect 31588 35222 31616 36110
rect 31668 36100 31720 36106
rect 31668 36042 31720 36048
rect 31576 35216 31628 35222
rect 31576 35158 31628 35164
rect 31680 35154 31708 36042
rect 31668 35148 31720 35154
rect 31668 35090 31720 35096
rect 31574 35048 31630 35057
rect 31574 34983 31576 34992
rect 31628 34983 31630 34992
rect 31668 35012 31720 35018
rect 31576 34954 31628 34960
rect 31668 34954 31720 34960
rect 31680 32026 31708 34954
rect 31668 32020 31720 32026
rect 31668 31962 31720 31968
rect 31772 29510 31800 36536
rect 31852 36236 31904 36242
rect 31852 36178 31904 36184
rect 31864 35766 31892 36178
rect 32036 36032 32088 36038
rect 32036 35974 32088 35980
rect 32048 35766 32076 35974
rect 32864 35828 32916 35834
rect 32864 35770 32916 35776
rect 31852 35760 31904 35766
rect 31852 35702 31904 35708
rect 32036 35760 32088 35766
rect 32036 35702 32088 35708
rect 32876 35494 32904 35770
rect 32496 35488 32548 35494
rect 32496 35430 32548 35436
rect 32864 35488 32916 35494
rect 32864 35430 32916 35436
rect 32508 35086 32536 35430
rect 32496 35080 32548 35086
rect 32496 35022 32548 35028
rect 32508 33454 32536 35022
rect 32312 33448 32364 33454
rect 32312 33390 32364 33396
rect 32496 33448 32548 33454
rect 32496 33390 32548 33396
rect 32324 32842 32352 33390
rect 32404 33108 32456 33114
rect 32404 33050 32456 33056
rect 32312 32836 32364 32842
rect 32312 32778 32364 32784
rect 32324 31890 32352 32778
rect 32312 31884 32364 31890
rect 32312 31826 32364 31832
rect 32416 31822 32444 33050
rect 32508 32434 32536 33390
rect 32588 32768 32640 32774
rect 32588 32710 32640 32716
rect 32496 32428 32548 32434
rect 32496 32370 32548 32376
rect 31852 31816 31904 31822
rect 31852 31758 31904 31764
rect 32220 31816 32272 31822
rect 32220 31758 32272 31764
rect 32404 31816 32456 31822
rect 32404 31758 32456 31764
rect 31576 29504 31628 29510
rect 31576 29446 31628 29452
rect 31760 29504 31812 29510
rect 31760 29446 31812 29452
rect 31588 29306 31616 29446
rect 31576 29300 31628 29306
rect 31576 29242 31628 29248
rect 31760 29300 31812 29306
rect 31760 29242 31812 29248
rect 31772 28490 31800 29242
rect 31760 28484 31812 28490
rect 31760 28426 31812 28432
rect 31680 26206 31800 26234
rect 31484 25288 31536 25294
rect 31484 25230 31536 25236
rect 31496 24886 31524 25230
rect 31680 25226 31708 26206
rect 31772 26042 31800 26206
rect 31760 26036 31812 26042
rect 31760 25978 31812 25984
rect 31668 25220 31720 25226
rect 31668 25162 31720 25168
rect 31484 24880 31536 24886
rect 31484 24822 31536 24828
rect 31484 22160 31536 22166
rect 31576 22160 31628 22166
rect 31484 22102 31536 22108
rect 31574 22128 31576 22137
rect 31628 22128 31630 22137
rect 31128 22066 31248 22094
rect 31024 16176 31076 16182
rect 31024 16118 31076 16124
rect 31024 16040 31076 16046
rect 31024 15982 31076 15988
rect 31036 15094 31064 15982
rect 31116 15496 31168 15502
rect 31116 15438 31168 15444
rect 31024 15088 31076 15094
rect 31024 15030 31076 15036
rect 31036 14074 31064 15030
rect 31024 14068 31076 14074
rect 31024 14010 31076 14016
rect 31036 12850 31064 14010
rect 31128 13394 31156 15438
rect 31116 13388 31168 13394
rect 31116 13330 31168 13336
rect 31024 12844 31076 12850
rect 31024 12786 31076 12792
rect 31220 7546 31248 22066
rect 31312 22066 31432 22094
rect 31312 12434 31340 22066
rect 31496 22012 31524 22102
rect 31574 22063 31630 22072
rect 31496 21984 31616 22012
rect 31484 21888 31536 21894
rect 31484 21830 31536 21836
rect 31496 21622 31524 21830
rect 31484 21616 31536 21622
rect 31484 21558 31536 21564
rect 31588 21554 31616 21984
rect 31392 21548 31444 21554
rect 31392 21490 31444 21496
rect 31576 21548 31628 21554
rect 31576 21490 31628 21496
rect 31404 21146 31432 21490
rect 31484 21480 31536 21486
rect 31484 21422 31536 21428
rect 31392 21140 31444 21146
rect 31392 21082 31444 21088
rect 31496 20942 31524 21422
rect 31484 20936 31536 20942
rect 31484 20878 31536 20884
rect 31588 20788 31616 21490
rect 31496 20760 31616 20788
rect 31496 19786 31524 20760
rect 31484 19780 31536 19786
rect 31484 19722 31536 19728
rect 31576 19712 31628 19718
rect 31576 19654 31628 19660
rect 31588 18766 31616 19654
rect 31576 18760 31628 18766
rect 31576 18702 31628 18708
rect 31680 16674 31708 25162
rect 31864 22094 31892 31758
rect 32232 31482 32260 31758
rect 32220 31476 32272 31482
rect 32220 31418 32272 31424
rect 32128 31340 32180 31346
rect 32128 31282 32180 31288
rect 31944 30728 31996 30734
rect 31944 30670 31996 30676
rect 31956 28558 31984 30670
rect 32140 30394 32168 31282
rect 32312 30592 32364 30598
rect 32312 30534 32364 30540
rect 32128 30388 32180 30394
rect 32128 30330 32180 30336
rect 32324 29646 32352 30534
rect 32600 30326 32628 32710
rect 32772 32428 32824 32434
rect 32772 32370 32824 32376
rect 32784 32026 32812 32370
rect 32772 32020 32824 32026
rect 32772 31962 32824 31968
rect 32876 31754 32904 35430
rect 33046 35048 33102 35057
rect 33046 34983 33048 34992
rect 33100 34983 33102 34992
rect 33048 34954 33100 34960
rect 32956 33652 33008 33658
rect 32956 33594 33008 33600
rect 32692 31726 32904 31754
rect 32588 30320 32640 30326
rect 32588 30262 32640 30268
rect 32036 29640 32088 29646
rect 32036 29582 32088 29588
rect 32312 29640 32364 29646
rect 32312 29582 32364 29588
rect 32048 28762 32076 29582
rect 32404 29572 32456 29578
rect 32404 29514 32456 29520
rect 32128 29504 32180 29510
rect 32128 29446 32180 29452
rect 32036 28756 32088 28762
rect 32036 28698 32088 28704
rect 31944 28552 31996 28558
rect 31944 28494 31996 28500
rect 32036 28076 32088 28082
rect 32036 28018 32088 28024
rect 32048 27674 32076 28018
rect 32036 27668 32088 27674
rect 32036 27610 32088 27616
rect 32140 26042 32168 29446
rect 32416 27448 32444 29514
rect 32588 28552 32640 28558
rect 32588 28494 32640 28500
rect 32600 28014 32628 28494
rect 32588 28008 32640 28014
rect 32588 27950 32640 27956
rect 32404 27442 32456 27448
rect 32404 27384 32456 27390
rect 32218 26888 32274 26897
rect 32218 26823 32274 26832
rect 32232 26790 32260 26823
rect 32220 26784 32272 26790
rect 32220 26726 32272 26732
rect 32404 26784 32456 26790
rect 32404 26726 32456 26732
rect 32128 26036 32180 26042
rect 32128 25978 32180 25984
rect 32416 25906 32444 26726
rect 32600 26042 32628 27950
rect 32692 26994 32720 31726
rect 32772 29640 32824 29646
rect 32772 29582 32824 29588
rect 32784 27470 32812 29582
rect 32968 29306 32996 33594
rect 33048 33516 33100 33522
rect 33048 33458 33100 33464
rect 33060 33114 33088 33458
rect 33048 33108 33100 33114
rect 33048 33050 33100 33056
rect 33324 32904 33376 32910
rect 33324 32846 33376 32852
rect 33336 32434 33364 32846
rect 33324 32428 33376 32434
rect 33324 32370 33376 32376
rect 33324 30592 33376 30598
rect 33324 30534 33376 30540
rect 33048 30320 33100 30326
rect 33048 30262 33100 30268
rect 32956 29300 33008 29306
rect 32956 29242 33008 29248
rect 33060 28150 33088 30262
rect 33336 30258 33364 30534
rect 33324 30252 33376 30258
rect 33324 30194 33376 30200
rect 33324 30048 33376 30054
rect 33324 29990 33376 29996
rect 33336 29238 33364 29990
rect 33232 29232 33284 29238
rect 33232 29174 33284 29180
rect 33324 29232 33376 29238
rect 33324 29174 33376 29180
rect 33244 28762 33272 29174
rect 33232 28756 33284 28762
rect 33232 28698 33284 28704
rect 33048 28144 33100 28150
rect 33048 28086 33100 28092
rect 32772 27464 32824 27470
rect 33060 27418 33088 28086
rect 33140 27668 33192 27674
rect 33140 27610 33192 27616
rect 32772 27406 32824 27412
rect 32968 27390 33088 27418
rect 32680 26988 32732 26994
rect 32680 26930 32732 26936
rect 32864 26988 32916 26994
rect 32864 26930 32916 26936
rect 32876 26790 32904 26930
rect 32968 26926 32996 27390
rect 33152 26994 33180 27610
rect 33140 26988 33192 26994
rect 33140 26930 33192 26936
rect 32956 26920 33008 26926
rect 32956 26862 33008 26868
rect 33244 26858 33272 28698
rect 33324 27396 33376 27402
rect 33324 27338 33376 27344
rect 33232 26852 33284 26858
rect 33232 26794 33284 26800
rect 32772 26784 32824 26790
rect 32772 26726 32824 26732
rect 32864 26784 32916 26790
rect 32864 26726 32916 26732
rect 32784 26330 32812 26726
rect 32876 26450 32904 26726
rect 32864 26444 32916 26450
rect 32864 26386 32916 26392
rect 32784 26302 32904 26330
rect 32588 26036 32640 26042
rect 32588 25978 32640 25984
rect 32220 25900 32272 25906
rect 32220 25842 32272 25848
rect 32404 25900 32456 25906
rect 32404 25842 32456 25848
rect 32128 25832 32180 25838
rect 32128 25774 32180 25780
rect 32140 23322 32168 25774
rect 32232 24818 32260 25842
rect 32772 25152 32824 25158
rect 32772 25094 32824 25100
rect 32220 24812 32272 24818
rect 32220 24754 32272 24760
rect 32784 24614 32812 25094
rect 32496 24608 32548 24614
rect 32496 24550 32548 24556
rect 32772 24608 32824 24614
rect 32772 24550 32824 24556
rect 32508 24274 32536 24550
rect 32678 24440 32734 24449
rect 32784 24410 32812 24550
rect 32678 24375 32734 24384
rect 32772 24404 32824 24410
rect 32692 24342 32720 24375
rect 32772 24346 32824 24352
rect 32680 24336 32732 24342
rect 32680 24278 32732 24284
rect 32496 24268 32548 24274
rect 32496 24210 32548 24216
rect 32312 24200 32364 24206
rect 32312 24142 32364 24148
rect 32402 24168 32458 24177
rect 32324 23905 32352 24142
rect 32402 24103 32458 24112
rect 32310 23896 32366 23905
rect 32310 23831 32366 23840
rect 32416 23798 32444 24103
rect 32404 23792 32456 23798
rect 32404 23734 32456 23740
rect 32128 23316 32180 23322
rect 32128 23258 32180 23264
rect 32140 22642 32168 23258
rect 32128 22636 32180 22642
rect 32128 22578 32180 22584
rect 31772 22066 31892 22094
rect 32036 22092 32088 22098
rect 31772 21842 31800 22066
rect 32876 22094 32904 26302
rect 33336 26042 33364 27338
rect 33428 26874 33456 48554
rect 33520 48498 33548 51200
rect 33888 48618 33916 51326
rect 34150 51200 34206 51326
rect 34716 51326 34850 51354
rect 33876 48612 33928 48618
rect 33876 48554 33928 48560
rect 33520 48470 34468 48498
rect 33508 48000 33560 48006
rect 33508 47942 33560 47948
rect 33520 47734 33548 47942
rect 33508 47728 33560 47734
rect 33508 47670 33560 47676
rect 34440 41414 34468 48470
rect 34716 47598 34744 51326
rect 34794 51200 34850 51326
rect 35438 51200 35494 52000
rect 36082 51200 36138 52000
rect 36726 51200 36782 52000
rect 37370 51354 37426 52000
rect 38014 51354 38070 52000
rect 37370 51326 37688 51354
rect 37370 51200 37426 51326
rect 34934 49532 35242 49552
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49456 35242 49476
rect 35808 49224 35860 49230
rect 35808 49166 35860 49172
rect 34888 49156 34940 49162
rect 34888 49098 34940 49104
rect 34900 48754 34928 49098
rect 34888 48748 34940 48754
rect 34888 48690 34940 48696
rect 34934 48444 35242 48464
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48368 35242 48388
rect 35820 48210 35848 49166
rect 36096 48686 36124 51200
rect 35900 48680 35952 48686
rect 35900 48622 35952 48628
rect 36084 48680 36136 48686
rect 36084 48622 36136 48628
rect 35808 48204 35860 48210
rect 35808 48146 35860 48152
rect 34796 48136 34848 48142
rect 34796 48078 34848 48084
rect 34704 47592 34756 47598
rect 34704 47534 34756 47540
rect 34520 47456 34572 47462
rect 34520 47398 34572 47404
rect 34532 45898 34560 47398
rect 34520 45892 34572 45898
rect 34520 45834 34572 45840
rect 34164 41386 34468 41414
rect 33508 32904 33560 32910
rect 33508 32846 33560 32852
rect 33520 32570 33548 32846
rect 33508 32564 33560 32570
rect 33508 32506 33560 32512
rect 33876 32428 33928 32434
rect 33876 32370 33928 32376
rect 33508 31884 33560 31890
rect 33508 31826 33560 31832
rect 33520 30190 33548 31826
rect 33508 30184 33560 30190
rect 33508 30126 33560 30132
rect 33520 29102 33548 30126
rect 33508 29096 33560 29102
rect 33508 29038 33560 29044
rect 33692 29028 33744 29034
rect 33692 28970 33744 28976
rect 33704 28558 33732 28970
rect 33692 28552 33744 28558
rect 33692 28494 33744 28500
rect 33692 27056 33744 27062
rect 33692 26998 33744 27004
rect 33704 26897 33732 26998
rect 33690 26888 33746 26897
rect 33428 26846 33640 26874
rect 33324 26036 33376 26042
rect 33324 25978 33376 25984
rect 33336 24818 33364 25978
rect 33140 24812 33192 24818
rect 33140 24754 33192 24760
rect 33324 24812 33376 24818
rect 33324 24754 33376 24760
rect 33152 24274 33180 24754
rect 33140 24268 33192 24274
rect 33140 24210 33192 24216
rect 33152 23118 33180 24210
rect 33232 23656 33284 23662
rect 33232 23598 33284 23604
rect 33416 23656 33468 23662
rect 33416 23598 33468 23604
rect 33140 23112 33192 23118
rect 33140 23054 33192 23060
rect 33244 22506 33272 23598
rect 33428 23322 33456 23598
rect 33416 23316 33468 23322
rect 33416 23258 33468 23264
rect 33232 22500 33284 22506
rect 33232 22442 33284 22448
rect 33508 22500 33560 22506
rect 33508 22442 33560 22448
rect 32876 22066 32996 22094
rect 32036 22034 32088 22040
rect 32048 22001 32076 22034
rect 32128 22024 32180 22030
rect 32034 21992 32090 22001
rect 32128 21966 32180 21972
rect 32588 22024 32640 22030
rect 32588 21966 32640 21972
rect 32034 21927 32090 21936
rect 31772 21814 31892 21842
rect 31760 20324 31812 20330
rect 31760 20266 31812 20272
rect 31772 19514 31800 20266
rect 31760 19508 31812 19514
rect 31760 19450 31812 19456
rect 31760 19372 31812 19378
rect 31760 19314 31812 19320
rect 31772 18630 31800 19314
rect 31760 18624 31812 18630
rect 31760 18566 31812 18572
rect 31772 17746 31800 18566
rect 31760 17740 31812 17746
rect 31760 17682 31812 17688
rect 31496 16646 31708 16674
rect 31496 16522 31524 16646
rect 31484 16516 31536 16522
rect 31484 16458 31536 16464
rect 31668 16516 31720 16522
rect 31668 16458 31720 16464
rect 31576 16108 31628 16114
rect 31576 16050 31628 16056
rect 31484 16040 31536 16046
rect 31484 15982 31536 15988
rect 31496 15502 31524 15982
rect 31484 15496 31536 15502
rect 31484 15438 31536 15444
rect 31588 15026 31616 16050
rect 31680 15026 31708 16458
rect 31760 15904 31812 15910
rect 31760 15846 31812 15852
rect 31772 15502 31800 15846
rect 31760 15496 31812 15502
rect 31760 15438 31812 15444
rect 31576 15020 31628 15026
rect 31576 14962 31628 14968
rect 31668 15020 31720 15026
rect 31668 14962 31720 14968
rect 31484 14408 31536 14414
rect 31484 14350 31536 14356
rect 31312 12406 31432 12434
rect 31300 11620 31352 11626
rect 31300 11562 31352 11568
rect 31312 11082 31340 11562
rect 31300 11076 31352 11082
rect 31300 11018 31352 11024
rect 31208 7540 31260 7546
rect 31208 7482 31260 7488
rect 31300 3936 31352 3942
rect 31300 3878 31352 3884
rect 31312 3602 31340 3878
rect 31300 3596 31352 3602
rect 31300 3538 31352 3544
rect 30668 2746 30972 2774
rect 30668 2038 30696 2746
rect 30932 2508 30984 2514
rect 30932 2450 30984 2456
rect 30656 2032 30708 2038
rect 30656 1974 30708 1980
rect 30944 800 30972 2450
rect 31404 2310 31432 12406
rect 31496 9586 31524 14350
rect 31588 13938 31616 14962
rect 31576 13932 31628 13938
rect 31576 13874 31628 13880
rect 31588 12170 31616 13874
rect 31680 13190 31708 14962
rect 31864 14074 31892 21814
rect 32140 21554 32168 21966
rect 32128 21548 32180 21554
rect 32128 21490 32180 21496
rect 32128 20936 32180 20942
rect 32128 20878 32180 20884
rect 32140 19378 32168 20878
rect 32600 20806 32628 21966
rect 32772 21344 32824 21350
rect 32772 21286 32824 21292
rect 32784 20942 32812 21286
rect 32772 20936 32824 20942
rect 32772 20878 32824 20884
rect 32220 20800 32272 20806
rect 32220 20742 32272 20748
rect 32588 20800 32640 20806
rect 32588 20742 32640 20748
rect 32232 20466 32260 20742
rect 32864 20596 32916 20602
rect 32864 20538 32916 20544
rect 32220 20460 32272 20466
rect 32220 20402 32272 20408
rect 32588 20460 32640 20466
rect 32588 20402 32640 20408
rect 32312 19916 32364 19922
rect 32312 19858 32364 19864
rect 32324 19514 32352 19858
rect 32600 19514 32628 20402
rect 32876 19786 32904 20538
rect 32864 19780 32916 19786
rect 32864 19722 32916 19728
rect 32680 19712 32732 19718
rect 32680 19654 32732 19660
rect 32312 19508 32364 19514
rect 32312 19450 32364 19456
rect 32588 19508 32640 19514
rect 32588 19450 32640 19456
rect 32128 19372 32180 19378
rect 32128 19314 32180 19320
rect 31944 16448 31996 16454
rect 31944 16390 31996 16396
rect 31956 16182 31984 16390
rect 31944 16176 31996 16182
rect 31944 16118 31996 16124
rect 32140 16114 32168 19314
rect 32128 16108 32180 16114
rect 32128 16050 32180 16056
rect 32220 16108 32272 16114
rect 32220 16050 32272 16056
rect 32232 15162 32260 16050
rect 32220 15156 32272 15162
rect 32220 15098 32272 15104
rect 32404 14272 32456 14278
rect 32404 14214 32456 14220
rect 31852 14068 31904 14074
rect 31852 14010 31904 14016
rect 32416 14006 32444 14214
rect 32404 14000 32456 14006
rect 32404 13942 32456 13948
rect 32036 13864 32088 13870
rect 32036 13806 32088 13812
rect 32220 13864 32272 13870
rect 32220 13806 32272 13812
rect 31668 13184 31720 13190
rect 31668 13126 31720 13132
rect 31680 12918 31708 13126
rect 32048 12986 32076 13806
rect 32232 13530 32260 13806
rect 32220 13524 32272 13530
rect 32220 13466 32272 13472
rect 32036 12980 32088 12986
rect 32036 12922 32088 12928
rect 32232 12918 32260 13466
rect 31668 12912 31720 12918
rect 31668 12854 31720 12860
rect 32220 12912 32272 12918
rect 32220 12854 32272 12860
rect 31852 12232 31904 12238
rect 31852 12174 31904 12180
rect 31576 12164 31628 12170
rect 31576 12106 31628 12112
rect 31864 11898 31892 12174
rect 31852 11892 31904 11898
rect 31852 11834 31904 11840
rect 31484 9580 31536 9586
rect 31484 9522 31536 9528
rect 32600 5166 32628 19450
rect 32692 19446 32720 19654
rect 32680 19440 32732 19446
rect 32680 19382 32732 19388
rect 32864 18216 32916 18222
rect 32864 18158 32916 18164
rect 32876 16590 32904 18158
rect 32864 16584 32916 16590
rect 32864 16526 32916 16532
rect 32876 15638 32904 16526
rect 32864 15632 32916 15638
rect 32864 15574 32916 15580
rect 32588 5160 32640 5166
rect 32588 5102 32640 5108
rect 32968 4826 32996 22066
rect 33520 22030 33548 22442
rect 33508 22024 33560 22030
rect 33508 21966 33560 21972
rect 33324 21956 33376 21962
rect 33324 21898 33376 21904
rect 33336 21690 33364 21898
rect 33324 21684 33376 21690
rect 33324 21626 33376 21632
rect 33140 20256 33192 20262
rect 33140 20198 33192 20204
rect 33152 19854 33180 20198
rect 33140 19848 33192 19854
rect 33140 19790 33192 19796
rect 33048 17740 33100 17746
rect 33048 17682 33100 17688
rect 32220 4820 32272 4826
rect 32220 4762 32272 4768
rect 32956 4820 33008 4826
rect 32956 4762 33008 4768
rect 32036 4004 32088 4010
rect 32036 3946 32088 3952
rect 32128 4004 32180 4010
rect 32128 3946 32180 3952
rect 31576 3596 31628 3602
rect 31576 3538 31628 3544
rect 31392 2304 31444 2310
rect 31392 2246 31444 2252
rect 31588 800 31616 3538
rect 32048 2922 32076 3946
rect 32140 3058 32168 3946
rect 32128 3052 32180 3058
rect 32128 2994 32180 3000
rect 32036 2916 32088 2922
rect 32036 2858 32088 2864
rect 32232 800 32260 4762
rect 32312 3936 32364 3942
rect 32312 3878 32364 3884
rect 32324 3126 32352 3878
rect 32312 3120 32364 3126
rect 32312 3062 32364 3068
rect 33060 2854 33088 17682
rect 33508 17536 33560 17542
rect 33508 17478 33560 17484
rect 33520 17270 33548 17478
rect 33508 17264 33560 17270
rect 33508 17206 33560 17212
rect 33612 17134 33640 26846
rect 33690 26823 33746 26832
rect 33508 17128 33560 17134
rect 33508 17070 33560 17076
rect 33600 17128 33652 17134
rect 33600 17070 33652 17076
rect 33520 15910 33548 17070
rect 33508 15904 33560 15910
rect 33508 15846 33560 15852
rect 33520 15094 33548 15846
rect 33508 15088 33560 15094
rect 33508 15030 33560 15036
rect 33508 2984 33560 2990
rect 33508 2926 33560 2932
rect 33048 2848 33100 2854
rect 33048 2790 33100 2796
rect 32864 2440 32916 2446
rect 32864 2382 32916 2388
rect 32876 800 32904 2382
rect 33520 800 33548 2926
rect 33888 2514 33916 32370
rect 34060 32224 34112 32230
rect 34060 32166 34112 32172
rect 34072 31822 34100 32166
rect 34060 31816 34112 31822
rect 34060 31758 34112 31764
rect 33968 29164 34020 29170
rect 33968 29106 34020 29112
rect 33980 27946 34008 29106
rect 34060 28416 34112 28422
rect 34060 28358 34112 28364
rect 33968 27940 34020 27946
rect 33968 27882 34020 27888
rect 34072 27538 34100 28358
rect 34060 27532 34112 27538
rect 34060 27474 34112 27480
rect 34164 22094 34192 41386
rect 34808 35698 34836 48078
rect 35912 47802 35940 48622
rect 36740 48210 36768 51200
rect 36728 48204 36780 48210
rect 36728 48146 36780 48152
rect 35900 47796 35952 47802
rect 35900 47738 35952 47744
rect 34934 47356 35242 47376
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47280 35242 47300
rect 34934 46268 35242 46288
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46192 35242 46212
rect 34934 45180 35242 45200
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45104 35242 45124
rect 34934 44092 35242 44112
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44016 35242 44036
rect 34934 43004 35242 43024
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42928 35242 42948
rect 34934 41916 35242 41936
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41840 35242 41860
rect 34934 40828 35242 40848
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40752 35242 40772
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 35164 38480 35216 38486
rect 35162 38448 35164 38457
rect 35216 38448 35218 38457
rect 35162 38383 35218 38392
rect 35624 37664 35676 37670
rect 35624 37606 35676 37612
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 34796 35692 34848 35698
rect 34796 35634 34848 35640
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 34244 34944 34296 34950
rect 34244 34886 34296 34892
rect 34256 31686 34284 34886
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 34244 31680 34296 31686
rect 34244 31622 34296 31628
rect 34256 26926 34284 31622
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 35348 30728 35400 30734
rect 35348 30670 35400 30676
rect 34520 30660 34572 30666
rect 34520 30602 34572 30608
rect 34532 30054 34560 30602
rect 34612 30252 34664 30258
rect 34612 30194 34664 30200
rect 34520 30048 34572 30054
rect 34520 29990 34572 29996
rect 34624 29866 34652 30194
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 34532 29838 34652 29866
rect 34532 28558 34560 29838
rect 34794 29744 34850 29753
rect 34794 29679 34796 29688
rect 34848 29679 34850 29688
rect 34796 29650 34848 29656
rect 35072 29640 35124 29646
rect 35072 29582 35124 29588
rect 34796 29504 34848 29510
rect 34796 29446 34848 29452
rect 34702 29336 34758 29345
rect 34702 29271 34704 29280
rect 34756 29271 34758 29280
rect 34704 29242 34756 29248
rect 34808 29170 34836 29446
rect 34704 29164 34756 29170
rect 34704 29106 34756 29112
rect 34796 29164 34848 29170
rect 34796 29106 34848 29112
rect 34716 28626 34744 29106
rect 35084 28994 35112 29582
rect 35256 29164 35308 29170
rect 35256 29106 35308 29112
rect 35268 29050 35296 29106
rect 35360 29050 35388 30670
rect 35530 29744 35586 29753
rect 35530 29679 35532 29688
rect 35584 29679 35586 29688
rect 35532 29650 35584 29656
rect 35636 29578 35664 37606
rect 37660 34066 37688 51326
rect 38014 51326 38240 51354
rect 38014 51200 38070 51326
rect 38212 49230 38240 51326
rect 38658 51200 38714 52000
rect 39302 51354 39358 52000
rect 38764 51326 39358 51354
rect 38200 49224 38252 49230
rect 38200 49166 38252 49172
rect 38016 49088 38068 49094
rect 38016 49030 38068 49036
rect 37648 34060 37700 34066
rect 37648 34002 37700 34008
rect 35992 33924 36044 33930
rect 35992 33866 36044 33872
rect 36004 33658 36032 33866
rect 35992 33652 36044 33658
rect 35992 33594 36044 33600
rect 35900 33516 35952 33522
rect 35900 33458 35952 33464
rect 35912 31346 35940 33458
rect 35992 31816 36044 31822
rect 35992 31758 36044 31764
rect 35900 31340 35952 31346
rect 35900 31282 35952 31288
rect 35808 30116 35860 30122
rect 35808 30058 35860 30064
rect 35820 29782 35848 30058
rect 35808 29776 35860 29782
rect 35808 29718 35860 29724
rect 35716 29640 35768 29646
rect 35716 29582 35768 29588
rect 35624 29572 35676 29578
rect 35624 29514 35676 29520
rect 35440 29504 35492 29510
rect 35440 29446 35492 29452
rect 35268 29022 35388 29050
rect 34808 28966 35112 28994
rect 34704 28620 34756 28626
rect 34704 28562 34756 28568
rect 34520 28552 34572 28558
rect 34520 28494 34572 28500
rect 34532 27538 34560 28494
rect 34520 27532 34572 27538
rect 34520 27474 34572 27480
rect 34336 26988 34388 26994
rect 34336 26930 34388 26936
rect 34244 26920 34296 26926
rect 34244 26862 34296 26868
rect 34348 26586 34376 26930
rect 34336 26580 34388 26586
rect 34336 26522 34388 26528
rect 34532 26466 34560 27474
rect 34716 27334 34744 28562
rect 34808 28082 34836 28966
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 34796 28076 34848 28082
rect 34796 28018 34848 28024
rect 34808 27606 34836 28018
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 34796 27600 34848 27606
rect 34796 27542 34848 27548
rect 35072 27600 35124 27606
rect 35072 27542 35124 27548
rect 34704 27328 34756 27334
rect 34704 27270 34756 27276
rect 34716 27130 34744 27270
rect 34704 27124 34756 27130
rect 34704 27066 34756 27072
rect 35084 26994 35112 27542
rect 35360 27470 35388 29022
rect 35452 28082 35480 29446
rect 35728 29345 35756 29582
rect 35714 29336 35770 29345
rect 35714 29271 35770 29280
rect 35912 28558 35940 31282
rect 36004 30938 36032 31758
rect 36176 31748 36228 31754
rect 36176 31690 36228 31696
rect 36188 31482 36216 31690
rect 36176 31476 36228 31482
rect 36176 31418 36228 31424
rect 35992 30932 36044 30938
rect 35992 30874 36044 30880
rect 36004 30326 36032 30874
rect 35992 30320 36044 30326
rect 35992 30262 36044 30268
rect 36636 29300 36688 29306
rect 36636 29242 36688 29248
rect 36648 28626 36676 29242
rect 36636 28620 36688 28626
rect 36636 28562 36688 28568
rect 35900 28552 35952 28558
rect 35900 28494 35952 28500
rect 35440 28076 35492 28082
rect 35440 28018 35492 28024
rect 35624 28076 35676 28082
rect 35624 28018 35676 28024
rect 35452 27614 35480 28018
rect 35636 27674 35664 28018
rect 35912 27946 35940 28494
rect 35900 27940 35952 27946
rect 35900 27882 35952 27888
rect 35992 27872 36044 27878
rect 35992 27814 36044 27820
rect 35624 27668 35676 27674
rect 35452 27586 35572 27614
rect 35624 27610 35676 27616
rect 35348 27464 35400 27470
rect 35348 27406 35400 27412
rect 35072 26988 35124 26994
rect 35072 26930 35124 26936
rect 34612 26784 34664 26790
rect 34612 26726 34664 26732
rect 34348 26438 34560 26466
rect 34348 26314 34376 26438
rect 34520 26376 34572 26382
rect 34520 26318 34572 26324
rect 34336 26308 34388 26314
rect 34336 26250 34388 26256
rect 34532 26042 34560 26318
rect 34520 26036 34572 26042
rect 34520 25978 34572 25984
rect 34624 25974 34652 26726
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 35360 26382 35388 27406
rect 35544 26858 35572 27586
rect 36004 27470 36032 27814
rect 35992 27464 36044 27470
rect 35992 27406 36044 27412
rect 36084 27124 36136 27130
rect 36084 27066 36136 27072
rect 36096 26994 36124 27066
rect 35992 26988 36044 26994
rect 35992 26930 36044 26936
rect 36084 26988 36136 26994
rect 36084 26930 36136 26936
rect 35532 26852 35584 26858
rect 35532 26794 35584 26800
rect 35440 26784 35492 26790
rect 35440 26726 35492 26732
rect 35452 26382 35480 26726
rect 36004 26586 36032 26930
rect 35992 26580 36044 26586
rect 35992 26522 36044 26528
rect 37280 26512 37332 26518
rect 37280 26454 37332 26460
rect 35348 26376 35400 26382
rect 35348 26318 35400 26324
rect 35440 26376 35492 26382
rect 35440 26318 35492 26324
rect 35256 26308 35308 26314
rect 35256 26250 35308 26256
rect 35268 26042 35296 26250
rect 36544 26240 36596 26246
rect 36544 26182 36596 26188
rect 36556 26042 36584 26182
rect 35256 26036 35308 26042
rect 35256 25978 35308 25984
rect 35624 26036 35676 26042
rect 35624 25978 35676 25984
rect 36544 26036 36596 26042
rect 36544 25978 36596 25984
rect 34612 25968 34664 25974
rect 34612 25910 34664 25916
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 35636 24750 35664 25978
rect 36544 25696 36596 25702
rect 36544 25638 36596 25644
rect 36556 25430 36584 25638
rect 36544 25424 36596 25430
rect 36544 25366 36596 25372
rect 36544 24812 36596 24818
rect 36544 24754 36596 24760
rect 34796 24744 34848 24750
rect 34796 24686 34848 24692
rect 35440 24744 35492 24750
rect 35440 24686 35492 24692
rect 35624 24744 35676 24750
rect 35624 24686 35676 24692
rect 34808 24410 34836 24686
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 34796 24404 34848 24410
rect 34796 24346 34848 24352
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 34164 22066 34376 22094
rect 34244 20936 34296 20942
rect 34244 20878 34296 20884
rect 34256 20466 34284 20878
rect 34244 20460 34296 20466
rect 34244 20402 34296 20408
rect 34256 17678 34284 20402
rect 34348 18290 34376 22066
rect 34796 21888 34848 21894
rect 34796 21830 34848 21836
rect 34520 21480 34572 21486
rect 34520 21422 34572 21428
rect 34704 21480 34756 21486
rect 34704 21422 34756 21428
rect 34532 20874 34560 21422
rect 34520 20868 34572 20874
rect 34520 20810 34572 20816
rect 34716 20602 34744 21422
rect 34808 21146 34836 21830
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 34796 21140 34848 21146
rect 34796 21082 34848 21088
rect 34704 20596 34756 20602
rect 34704 20538 34756 20544
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 34336 18284 34388 18290
rect 34336 18226 34388 18232
rect 34428 18216 34480 18222
rect 34428 18158 34480 18164
rect 34440 17882 34468 18158
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 34428 17876 34480 17882
rect 34428 17818 34480 17824
rect 34244 17672 34296 17678
rect 34244 17614 34296 17620
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 34520 5636 34572 5642
rect 34520 5578 34572 5584
rect 33876 2508 33928 2514
rect 33876 2450 33928 2456
rect 34152 2372 34204 2378
rect 34152 2314 34204 2320
rect 34060 2304 34112 2310
rect 34060 2246 34112 2252
rect 34072 2106 34100 2246
rect 34060 2100 34112 2106
rect 34060 2042 34112 2048
rect 34164 800 34192 2314
rect 34532 2310 34560 5578
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 35452 4078 35480 24686
rect 36556 24614 36584 24754
rect 36544 24608 36596 24614
rect 36544 24550 36596 24556
rect 37292 24274 37320 26454
rect 37372 26376 37424 26382
rect 37372 26318 37424 26324
rect 37384 24614 37412 26318
rect 38028 25294 38056 49030
rect 38476 28484 38528 28490
rect 38476 28426 38528 28432
rect 38108 27600 38160 27606
rect 38108 27542 38160 27548
rect 38120 25906 38148 27542
rect 38292 26240 38344 26246
rect 38292 26182 38344 26188
rect 38304 25974 38332 26182
rect 38292 25968 38344 25974
rect 38292 25910 38344 25916
rect 38108 25900 38160 25906
rect 38108 25842 38160 25848
rect 38108 25492 38160 25498
rect 38108 25434 38160 25440
rect 38016 25288 38068 25294
rect 38016 25230 38068 25236
rect 37372 24608 37424 24614
rect 37372 24550 37424 24556
rect 37280 24268 37332 24274
rect 37280 24210 37332 24216
rect 37384 23730 37412 24550
rect 37464 24132 37516 24138
rect 37464 24074 37516 24080
rect 37476 23866 37504 24074
rect 37464 23860 37516 23866
rect 37464 23802 37516 23808
rect 37372 23724 37424 23730
rect 37372 23666 37424 23672
rect 36544 16448 36596 16454
rect 36544 16390 36596 16396
rect 36556 16250 36584 16390
rect 36544 16244 36596 16250
rect 36544 16186 36596 16192
rect 37464 11688 37516 11694
rect 37464 11630 37516 11636
rect 37280 11620 37332 11626
rect 37280 11562 37332 11568
rect 37292 11150 37320 11562
rect 37476 11354 37504 11630
rect 37464 11348 37516 11354
rect 37464 11290 37516 11296
rect 37280 11144 37332 11150
rect 37280 11086 37332 11092
rect 37292 7970 37320 11086
rect 37292 7942 37412 7970
rect 37280 7880 37332 7886
rect 37280 7822 37332 7828
rect 35900 7812 35952 7818
rect 35900 7754 35952 7760
rect 35440 4072 35492 4078
rect 35440 4014 35492 4020
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 35912 2514 35940 7754
rect 37292 7410 37320 7822
rect 37280 7404 37332 7410
rect 37280 7346 37332 7352
rect 37384 7274 37412 7942
rect 38016 7336 38068 7342
rect 38016 7278 38068 7284
rect 37372 7268 37424 7274
rect 37372 7210 37424 7216
rect 37384 4706 37412 7210
rect 37384 4678 37504 4706
rect 37476 4078 37504 4678
rect 37924 4140 37976 4146
rect 37924 4082 37976 4088
rect 37372 4072 37424 4078
rect 37372 4014 37424 4020
rect 37464 4072 37516 4078
rect 37464 4014 37516 4020
rect 36176 4004 36228 4010
rect 36176 3946 36228 3952
rect 36188 3670 36216 3946
rect 36544 3936 36596 3942
rect 36544 3878 36596 3884
rect 36176 3664 36228 3670
rect 36176 3606 36228 3612
rect 36556 3602 36584 3878
rect 36544 3596 36596 3602
rect 36544 3538 36596 3544
rect 36728 3596 36780 3602
rect 36728 3538 36780 3544
rect 36360 3528 36412 3534
rect 36360 3470 36412 3476
rect 36372 3058 36400 3470
rect 36360 3052 36412 3058
rect 36360 2994 36412 3000
rect 35900 2508 35952 2514
rect 35900 2450 35952 2456
rect 34796 2440 34848 2446
rect 34796 2382 34848 2388
rect 36084 2440 36136 2446
rect 36084 2382 36136 2388
rect 34520 2304 34572 2310
rect 34520 2246 34572 2252
rect 34808 800 34836 2382
rect 36096 800 36124 2382
rect 36740 800 36768 3538
rect 37384 800 37412 4014
rect 37936 2854 37964 4082
rect 37924 2848 37976 2854
rect 37924 2790 37976 2796
rect 38028 800 38056 7278
rect 38120 3602 38148 25434
rect 38292 25288 38344 25294
rect 38292 25230 38344 25236
rect 38304 8838 38332 25230
rect 38488 12442 38516 28426
rect 38568 24608 38620 24614
rect 38568 24550 38620 24556
rect 38476 12436 38528 12442
rect 38476 12378 38528 12384
rect 38580 9654 38608 24550
rect 38672 24070 38700 51200
rect 38764 38554 38792 51326
rect 39302 51200 39358 51326
rect 39946 51200 40002 52000
rect 40590 51354 40646 52000
rect 41234 51354 41290 52000
rect 41878 51354 41934 52000
rect 40590 51326 40724 51354
rect 40590 51200 40646 51326
rect 39304 49224 39356 49230
rect 39304 49166 39356 49172
rect 38752 38548 38804 38554
rect 38752 38490 38804 38496
rect 39316 38486 39344 49166
rect 39672 48884 39724 48890
rect 39672 48826 39724 48832
rect 39684 48346 39712 48826
rect 39764 48680 39816 48686
rect 39960 48668 39988 51200
rect 40696 49298 40724 51326
rect 40880 51326 41290 51354
rect 40684 49292 40736 49298
rect 40684 49234 40736 49240
rect 40040 48680 40092 48686
rect 39960 48640 40040 48668
rect 39764 48622 39816 48628
rect 40040 48622 40092 48628
rect 39776 48346 39804 48622
rect 39672 48340 39724 48346
rect 39672 48282 39724 48288
rect 39764 48340 39816 48346
rect 39764 48282 39816 48288
rect 40684 47524 40736 47530
rect 40684 47466 40736 47472
rect 40696 47258 40724 47466
rect 40684 47252 40736 47258
rect 40684 47194 40736 47200
rect 39856 47116 39908 47122
rect 39856 47058 39908 47064
rect 39304 38480 39356 38486
rect 39304 38422 39356 38428
rect 38936 38276 38988 38282
rect 38936 38218 38988 38224
rect 38948 26586 38976 38218
rect 38936 26580 38988 26586
rect 38936 26522 38988 26528
rect 39120 24812 39172 24818
rect 39120 24754 39172 24760
rect 39132 24614 39160 24754
rect 39120 24608 39172 24614
rect 39120 24550 39172 24556
rect 39120 24132 39172 24138
rect 39120 24074 39172 24080
rect 38660 24064 38712 24070
rect 38660 24006 38712 24012
rect 38568 9648 38620 9654
rect 38568 9590 38620 9596
rect 38292 8832 38344 8838
rect 38292 8774 38344 8780
rect 39132 5574 39160 24074
rect 39120 5568 39172 5574
rect 39120 5510 39172 5516
rect 38752 4072 38804 4078
rect 38752 4014 38804 4020
rect 39764 4072 39816 4078
rect 39764 4014 39816 4020
rect 38764 3738 38792 4014
rect 38752 3732 38804 3738
rect 38752 3674 38804 3680
rect 38844 3664 38896 3670
rect 38844 3606 38896 3612
rect 38108 3596 38160 3602
rect 38108 3538 38160 3544
rect 38856 3534 38884 3606
rect 39028 3596 39080 3602
rect 39028 3538 39080 3544
rect 38844 3528 38896 3534
rect 38844 3470 38896 3476
rect 39040 3369 39068 3538
rect 39026 3360 39082 3369
rect 39026 3295 39082 3304
rect 38660 2440 38712 2446
rect 38660 2382 38712 2388
rect 38672 800 38700 2382
rect 39776 2122 39804 4014
rect 39868 3534 39896 47058
rect 40880 45554 40908 51326
rect 41234 51200 41290 51326
rect 41800 51326 41934 51354
rect 41800 48142 41828 51326
rect 41878 51200 41934 51326
rect 42522 51354 42578 52000
rect 42522 51326 42748 51354
rect 42522 51200 42578 51326
rect 42340 49224 42392 49230
rect 42340 49166 42392 49172
rect 41052 48136 41104 48142
rect 41052 48078 41104 48084
rect 41788 48136 41840 48142
rect 41788 48078 41840 48084
rect 40052 45526 40908 45554
rect 40052 23662 40080 45526
rect 41064 34746 41092 48078
rect 42064 48068 42116 48074
rect 42064 48010 42116 48016
rect 41880 48000 41932 48006
rect 41880 47942 41932 47948
rect 41696 47660 41748 47666
rect 41696 47602 41748 47608
rect 41708 47190 41736 47602
rect 41696 47184 41748 47190
rect 41696 47126 41748 47132
rect 41052 34740 41104 34746
rect 41052 34682 41104 34688
rect 40040 23656 40092 23662
rect 40040 23598 40092 23604
rect 41892 22778 41920 47942
rect 42076 47802 42104 48010
rect 42064 47796 42116 47802
rect 42064 47738 42116 47744
rect 42352 45490 42380 49166
rect 42720 48770 42748 51326
rect 43166 51200 43222 52000
rect 43810 51354 43866 52000
rect 44454 51354 44510 52000
rect 43810 51326 43944 51354
rect 43810 51200 43866 51326
rect 42720 48742 42840 48770
rect 42812 48686 42840 48742
rect 42432 48680 42484 48686
rect 42432 48622 42484 48628
rect 42616 48680 42668 48686
rect 42616 48622 42668 48628
rect 42800 48680 42852 48686
rect 42800 48622 42852 48628
rect 42444 47258 42472 48622
rect 42628 48278 42656 48622
rect 42616 48272 42668 48278
rect 42616 48214 42668 48220
rect 43180 48210 43208 51200
rect 42524 48204 42576 48210
rect 42524 48146 42576 48152
rect 42800 48204 42852 48210
rect 42800 48146 42852 48152
rect 43168 48204 43220 48210
rect 43168 48146 43220 48152
rect 42536 47802 42564 48146
rect 42524 47796 42576 47802
rect 42524 47738 42576 47744
rect 42432 47252 42484 47258
rect 42432 47194 42484 47200
rect 42812 46578 42840 48146
rect 43444 47592 43496 47598
rect 43444 47534 43496 47540
rect 43456 47258 43484 47534
rect 43444 47252 43496 47258
rect 43444 47194 43496 47200
rect 43916 47054 43944 51326
rect 44454 51326 44772 51354
rect 44454 51200 44510 51326
rect 44088 49224 44140 49230
rect 44088 49166 44140 49172
rect 43996 47184 44048 47190
rect 43996 47126 44048 47132
rect 43904 47048 43956 47054
rect 43904 46990 43956 46996
rect 42800 46572 42852 46578
rect 42800 46514 42852 46520
rect 42340 45484 42392 45490
rect 42340 45426 42392 45432
rect 44008 24342 44036 47126
rect 44100 46578 44128 49166
rect 44640 49156 44692 49162
rect 44640 49098 44692 49104
rect 44180 48000 44232 48006
rect 44180 47942 44232 47948
rect 44088 46572 44140 46578
rect 44088 46514 44140 46520
rect 44192 45966 44220 47942
rect 44548 47456 44600 47462
rect 44548 47398 44600 47404
rect 44560 46578 44588 47398
rect 44652 46714 44680 49098
rect 44744 48142 44772 51326
rect 45098 51200 45154 52000
rect 45742 51200 45798 52000
rect 46386 51200 46442 52000
rect 46662 51776 46718 51785
rect 46662 51711 46718 51720
rect 44732 48136 44784 48142
rect 45112 48124 45140 51200
rect 45756 48686 45784 51200
rect 46570 51096 46626 51105
rect 46570 51031 46626 51040
rect 46204 49360 46256 49366
rect 46204 49302 46256 49308
rect 45376 48680 45428 48686
rect 45376 48622 45428 48628
rect 45744 48680 45796 48686
rect 45744 48622 45796 48628
rect 45112 48096 45324 48124
rect 44732 48078 44784 48084
rect 45100 48000 45152 48006
rect 45100 47942 45152 47948
rect 45008 47048 45060 47054
rect 45008 46990 45060 46996
rect 44640 46708 44692 46714
rect 44640 46650 44692 46656
rect 44548 46572 44600 46578
rect 44548 46514 44600 46520
rect 44180 45960 44232 45966
rect 44180 45902 44232 45908
rect 44560 40050 44588 46514
rect 45020 46170 45048 46990
rect 45008 46164 45060 46170
rect 45008 46106 45060 46112
rect 44548 40044 44600 40050
rect 44548 39986 44600 39992
rect 45112 35894 45140 47942
rect 45192 47456 45244 47462
rect 45192 47398 45244 47404
rect 45204 47122 45232 47398
rect 45296 47122 45324 48096
rect 45192 47116 45244 47122
rect 45192 47058 45244 47064
rect 45284 47116 45336 47122
rect 45284 47058 45336 47064
rect 45388 46170 45416 48622
rect 45468 48612 45520 48618
rect 45468 48554 45520 48560
rect 45376 46164 45428 46170
rect 45376 46106 45428 46112
rect 45480 45490 45508 48554
rect 46216 47802 46244 49302
rect 46296 48136 46348 48142
rect 46296 48078 46348 48084
rect 46204 47796 46256 47802
rect 46204 47738 46256 47744
rect 46020 47592 46072 47598
rect 46020 47534 46072 47540
rect 45928 45960 45980 45966
rect 45928 45902 45980 45908
rect 45468 45484 45520 45490
rect 45468 45426 45520 45432
rect 45192 44872 45244 44878
rect 45192 44814 45244 44820
rect 45204 44402 45232 44814
rect 45192 44396 45244 44402
rect 45192 44338 45244 44344
rect 45744 41132 45796 41138
rect 45744 41074 45796 41080
rect 45112 35866 45232 35894
rect 45204 25702 45232 35866
rect 45466 26616 45522 26625
rect 45466 26551 45522 26560
rect 45192 25696 45244 25702
rect 45192 25638 45244 25644
rect 43996 24336 44048 24342
rect 43996 24278 44048 24284
rect 41880 22772 41932 22778
rect 41880 22714 41932 22720
rect 45480 22030 45508 26551
rect 45756 23186 45784 41074
rect 45836 36848 45888 36854
rect 45836 36790 45888 36796
rect 45744 23180 45796 23186
rect 45744 23122 45796 23128
rect 45468 22024 45520 22030
rect 45468 21966 45520 21972
rect 42800 12708 42852 12714
rect 42800 12650 42852 12656
rect 42812 11830 42840 12650
rect 42800 11824 42852 11830
rect 42800 11766 42852 11772
rect 45652 7404 45704 7410
rect 45652 7346 45704 7352
rect 45008 4616 45060 4622
rect 45008 4558 45060 4564
rect 41696 4140 41748 4146
rect 41696 4082 41748 4088
rect 41512 3936 41564 3942
rect 41512 3878 41564 3884
rect 41524 3602 41552 3878
rect 41708 3738 41736 4082
rect 42432 4072 42484 4078
rect 42708 4072 42760 4078
rect 42432 4014 42484 4020
rect 42536 4032 42708 4060
rect 41696 3732 41748 3738
rect 41696 3674 41748 3680
rect 41512 3596 41564 3602
rect 41512 3538 41564 3544
rect 41880 3596 41932 3602
rect 41880 3538 41932 3544
rect 39856 3528 39908 3534
rect 39856 3470 39908 3476
rect 40132 3392 40184 3398
rect 40132 3334 40184 3340
rect 40144 3126 40172 3334
rect 40132 3120 40184 3126
rect 40132 3062 40184 3068
rect 39948 2984 40000 2990
rect 39948 2926 40000 2932
rect 41144 2984 41196 2990
rect 41144 2926 41196 2932
rect 39960 2514 39988 2926
rect 39948 2508 40000 2514
rect 39948 2450 40000 2456
rect 39776 2094 39988 2122
rect 39960 800 39988 2094
rect 41156 1578 41184 2926
rect 41156 1550 41276 1578
rect 41248 800 41276 1550
rect 41892 800 41920 3538
rect 42444 3058 42472 4014
rect 42432 3052 42484 3058
rect 42432 2994 42484 3000
rect 42536 800 42564 4032
rect 42708 4014 42760 4020
rect 44180 3392 44232 3398
rect 44180 3334 44232 3340
rect 44192 3126 44220 3334
rect 44180 3120 44232 3126
rect 44180 3062 44232 3068
rect 44364 3120 44416 3126
rect 44364 3062 44416 3068
rect 44272 2984 44324 2990
rect 44272 2926 44324 2932
rect 44284 2514 44312 2926
rect 44376 2854 44404 3062
rect 44456 2984 44508 2990
rect 44456 2926 44508 2932
rect 44364 2848 44416 2854
rect 44364 2790 44416 2796
rect 44272 2508 44324 2514
rect 44272 2450 44324 2456
rect 43168 2372 43220 2378
rect 43168 2314 43220 2320
rect 43180 800 43208 2314
rect 43444 2304 43496 2310
rect 43444 2246 43496 2252
rect 43456 1970 43484 2246
rect 43444 1964 43496 1970
rect 43444 1906 43496 1912
rect 44468 800 44496 2926
rect 45020 2514 45048 4558
rect 45376 3936 45428 3942
rect 45376 3878 45428 3884
rect 45388 3602 45416 3878
rect 45664 3670 45692 7346
rect 45848 6322 45876 36790
rect 45940 35698 45968 45902
rect 45928 35692 45980 35698
rect 45928 35634 45980 35640
rect 45940 35290 45968 35634
rect 45928 35284 45980 35290
rect 45928 35226 45980 35232
rect 46032 30122 46060 47534
rect 46308 45490 46336 48078
rect 46388 47456 46440 47462
rect 46388 47398 46440 47404
rect 46400 46510 46428 47398
rect 46388 46504 46440 46510
rect 46388 46446 46440 46452
rect 46584 45914 46612 51031
rect 46676 49298 46704 51711
rect 47030 51200 47086 52000
rect 47674 51354 47730 52000
rect 47674 51326 47808 51354
rect 47674 51200 47730 51326
rect 46754 50416 46810 50425
rect 46754 50351 46810 50360
rect 46664 49292 46716 49298
rect 46664 49234 46716 49240
rect 46768 48210 46796 50351
rect 46846 49736 46902 49745
rect 46846 49671 46902 49680
rect 46860 49298 46888 49671
rect 46848 49292 46900 49298
rect 46848 49234 46900 49240
rect 47780 49230 47808 51326
rect 48318 51200 48374 52000
rect 48962 51200 49018 52000
rect 49606 51200 49662 52000
rect 47768 49224 47820 49230
rect 47768 49166 47820 49172
rect 47766 49056 47822 49065
rect 47766 48991 47822 49000
rect 47780 48822 47808 48991
rect 47768 48816 47820 48822
rect 47768 48758 47820 48764
rect 47766 48376 47822 48385
rect 47766 48311 47822 48320
rect 47032 48272 47084 48278
rect 47032 48214 47084 48220
rect 46756 48204 46808 48210
rect 46756 48146 46808 48152
rect 46846 47016 46902 47025
rect 46846 46951 46902 46960
rect 46584 45886 46704 45914
rect 46296 45484 46348 45490
rect 46296 45426 46348 45432
rect 46480 45280 46532 45286
rect 46480 45222 46532 45228
rect 46492 44946 46520 45222
rect 46570 44976 46626 44985
rect 46480 44940 46532 44946
rect 46570 44911 46626 44920
rect 46480 44882 46532 44888
rect 46110 44296 46166 44305
rect 46110 44231 46166 44240
rect 46124 31890 46152 44231
rect 46480 42016 46532 42022
rect 46480 41958 46532 41964
rect 46492 41682 46520 41958
rect 46480 41676 46532 41682
rect 46480 41618 46532 41624
rect 46204 41064 46256 41070
rect 46204 41006 46256 41012
rect 46216 40905 46244 41006
rect 46296 40928 46348 40934
rect 46202 40896 46258 40905
rect 46296 40870 46348 40876
rect 46202 40831 46258 40840
rect 46308 40594 46336 40870
rect 46296 40588 46348 40594
rect 46296 40530 46348 40536
rect 46202 37496 46258 37505
rect 46202 37431 46258 37440
rect 46112 31884 46164 31890
rect 46112 31826 46164 31832
rect 46020 30116 46072 30122
rect 46020 30058 46072 30064
rect 46032 29238 46060 30058
rect 46020 29232 46072 29238
rect 46020 29174 46072 29180
rect 46216 13938 46244 37431
rect 46480 37120 46532 37126
rect 46480 37062 46532 37068
rect 46492 36242 46520 37062
rect 46480 36236 46532 36242
rect 46480 36178 46532 36184
rect 46388 34536 46440 34542
rect 46388 34478 46440 34484
rect 46400 33658 46428 34478
rect 46388 33652 46440 33658
rect 46388 33594 46440 33600
rect 46296 28960 46348 28966
rect 46296 28902 46348 28908
rect 46480 28960 46532 28966
rect 46480 28902 46532 28908
rect 46308 28626 46336 28902
rect 46492 28626 46520 28902
rect 46296 28620 46348 28626
rect 46296 28562 46348 28568
rect 46480 28620 46532 28626
rect 46480 28562 46532 28568
rect 46388 27056 46440 27062
rect 46388 26998 46440 27004
rect 46296 20256 46348 20262
rect 46296 20198 46348 20204
rect 46308 19922 46336 20198
rect 46296 19916 46348 19922
rect 46296 19858 46348 19864
rect 46400 17785 46428 26998
rect 46480 25968 46532 25974
rect 46480 25910 46532 25916
rect 46492 25226 46520 25910
rect 46480 25220 46532 25226
rect 46480 25162 46532 25168
rect 46584 21486 46612 44911
rect 46676 38214 46704 45886
rect 46756 45416 46808 45422
rect 46756 45358 46808 45364
rect 46768 44010 46796 45358
rect 46860 44334 46888 46951
rect 47044 46578 47072 48214
rect 47676 48068 47728 48074
rect 47676 48010 47728 48016
rect 47688 46714 47716 48010
rect 47780 47734 47808 48311
rect 48332 47802 48360 51200
rect 48320 47796 48372 47802
rect 48320 47738 48372 47744
rect 47768 47728 47820 47734
rect 47768 47670 47820 47676
rect 48976 47054 49004 51200
rect 49620 48278 49648 51200
rect 49608 48272 49660 48278
rect 49608 48214 49660 48220
rect 48964 47048 49016 47054
rect 48964 46990 49016 46996
rect 47952 46912 48004 46918
rect 47952 46854 48004 46860
rect 47676 46708 47728 46714
rect 47676 46650 47728 46656
rect 47032 46572 47084 46578
rect 47032 46514 47084 46520
rect 47768 46028 47820 46034
rect 47768 45970 47820 45976
rect 47676 45892 47728 45898
rect 47676 45834 47728 45840
rect 47688 45558 47716 45834
rect 47676 45552 47728 45558
rect 47676 45494 47728 45500
rect 47124 45484 47176 45490
rect 47124 45426 47176 45432
rect 46848 44328 46900 44334
rect 46848 44270 46900 44276
rect 46768 43982 46888 44010
rect 46756 42220 46808 42226
rect 46756 42162 46808 42168
rect 46664 38208 46716 38214
rect 46664 38150 46716 38156
rect 46768 36854 46796 42162
rect 46860 37262 46888 43982
rect 46940 43716 46992 43722
rect 46940 43658 46992 43664
rect 46952 43450 46980 43658
rect 46940 43444 46992 43450
rect 46940 43386 46992 43392
rect 47032 37936 47084 37942
rect 47032 37878 47084 37884
rect 46848 37256 46900 37262
rect 46848 37198 46900 37204
rect 46756 36848 46808 36854
rect 46756 36790 46808 36796
rect 46848 36576 46900 36582
rect 46848 36518 46900 36524
rect 46860 35894 46888 36518
rect 46768 35866 46888 35894
rect 46664 35692 46716 35698
rect 46664 35634 46716 35640
rect 46676 33522 46704 35634
rect 46768 34134 46796 35866
rect 46940 35488 46992 35494
rect 46940 35430 46992 35436
rect 46848 34400 46900 34406
rect 46848 34342 46900 34348
rect 46756 34128 46808 34134
rect 46860 34105 46888 34342
rect 46756 34070 46808 34076
rect 46846 34096 46902 34105
rect 46952 34066 46980 35430
rect 46846 34031 46902 34040
rect 46940 34060 46992 34066
rect 46940 34002 46992 34008
rect 46664 33516 46716 33522
rect 46664 33458 46716 33464
rect 46940 33312 46992 33318
rect 46940 33254 46992 33260
rect 46848 32360 46900 32366
rect 46848 32302 46900 32308
rect 46756 29164 46808 29170
rect 46756 29106 46808 29112
rect 46664 29028 46716 29034
rect 46664 28970 46716 28976
rect 46676 27402 46704 28970
rect 46664 27396 46716 27402
rect 46664 27338 46716 27344
rect 46664 23044 46716 23050
rect 46664 22986 46716 22992
rect 46572 21480 46624 21486
rect 46572 21422 46624 21428
rect 46386 17776 46442 17785
rect 46386 17711 46442 17720
rect 46296 17672 46348 17678
rect 46296 17614 46348 17620
rect 46308 16658 46336 17614
rect 46296 16652 46348 16658
rect 46296 16594 46348 16600
rect 46296 15904 46348 15910
rect 46296 15846 46348 15852
rect 46308 15570 46336 15846
rect 46296 15564 46348 15570
rect 46296 15506 46348 15512
rect 46676 15162 46704 22986
rect 46768 19378 46796 29106
rect 46860 26042 46888 32302
rect 46952 29850 46980 33254
rect 46940 29844 46992 29850
rect 46940 29786 46992 29792
rect 47044 27962 47072 37878
rect 47136 28082 47164 45426
rect 47308 44464 47360 44470
rect 47308 44406 47360 44412
rect 47320 42770 47348 44406
rect 47780 44402 47808 45970
rect 47768 44396 47820 44402
rect 47768 44338 47820 44344
rect 47860 43308 47912 43314
rect 47860 43250 47912 43256
rect 47872 42945 47900 43250
rect 47858 42936 47914 42945
rect 47858 42871 47914 42880
rect 47964 42786 47992 46854
rect 48134 46336 48190 46345
rect 48134 46271 48190 46280
rect 48148 46034 48176 46271
rect 48136 46028 48188 46034
rect 48136 45970 48188 45976
rect 48134 45656 48190 45665
rect 48134 45591 48190 45600
rect 48148 44946 48176 45591
rect 48136 44940 48188 44946
rect 48136 44882 48188 44888
rect 48136 43716 48188 43722
rect 48136 43658 48188 43664
rect 48148 43625 48176 43658
rect 48134 43616 48190 43625
rect 48134 43551 48190 43560
rect 48228 43104 48280 43110
rect 48228 43046 48280 43052
rect 47308 42764 47360 42770
rect 47308 42706 47360 42712
rect 47872 42758 47992 42786
rect 47216 42696 47268 42702
rect 47216 42638 47268 42644
rect 47228 37942 47256 42638
rect 47768 42016 47820 42022
rect 47768 41958 47820 41964
rect 47780 41750 47808 41958
rect 47768 41744 47820 41750
rect 47768 41686 47820 41692
rect 47872 40746 47900 42758
rect 47952 42628 48004 42634
rect 47952 42570 48004 42576
rect 47964 42265 47992 42570
rect 47950 42256 48006 42265
rect 47950 42191 48006 42200
rect 48134 41576 48190 41585
rect 48134 41511 48136 41520
rect 48188 41511 48190 41520
rect 48136 41482 48188 41488
rect 47780 40718 47900 40746
rect 47676 40452 47728 40458
rect 47676 40394 47728 40400
rect 47688 40050 47716 40394
rect 47308 40044 47360 40050
rect 47308 39986 47360 39992
rect 47676 40044 47728 40050
rect 47676 39986 47728 39992
rect 47216 37936 47268 37942
rect 47216 37878 47268 37884
rect 47320 31754 47348 39986
rect 47676 39432 47728 39438
rect 47676 39374 47728 39380
rect 47688 38418 47716 39374
rect 47676 38412 47728 38418
rect 47676 38354 47728 38360
rect 47492 37664 47544 37670
rect 47492 37606 47544 37612
rect 47400 34672 47452 34678
rect 47400 34614 47452 34620
rect 47412 33114 47440 34614
rect 47400 33108 47452 33114
rect 47400 33050 47452 33056
rect 47320 31726 47440 31754
rect 47306 30016 47362 30025
rect 47306 29951 47362 29960
rect 47320 29646 47348 29951
rect 47308 29640 47360 29646
rect 47308 29582 47360 29588
rect 47124 28076 47176 28082
rect 47124 28018 47176 28024
rect 47044 27934 47256 27962
rect 47032 27872 47084 27878
rect 47032 27814 47084 27820
rect 47124 27872 47176 27878
rect 47124 27814 47176 27820
rect 47044 27538 47072 27814
rect 47032 27532 47084 27538
rect 47032 27474 47084 27480
rect 46940 27328 46992 27334
rect 46940 27270 46992 27276
rect 46848 26036 46900 26042
rect 46848 25978 46900 25984
rect 46860 25906 46888 25978
rect 46848 25900 46900 25906
rect 46848 25842 46900 25848
rect 46952 24274 46980 27270
rect 46940 24268 46992 24274
rect 46940 24210 46992 24216
rect 46940 19780 46992 19786
rect 46940 19722 46992 19728
rect 46952 19514 46980 19722
rect 46940 19508 46992 19514
rect 46940 19450 46992 19456
rect 46756 19372 46808 19378
rect 46756 19314 46808 19320
rect 46768 15978 46796 19314
rect 46756 15972 46808 15978
rect 46756 15914 46808 15920
rect 46664 15156 46716 15162
rect 46664 15098 46716 15104
rect 46846 15056 46902 15065
rect 46846 14991 46848 15000
rect 46900 14991 46902 15000
rect 46848 14962 46900 14968
rect 46480 14816 46532 14822
rect 46480 14758 46532 14764
rect 46492 14482 46520 14758
rect 46480 14476 46532 14482
rect 46480 14418 46532 14424
rect 46204 13932 46256 13938
rect 46204 13874 46256 13880
rect 46846 13016 46902 13025
rect 46846 12951 46902 12960
rect 46860 12714 46888 12951
rect 46848 12708 46900 12714
rect 46848 12650 46900 12656
rect 46848 12436 46900 12442
rect 46848 12378 46900 12384
rect 46860 12345 46888 12378
rect 46846 12336 46902 12345
rect 46846 12271 46902 12280
rect 47136 11150 47164 27814
rect 47228 16574 47256 27934
rect 47308 24200 47360 24206
rect 47308 24142 47360 24148
rect 47320 23905 47348 24142
rect 47306 23896 47362 23905
rect 47306 23831 47362 23840
rect 47412 17202 47440 31726
rect 47504 28626 47532 37606
rect 47584 35488 47636 35494
rect 47584 35430 47636 35436
rect 47492 28620 47544 28626
rect 47492 28562 47544 28568
rect 47596 28506 47624 35430
rect 47676 35012 47728 35018
rect 47676 34954 47728 34960
rect 47688 34746 47716 34954
rect 47676 34740 47728 34746
rect 47676 34682 47728 34688
rect 47676 32428 47728 32434
rect 47676 32370 47728 32376
rect 47688 32065 47716 32370
rect 47674 32056 47730 32065
rect 47674 31991 47730 32000
rect 47676 28620 47728 28626
rect 47676 28562 47728 28568
rect 47504 28478 47624 28506
rect 47504 24954 47532 28478
rect 47584 28416 47636 28422
rect 47584 28358 47636 28364
rect 47492 24948 47544 24954
rect 47492 24890 47544 24896
rect 47492 23112 47544 23118
rect 47492 23054 47544 23060
rect 47504 22778 47532 23054
rect 47492 22772 47544 22778
rect 47492 22714 47544 22720
rect 47596 22094 47624 28358
rect 47688 23526 47716 28562
rect 47780 27554 47808 40718
rect 48136 40452 48188 40458
rect 48136 40394 48188 40400
rect 48148 40225 48176 40394
rect 48134 40216 48190 40225
rect 48134 40151 48190 40160
rect 48134 39536 48190 39545
rect 48134 39471 48190 39480
rect 47952 38956 48004 38962
rect 47952 38898 48004 38904
rect 47964 38865 47992 38898
rect 47950 38856 48006 38865
rect 47950 38791 48006 38800
rect 48148 38418 48176 39471
rect 48136 38412 48188 38418
rect 48136 38354 48188 38360
rect 47858 38176 47914 38185
rect 47858 38111 47914 38120
rect 47872 37874 47900 38111
rect 47860 37868 47912 37874
rect 47860 37810 47912 37816
rect 47952 37256 48004 37262
rect 47952 37198 48004 37204
rect 47964 36310 47992 37198
rect 48134 36816 48190 36825
rect 48134 36751 48190 36760
rect 47952 36304 48004 36310
rect 47952 36246 48004 36252
rect 48148 36242 48176 36751
rect 48136 36236 48188 36242
rect 48136 36178 48188 36184
rect 47858 36136 47914 36145
rect 47858 36071 47914 36080
rect 47872 35698 47900 36071
rect 48240 35894 48268 43046
rect 48056 35866 48268 35894
rect 47860 35692 47912 35698
rect 47860 35634 47912 35640
rect 47860 34604 47912 34610
rect 47860 34546 47912 34552
rect 47872 28422 47900 34546
rect 47952 33516 48004 33522
rect 47952 33458 48004 33464
rect 47964 33425 47992 33458
rect 47950 33416 48006 33425
rect 47950 33351 48006 33360
rect 47952 31816 48004 31822
rect 47952 31758 48004 31764
rect 48056 31770 48084 35866
rect 48226 35456 48282 35465
rect 48226 35391 48282 35400
rect 48136 35012 48188 35018
rect 48136 34954 48188 34960
rect 48148 34785 48176 34954
rect 48134 34776 48190 34785
rect 48134 34711 48190 34720
rect 48240 34066 48268 35391
rect 48228 34060 48280 34066
rect 48228 34002 48280 34008
rect 47964 31385 47992 31758
rect 48056 31742 48176 31770
rect 48044 31680 48096 31686
rect 48044 31622 48096 31628
rect 48056 31414 48084 31622
rect 48044 31408 48096 31414
rect 47950 31376 48006 31385
rect 48044 31350 48096 31356
rect 47950 31311 48006 31320
rect 48148 29458 48176 31742
rect 48056 29430 48176 29458
rect 47860 28416 47912 28422
rect 47860 28358 47912 28364
rect 47860 28076 47912 28082
rect 47860 28018 47912 28024
rect 47872 27985 47900 28018
rect 47858 27976 47914 27985
rect 47858 27911 47914 27920
rect 47780 27526 47900 27554
rect 47768 25696 47820 25702
rect 47768 25638 47820 25644
rect 47780 25362 47808 25638
rect 47768 25356 47820 25362
rect 47768 25298 47820 25304
rect 47676 23520 47728 23526
rect 47676 23462 47728 23468
rect 47872 23322 47900 27526
rect 48056 26466 48084 29430
rect 48134 29336 48190 29345
rect 48134 29271 48190 29280
rect 48148 28626 48176 29271
rect 48226 28656 48282 28665
rect 48136 28620 48188 28626
rect 48226 28591 48282 28600
rect 48136 28562 48188 28568
rect 48240 27538 48268 28591
rect 48228 27532 48280 27538
rect 48228 27474 48280 27480
rect 48056 26438 48268 26466
rect 47952 26308 48004 26314
rect 47952 26250 48004 26256
rect 48044 26308 48096 26314
rect 48044 26250 48096 26256
rect 47964 25945 47992 26250
rect 47950 25936 48006 25945
rect 47950 25871 48006 25880
rect 47950 25256 48006 25265
rect 47950 25191 48006 25200
rect 47964 24818 47992 25191
rect 47952 24812 48004 24818
rect 47952 24754 48004 24760
rect 48056 23798 48084 26250
rect 48136 25220 48188 25226
rect 48136 25162 48188 25168
rect 48148 24585 48176 25162
rect 48134 24576 48190 24585
rect 48134 24511 48190 24520
rect 48044 23792 48096 23798
rect 48044 23734 48096 23740
rect 47860 23316 47912 23322
rect 47860 23258 47912 23264
rect 48240 23254 48268 26438
rect 48504 25832 48556 25838
rect 48504 25774 48556 25780
rect 48228 23248 48280 23254
rect 48228 23190 48280 23196
rect 48044 22976 48096 22982
rect 48044 22918 48096 22924
rect 48056 22166 48084 22918
rect 48136 22636 48188 22642
rect 48136 22578 48188 22584
rect 48148 22545 48176 22578
rect 48134 22536 48190 22545
rect 48134 22471 48190 22480
rect 48044 22160 48096 22166
rect 48044 22102 48096 22108
rect 47504 22066 47624 22094
rect 47400 17196 47452 17202
rect 47400 17138 47452 17144
rect 47228 16546 47348 16574
rect 47124 11144 47176 11150
rect 47124 11086 47176 11092
rect 46848 9648 46900 9654
rect 46846 9616 46848 9625
rect 46900 9616 46902 9625
rect 46846 9551 46902 9560
rect 46296 7880 46348 7886
rect 46296 7822 46348 7828
rect 46308 7478 46336 7822
rect 46756 7812 46808 7818
rect 46756 7754 46808 7760
rect 46768 7546 46796 7754
rect 46756 7540 46808 7546
rect 46756 7482 46808 7488
rect 46296 7472 46348 7478
rect 46296 7414 46348 7420
rect 46020 6724 46072 6730
rect 46020 6666 46072 6672
rect 46032 6458 46060 6666
rect 46020 6452 46072 6458
rect 46020 6394 46072 6400
rect 45836 6316 45888 6322
rect 45836 6258 45888 6264
rect 45848 4146 45876 6258
rect 46296 6112 46348 6118
rect 46296 6054 46348 6060
rect 46308 5778 46336 6054
rect 46296 5772 46348 5778
rect 46296 5714 46348 5720
rect 46940 5636 46992 5642
rect 46940 5578 46992 5584
rect 46952 5370 46980 5578
rect 47032 5568 47084 5574
rect 47032 5510 47084 5516
rect 46940 5364 46992 5370
rect 46940 5306 46992 5312
rect 46664 5228 46716 5234
rect 46664 5170 46716 5176
rect 45836 4140 45888 4146
rect 45836 4082 45888 4088
rect 45928 4140 45980 4146
rect 45928 4082 45980 4088
rect 45652 3664 45704 3670
rect 45652 3606 45704 3612
rect 45376 3596 45428 3602
rect 45376 3538 45428 3544
rect 45940 3534 45968 4082
rect 46204 3936 46256 3942
rect 46204 3878 46256 3884
rect 46216 3602 46244 3878
rect 46204 3596 46256 3602
rect 46204 3538 46256 3544
rect 46388 3596 46440 3602
rect 46388 3538 46440 3544
rect 45928 3528 45980 3534
rect 45928 3470 45980 3476
rect 45192 3392 45244 3398
rect 45192 3334 45244 3340
rect 45204 2514 45232 3334
rect 45744 3052 45796 3058
rect 45744 2994 45796 3000
rect 45008 2508 45060 2514
rect 45008 2450 45060 2456
rect 45192 2508 45244 2514
rect 45192 2450 45244 2456
rect 45376 2508 45428 2514
rect 45376 2450 45428 2456
rect 45112 870 45232 898
rect 45112 800 45140 870
rect 21376 734 21680 762
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 23846 0 23902 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 25778 0 25834 800
rect 26422 0 26478 800
rect 27066 0 27122 800
rect 27710 0 27766 800
rect 28354 0 28410 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30286 0 30342 800
rect 30930 0 30986 800
rect 31574 0 31630 800
rect 32218 0 32274 800
rect 32862 0 32918 800
rect 33506 0 33562 800
rect 34150 0 34206 800
rect 34794 0 34850 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 36726 0 36782 800
rect 37370 0 37426 800
rect 38014 0 38070 800
rect 38658 0 38714 800
rect 39946 0 40002 800
rect 40590 0 40646 800
rect 41234 0 41290 800
rect 41878 0 41934 800
rect 42522 0 42578 800
rect 43166 0 43222 800
rect 43810 0 43866 800
rect 44454 0 44510 800
rect 45098 0 45154 800
rect 45204 762 45232 870
rect 45388 762 45416 2450
rect 45756 800 45784 2994
rect 46400 800 46428 3538
rect 46570 3360 46626 3369
rect 46570 3295 46626 3304
rect 46584 3058 46612 3295
rect 46676 3126 46704 5170
rect 46756 5160 46808 5166
rect 46756 5102 46808 5108
rect 46768 4185 46796 5102
rect 46848 4820 46900 4826
rect 46848 4762 46900 4768
rect 46754 4176 46810 4185
rect 46754 4111 46810 4120
rect 46756 4072 46808 4078
rect 46756 4014 46808 4020
rect 46664 3120 46716 3126
rect 46664 3062 46716 3068
rect 46572 3052 46624 3058
rect 46572 2994 46624 3000
rect 45204 734 45416 762
rect 45742 0 45798 800
rect 46386 0 46442 800
rect 46768 105 46796 4014
rect 46860 3505 46888 4762
rect 46940 4548 46992 4554
rect 46940 4490 46992 4496
rect 46952 4146 46980 4490
rect 46940 4140 46992 4146
rect 46940 4082 46992 4088
rect 46846 3496 46902 3505
rect 46846 3431 46902 3440
rect 46848 2644 46900 2650
rect 46848 2586 46900 2592
rect 46860 1465 46888 2586
rect 46846 1456 46902 1465
rect 46846 1391 46902 1400
rect 47044 800 47072 5510
rect 47136 3738 47164 11086
rect 47216 11008 47268 11014
rect 47216 10950 47268 10956
rect 47228 10130 47256 10950
rect 47216 10124 47268 10130
rect 47216 10066 47268 10072
rect 47320 6914 47348 16546
rect 47504 16454 47532 22066
rect 47952 21956 48004 21962
rect 47952 21898 48004 21904
rect 47964 21865 47992 21898
rect 47950 21856 48006 21865
rect 47950 21791 48006 21800
rect 48136 19848 48188 19854
rect 48134 19816 48136 19825
rect 48188 19816 48190 19825
rect 48134 19751 48190 19760
rect 47952 19372 48004 19378
rect 47952 19314 48004 19320
rect 47964 19145 47992 19314
rect 48044 19168 48096 19174
rect 47950 19136 48006 19145
rect 48044 19110 48096 19116
rect 47950 19071 48006 19080
rect 47676 16992 47728 16998
rect 47676 16934 47728 16940
rect 47688 16522 47716 16934
rect 47676 16516 47728 16522
rect 47676 16458 47728 16464
rect 47492 16448 47544 16454
rect 47492 16390 47544 16396
rect 47584 15020 47636 15026
rect 47584 14962 47636 14968
rect 47228 6886 47348 6914
rect 47228 5234 47256 6886
rect 47216 5228 47268 5234
rect 47216 5170 47268 5176
rect 47596 4010 47624 14962
rect 47676 14340 47728 14346
rect 47676 14282 47728 14288
rect 47688 13530 47716 14282
rect 47860 13932 47912 13938
rect 47860 13874 47912 13880
rect 47872 13705 47900 13874
rect 47858 13696 47914 13705
rect 47858 13631 47914 13640
rect 47676 13524 47728 13530
rect 47676 13466 47728 13472
rect 47952 11144 48004 11150
rect 47952 11086 48004 11092
rect 47768 10668 47820 10674
rect 47768 10610 47820 10616
rect 47780 10305 47808 10610
rect 47766 10296 47822 10305
rect 47766 10231 47822 10240
rect 47964 10198 47992 11086
rect 47952 10192 48004 10198
rect 47952 10134 48004 10140
rect 48056 9110 48084 19110
rect 48134 17096 48190 17105
rect 48134 17031 48190 17040
rect 48148 16658 48176 17031
rect 48136 16652 48188 16658
rect 48136 16594 48188 16600
rect 48134 16416 48190 16425
rect 48134 16351 48190 16360
rect 48148 15570 48176 16351
rect 48136 15564 48188 15570
rect 48136 15506 48188 15512
rect 48134 14376 48190 14385
rect 48134 14311 48136 14320
rect 48188 14311 48190 14320
rect 48136 14282 48188 14288
rect 48134 10976 48190 10985
rect 48134 10911 48190 10920
rect 48148 10130 48176 10911
rect 48136 10124 48188 10130
rect 48136 10066 48188 10072
rect 48044 9104 48096 9110
rect 48044 9046 48096 9052
rect 47950 8936 48006 8945
rect 47950 8871 47952 8880
rect 48004 8871 48006 8880
rect 47952 8842 48004 8848
rect 47768 8492 47820 8498
rect 47768 8434 47820 8440
rect 47780 8265 47808 8434
rect 47766 8256 47822 8265
rect 47766 8191 47822 8200
rect 48136 7812 48188 7818
rect 48136 7754 48188 7760
rect 48148 7585 48176 7754
rect 48134 7576 48190 7585
rect 48134 7511 48190 7520
rect 47676 6724 47728 6730
rect 47676 6666 47728 6672
rect 47688 6225 47716 6666
rect 47674 6216 47730 6225
rect 47674 6151 47730 6160
rect 48136 5636 48188 5642
rect 48136 5578 48188 5584
rect 47950 5536 48006 5545
rect 47950 5471 48006 5480
rect 47964 5302 47992 5471
rect 47952 5296 48004 5302
rect 47952 5238 48004 5244
rect 48148 4865 48176 5578
rect 48134 4856 48190 4865
rect 48134 4791 48190 4800
rect 48320 4548 48372 4554
rect 48320 4490 48372 4496
rect 47584 4004 47636 4010
rect 47584 3946 47636 3952
rect 48044 3936 48096 3942
rect 48044 3878 48096 3884
rect 47124 3732 47176 3738
rect 47124 3674 47176 3680
rect 48056 3194 48084 3878
rect 48044 3188 48096 3194
rect 48044 3130 48096 3136
rect 47768 2372 47820 2378
rect 47768 2314 47820 2320
rect 46754 96 46810 105
rect 46754 31 46810 40
rect 47030 0 47086 800
rect 47674 0 47730 800
rect 47780 785 47808 2314
rect 48332 800 48360 4490
rect 47766 776 47822 785
rect 47766 711 47822 720
rect 48318 0 48374 800
rect 48516 762 48544 25774
rect 49608 3052 49660 3058
rect 49608 2994 49660 3000
rect 48884 870 49004 898
rect 48884 762 48912 870
rect 48976 800 49004 870
rect 49620 800 49648 2994
rect 48516 734 48912 762
rect 48962 0 49018 800
rect 49606 0 49662 800
<< via2 >>
rect 3790 51720 3846 51776
rect 1398 47640 1454 47696
rect 1398 45600 1454 45656
rect 1398 40160 1454 40216
rect 1398 36760 1454 36816
rect 1398 23840 1454 23896
rect 1398 22480 1454 22536
rect 1398 12280 1454 12336
rect 1398 7520 1454 7576
rect 2870 50360 2926 50416
rect 1858 44240 1914 44296
rect 1858 43560 1914 43616
rect 1858 41520 1914 41576
rect 1858 40840 1914 40896
rect 1858 37440 1914 37496
rect 1582 25900 1638 25936
rect 1582 25880 1584 25900
rect 1584 25880 1636 25900
rect 1636 25880 1638 25900
rect 1858 34720 1914 34776
rect 1858 31320 1914 31376
rect 1858 27240 1914 27296
rect 1858 17040 1914 17096
rect 1858 10920 1914 10976
rect 1858 8200 1914 8256
rect 2778 46280 2834 46336
rect 2870 44920 2926 44976
rect 3054 49000 3110 49056
rect 3422 48340 3478 48376
rect 3422 48320 3424 48340
rect 3424 48320 3476 48340
rect 3476 48320 3478 48340
rect 3054 39480 3110 39536
rect 4066 51040 4122 51096
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4066 46960 4122 47016
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4066 38120 4122 38176
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 2778 36080 2834 36136
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 2778 34060 2834 34096
rect 2778 34040 2780 34060
rect 2780 34040 2832 34060
rect 2832 34040 2834 34060
rect 2778 33396 2780 33416
rect 2780 33396 2832 33416
rect 2832 33396 2834 33416
rect 2778 33360 2834 33396
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 2870 32680 2926 32736
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 3054 32000 3110 32056
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 2870 29960 2926 30016
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 2778 28620 2834 28656
rect 2778 28600 2780 28620
rect 2780 28600 2832 28620
rect 2832 28600 2834 28620
rect 2778 26560 2834 26616
rect 2778 23180 2834 23216
rect 2778 23160 2780 23180
rect 2780 23160 2832 23180
rect 2832 23160 2834 23180
rect 2778 19080 2834 19136
rect 2778 17720 2834 17776
rect 2778 16360 2834 16416
rect 4066 29280 4122 29336
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 2778 13640 2834 13696
rect 2870 10240 2926 10296
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 3974 21800 4030 21856
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4066 21120 4122 21176
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4066 19760 4122 19816
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4066 18400 4122 18456
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4066 12960 4122 13016
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 2962 9560 3018 9616
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4066 8880 4122 8936
rect 2778 6860 2834 6896
rect 2778 6840 2780 6860
rect 2780 6840 2832 6860
rect 2832 6840 2834 6860
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 3606 6160 3662 6216
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 2778 5480 2834 5536
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 2778 4800 2834 4856
rect 1858 3440 1914 3496
rect 3698 4120 3754 4176
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 3422 2080 3478 2136
rect 9402 29164 9458 29200
rect 9402 29144 9404 29164
rect 9404 29144 9456 29164
rect 9456 29144 9458 29164
rect 8666 26988 8722 27024
rect 9494 27920 9550 27976
rect 8666 26968 8668 26988
rect 8668 26968 8720 26988
rect 8720 26968 8722 26988
rect 8850 26560 8906 26616
rect 8390 23044 8446 23080
rect 8390 23024 8392 23044
rect 8392 23024 8444 23044
rect 8444 23024 8446 23044
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4802 2352 4858 2408
rect 2778 720 2834 776
rect 9218 26444 9274 26480
rect 9218 26424 9220 26444
rect 9220 26424 9272 26444
rect 9272 26424 9274 26444
rect 9126 24792 9182 24848
rect 9678 27784 9734 27840
rect 9678 26852 9734 26888
rect 9678 26832 9680 26852
rect 9680 26832 9732 26852
rect 9732 26832 9734 26852
rect 9954 27920 10010 27976
rect 9954 27820 9956 27840
rect 9956 27820 10008 27840
rect 10008 27820 10010 27840
rect 9954 27784 10010 27820
rect 10046 26852 10102 26888
rect 10046 26832 10048 26852
rect 10048 26832 10100 26852
rect 10100 26832 10102 26852
rect 10414 27004 10416 27024
rect 10416 27004 10468 27024
rect 10468 27004 10470 27024
rect 10414 26968 10470 27004
rect 10598 26560 10654 26616
rect 9954 25492 10010 25528
rect 9954 25472 9956 25492
rect 9956 25472 10008 25492
rect 10008 25472 10010 25492
rect 12254 24132 12310 24168
rect 12254 24112 12256 24132
rect 12256 24112 12308 24132
rect 12308 24112 12310 24132
rect 9862 23044 9918 23080
rect 9862 23024 9864 23044
rect 9864 23024 9916 23044
rect 9916 23024 9918 23044
rect 12346 22616 12402 22672
rect 10414 17312 10470 17368
rect 14554 25492 14610 25528
rect 14554 25472 14556 25492
rect 14556 25472 14608 25492
rect 14608 25472 14610 25492
rect 14554 22616 14610 22672
rect 15014 22636 15070 22672
rect 15014 22616 15016 22636
rect 15016 22616 15068 22636
rect 15068 22616 15070 22636
rect 14922 18128 14978 18184
rect 14646 17856 14702 17912
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 16210 22636 16266 22672
rect 16210 22616 16212 22636
rect 16212 22616 16264 22636
rect 16264 22616 16266 22636
rect 17774 29164 17830 29200
rect 17774 29144 17776 29164
rect 17776 29144 17828 29164
rect 17828 29144 17830 29164
rect 17590 26424 17646 26480
rect 17682 26288 17738 26344
rect 17406 24812 17462 24848
rect 18142 26288 18198 26344
rect 17958 25200 18014 25256
rect 17406 24792 17408 24812
rect 17408 24792 17460 24812
rect 17460 24792 17462 24812
rect 16854 24112 16910 24168
rect 15382 17584 15438 17640
rect 16026 17312 16082 17368
rect 16946 17584 17002 17640
rect 17406 18164 17408 18184
rect 17408 18164 17460 18184
rect 17460 18164 17462 18184
rect 17406 18128 17462 18164
rect 14738 2508 14794 2544
rect 14738 2488 14740 2508
rect 14740 2488 14792 2508
rect 14792 2488 14794 2508
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19706 37884 19708 37904
rect 19708 37884 19760 37904
rect 19760 37884 19762 37904
rect 19706 37848 19762 37884
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 20350 37032 20406 37088
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19706 30096 19762 30152
rect 19982 29688 20038 29744
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19982 28192 20038 28248
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 18418 17856 18474 17912
rect 20994 35692 21050 35728
rect 20994 35672 20996 35692
rect 20996 35672 21048 35692
rect 21048 35672 21050 35692
rect 20534 30368 20590 30424
rect 20350 30232 20406 30288
rect 20350 29280 20406 29336
rect 20350 26968 20406 27024
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19982 25472 20038 25528
rect 20258 25608 20314 25664
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19890 24828 19892 24848
rect 19892 24828 19944 24848
rect 19944 24828 19946 24848
rect 19890 24792 19946 24828
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19522 22616 19578 22672
rect 19798 22228 19854 22264
rect 19798 22208 19800 22228
rect 19800 22208 19852 22228
rect 19852 22208 19854 22228
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19890 19352 19946 19408
rect 19890 18672 19946 18728
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19430 15408 19486 15464
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19614 15000 19670 15056
rect 19614 14340 19670 14376
rect 19614 14320 19616 14340
rect 19616 14320 19668 14340
rect 19668 14320 19670 14340
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19338 12144 19394 12200
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19890 11756 19946 11792
rect 19890 11736 19892 11756
rect 19892 11736 19944 11756
rect 19944 11736 19946 11756
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19338 9560 19394 9616
rect 20258 23024 20314 23080
rect 20166 14320 20222 14376
rect 20074 12688 20130 12744
rect 20994 29688 21050 29744
rect 20350 19624 20406 19680
rect 20350 17312 20406 17368
rect 21178 25200 21234 25256
rect 20626 19760 20682 19816
rect 20074 9968 20130 10024
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19614 9580 19670 9616
rect 19614 9560 19616 9580
rect 19616 9560 19668 9580
rect 19668 9560 19670 9580
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19430 7384 19486 7440
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 20350 10376 20406 10432
rect 20626 16904 20682 16960
rect 21086 17720 21142 17776
rect 20534 11600 20590 11656
rect 21270 11600 21326 11656
rect 20350 3576 20406 3632
rect 19890 3476 19892 3496
rect 19892 3476 19944 3496
rect 19944 3476 19946 3496
rect 19890 3440 19946 3476
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 21822 24656 21878 24712
rect 21914 24112 21970 24168
rect 22098 21292 22100 21312
rect 22100 21292 22152 21312
rect 22152 21292 22154 21312
rect 22098 21256 22154 21292
rect 22098 19352 22154 19408
rect 22282 17720 22338 17776
rect 21822 13368 21878 13424
rect 23478 39092 23534 39128
rect 23478 39072 23480 39092
rect 23480 39072 23532 39092
rect 23532 39072 23534 39092
rect 23386 29452 23388 29472
rect 23388 29452 23440 29472
rect 23440 29452 23442 29472
rect 23386 29416 23442 29452
rect 24766 33940 24768 33960
rect 24768 33940 24820 33960
rect 24820 33940 24822 33960
rect 23754 25492 23810 25528
rect 23754 25472 23756 25492
rect 23756 25472 23808 25492
rect 23808 25472 23810 25492
rect 23110 24928 23166 24984
rect 23386 23468 23388 23488
rect 23388 23468 23440 23488
rect 23440 23468 23442 23488
rect 23386 23432 23442 23468
rect 23846 24928 23902 24984
rect 23754 20848 23810 20904
rect 23662 20304 23718 20360
rect 23386 7928 23442 7984
rect 23294 7792 23350 7848
rect 24122 25744 24178 25800
rect 24766 33904 24822 33940
rect 24582 30368 24638 30424
rect 24858 29452 24860 29472
rect 24860 29452 24912 29472
rect 24912 29452 24914 29472
rect 24858 29416 24914 29452
rect 24122 22344 24178 22400
rect 24122 20712 24178 20768
rect 24122 17584 24178 17640
rect 24122 17176 24178 17232
rect 25042 29824 25098 29880
rect 26330 37848 26386 37904
rect 26054 34060 26110 34096
rect 26054 34040 26056 34060
rect 26056 34040 26108 34060
rect 26108 34040 26110 34060
rect 26790 39072 26846 39128
rect 26054 30368 26110 30424
rect 25134 24792 25190 24848
rect 24122 9696 24178 9752
rect 24674 23468 24676 23488
rect 24676 23468 24728 23488
rect 24728 23468 24730 23488
rect 24674 23432 24730 23468
rect 24950 20712 25006 20768
rect 24766 17176 24822 17232
rect 25686 25608 25742 25664
rect 25502 22616 25558 22672
rect 25042 14340 25098 14376
rect 25042 14320 25044 14340
rect 25044 14320 25096 14340
rect 25096 14320 25098 14340
rect 25042 7828 25044 7848
rect 25044 7828 25096 7848
rect 25096 7828 25098 7848
rect 25042 7792 25098 7828
rect 25318 7928 25374 7984
rect 25686 21256 25742 21312
rect 25870 29280 25926 29336
rect 26330 24248 26386 24304
rect 26146 22636 26202 22672
rect 26146 22616 26148 22636
rect 26148 22616 26200 22636
rect 26200 22616 26202 22636
rect 26238 13368 26294 13424
rect 26238 3576 26294 3632
rect 27066 34076 27068 34096
rect 27068 34076 27120 34096
rect 27120 34076 27122 34096
rect 27066 34040 27122 34076
rect 27710 35692 27766 35728
rect 27710 35672 27712 35692
rect 27712 35672 27764 35692
rect 27764 35672 27766 35692
rect 27342 30096 27398 30152
rect 27986 29844 28042 29880
rect 27986 29824 27988 29844
rect 27988 29824 28040 29844
rect 28040 29824 28042 29844
rect 28354 33924 28410 33960
rect 28354 33904 28356 33924
rect 28356 33904 28408 33924
rect 28408 33904 28410 33924
rect 27618 24248 27674 24304
rect 28630 24656 28686 24712
rect 27158 16244 27214 16280
rect 27158 16224 27160 16244
rect 27160 16224 27212 16244
rect 27212 16224 27214 16244
rect 26974 14320 27030 14376
rect 26606 11736 26662 11792
rect 27618 17584 27674 17640
rect 27894 11872 27950 11928
rect 28078 11872 28134 11928
rect 28078 11600 28134 11656
rect 27250 7828 27252 7848
rect 27252 7828 27304 7848
rect 27304 7828 27306 7848
rect 27250 7792 27306 7828
rect 27986 3476 27988 3496
rect 27988 3476 28040 3496
rect 28040 3476 28042 3496
rect 27986 3440 28042 3476
rect 28998 23840 29054 23896
rect 29642 38664 29698 38720
rect 29918 38156 29920 38176
rect 29920 38156 29972 38176
rect 29972 38156 29974 38176
rect 29918 38120 29974 38156
rect 31666 38392 31722 38448
rect 29366 24384 29422 24440
rect 28998 23060 29000 23080
rect 29000 23060 29052 23080
rect 29052 23060 29054 23080
rect 28998 23024 29054 23060
rect 30194 23060 30196 23080
rect 30196 23060 30248 23080
rect 30248 23060 30250 23080
rect 30194 23024 30250 23060
rect 30378 21956 30434 21992
rect 30378 21936 30380 21956
rect 30380 21936 30432 21956
rect 30432 21936 30434 21956
rect 28354 14356 28356 14376
rect 28356 14356 28408 14376
rect 28408 14356 28410 14376
rect 28354 14320 28410 14356
rect 30654 22108 30656 22128
rect 30656 22108 30708 22128
rect 30708 22108 30710 22128
rect 30654 22072 30710 22108
rect 30378 16224 30434 16280
rect 32034 38156 32036 38176
rect 32036 38156 32088 38176
rect 32088 38156 32090 38176
rect 32034 38120 32090 38156
rect 31574 35012 31630 35048
rect 31574 34992 31576 35012
rect 31576 34992 31628 35012
rect 31628 34992 31630 35012
rect 31574 22108 31576 22128
rect 31576 22108 31628 22128
rect 31628 22108 31630 22128
rect 31574 22072 31630 22108
rect 33046 35012 33102 35048
rect 33046 34992 33048 35012
rect 33048 34992 33100 35012
rect 33100 34992 33102 35012
rect 32218 26832 32274 26888
rect 32678 24384 32734 24440
rect 32402 24112 32458 24168
rect 32310 23840 32366 23896
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 32034 21936 32090 21992
rect 33690 26832 33746 26888
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 35162 38428 35164 38448
rect 35164 38428 35216 38448
rect 35216 38428 35218 38448
rect 35162 38392 35218 38428
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34794 29708 34850 29744
rect 34794 29688 34796 29708
rect 34796 29688 34848 29708
rect 34848 29688 34850 29708
rect 34702 29300 34758 29336
rect 34702 29280 34704 29300
rect 34704 29280 34756 29300
rect 34756 29280 34758 29300
rect 35530 29708 35586 29744
rect 35530 29688 35532 29708
rect 35532 29688 35584 29708
rect 35584 29688 35586 29708
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 35714 29280 35770 29336
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 39026 3304 39082 3360
rect 46662 51720 46718 51776
rect 46570 51040 46626 51096
rect 45466 26560 45522 26616
rect 46754 50360 46810 50416
rect 46846 49680 46902 49736
rect 47766 49000 47822 49056
rect 47766 48320 47822 48376
rect 46846 46960 46902 47016
rect 46570 44920 46626 44976
rect 46110 44240 46166 44296
rect 46202 40840 46258 40896
rect 46202 37440 46258 37496
rect 46846 34040 46902 34096
rect 46386 17720 46442 17776
rect 47858 42880 47914 42936
rect 48134 46280 48190 46336
rect 48134 45600 48190 45656
rect 48134 43560 48190 43616
rect 47950 42200 48006 42256
rect 48134 41540 48190 41576
rect 48134 41520 48136 41540
rect 48136 41520 48188 41540
rect 48188 41520 48190 41540
rect 47306 29960 47362 30016
rect 46846 15020 46902 15056
rect 46846 15000 46848 15020
rect 46848 15000 46900 15020
rect 46900 15000 46902 15020
rect 46846 12960 46902 13016
rect 46846 12280 46902 12336
rect 47306 23840 47362 23896
rect 47674 32000 47730 32056
rect 48134 40160 48190 40216
rect 48134 39480 48190 39536
rect 47950 38800 48006 38856
rect 47858 38120 47914 38176
rect 48134 36760 48190 36816
rect 47858 36080 47914 36136
rect 47950 33360 48006 33416
rect 48226 35400 48282 35456
rect 48134 34720 48190 34776
rect 47950 31320 48006 31376
rect 47858 27920 47914 27976
rect 48134 29280 48190 29336
rect 48226 28600 48282 28656
rect 47950 25880 48006 25936
rect 47950 25200 48006 25256
rect 48134 24520 48190 24576
rect 48134 22480 48190 22536
rect 46846 9596 46848 9616
rect 46848 9596 46900 9616
rect 46900 9596 46902 9616
rect 46846 9560 46902 9596
rect 46570 3304 46626 3360
rect 46754 4120 46810 4176
rect 46846 3440 46902 3496
rect 46846 1400 46902 1456
rect 47950 21800 48006 21856
rect 48134 19796 48136 19816
rect 48136 19796 48188 19816
rect 48188 19796 48190 19816
rect 48134 19760 48190 19796
rect 47950 19080 48006 19136
rect 47858 13640 47914 13696
rect 47766 10240 47822 10296
rect 48134 17040 48190 17096
rect 48134 16360 48190 16416
rect 48134 14340 48190 14376
rect 48134 14320 48136 14340
rect 48136 14320 48188 14340
rect 48188 14320 48190 14340
rect 48134 10920 48190 10976
rect 47950 8900 48006 8936
rect 47950 8880 47952 8900
rect 47952 8880 48004 8900
rect 48004 8880 48006 8900
rect 47766 8200 47822 8256
rect 48134 7520 48190 7576
rect 47674 6160 47730 6216
rect 47950 5480 48006 5536
rect 48134 4800 48190 4856
rect 46754 40 46810 96
rect 47766 720 47822 776
<< metal3 >>
rect 0 51778 800 51808
rect 3785 51778 3851 51781
rect 0 51776 3851 51778
rect 0 51720 3790 51776
rect 3846 51720 3851 51776
rect 0 51718 3851 51720
rect 0 51688 800 51718
rect 3785 51715 3851 51718
rect 46657 51778 46723 51781
rect 49200 51778 50000 51808
rect 46657 51776 50000 51778
rect 46657 51720 46662 51776
rect 46718 51720 50000 51776
rect 46657 51718 50000 51720
rect 46657 51715 46723 51718
rect 49200 51688 50000 51718
rect 0 51098 800 51128
rect 4061 51098 4127 51101
rect 0 51096 4127 51098
rect 0 51040 4066 51096
rect 4122 51040 4127 51096
rect 0 51038 4127 51040
rect 0 51008 800 51038
rect 4061 51035 4127 51038
rect 46565 51098 46631 51101
rect 49200 51098 50000 51128
rect 46565 51096 50000 51098
rect 46565 51040 46570 51096
rect 46626 51040 50000 51096
rect 46565 51038 50000 51040
rect 46565 51035 46631 51038
rect 49200 51008 50000 51038
rect 0 50418 800 50448
rect 2865 50418 2931 50421
rect 0 50416 2931 50418
rect 0 50360 2870 50416
rect 2926 50360 2931 50416
rect 0 50358 2931 50360
rect 0 50328 800 50358
rect 2865 50355 2931 50358
rect 46749 50418 46815 50421
rect 49200 50418 50000 50448
rect 46749 50416 50000 50418
rect 46749 50360 46754 50416
rect 46810 50360 50000 50416
rect 46749 50358 50000 50360
rect 46749 50355 46815 50358
rect 49200 50328 50000 50358
rect 0 49648 800 49768
rect 46841 49738 46907 49741
rect 49200 49738 50000 49768
rect 46841 49736 50000 49738
rect 46841 49680 46846 49736
rect 46902 49680 50000 49736
rect 46841 49678 50000 49680
rect 46841 49675 46907 49678
rect 49200 49648 50000 49678
rect 4208 49536 4528 49537
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 49471 4528 49472
rect 34928 49536 35248 49537
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 49471 35248 49472
rect 0 49058 800 49088
rect 3049 49058 3115 49061
rect 0 49056 3115 49058
rect 0 49000 3054 49056
rect 3110 49000 3115 49056
rect 0 48998 3115 49000
rect 0 48968 800 48998
rect 3049 48995 3115 48998
rect 47761 49058 47827 49061
rect 49200 49058 50000 49088
rect 47761 49056 50000 49058
rect 47761 49000 47766 49056
rect 47822 49000 50000 49056
rect 47761 48998 50000 49000
rect 47761 48995 47827 48998
rect 19568 48992 19888 48993
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 49200 48968 50000 48998
rect 19568 48927 19888 48928
rect 4208 48448 4528 48449
rect 0 48378 800 48408
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 48383 4528 48384
rect 34928 48448 35248 48449
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 48383 35248 48384
rect 3417 48378 3483 48381
rect 0 48376 3483 48378
rect 0 48320 3422 48376
rect 3478 48320 3483 48376
rect 0 48318 3483 48320
rect 0 48288 800 48318
rect 3417 48315 3483 48318
rect 47761 48378 47827 48381
rect 49200 48378 50000 48408
rect 47761 48376 50000 48378
rect 47761 48320 47766 48376
rect 47822 48320 50000 48376
rect 47761 48318 50000 48320
rect 47761 48315 47827 48318
rect 49200 48288 50000 48318
rect 19568 47904 19888 47905
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 47839 19888 47840
rect 0 47698 800 47728
rect 1393 47698 1459 47701
rect 0 47696 1459 47698
rect 0 47640 1398 47696
rect 1454 47640 1459 47696
rect 0 47638 1459 47640
rect 0 47608 800 47638
rect 1393 47635 1459 47638
rect 49200 47608 50000 47728
rect 4208 47360 4528 47361
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 47295 4528 47296
rect 34928 47360 35248 47361
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 47295 35248 47296
rect 0 47018 800 47048
rect 4061 47018 4127 47021
rect 0 47016 4127 47018
rect 0 46960 4066 47016
rect 4122 46960 4127 47016
rect 0 46958 4127 46960
rect 0 46928 800 46958
rect 4061 46955 4127 46958
rect 46841 47018 46907 47021
rect 49200 47018 50000 47048
rect 46841 47016 50000 47018
rect 46841 46960 46846 47016
rect 46902 46960 50000 47016
rect 46841 46958 50000 46960
rect 46841 46955 46907 46958
rect 49200 46928 50000 46958
rect 19568 46816 19888 46817
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 46751 19888 46752
rect 0 46338 800 46368
rect 2773 46338 2839 46341
rect 0 46336 2839 46338
rect 0 46280 2778 46336
rect 2834 46280 2839 46336
rect 0 46278 2839 46280
rect 0 46248 800 46278
rect 2773 46275 2839 46278
rect 48129 46338 48195 46341
rect 49200 46338 50000 46368
rect 48129 46336 50000 46338
rect 48129 46280 48134 46336
rect 48190 46280 50000 46336
rect 48129 46278 50000 46280
rect 48129 46275 48195 46278
rect 4208 46272 4528 46273
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 46207 4528 46208
rect 34928 46272 35248 46273
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 49200 46248 50000 46278
rect 34928 46207 35248 46208
rect 19568 45728 19888 45729
rect 0 45658 800 45688
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 45663 19888 45664
rect 1393 45658 1459 45661
rect 0 45656 1459 45658
rect 0 45600 1398 45656
rect 1454 45600 1459 45656
rect 0 45598 1459 45600
rect 0 45568 800 45598
rect 1393 45595 1459 45598
rect 48129 45658 48195 45661
rect 49200 45658 50000 45688
rect 48129 45656 50000 45658
rect 48129 45600 48134 45656
rect 48190 45600 50000 45656
rect 48129 45598 50000 45600
rect 48129 45595 48195 45598
rect 49200 45568 50000 45598
rect 4208 45184 4528 45185
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 45119 4528 45120
rect 34928 45184 35248 45185
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 45119 35248 45120
rect 0 44978 800 45008
rect 2865 44978 2931 44981
rect 0 44976 2931 44978
rect 0 44920 2870 44976
rect 2926 44920 2931 44976
rect 0 44918 2931 44920
rect 0 44888 800 44918
rect 2865 44915 2931 44918
rect 46565 44978 46631 44981
rect 49200 44978 50000 45008
rect 46565 44976 50000 44978
rect 46565 44920 46570 44976
rect 46626 44920 50000 44976
rect 46565 44918 50000 44920
rect 46565 44915 46631 44918
rect 49200 44888 50000 44918
rect 19568 44640 19888 44641
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 44575 19888 44576
rect 0 44298 800 44328
rect 1853 44298 1919 44301
rect 0 44296 1919 44298
rect 0 44240 1858 44296
rect 1914 44240 1919 44296
rect 0 44238 1919 44240
rect 0 44208 800 44238
rect 1853 44235 1919 44238
rect 46105 44298 46171 44301
rect 49200 44298 50000 44328
rect 46105 44296 50000 44298
rect 46105 44240 46110 44296
rect 46166 44240 50000 44296
rect 46105 44238 50000 44240
rect 46105 44235 46171 44238
rect 49200 44208 50000 44238
rect 4208 44096 4528 44097
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 44031 4528 44032
rect 34928 44096 35248 44097
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 44031 35248 44032
rect 0 43618 800 43648
rect 1853 43618 1919 43621
rect 0 43616 1919 43618
rect 0 43560 1858 43616
rect 1914 43560 1919 43616
rect 0 43558 1919 43560
rect 0 43528 800 43558
rect 1853 43555 1919 43558
rect 48129 43618 48195 43621
rect 49200 43618 50000 43648
rect 48129 43616 50000 43618
rect 48129 43560 48134 43616
rect 48190 43560 50000 43616
rect 48129 43558 50000 43560
rect 48129 43555 48195 43558
rect 19568 43552 19888 43553
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 49200 43528 50000 43558
rect 19568 43487 19888 43488
rect 4208 43008 4528 43009
rect 0 42848 800 42968
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 42943 4528 42944
rect 34928 43008 35248 43009
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 42943 35248 42944
rect 47853 42938 47919 42941
rect 49200 42938 50000 42968
rect 47853 42936 50000 42938
rect 47853 42880 47858 42936
rect 47914 42880 50000 42936
rect 47853 42878 50000 42880
rect 47853 42875 47919 42878
rect 49200 42848 50000 42878
rect 19568 42464 19888 42465
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 42399 19888 42400
rect 47945 42258 48011 42261
rect 49200 42258 50000 42288
rect 47945 42256 50000 42258
rect 47945 42200 47950 42256
rect 48006 42200 50000 42256
rect 47945 42198 50000 42200
rect 47945 42195 48011 42198
rect 49200 42168 50000 42198
rect 4208 41920 4528 41921
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 41855 4528 41856
rect 34928 41920 35248 41921
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 41855 35248 41856
rect 0 41578 800 41608
rect 1853 41578 1919 41581
rect 0 41576 1919 41578
rect 0 41520 1858 41576
rect 1914 41520 1919 41576
rect 0 41518 1919 41520
rect 0 41488 800 41518
rect 1853 41515 1919 41518
rect 48129 41578 48195 41581
rect 49200 41578 50000 41608
rect 48129 41576 50000 41578
rect 48129 41520 48134 41576
rect 48190 41520 50000 41576
rect 48129 41518 50000 41520
rect 48129 41515 48195 41518
rect 49200 41488 50000 41518
rect 19568 41376 19888 41377
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 41311 19888 41312
rect 0 40898 800 40928
rect 1853 40898 1919 40901
rect 0 40896 1919 40898
rect 0 40840 1858 40896
rect 1914 40840 1919 40896
rect 0 40838 1919 40840
rect 0 40808 800 40838
rect 1853 40835 1919 40838
rect 46197 40898 46263 40901
rect 49200 40898 50000 40928
rect 46197 40896 50000 40898
rect 46197 40840 46202 40896
rect 46258 40840 50000 40896
rect 46197 40838 50000 40840
rect 46197 40835 46263 40838
rect 4208 40832 4528 40833
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 40767 4528 40768
rect 34928 40832 35248 40833
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 49200 40808 50000 40838
rect 34928 40767 35248 40768
rect 19568 40288 19888 40289
rect 0 40218 800 40248
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 40223 19888 40224
rect 1393 40218 1459 40221
rect 0 40216 1459 40218
rect 0 40160 1398 40216
rect 1454 40160 1459 40216
rect 0 40158 1459 40160
rect 0 40128 800 40158
rect 1393 40155 1459 40158
rect 48129 40218 48195 40221
rect 49200 40218 50000 40248
rect 48129 40216 50000 40218
rect 48129 40160 48134 40216
rect 48190 40160 50000 40216
rect 48129 40158 50000 40160
rect 48129 40155 48195 40158
rect 49200 40128 50000 40158
rect 4208 39744 4528 39745
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 0 39538 800 39568
rect 3049 39538 3115 39541
rect 0 39536 3115 39538
rect 0 39480 3054 39536
rect 3110 39480 3115 39536
rect 0 39478 3115 39480
rect 0 39448 800 39478
rect 3049 39475 3115 39478
rect 48129 39538 48195 39541
rect 49200 39538 50000 39568
rect 48129 39536 50000 39538
rect 48129 39480 48134 39536
rect 48190 39480 50000 39536
rect 48129 39478 50000 39480
rect 48129 39475 48195 39478
rect 49200 39448 50000 39478
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 39135 19888 39136
rect 23473 39130 23539 39133
rect 26785 39130 26851 39133
rect 23473 39128 26851 39130
rect 23473 39072 23478 39128
rect 23534 39072 26790 39128
rect 26846 39072 26851 39128
rect 23473 39070 26851 39072
rect 23473 39067 23539 39070
rect 26785 39067 26851 39070
rect 0 38768 800 38888
rect 47945 38858 48011 38861
rect 49200 38858 50000 38888
rect 47945 38856 50000 38858
rect 47945 38800 47950 38856
rect 48006 38800 50000 38856
rect 47945 38798 50000 38800
rect 47945 38795 48011 38798
rect 49200 38768 50000 38798
rect 24158 38660 24164 38724
rect 24228 38722 24234 38724
rect 29637 38722 29703 38725
rect 24228 38720 29703 38722
rect 24228 38664 29642 38720
rect 29698 38664 29703 38720
rect 24228 38662 29703 38664
rect 24228 38660 24234 38662
rect 29637 38659 29703 38662
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 38591 35248 38592
rect 31661 38450 31727 38453
rect 35157 38450 35223 38453
rect 31661 38448 35223 38450
rect 31661 38392 31666 38448
rect 31722 38392 35162 38448
rect 35218 38392 35223 38448
rect 31661 38390 35223 38392
rect 31661 38387 31727 38390
rect 35157 38387 35223 38390
rect 0 38178 800 38208
rect 4061 38178 4127 38181
rect 0 38176 4127 38178
rect 0 38120 4066 38176
rect 4122 38120 4127 38176
rect 0 38118 4127 38120
rect 0 38088 800 38118
rect 4061 38115 4127 38118
rect 29913 38178 29979 38181
rect 32029 38178 32095 38181
rect 29913 38176 32095 38178
rect 29913 38120 29918 38176
rect 29974 38120 32034 38176
rect 32090 38120 32095 38176
rect 29913 38118 32095 38120
rect 29913 38115 29979 38118
rect 32029 38115 32095 38118
rect 47853 38178 47919 38181
rect 49200 38178 50000 38208
rect 47853 38176 50000 38178
rect 47853 38120 47858 38176
rect 47914 38120 50000 38176
rect 47853 38118 50000 38120
rect 47853 38115 47919 38118
rect 19568 38112 19888 38113
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 49200 38088 50000 38118
rect 19568 38047 19888 38048
rect 19701 37906 19767 37909
rect 26325 37906 26391 37909
rect 19701 37904 26391 37906
rect 19701 37848 19706 37904
rect 19762 37848 26330 37904
rect 26386 37848 26391 37904
rect 19701 37846 26391 37848
rect 19701 37843 19767 37846
rect 26325 37843 26391 37846
rect 4208 37568 4528 37569
rect 0 37498 800 37528
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 1853 37498 1919 37501
rect 0 37496 1919 37498
rect 0 37440 1858 37496
rect 1914 37440 1919 37496
rect 0 37438 1919 37440
rect 0 37408 800 37438
rect 1853 37435 1919 37438
rect 46197 37498 46263 37501
rect 49200 37498 50000 37528
rect 46197 37496 50000 37498
rect 46197 37440 46202 37496
rect 46258 37440 50000 37496
rect 46197 37438 50000 37440
rect 46197 37435 46263 37438
rect 49200 37408 50000 37438
rect 20345 37092 20411 37093
rect 20294 37028 20300 37092
rect 20364 37090 20411 37092
rect 20364 37088 20456 37090
rect 20406 37032 20456 37088
rect 20364 37030 20456 37032
rect 20364 37028 20411 37030
rect 20345 37027 20411 37028
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 0 36818 800 36848
rect 1393 36818 1459 36821
rect 0 36816 1459 36818
rect 0 36760 1398 36816
rect 1454 36760 1459 36816
rect 0 36758 1459 36760
rect 0 36728 800 36758
rect 1393 36755 1459 36758
rect 48129 36818 48195 36821
rect 49200 36818 50000 36848
rect 48129 36816 50000 36818
rect 48129 36760 48134 36816
rect 48190 36760 50000 36816
rect 48129 36758 50000 36760
rect 48129 36755 48195 36758
rect 49200 36728 50000 36758
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 0 36138 800 36168
rect 2773 36138 2839 36141
rect 0 36136 2839 36138
rect 0 36080 2778 36136
rect 2834 36080 2839 36136
rect 0 36078 2839 36080
rect 0 36048 800 36078
rect 2773 36075 2839 36078
rect 47853 36138 47919 36141
rect 49200 36138 50000 36168
rect 47853 36136 50000 36138
rect 47853 36080 47858 36136
rect 47914 36080 50000 36136
rect 47853 36078 50000 36080
rect 47853 36075 47919 36078
rect 49200 36048 50000 36078
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 20989 35730 21055 35733
rect 27705 35730 27771 35733
rect 20989 35728 27771 35730
rect 20989 35672 20994 35728
rect 21050 35672 27710 35728
rect 27766 35672 27771 35728
rect 20989 35670 27771 35672
rect 20989 35667 21055 35670
rect 27705 35667 27771 35670
rect 0 35368 800 35488
rect 48221 35458 48287 35461
rect 49200 35458 50000 35488
rect 48221 35456 50000 35458
rect 48221 35400 48226 35456
rect 48282 35400 50000 35456
rect 48221 35398 50000 35400
rect 48221 35395 48287 35398
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 49200 35368 50000 35398
rect 34928 35327 35248 35328
rect 31569 35050 31635 35053
rect 33041 35050 33107 35053
rect 31569 35048 33107 35050
rect 31569 34992 31574 35048
rect 31630 34992 33046 35048
rect 33102 34992 33107 35048
rect 31569 34990 33107 34992
rect 31569 34987 31635 34990
rect 33041 34987 33107 34990
rect 19568 34848 19888 34849
rect 0 34778 800 34808
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 1853 34778 1919 34781
rect 0 34776 1919 34778
rect 0 34720 1858 34776
rect 1914 34720 1919 34776
rect 0 34718 1919 34720
rect 0 34688 800 34718
rect 1853 34715 1919 34718
rect 48129 34778 48195 34781
rect 49200 34778 50000 34808
rect 48129 34776 50000 34778
rect 48129 34720 48134 34776
rect 48190 34720 50000 34776
rect 48129 34718 50000 34720
rect 48129 34715 48195 34718
rect 49200 34688 50000 34718
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 0 34098 800 34128
rect 2773 34098 2839 34101
rect 0 34096 2839 34098
rect 0 34040 2778 34096
rect 2834 34040 2839 34096
rect 0 34038 2839 34040
rect 0 34008 800 34038
rect 2773 34035 2839 34038
rect 26049 34098 26115 34101
rect 27061 34098 27127 34101
rect 26049 34096 27127 34098
rect 26049 34040 26054 34096
rect 26110 34040 27066 34096
rect 27122 34040 27127 34096
rect 26049 34038 27127 34040
rect 26049 34035 26115 34038
rect 27061 34035 27127 34038
rect 46841 34098 46907 34101
rect 49200 34098 50000 34128
rect 46841 34096 50000 34098
rect 46841 34040 46846 34096
rect 46902 34040 50000 34096
rect 46841 34038 50000 34040
rect 46841 34035 46907 34038
rect 49200 34008 50000 34038
rect 24761 33962 24827 33965
rect 28349 33962 28415 33965
rect 24761 33960 28415 33962
rect 24761 33904 24766 33960
rect 24822 33904 28354 33960
rect 28410 33904 28415 33960
rect 24761 33902 28415 33904
rect 24761 33899 24827 33902
rect 28349 33899 28415 33902
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 0 33418 800 33448
rect 2773 33418 2839 33421
rect 0 33416 2839 33418
rect 0 33360 2778 33416
rect 2834 33360 2839 33416
rect 0 33358 2839 33360
rect 0 33328 800 33358
rect 2773 33355 2839 33358
rect 47945 33418 48011 33421
rect 49200 33418 50000 33448
rect 47945 33416 50000 33418
rect 47945 33360 47950 33416
rect 48006 33360 50000 33416
rect 47945 33358 50000 33360
rect 47945 33355 48011 33358
rect 49200 33328 50000 33358
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 0 32738 800 32768
rect 2865 32738 2931 32741
rect 0 32736 2931 32738
rect 0 32680 2870 32736
rect 2926 32680 2931 32736
rect 0 32678 2931 32680
rect 0 32648 800 32678
rect 2865 32675 2931 32678
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 49200 32648 50000 32768
rect 19568 32607 19888 32608
rect 4208 32128 4528 32129
rect 0 32058 800 32088
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 3049 32058 3115 32061
rect 0 32056 3115 32058
rect 0 32000 3054 32056
rect 3110 32000 3115 32056
rect 0 31998 3115 32000
rect 0 31968 800 31998
rect 3049 31995 3115 31998
rect 47669 32058 47735 32061
rect 49200 32058 50000 32088
rect 47669 32056 50000 32058
rect 47669 32000 47674 32056
rect 47730 32000 50000 32056
rect 47669 31998 50000 32000
rect 47669 31995 47735 31998
rect 49200 31968 50000 31998
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 0 31378 800 31408
rect 1853 31378 1919 31381
rect 0 31376 1919 31378
rect 0 31320 1858 31376
rect 1914 31320 1919 31376
rect 0 31318 1919 31320
rect 0 31288 800 31318
rect 1853 31315 1919 31318
rect 47945 31378 48011 31381
rect 49200 31378 50000 31408
rect 47945 31376 50000 31378
rect 47945 31320 47950 31376
rect 48006 31320 50000 31376
rect 47945 31318 50000 31320
rect 47945 31315 48011 31318
rect 49200 31288 50000 31318
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 0 30608 800 30728
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 20529 30426 20595 30429
rect 21214 30426 21220 30428
rect 20529 30424 21220 30426
rect 20529 30368 20534 30424
rect 20590 30368 21220 30424
rect 20529 30366 21220 30368
rect 20529 30363 20595 30366
rect 21214 30364 21220 30366
rect 21284 30364 21290 30428
rect 24577 30426 24643 30429
rect 26049 30426 26115 30429
rect 24577 30424 26115 30426
rect 24577 30368 24582 30424
rect 24638 30368 26054 30424
rect 26110 30368 26115 30424
rect 24577 30366 26115 30368
rect 24577 30363 24643 30366
rect 26049 30363 26115 30366
rect 20345 30290 20411 30293
rect 20302 30288 20411 30290
rect 20302 30232 20350 30288
rect 20406 30232 20411 30288
rect 20302 30227 20411 30232
rect 19701 30154 19767 30157
rect 20302 30154 20362 30227
rect 27337 30154 27403 30157
rect 19701 30152 27403 30154
rect 19701 30096 19706 30152
rect 19762 30096 27342 30152
rect 27398 30096 27403 30152
rect 19701 30094 27403 30096
rect 19701 30091 19767 30094
rect 27337 30091 27403 30094
rect 0 30018 800 30048
rect 2865 30018 2931 30021
rect 0 30016 2931 30018
rect 0 29960 2870 30016
rect 2926 29960 2931 30016
rect 0 29958 2931 29960
rect 0 29928 800 29958
rect 2865 29955 2931 29958
rect 47301 30018 47367 30021
rect 49200 30018 50000 30048
rect 47301 30016 50000 30018
rect 47301 29960 47306 30016
rect 47362 29960 50000 30016
rect 47301 29958 50000 29960
rect 47301 29955 47367 29958
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 49200 29928 50000 29958
rect 34928 29887 35248 29888
rect 25037 29882 25103 29885
rect 27981 29882 28047 29885
rect 25037 29880 28047 29882
rect 25037 29824 25042 29880
rect 25098 29824 27986 29880
rect 28042 29824 28047 29880
rect 25037 29822 28047 29824
rect 25037 29819 25103 29822
rect 27981 29819 28047 29822
rect 19977 29746 20043 29749
rect 20989 29746 21055 29749
rect 19977 29744 21055 29746
rect 19977 29688 19982 29744
rect 20038 29688 20994 29744
rect 21050 29688 21055 29744
rect 19977 29686 21055 29688
rect 19977 29683 20043 29686
rect 20989 29683 21055 29686
rect 34789 29746 34855 29749
rect 35525 29746 35591 29749
rect 34789 29744 35591 29746
rect 34789 29688 34794 29744
rect 34850 29688 35530 29744
rect 35586 29688 35591 29744
rect 34789 29686 35591 29688
rect 34789 29683 34855 29686
rect 35525 29683 35591 29686
rect 23381 29474 23447 29477
rect 24853 29474 24919 29477
rect 23381 29472 24919 29474
rect 23381 29416 23386 29472
rect 23442 29416 24858 29472
rect 24914 29416 24919 29472
rect 23381 29414 24919 29416
rect 23381 29411 23447 29414
rect 24853 29411 24919 29414
rect 19568 29408 19888 29409
rect 0 29338 800 29368
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 4061 29338 4127 29341
rect 20345 29340 20411 29341
rect 20294 29338 20300 29340
rect 0 29336 4127 29338
rect 0 29280 4066 29336
rect 4122 29280 4127 29336
rect 0 29278 4127 29280
rect 20218 29278 20300 29338
rect 20364 29338 20411 29340
rect 25865 29338 25931 29341
rect 20364 29336 25931 29338
rect 20406 29280 25870 29336
rect 25926 29280 25931 29336
rect 0 29248 800 29278
rect 4061 29275 4127 29278
rect 20294 29276 20300 29278
rect 20364 29278 25931 29280
rect 20364 29276 20411 29278
rect 20345 29275 20411 29276
rect 25865 29275 25931 29278
rect 34697 29338 34763 29341
rect 35709 29338 35775 29341
rect 34697 29336 35775 29338
rect 34697 29280 34702 29336
rect 34758 29280 35714 29336
rect 35770 29280 35775 29336
rect 34697 29278 35775 29280
rect 34697 29275 34763 29278
rect 35709 29275 35775 29278
rect 48129 29338 48195 29341
rect 49200 29338 50000 29368
rect 48129 29336 50000 29338
rect 48129 29280 48134 29336
rect 48190 29280 50000 29336
rect 48129 29278 50000 29280
rect 48129 29275 48195 29278
rect 49200 29248 50000 29278
rect 9397 29202 9463 29205
rect 17769 29202 17835 29205
rect 9397 29200 17835 29202
rect 9397 29144 9402 29200
rect 9458 29144 17774 29200
rect 17830 29144 17835 29200
rect 9397 29142 17835 29144
rect 9397 29139 9463 29142
rect 17769 29139 17835 29142
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 0 28658 800 28688
rect 2773 28658 2839 28661
rect 0 28656 2839 28658
rect 0 28600 2778 28656
rect 2834 28600 2839 28656
rect 0 28598 2839 28600
rect 0 28568 800 28598
rect 2773 28595 2839 28598
rect 48221 28658 48287 28661
rect 49200 28658 50000 28688
rect 48221 28656 50000 28658
rect 48221 28600 48226 28656
rect 48282 28600 50000 28656
rect 48221 28598 50000 28600
rect 48221 28595 48287 28598
rect 49200 28568 50000 28598
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 19977 28250 20043 28253
rect 20110 28250 20116 28252
rect 19977 28248 20116 28250
rect 19977 28192 19982 28248
rect 20038 28192 20116 28248
rect 19977 28190 20116 28192
rect 19977 28187 20043 28190
rect 20110 28188 20116 28190
rect 20180 28188 20186 28252
rect 0 27888 800 28008
rect 9489 27978 9555 27981
rect 9949 27978 10015 27981
rect 9489 27976 10015 27978
rect 9489 27920 9494 27976
rect 9550 27920 9954 27976
rect 10010 27920 10015 27976
rect 9489 27918 10015 27920
rect 9489 27915 9555 27918
rect 9949 27915 10015 27918
rect 47853 27978 47919 27981
rect 49200 27978 50000 28008
rect 47853 27976 50000 27978
rect 47853 27920 47858 27976
rect 47914 27920 50000 27976
rect 47853 27918 50000 27920
rect 47853 27915 47919 27918
rect 49200 27888 50000 27918
rect 9673 27842 9739 27845
rect 9949 27842 10015 27845
rect 9673 27840 10015 27842
rect 9673 27784 9678 27840
rect 9734 27784 9954 27840
rect 10010 27784 10015 27840
rect 9673 27782 10015 27784
rect 9673 27779 9739 27782
rect 9949 27779 10015 27782
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 0 27298 800 27328
rect 1853 27298 1919 27301
rect 0 27296 1919 27298
rect 0 27240 1858 27296
rect 1914 27240 1919 27296
rect 0 27238 1919 27240
rect 0 27208 800 27238
rect 1853 27235 1919 27238
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 49200 27208 50000 27328
rect 19568 27167 19888 27168
rect 8661 27026 8727 27029
rect 10409 27026 10475 27029
rect 20345 27028 20411 27029
rect 20294 27026 20300 27028
rect 8661 27024 10475 27026
rect 8661 26968 8666 27024
rect 8722 26968 10414 27024
rect 10470 26968 10475 27024
rect 8661 26966 10475 26968
rect 20254 26966 20300 27026
rect 20364 27024 20411 27028
rect 20406 26968 20411 27024
rect 8661 26963 8727 26966
rect 10409 26963 10475 26966
rect 20294 26964 20300 26966
rect 20364 26964 20411 26968
rect 20345 26963 20411 26964
rect 9673 26890 9739 26893
rect 10041 26890 10107 26893
rect 9673 26888 10107 26890
rect 9673 26832 9678 26888
rect 9734 26832 10046 26888
rect 10102 26832 10107 26888
rect 9673 26830 10107 26832
rect 9673 26827 9739 26830
rect 10041 26827 10107 26830
rect 32213 26890 32279 26893
rect 33685 26890 33751 26893
rect 32213 26888 33751 26890
rect 32213 26832 32218 26888
rect 32274 26832 33690 26888
rect 33746 26832 33751 26888
rect 32213 26830 33751 26832
rect 32213 26827 32279 26830
rect 33685 26827 33751 26830
rect 4208 26688 4528 26689
rect 0 26618 800 26648
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 2773 26618 2839 26621
rect 0 26616 2839 26618
rect 0 26560 2778 26616
rect 2834 26560 2839 26616
rect 0 26558 2839 26560
rect 0 26528 800 26558
rect 2773 26555 2839 26558
rect 8845 26618 8911 26621
rect 10593 26618 10659 26621
rect 8845 26616 10659 26618
rect 8845 26560 8850 26616
rect 8906 26560 10598 26616
rect 10654 26560 10659 26616
rect 8845 26558 10659 26560
rect 8845 26555 8911 26558
rect 10593 26555 10659 26558
rect 45461 26618 45527 26621
rect 49200 26618 50000 26648
rect 45461 26616 50000 26618
rect 45461 26560 45466 26616
rect 45522 26560 50000 26616
rect 45461 26558 50000 26560
rect 45461 26555 45527 26558
rect 49200 26528 50000 26558
rect 9213 26482 9279 26485
rect 17585 26482 17651 26485
rect 9213 26480 17651 26482
rect 9213 26424 9218 26480
rect 9274 26424 17590 26480
rect 17646 26424 17651 26480
rect 9213 26422 17651 26424
rect 9213 26419 9279 26422
rect 17585 26419 17651 26422
rect 17677 26346 17743 26349
rect 18137 26346 18203 26349
rect 17677 26344 18203 26346
rect 17677 26288 17682 26344
rect 17738 26288 18142 26344
rect 18198 26288 18203 26344
rect 17677 26286 18203 26288
rect 17677 26283 17743 26286
rect 18137 26283 18203 26286
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 0 25938 800 25968
rect 1577 25938 1643 25941
rect 0 25936 1643 25938
rect 0 25880 1582 25936
rect 1638 25880 1643 25936
rect 0 25878 1643 25880
rect 0 25848 800 25878
rect 1577 25875 1643 25878
rect 47945 25938 48011 25941
rect 49200 25938 50000 25968
rect 47945 25936 50000 25938
rect 47945 25880 47950 25936
rect 48006 25880 50000 25936
rect 47945 25878 50000 25880
rect 47945 25875 48011 25878
rect 49200 25848 50000 25878
rect 24117 25804 24183 25805
rect 24117 25802 24164 25804
rect 24072 25800 24164 25802
rect 24072 25744 24122 25800
rect 24072 25742 24164 25744
rect 24117 25740 24164 25742
rect 24228 25740 24234 25804
rect 24117 25739 24183 25740
rect 20253 25666 20319 25669
rect 25681 25666 25747 25669
rect 20253 25664 25747 25666
rect 20253 25608 20258 25664
rect 20314 25608 25686 25664
rect 25742 25608 25747 25664
rect 20253 25606 25747 25608
rect 20253 25603 20319 25606
rect 25681 25603 25747 25606
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 9949 25530 10015 25533
rect 14549 25530 14615 25533
rect 9949 25528 14615 25530
rect 9949 25472 9954 25528
rect 10010 25472 14554 25528
rect 14610 25472 14615 25528
rect 9949 25470 14615 25472
rect 9949 25467 10015 25470
rect 14549 25467 14615 25470
rect 19977 25530 20043 25533
rect 23749 25530 23815 25533
rect 19977 25528 23815 25530
rect 19977 25472 19982 25528
rect 20038 25472 23754 25528
rect 23810 25472 23815 25528
rect 19977 25470 23815 25472
rect 19977 25467 20043 25470
rect 23749 25467 23815 25470
rect 0 25168 800 25288
rect 17953 25258 18019 25261
rect 21173 25258 21239 25261
rect 17953 25256 21239 25258
rect 17953 25200 17958 25256
rect 18014 25200 21178 25256
rect 21234 25200 21239 25256
rect 17953 25198 21239 25200
rect 17953 25195 18019 25198
rect 21173 25195 21239 25198
rect 47945 25258 48011 25261
rect 49200 25258 50000 25288
rect 47945 25256 50000 25258
rect 47945 25200 47950 25256
rect 48006 25200 50000 25256
rect 47945 25198 50000 25200
rect 47945 25195 48011 25198
rect 49200 25168 50000 25198
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 23105 24988 23171 24989
rect 23054 24986 23060 24988
rect 23014 24926 23060 24986
rect 23124 24984 23171 24988
rect 23166 24928 23171 24984
rect 23054 24924 23060 24926
rect 23124 24924 23171 24928
rect 23105 24923 23171 24924
rect 23841 24986 23907 24989
rect 23974 24986 23980 24988
rect 23841 24984 23980 24986
rect 23841 24928 23846 24984
rect 23902 24928 23980 24984
rect 23841 24926 23980 24928
rect 23841 24923 23907 24926
rect 23974 24924 23980 24926
rect 24044 24924 24050 24988
rect 9121 24850 9187 24853
rect 17401 24850 17467 24853
rect 9121 24848 17467 24850
rect 9121 24792 9126 24848
rect 9182 24792 17406 24848
rect 17462 24792 17467 24848
rect 9121 24790 17467 24792
rect 9121 24787 9187 24790
rect 17401 24787 17467 24790
rect 19885 24850 19951 24853
rect 25129 24850 25195 24853
rect 19885 24848 25195 24850
rect 19885 24792 19890 24848
rect 19946 24792 25134 24848
rect 25190 24792 25195 24848
rect 19885 24790 25195 24792
rect 19885 24787 19951 24790
rect 25129 24787 25195 24790
rect 21817 24714 21883 24717
rect 28625 24714 28691 24717
rect 21817 24712 28691 24714
rect 21817 24656 21822 24712
rect 21878 24656 28630 24712
rect 28686 24656 28691 24712
rect 21817 24654 28691 24656
rect 21817 24651 21883 24654
rect 28625 24651 28691 24654
rect 0 24488 800 24608
rect 48129 24578 48195 24581
rect 49200 24578 50000 24608
rect 48129 24576 50000 24578
rect 48129 24520 48134 24576
rect 48190 24520 50000 24576
rect 48129 24518 50000 24520
rect 48129 24515 48195 24518
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 49200 24488 50000 24518
rect 34928 24447 35248 24448
rect 29361 24442 29427 24445
rect 32673 24442 32739 24445
rect 29361 24440 32739 24442
rect 29361 24384 29366 24440
rect 29422 24384 32678 24440
rect 32734 24384 32739 24440
rect 29361 24382 32739 24384
rect 29361 24379 29427 24382
rect 32673 24379 32739 24382
rect 26325 24306 26391 24309
rect 27613 24306 27679 24309
rect 26325 24304 27679 24306
rect 26325 24248 26330 24304
rect 26386 24248 27618 24304
rect 27674 24248 27679 24304
rect 26325 24246 27679 24248
rect 26325 24243 26391 24246
rect 27613 24243 27679 24246
rect 12249 24170 12315 24173
rect 16849 24170 16915 24173
rect 12249 24168 16915 24170
rect 12249 24112 12254 24168
rect 12310 24112 16854 24168
rect 16910 24112 16915 24168
rect 12249 24110 16915 24112
rect 12249 24107 12315 24110
rect 16849 24107 16915 24110
rect 21909 24170 21975 24173
rect 32397 24170 32463 24173
rect 21909 24168 32463 24170
rect 21909 24112 21914 24168
rect 21970 24112 32402 24168
rect 32458 24112 32463 24168
rect 21909 24110 32463 24112
rect 21909 24107 21975 24110
rect 32397 24107 32463 24110
rect 19568 23968 19888 23969
rect 0 23898 800 23928
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 1393 23898 1459 23901
rect 0 23896 1459 23898
rect 0 23840 1398 23896
rect 1454 23840 1459 23896
rect 0 23838 1459 23840
rect 0 23808 800 23838
rect 1393 23835 1459 23838
rect 28993 23898 29059 23901
rect 32305 23898 32371 23901
rect 28993 23896 32371 23898
rect 28993 23840 28998 23896
rect 29054 23840 32310 23896
rect 32366 23840 32371 23896
rect 28993 23838 32371 23840
rect 28993 23835 29059 23838
rect 32305 23835 32371 23838
rect 47301 23898 47367 23901
rect 49200 23898 50000 23928
rect 47301 23896 50000 23898
rect 47301 23840 47306 23896
rect 47362 23840 50000 23896
rect 47301 23838 50000 23840
rect 47301 23835 47367 23838
rect 49200 23808 50000 23838
rect 23381 23490 23447 23493
rect 24669 23490 24735 23493
rect 23381 23488 24735 23490
rect 23381 23432 23386 23488
rect 23442 23432 24674 23488
rect 24730 23432 24735 23488
rect 23381 23430 24735 23432
rect 23381 23427 23447 23430
rect 24669 23427 24735 23430
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 0 23218 800 23248
rect 2773 23218 2839 23221
rect 0 23216 2839 23218
rect 0 23160 2778 23216
rect 2834 23160 2839 23216
rect 0 23158 2839 23160
rect 0 23128 800 23158
rect 2773 23155 2839 23158
rect 49200 23128 50000 23248
rect 8385 23082 8451 23085
rect 9857 23082 9923 23085
rect 8385 23080 9923 23082
rect 8385 23024 8390 23080
rect 8446 23024 9862 23080
rect 9918 23024 9923 23080
rect 8385 23022 9923 23024
rect 8385 23019 8451 23022
rect 9857 23019 9923 23022
rect 20110 23020 20116 23084
rect 20180 23082 20186 23084
rect 20253 23082 20319 23085
rect 20180 23080 20319 23082
rect 20180 23024 20258 23080
rect 20314 23024 20319 23080
rect 20180 23022 20319 23024
rect 20180 23020 20186 23022
rect 20253 23019 20319 23022
rect 28993 23082 29059 23085
rect 30189 23082 30255 23085
rect 28993 23080 30255 23082
rect 28993 23024 28998 23080
rect 29054 23024 30194 23080
rect 30250 23024 30255 23080
rect 28993 23022 30255 23024
rect 28993 23019 29059 23022
rect 30189 23019 30255 23022
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 12341 22674 12407 22677
rect 14549 22674 14615 22677
rect 15009 22674 15075 22677
rect 16205 22674 16271 22677
rect 12341 22672 16271 22674
rect 12341 22616 12346 22672
rect 12402 22616 14554 22672
rect 14610 22616 15014 22672
rect 15070 22616 16210 22672
rect 16266 22616 16271 22672
rect 12341 22614 16271 22616
rect 12341 22611 12407 22614
rect 14549 22611 14615 22614
rect 15009 22611 15075 22614
rect 16205 22611 16271 22614
rect 19517 22674 19583 22677
rect 25497 22674 25563 22677
rect 26141 22674 26207 22677
rect 19517 22672 26207 22674
rect 19517 22616 19522 22672
rect 19578 22616 25502 22672
rect 25558 22616 26146 22672
rect 26202 22616 26207 22672
rect 19517 22614 26207 22616
rect 19517 22611 19583 22614
rect 25497 22611 25563 22614
rect 26141 22611 26207 22614
rect 0 22538 800 22568
rect 1393 22538 1459 22541
rect 0 22536 1459 22538
rect 0 22480 1398 22536
rect 1454 22480 1459 22536
rect 0 22478 1459 22480
rect 0 22448 800 22478
rect 1393 22475 1459 22478
rect 48129 22538 48195 22541
rect 49200 22538 50000 22568
rect 48129 22536 50000 22538
rect 48129 22480 48134 22536
rect 48190 22480 50000 22536
rect 48129 22478 50000 22480
rect 48129 22475 48195 22478
rect 49200 22448 50000 22478
rect 24117 22404 24183 22405
rect 24117 22400 24164 22404
rect 24228 22402 24234 22404
rect 24117 22344 24122 22400
rect 24117 22340 24164 22344
rect 24228 22342 24274 22402
rect 24228 22340 24234 22342
rect 24117 22339 24183 22340
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 19793 22266 19859 22269
rect 20294 22266 20300 22268
rect 19793 22264 20300 22266
rect 19793 22208 19798 22264
rect 19854 22208 20300 22264
rect 19793 22206 20300 22208
rect 19793 22203 19859 22206
rect 20294 22204 20300 22206
rect 20364 22204 20370 22268
rect 30649 22130 30715 22133
rect 31569 22130 31635 22133
rect 30649 22128 31635 22130
rect 30649 22072 30654 22128
rect 30710 22072 31574 22128
rect 31630 22072 31635 22128
rect 30649 22070 31635 22072
rect 30649 22067 30715 22070
rect 31569 22067 31635 22070
rect 30373 21994 30439 21997
rect 32029 21994 32095 21997
rect 30373 21992 32095 21994
rect 30373 21936 30378 21992
rect 30434 21936 32034 21992
rect 32090 21936 32095 21992
rect 30373 21934 32095 21936
rect 30373 21931 30439 21934
rect 32029 21931 32095 21934
rect 0 21858 800 21888
rect 3969 21858 4035 21861
rect 0 21856 4035 21858
rect 0 21800 3974 21856
rect 4030 21800 4035 21856
rect 0 21798 4035 21800
rect 0 21768 800 21798
rect 3969 21795 4035 21798
rect 47945 21858 48011 21861
rect 49200 21858 50000 21888
rect 47945 21856 50000 21858
rect 47945 21800 47950 21856
rect 48006 21800 50000 21856
rect 47945 21798 50000 21800
rect 47945 21795 48011 21798
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 49200 21768 50000 21798
rect 19568 21727 19888 21728
rect 22093 21314 22159 21317
rect 25681 21314 25747 21317
rect 22093 21312 25747 21314
rect 22093 21256 22098 21312
rect 22154 21256 25686 21312
rect 25742 21256 25747 21312
rect 22093 21254 25747 21256
rect 22093 21251 22159 21254
rect 25681 21251 25747 21254
rect 4208 21248 4528 21249
rect 0 21178 800 21208
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 4061 21178 4127 21181
rect 0 21176 4127 21178
rect 0 21120 4066 21176
rect 4122 21120 4127 21176
rect 0 21118 4127 21120
rect 0 21088 800 21118
rect 4061 21115 4127 21118
rect 49200 21088 50000 21208
rect 23749 20906 23815 20909
rect 23614 20904 23815 20906
rect 23614 20848 23754 20904
rect 23810 20848 23815 20904
rect 23614 20846 23815 20848
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 0 20408 800 20528
rect 23614 20365 23674 20846
rect 23749 20843 23815 20846
rect 24117 20770 24183 20773
rect 24945 20770 25011 20773
rect 24117 20768 25011 20770
rect 24117 20712 24122 20768
rect 24178 20712 24950 20768
rect 25006 20712 25011 20768
rect 24117 20710 25011 20712
rect 24117 20707 24183 20710
rect 24945 20707 25011 20710
rect 49200 20408 50000 20528
rect 23614 20360 23723 20365
rect 23614 20304 23662 20360
rect 23718 20304 23723 20360
rect 23614 20302 23723 20304
rect 23657 20299 23723 20302
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 0 19818 800 19848
rect 4061 19818 4127 19821
rect 20621 19818 20687 19821
rect 0 19816 4127 19818
rect 0 19760 4066 19816
rect 4122 19760 4127 19816
rect 0 19758 4127 19760
rect 0 19728 800 19758
rect 4061 19755 4127 19758
rect 20348 19816 20687 19818
rect 20348 19760 20626 19816
rect 20682 19760 20687 19816
rect 20348 19758 20687 19760
rect 20348 19685 20408 19758
rect 20621 19755 20687 19758
rect 48129 19818 48195 19821
rect 49200 19818 50000 19848
rect 48129 19816 50000 19818
rect 48129 19760 48134 19816
rect 48190 19760 50000 19816
rect 48129 19758 50000 19760
rect 48129 19755 48195 19758
rect 49200 19728 50000 19758
rect 20345 19680 20411 19685
rect 20345 19624 20350 19680
rect 20406 19624 20411 19680
rect 20345 19619 20411 19624
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 19885 19410 19951 19413
rect 22093 19410 22159 19413
rect 19885 19408 22159 19410
rect 19885 19352 19890 19408
rect 19946 19352 22098 19408
rect 22154 19352 22159 19408
rect 19885 19350 22159 19352
rect 19885 19347 19951 19350
rect 22093 19347 22159 19350
rect 0 19138 800 19168
rect 2773 19138 2839 19141
rect 0 19136 2839 19138
rect 0 19080 2778 19136
rect 2834 19080 2839 19136
rect 0 19078 2839 19080
rect 0 19048 800 19078
rect 2773 19075 2839 19078
rect 47945 19138 48011 19141
rect 49200 19138 50000 19168
rect 47945 19136 50000 19138
rect 47945 19080 47950 19136
rect 48006 19080 50000 19136
rect 47945 19078 50000 19080
rect 47945 19075 48011 19078
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 49200 19048 50000 19078
rect 34928 19007 35248 19008
rect 19885 18730 19951 18733
rect 20110 18730 20116 18732
rect 19885 18728 20116 18730
rect 19885 18672 19890 18728
rect 19946 18672 20116 18728
rect 19885 18670 20116 18672
rect 19885 18667 19951 18670
rect 20110 18668 20116 18670
rect 20180 18668 20186 18732
rect 19568 18528 19888 18529
rect 0 18458 800 18488
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 4061 18458 4127 18461
rect 0 18456 4127 18458
rect 0 18400 4066 18456
rect 4122 18400 4127 18456
rect 0 18398 4127 18400
rect 0 18368 800 18398
rect 4061 18395 4127 18398
rect 49200 18368 50000 18488
rect 14917 18186 14983 18189
rect 17401 18186 17467 18189
rect 14917 18184 17467 18186
rect 14917 18128 14922 18184
rect 14978 18128 17406 18184
rect 17462 18128 17467 18184
rect 14917 18126 17467 18128
rect 14917 18123 14983 18126
rect 17401 18123 17467 18126
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 14641 17914 14707 17917
rect 18413 17914 18479 17917
rect 14641 17912 18479 17914
rect 14641 17856 14646 17912
rect 14702 17856 18418 17912
rect 18474 17856 18479 17912
rect 14641 17854 18479 17856
rect 14641 17851 14707 17854
rect 18413 17851 18479 17854
rect 0 17778 800 17808
rect 2773 17778 2839 17781
rect 0 17776 2839 17778
rect 0 17720 2778 17776
rect 2834 17720 2839 17776
rect 0 17718 2839 17720
rect 0 17688 800 17718
rect 2773 17715 2839 17718
rect 21081 17778 21147 17781
rect 22277 17778 22343 17781
rect 21081 17776 22343 17778
rect 21081 17720 21086 17776
rect 21142 17720 22282 17776
rect 22338 17720 22343 17776
rect 21081 17718 22343 17720
rect 21081 17715 21147 17718
rect 22277 17715 22343 17718
rect 46381 17778 46447 17781
rect 49200 17778 50000 17808
rect 46381 17776 50000 17778
rect 46381 17720 46386 17776
rect 46442 17720 50000 17776
rect 46381 17718 50000 17720
rect 46381 17715 46447 17718
rect 49200 17688 50000 17718
rect 15377 17642 15443 17645
rect 16941 17642 17007 17645
rect 15377 17640 17007 17642
rect 15377 17584 15382 17640
rect 15438 17584 16946 17640
rect 17002 17584 17007 17640
rect 15377 17582 17007 17584
rect 15377 17579 15443 17582
rect 16941 17579 17007 17582
rect 24117 17642 24183 17645
rect 27613 17642 27679 17645
rect 24117 17640 27679 17642
rect 24117 17584 24122 17640
rect 24178 17584 27618 17640
rect 27674 17584 27679 17640
rect 24117 17582 27679 17584
rect 24117 17579 24183 17582
rect 27613 17579 27679 17582
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 10409 17370 10475 17373
rect 16021 17370 16087 17373
rect 10409 17368 16087 17370
rect 10409 17312 10414 17368
rect 10470 17312 16026 17368
rect 16082 17312 16087 17368
rect 10409 17310 16087 17312
rect 10409 17307 10475 17310
rect 16021 17307 16087 17310
rect 20345 17370 20411 17373
rect 20345 17368 20546 17370
rect 20345 17312 20350 17368
rect 20406 17312 20546 17368
rect 20345 17310 20546 17312
rect 20345 17307 20411 17310
rect 0 17098 800 17128
rect 1853 17098 1919 17101
rect 0 17096 1919 17098
rect 0 17040 1858 17096
rect 1914 17040 1919 17096
rect 0 17038 1919 17040
rect 0 17008 800 17038
rect 1853 17035 1919 17038
rect 20486 16962 20546 17310
rect 24117 17234 24183 17237
rect 24761 17234 24827 17237
rect 24117 17232 24827 17234
rect 24117 17176 24122 17232
rect 24178 17176 24766 17232
rect 24822 17176 24827 17232
rect 24117 17174 24827 17176
rect 24117 17171 24183 17174
rect 24761 17171 24827 17174
rect 48129 17098 48195 17101
rect 49200 17098 50000 17128
rect 48129 17096 50000 17098
rect 48129 17040 48134 17096
rect 48190 17040 50000 17096
rect 48129 17038 50000 17040
rect 48129 17035 48195 17038
rect 49200 17008 50000 17038
rect 20621 16962 20687 16965
rect 20486 16960 20687 16962
rect 20486 16904 20626 16960
rect 20682 16904 20687 16960
rect 20486 16902 20687 16904
rect 20621 16899 20687 16902
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 0 16418 800 16448
rect 2773 16418 2839 16421
rect 0 16416 2839 16418
rect 0 16360 2778 16416
rect 2834 16360 2839 16416
rect 0 16358 2839 16360
rect 0 16328 800 16358
rect 2773 16355 2839 16358
rect 48129 16418 48195 16421
rect 49200 16418 50000 16448
rect 48129 16416 50000 16418
rect 48129 16360 48134 16416
rect 48190 16360 50000 16416
rect 48129 16358 50000 16360
rect 48129 16355 48195 16358
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 49200 16328 50000 16358
rect 19568 16287 19888 16288
rect 27153 16282 27219 16285
rect 30373 16282 30439 16285
rect 27153 16280 30439 16282
rect 27153 16224 27158 16280
rect 27214 16224 30378 16280
rect 30434 16224 30439 16280
rect 27153 16222 30439 16224
rect 27153 16219 27219 16222
rect 30373 16219 30439 16222
rect 4208 15808 4528 15809
rect 0 15648 800 15768
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 49200 15648 50000 15768
rect 19425 15466 19491 15469
rect 19382 15464 19491 15466
rect 19382 15408 19430 15464
rect 19486 15408 19491 15464
rect 19382 15403 19491 15408
rect 0 14968 800 15088
rect 19382 15058 19442 15403
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 19609 15058 19675 15061
rect 19382 15056 19675 15058
rect 19382 15000 19614 15056
rect 19670 15000 19675 15056
rect 19382 14998 19675 15000
rect 19609 14995 19675 14998
rect 46841 15058 46907 15061
rect 49200 15058 50000 15088
rect 46841 15056 50000 15058
rect 46841 15000 46846 15056
rect 46902 15000 50000 15056
rect 46841 14998 50000 15000
rect 46841 14995 46907 14998
rect 49200 14968 50000 14998
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 0 14288 800 14408
rect 19609 14378 19675 14381
rect 20161 14378 20227 14381
rect 19609 14376 20227 14378
rect 19609 14320 19614 14376
rect 19670 14320 20166 14376
rect 20222 14320 20227 14376
rect 19609 14318 20227 14320
rect 19609 14315 19675 14318
rect 20161 14315 20227 14318
rect 25037 14378 25103 14381
rect 26969 14378 27035 14381
rect 28349 14378 28415 14381
rect 25037 14376 28415 14378
rect 25037 14320 25042 14376
rect 25098 14320 26974 14376
rect 27030 14320 28354 14376
rect 28410 14320 28415 14376
rect 25037 14318 28415 14320
rect 25037 14315 25103 14318
rect 26969 14315 27035 14318
rect 28349 14315 28415 14318
rect 48129 14378 48195 14381
rect 49200 14378 50000 14408
rect 48129 14376 50000 14378
rect 48129 14320 48134 14376
rect 48190 14320 50000 14376
rect 48129 14318 50000 14320
rect 48129 14315 48195 14318
rect 49200 14288 50000 14318
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 0 13698 800 13728
rect 2773 13698 2839 13701
rect 0 13696 2839 13698
rect 0 13640 2778 13696
rect 2834 13640 2839 13696
rect 0 13638 2839 13640
rect 0 13608 800 13638
rect 2773 13635 2839 13638
rect 47853 13698 47919 13701
rect 49200 13698 50000 13728
rect 47853 13696 50000 13698
rect 47853 13640 47858 13696
rect 47914 13640 50000 13696
rect 47853 13638 50000 13640
rect 47853 13635 47919 13638
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 49200 13608 50000 13638
rect 34928 13567 35248 13568
rect 21817 13426 21883 13429
rect 26233 13426 26299 13429
rect 21817 13424 26299 13426
rect 21817 13368 21822 13424
rect 21878 13368 26238 13424
rect 26294 13368 26299 13424
rect 21817 13366 26299 13368
rect 21817 13363 21883 13366
rect 26233 13363 26299 13366
rect 19568 13088 19888 13089
rect 0 13018 800 13048
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 4061 13018 4127 13021
rect 0 13016 4127 13018
rect 0 12960 4066 13016
rect 4122 12960 4127 13016
rect 0 12958 4127 12960
rect 0 12928 800 12958
rect 4061 12955 4127 12958
rect 46841 13018 46907 13021
rect 49200 13018 50000 13048
rect 46841 13016 50000 13018
rect 46841 12960 46846 13016
rect 46902 12960 50000 13016
rect 46841 12958 50000 12960
rect 46841 12955 46907 12958
rect 49200 12928 50000 12958
rect 20069 12748 20135 12749
rect 20069 12744 20116 12748
rect 20180 12746 20186 12748
rect 20069 12688 20074 12744
rect 20069 12684 20116 12688
rect 20180 12686 20226 12746
rect 20180 12684 20186 12686
rect 20069 12683 20135 12684
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 0 12338 800 12368
rect 1393 12338 1459 12341
rect 0 12336 1459 12338
rect 0 12280 1398 12336
rect 1454 12280 1459 12336
rect 0 12278 1459 12280
rect 0 12248 800 12278
rect 1393 12275 1459 12278
rect 46841 12338 46907 12341
rect 49200 12338 50000 12368
rect 46841 12336 50000 12338
rect 46841 12280 46846 12336
rect 46902 12280 50000 12336
rect 46841 12278 50000 12280
rect 46841 12275 46907 12278
rect 49200 12248 50000 12278
rect 19333 12204 19399 12205
rect 19333 12200 19380 12204
rect 19444 12202 19450 12204
rect 19333 12144 19338 12200
rect 19333 12140 19380 12144
rect 19444 12142 19490 12202
rect 19444 12140 19450 12142
rect 19333 12139 19399 12140
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 27889 11930 27955 11933
rect 28073 11930 28139 11933
rect 27889 11928 28139 11930
rect 27889 11872 27894 11928
rect 27950 11872 28078 11928
rect 28134 11872 28139 11928
rect 27889 11870 28139 11872
rect 27889 11867 27955 11870
rect 28073 11867 28139 11870
rect 19885 11794 19951 11797
rect 26601 11794 26667 11797
rect 19885 11792 26667 11794
rect 19885 11736 19890 11792
rect 19946 11736 26606 11792
rect 26662 11736 26667 11792
rect 19885 11734 26667 11736
rect 19885 11731 19951 11734
rect 26601 11731 26667 11734
rect 0 11568 800 11688
rect 20529 11658 20595 11661
rect 21265 11658 21331 11661
rect 28073 11658 28139 11661
rect 20529 11656 28139 11658
rect 20529 11600 20534 11656
rect 20590 11600 21270 11656
rect 21326 11600 28078 11656
rect 28134 11600 28139 11656
rect 20529 11598 28139 11600
rect 20529 11595 20595 11598
rect 21265 11595 21331 11598
rect 28073 11595 28139 11598
rect 49200 11568 50000 11688
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 0 10978 800 11008
rect 1853 10978 1919 10981
rect 0 10976 1919 10978
rect 0 10920 1858 10976
rect 1914 10920 1919 10976
rect 0 10918 1919 10920
rect 0 10888 800 10918
rect 1853 10915 1919 10918
rect 48129 10978 48195 10981
rect 49200 10978 50000 11008
rect 48129 10976 50000 10978
rect 48129 10920 48134 10976
rect 48190 10920 50000 10976
rect 48129 10918 50000 10920
rect 48129 10915 48195 10918
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 49200 10888 50000 10918
rect 19568 10847 19888 10848
rect 20345 10434 20411 10437
rect 20118 10432 20411 10434
rect 20118 10376 20350 10432
rect 20406 10376 20411 10432
rect 20118 10374 20411 10376
rect 4208 10368 4528 10369
rect 0 10298 800 10328
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 2865 10298 2931 10301
rect 0 10296 2931 10298
rect 0 10240 2870 10296
rect 2926 10240 2931 10296
rect 0 10238 2931 10240
rect 0 10208 800 10238
rect 2865 10235 2931 10238
rect 20118 10029 20178 10374
rect 20345 10371 20411 10374
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 47761 10298 47827 10301
rect 49200 10298 50000 10328
rect 47761 10296 50000 10298
rect 47761 10240 47766 10296
rect 47822 10240 50000 10296
rect 47761 10238 50000 10240
rect 47761 10235 47827 10238
rect 49200 10208 50000 10238
rect 20069 10024 20178 10029
rect 20069 9968 20074 10024
rect 20130 9968 20178 10024
rect 20069 9966 20178 9968
rect 20069 9963 20135 9966
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 23054 9692 23060 9756
rect 23124 9754 23130 9756
rect 24117 9754 24183 9757
rect 23124 9752 24183 9754
rect 23124 9696 24122 9752
rect 24178 9696 24183 9752
rect 23124 9694 24183 9696
rect 23124 9692 23130 9694
rect 24117 9691 24183 9694
rect 0 9618 800 9648
rect 2957 9618 3023 9621
rect 0 9616 3023 9618
rect 0 9560 2962 9616
rect 3018 9560 3023 9616
rect 0 9558 3023 9560
rect 0 9528 800 9558
rect 2957 9555 3023 9558
rect 19333 9618 19399 9621
rect 19609 9618 19675 9621
rect 19333 9616 19675 9618
rect 19333 9560 19338 9616
rect 19394 9560 19614 9616
rect 19670 9560 19675 9616
rect 19333 9558 19675 9560
rect 19333 9555 19399 9558
rect 19609 9555 19675 9558
rect 46841 9618 46907 9621
rect 49200 9618 50000 9648
rect 46841 9616 50000 9618
rect 46841 9560 46846 9616
rect 46902 9560 50000 9616
rect 46841 9558 50000 9560
rect 46841 9555 46907 9558
rect 49200 9528 50000 9558
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 0 8938 800 8968
rect 4061 8938 4127 8941
rect 0 8936 4127 8938
rect 0 8880 4066 8936
rect 4122 8880 4127 8936
rect 0 8878 4127 8880
rect 0 8848 800 8878
rect 4061 8875 4127 8878
rect 47945 8938 48011 8941
rect 49200 8938 50000 8968
rect 47945 8936 50000 8938
rect 47945 8880 47950 8936
rect 48006 8880 50000 8936
rect 47945 8878 50000 8880
rect 47945 8875 48011 8878
rect 49200 8848 50000 8878
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 0 8258 800 8288
rect 1853 8258 1919 8261
rect 0 8256 1919 8258
rect 0 8200 1858 8256
rect 1914 8200 1919 8256
rect 0 8198 1919 8200
rect 0 8168 800 8198
rect 1853 8195 1919 8198
rect 47761 8258 47827 8261
rect 49200 8258 50000 8288
rect 47761 8256 50000 8258
rect 47761 8200 47766 8256
rect 47822 8200 50000 8256
rect 47761 8198 50000 8200
rect 47761 8195 47827 8198
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 49200 8168 50000 8198
rect 34928 8127 35248 8128
rect 23381 7986 23447 7989
rect 25313 7986 25379 7989
rect 23381 7984 25379 7986
rect 23381 7928 23386 7984
rect 23442 7928 25318 7984
rect 25374 7928 25379 7984
rect 23381 7926 25379 7928
rect 23381 7923 23447 7926
rect 25313 7923 25379 7926
rect 23289 7850 23355 7853
rect 25037 7850 25103 7853
rect 27245 7850 27311 7853
rect 23289 7848 27311 7850
rect 23289 7792 23294 7848
rect 23350 7792 25042 7848
rect 25098 7792 27250 7848
rect 27306 7792 27311 7848
rect 23289 7790 27311 7792
rect 23289 7787 23355 7790
rect 25037 7787 25103 7790
rect 27245 7787 27311 7790
rect 19568 7648 19888 7649
rect 0 7578 800 7608
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 1393 7578 1459 7581
rect 0 7576 1459 7578
rect 0 7520 1398 7576
rect 1454 7520 1459 7576
rect 0 7518 1459 7520
rect 0 7488 800 7518
rect 1393 7515 1459 7518
rect 48129 7578 48195 7581
rect 49200 7578 50000 7608
rect 48129 7576 50000 7578
rect 48129 7520 48134 7576
rect 48190 7520 50000 7576
rect 48129 7518 50000 7520
rect 48129 7515 48195 7518
rect 49200 7488 50000 7518
rect 19425 7444 19491 7445
rect 19374 7380 19380 7444
rect 19444 7442 19491 7444
rect 19444 7440 19536 7442
rect 19486 7384 19536 7440
rect 19444 7382 19536 7384
rect 19444 7380 19491 7382
rect 19425 7379 19491 7380
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 0 6898 800 6928
rect 2773 6898 2839 6901
rect 49200 6898 50000 6928
rect 0 6896 2839 6898
rect 0 6840 2778 6896
rect 2834 6840 2839 6896
rect 0 6838 2839 6840
rect 0 6808 800 6838
rect 2773 6835 2839 6838
rect 45510 6838 50000 6898
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 0 6218 800 6248
rect 3601 6218 3667 6221
rect 0 6216 3667 6218
rect 0 6160 3606 6216
rect 3662 6160 3667 6216
rect 0 6158 3667 6160
rect 0 6128 800 6158
rect 3601 6155 3667 6158
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 21214 5748 21220 5812
rect 21284 5810 21290 5812
rect 45510 5810 45570 6838
rect 49200 6808 50000 6838
rect 47669 6218 47735 6221
rect 49200 6218 50000 6248
rect 47669 6216 50000 6218
rect 47669 6160 47674 6216
rect 47730 6160 50000 6216
rect 47669 6158 50000 6160
rect 47669 6155 47735 6158
rect 49200 6128 50000 6158
rect 21284 5750 45570 5810
rect 21284 5748 21290 5750
rect 0 5538 800 5568
rect 2773 5538 2839 5541
rect 0 5536 2839 5538
rect 0 5480 2778 5536
rect 2834 5480 2839 5536
rect 0 5478 2839 5480
rect 0 5448 800 5478
rect 2773 5475 2839 5478
rect 47945 5538 48011 5541
rect 49200 5538 50000 5568
rect 47945 5536 50000 5538
rect 47945 5480 47950 5536
rect 48006 5480 50000 5536
rect 47945 5478 50000 5480
rect 47945 5475 48011 5478
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 49200 5448 50000 5478
rect 19568 5407 19888 5408
rect 4208 4928 4528 4929
rect 0 4858 800 4888
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 2773 4858 2839 4861
rect 0 4856 2839 4858
rect 0 4800 2778 4856
rect 2834 4800 2839 4856
rect 0 4798 2839 4800
rect 0 4768 800 4798
rect 2773 4795 2839 4798
rect 48129 4858 48195 4861
rect 49200 4858 50000 4888
rect 48129 4856 50000 4858
rect 48129 4800 48134 4856
rect 48190 4800 50000 4856
rect 48129 4798 50000 4800
rect 48129 4795 48195 4798
rect 49200 4768 50000 4798
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 0 4178 800 4208
rect 3693 4178 3759 4181
rect 0 4176 3759 4178
rect 0 4120 3698 4176
rect 3754 4120 3759 4176
rect 0 4118 3759 4120
rect 0 4088 800 4118
rect 3693 4115 3759 4118
rect 46749 4178 46815 4181
rect 49200 4178 50000 4208
rect 46749 4176 50000 4178
rect 46749 4120 46754 4176
rect 46810 4120 50000 4176
rect 46749 4118 50000 4120
rect 46749 4115 46815 4118
rect 49200 4088 50000 4118
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 20345 3634 20411 3637
rect 26233 3634 26299 3637
rect 20345 3632 26299 3634
rect 20345 3576 20350 3632
rect 20406 3576 26238 3632
rect 26294 3576 26299 3632
rect 20345 3574 26299 3576
rect 20345 3571 20411 3574
rect 26233 3571 26299 3574
rect 0 3498 800 3528
rect 1853 3498 1919 3501
rect 0 3496 1919 3498
rect 0 3440 1858 3496
rect 1914 3440 1919 3496
rect 0 3438 1919 3440
rect 0 3408 800 3438
rect 1853 3435 1919 3438
rect 19885 3498 19951 3501
rect 27981 3498 28047 3501
rect 19885 3496 28047 3498
rect 19885 3440 19890 3496
rect 19946 3440 27986 3496
rect 28042 3440 28047 3496
rect 19885 3438 28047 3440
rect 19885 3435 19951 3438
rect 27981 3435 28047 3438
rect 46841 3498 46907 3501
rect 49200 3498 50000 3528
rect 46841 3496 50000 3498
rect 46841 3440 46846 3496
rect 46902 3440 50000 3496
rect 46841 3438 50000 3440
rect 46841 3435 46907 3438
rect 49200 3408 50000 3438
rect 39021 3362 39087 3365
rect 46565 3362 46631 3365
rect 39021 3360 46631 3362
rect 39021 3304 39026 3360
rect 39082 3304 46570 3360
rect 46626 3304 46631 3360
rect 39021 3302 46631 3304
rect 39021 3299 39087 3302
rect 46565 3299 46631 3302
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 0 2728 800 2848
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 49200 2728 50000 2848
rect 34928 2687 35248 2688
rect 14733 2546 14799 2549
rect 23974 2546 23980 2548
rect 14733 2544 23980 2546
rect 14733 2488 14738 2544
rect 14794 2488 23980 2544
rect 14733 2486 23980 2488
rect 14733 2483 14799 2486
rect 23974 2484 23980 2486
rect 24044 2484 24050 2548
rect 4797 2410 4863 2413
rect 24158 2410 24164 2412
rect 4797 2408 24164 2410
rect 4797 2352 4802 2408
rect 4858 2352 24164 2408
rect 4797 2350 24164 2352
rect 4797 2347 4863 2350
rect 24158 2348 24164 2350
rect 24228 2348 24234 2412
rect 19568 2208 19888 2209
rect 0 2138 800 2168
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 3417 2138 3483 2141
rect 0 2136 3483 2138
rect 0 2080 3422 2136
rect 3478 2080 3483 2136
rect 0 2078 3483 2080
rect 0 2048 800 2078
rect 3417 2075 3483 2078
rect 49200 2048 50000 2168
rect 0 1368 800 1488
rect 46841 1458 46907 1461
rect 49200 1458 50000 1488
rect 46841 1456 50000 1458
rect 46841 1400 46846 1456
rect 46902 1400 50000 1456
rect 46841 1398 50000 1400
rect 46841 1395 46907 1398
rect 49200 1368 50000 1398
rect 0 778 800 808
rect 2773 778 2839 781
rect 0 776 2839 778
rect 0 720 2778 776
rect 2834 720 2839 776
rect 0 718 2839 720
rect 0 688 800 718
rect 2773 715 2839 718
rect 47761 778 47827 781
rect 49200 778 50000 808
rect 47761 776 50000 778
rect 47761 720 47766 776
rect 47822 720 50000 776
rect 47761 718 50000 720
rect 47761 715 47827 718
rect 49200 688 50000 718
rect 46749 98 46815 101
rect 49200 98 50000 128
rect 46749 96 50000 98
rect 46749 40 46754 96
rect 46810 40 50000 96
rect 46749 38 50000 40
rect 46749 35 46815 38
rect 49200 8 50000 38
<< via3 >>
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 24164 38660 24228 38724
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 20300 37088 20364 37092
rect 20300 37032 20350 37088
rect 20350 37032 20364 37088
rect 20300 37028 20364 37032
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 21220 30364 21284 30428
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 20300 29336 20364 29340
rect 20300 29280 20350 29336
rect 20350 29280 20364 29336
rect 20300 29276 20364 29280
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 20116 28188 20180 28252
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 20300 27024 20364 27028
rect 20300 26968 20350 27024
rect 20350 26968 20364 27024
rect 20300 26964 20364 26968
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 24164 25800 24228 25804
rect 24164 25744 24178 25800
rect 24178 25744 24228 25800
rect 24164 25740 24228 25744
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 23060 24984 23124 24988
rect 23060 24928 23110 24984
rect 23110 24928 23124 24984
rect 23060 24924 23124 24928
rect 23980 24924 24044 24988
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 20116 23020 20180 23084
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 24164 22400 24228 22404
rect 24164 22344 24178 22400
rect 24178 22344 24228 22400
rect 24164 22340 24228 22344
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 20300 22204 20364 22268
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 20116 18668 20180 18732
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 20116 12744 20180 12748
rect 20116 12688 20130 12744
rect 20130 12688 20180 12744
rect 20116 12684 20180 12688
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19380 12200 19444 12204
rect 19380 12144 19394 12200
rect 19394 12144 19444 12200
rect 19380 12140 19444 12144
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 23060 9692 23124 9756
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 19380 7440 19444 7444
rect 19380 7384 19430 7440
rect 19430 7384 19444 7440
rect 19380 7380 19444 7384
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 21220 5748 21284 5812
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 23980 2484 24044 2548
rect 24164 2348 24228 2412
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 49536 4528 49552
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 19568 48992 19888 49552
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 34928 49536 35248 49552
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 24163 38724 24229 38725
rect 24163 38660 24164 38724
rect 24228 38660 24229 38724
rect 24163 38659 24229 38660
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 20299 37092 20365 37093
rect 20299 37028 20300 37092
rect 20364 37028 20365 37092
rect 20299 37027 20365 37028
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 20302 29341 20362 37027
rect 21219 30428 21285 30429
rect 21219 30364 21220 30428
rect 21284 30364 21285 30428
rect 21219 30363 21285 30364
rect 20299 29340 20365 29341
rect 20299 29276 20300 29340
rect 20364 29276 20365 29340
rect 20299 29275 20365 29276
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 20115 28252 20181 28253
rect 20115 28188 20116 28252
rect 20180 28188 20181 28252
rect 20115 28187 20181 28188
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 20118 23085 20178 28187
rect 20299 27028 20365 27029
rect 20299 26964 20300 27028
rect 20364 26964 20365 27028
rect 20299 26963 20365 26964
rect 20115 23084 20181 23085
rect 20115 23020 20116 23084
rect 20180 23020 20181 23084
rect 20115 23019 20181 23020
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 20302 22269 20362 26963
rect 20299 22268 20365 22269
rect 20299 22204 20300 22268
rect 20364 22204 20365 22268
rect 20299 22203 20365 22204
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 20115 18732 20181 18733
rect 20115 18668 20116 18732
rect 20180 18668 20181 18732
rect 20115 18667 20181 18668
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19379 12204 19445 12205
rect 19379 12140 19380 12204
rect 19444 12140 19445 12204
rect 19379 12139 19445 12140
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 19382 7445 19442 12139
rect 19568 12000 19888 13024
rect 20118 12749 20178 18667
rect 20115 12748 20181 12749
rect 20115 12684 20116 12748
rect 20180 12684 20181 12748
rect 20115 12683 20181 12684
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19379 7444 19445 7445
rect 19379 7380 19380 7444
rect 19444 7380 19445 7444
rect 19379 7379 19445 7380
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 21222 5813 21282 30363
rect 24166 25805 24226 38659
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 24163 25804 24229 25805
rect 24163 25740 24164 25804
rect 24228 25740 24229 25804
rect 24163 25739 24229 25740
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 23059 24988 23125 24989
rect 23059 24924 23060 24988
rect 23124 24924 23125 24988
rect 23059 24923 23125 24924
rect 23979 24988 24045 24989
rect 23979 24924 23980 24988
rect 24044 24924 24045 24988
rect 23979 24923 24045 24924
rect 23062 9757 23122 24923
rect 23059 9756 23125 9757
rect 23059 9692 23060 9756
rect 23124 9692 23125 9756
rect 23059 9691 23125 9692
rect 21219 5812 21285 5813
rect 21219 5748 21220 5812
rect 21284 5748 21285 5812
rect 21219 5747 21285 5748
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 23982 2549 24042 24923
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 24163 22404 24229 22405
rect 24163 22340 24164 22404
rect 24228 22340 24229 22404
rect 24163 22339 24229 22340
rect 23979 2548 24045 2549
rect 23979 2484 23980 2548
rect 24044 2484 24045 2548
rect 23979 2483 24045 2484
rect 24166 2413 24226 22339
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 24163 2412 24229 2413
rect 24163 2348 24164 2412
rect 24228 2348 24229 2412
rect 24163 2347 24229 2348
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 18584 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1644511149
transform -1 0 31004 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1644511149
transform 1 0 22540 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1644511149
transform 1 0 24104 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1644511149
transform 1 0 23644 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1644511149
transform 1 0 30452 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1644511149
transform 1 0 31188 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1644511149
transform 1 0 37628 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1644511149
transform 1 0 5796 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1644511149
transform 1 0 24656 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1644511149
transform 1 0 15088 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1644511149
transform 1 0 18400 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4048 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_42 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4968 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78
timestamp 1644511149
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_95
timestamp 1644511149
transform 1 0 9844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_103 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_134
timestamp 1644511149
transform 1 0 13432 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_149
timestamp 1644511149
transform 1 0 14812 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_161
timestamp 1644511149
transform 1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1644511149
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177
timestamp 1644511149
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_182
timestamp 1644511149
transform 1 0 17848 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1644511149
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_205
timestamp 1644511149
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_210
timestamp 1644511149
transform 1 0 20424 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1644511149
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_233
timestamp 1644511149
transform 1 0 22540 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_238
timestamp 1644511149
transform 1 0 23000 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_245
timestamp 1644511149
transform 1 0 23644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1644511149
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_265
timestamp 1644511149
transform 1 0 25484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_272
timestamp 1644511149
transform 1 0 26128 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_286
timestamp 1644511149
transform 1 0 27416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_300
timestamp 1644511149
transform 1 0 28704 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_330
timestamp 1644511149
transform 1 0 31464 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_345
timestamp 1644511149
transform 1 0 32844 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_350
timestamp 1644511149
transform 1 0 33304 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_360
timestamp 1644511149
transform 1 0 34224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_371
timestamp 1644511149
transform 1 0 35236 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_379
timestamp 1644511149
transform 1 0 35972 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_384
timestamp 1644511149
transform 1 0 36432 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_393
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_405
timestamp 1644511149
transform 1 0 38364 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_416
timestamp 1644511149
transform 1 0 39376 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_421
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_425
timestamp 1644511149
transform 1 0 40204 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_437
timestamp 1644511149
transform 1 0 41308 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_449
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_457
timestamp 1644511149
transform 1 0 43148 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_462
timestamp 1644511149
transform 1 0 43608 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_466
timestamp 1644511149
transform 1 0 43976 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_470
timestamp 1644511149
transform 1 0 44344 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_498
timestamp 1644511149
transform 1 0 46920 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_505
timestamp 1644511149
transform 1 0 47564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_512
timestamp 1644511149
transform 1 0 48208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_11
timestamp 1644511149
transform 1 0 2116 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_19
timestamp 1644511149
transform 1 0 2852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_23
timestamp 1644511149
transform 1 0 3220 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_45
timestamp 1644511149
transform 1 0 5244 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1644511149
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_81
timestamp 1644511149
transform 1 0 8556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_89
timestamp 1644511149
transform 1 0 9292 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_101
timestamp 1644511149
transform 1 0 10396 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_109
timestamp 1644511149
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_117
timestamp 1644511149
transform 1 0 11868 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_139
timestamp 1644511149
transform 1 0 13892 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1644511149
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_175
timestamp 1644511149
transform 1 0 17204 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_197
timestamp 1644511149
transform 1 0 19228 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_205
timestamp 1644511149
transform 1 0 19964 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_211
timestamp 1644511149
transform 1 0 20516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1644511149
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_237
timestamp 1644511149
transform 1 0 22908 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_261
timestamp 1644511149
transform 1 0 25116 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_269
timestamp 1644511149
transform 1 0 25852 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_274
timestamp 1644511149
transform 1 0 26312 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_293
timestamp 1644511149
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_305
timestamp 1644511149
transform 1 0 29164 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_332
timestamp 1644511149
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_358
timestamp 1644511149
transform 1 0 34040 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_370
timestamp 1644511149
transform 1 0 35144 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_382
timestamp 1644511149
transform 1 0 36248 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_386
timestamp 1644511149
transform 1 0 36616 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_405
timestamp 1644511149
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_417
timestamp 1644511149
transform 1 0 39468 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_421
timestamp 1644511149
transform 1 0 39836 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_443
timestamp 1644511149
transform 1 0 41860 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1644511149
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_452
timestamp 1644511149
transform 1 0 42688 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_464
timestamp 1644511149
transform 1 0 43792 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_487
timestamp 1644511149
transform 1 0 45908 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_495
timestamp 1644511149
transform 1 0 46644 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1644511149
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_505
timestamp 1644511149
transform 1 0 47564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_512
timestamp 1644511149
transform 1 0 48208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1644511149
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_32
timestamp 1644511149
transform 1 0 4048 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_57
timestamp 1644511149
transform 1 0 6348 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_65
timestamp 1644511149
transform 1 0 7084 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_70
timestamp 1644511149
transform 1 0 7544 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1644511149
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1644511149
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_97
timestamp 1644511149
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_109
timestamp 1644511149
transform 1 0 11132 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_113
timestamp 1644511149
transform 1 0 11500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_117
timestamp 1644511149
transform 1 0 11868 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_124
timestamp 1644511149
transform 1 0 12512 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1644511149
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_147
timestamp 1644511149
transform 1 0 14628 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1644511149
transform 1 0 15272 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_166
timestamp 1644511149
transform 1 0 16376 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_172
timestamp 1644511149
transform 1 0 16928 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_176
timestamp 1644511149
transform 1 0 17296 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_183
timestamp 1644511149
transform 1 0 17940 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1644511149
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_226
timestamp 1644511149
transform 1 0 21896 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_234
timestamp 1644511149
transform 1 0 22632 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_240
timestamp 1644511149
transform 1 0 23184 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_247
timestamp 1644511149
transform 1 0 23828 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1644511149
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_261
timestamp 1644511149
transform 1 0 25116 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_266
timestamp 1644511149
transform 1 0 25576 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_291
timestamp 1644511149
transform 1 0 27876 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_299
timestamp 1644511149
transform 1 0 28612 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_303
timestamp 1644511149
transform 1 0 28980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1644511149
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_314
timestamp 1644511149
transform 1 0 29992 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_318
timestamp 1644511149
transform 1 0 30360 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_322
timestamp 1644511149
transform 1 0 30728 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_347
timestamp 1644511149
transform 1 0 33028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_359
timestamp 1644511149
transform 1 0 34132 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1644511149
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_404
timestamp 1644511149
transform 1 0 38272 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_408
timestamp 1644511149
transform 1 0 38640 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_412
timestamp 1644511149
transform 1 0 39008 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_424
timestamp 1644511149
transform 1 0 40112 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_435
timestamp 1644511149
transform 1 0 41124 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_460
timestamp 1644511149
transform 1 0 43424 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_467
timestamp 1644511149
transform 1 0 44068 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1644511149
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_480
timestamp 1644511149
transform 1 0 45264 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_509
timestamp 1644511149
transform 1 0 47932 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_515
timestamp 1644511149
transform 1 0 48484 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_6
timestamp 1644511149
transform 1 0 1656 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_13
timestamp 1644511149
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_20
timestamp 1644511149
transform 1 0 2944 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_27
timestamp 1644511149
transform 1 0 3588 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_33
timestamp 1644511149
transform 1 0 4140 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_37
timestamp 1644511149
transform 1 0 4508 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_44
timestamp 1644511149
transform 1 0 5152 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_64
timestamp 1644511149
transform 1 0 6992 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_68
timestamp 1644511149
transform 1 0 7360 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_72
timestamp 1644511149
transform 1 0 7728 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_84
timestamp 1644511149
transform 1 0 8832 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_96
timestamp 1644511149
transform 1 0 9936 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1644511149
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_120
timestamp 1644511149
transform 1 0 12144 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_124
timestamp 1644511149
transform 1 0 12512 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_128
timestamp 1644511149
transform 1 0 12880 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_140
timestamp 1644511149
transform 1 0 13984 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_152
timestamp 1644511149
transform 1 0 15088 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1644511149
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_181
timestamp 1644511149
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_193
timestamp 1644511149
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1644511149
transform 1 0 20240 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_220
timestamp 1644511149
transform 1 0 21344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_237
timestamp 1644511149
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_249
timestamp 1644511149
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_261
timestamp 1644511149
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1644511149
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_310
timestamp 1644511149
transform 1 0 29624 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_317
timestamp 1644511149
transform 1 0 30268 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_321
timestamp 1644511149
transform 1 0 30636 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_325
timestamp 1644511149
transform 1 0 31004 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_333
timestamp 1644511149
transform 1 0 31740 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_340
timestamp 1644511149
transform 1 0 32384 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_347
timestamp 1644511149
transform 1 0 33028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_359
timestamp 1644511149
transform 1 0 34132 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_371
timestamp 1644511149
transform 1 0 35236 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_379
timestamp 1644511149
transform 1 0 35972 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_384
timestamp 1644511149
transform 1 0 36432 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_404
timestamp 1644511149
transform 1 0 38272 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_408
timestamp 1644511149
transform 1 0 38640 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_430
timestamp 1644511149
transform 1 0 40664 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_437
timestamp 1644511149
transform 1 0 41308 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_444
timestamp 1644511149
transform 1 0 41952 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_470
timestamp 1644511149
transform 1 0 44344 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_478
timestamp 1644511149
transform 1 0 45080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_482
timestamp 1644511149
transform 1 0 45448 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_489
timestamp 1644511149
transform 1 0 46092 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_500
timestamp 1644511149
transform 1 0 47104 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_505
timestamp 1644511149
transform 1 0 47564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_512
timestamp 1644511149
transform 1 0 48208 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1644511149
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_109
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_121
timestamp 1644511149
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1644511149
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_221
timestamp 1644511149
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_233
timestamp 1644511149
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1644511149
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1644511149
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1644511149
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_345
timestamp 1644511149
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1644511149
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_401
timestamp 1644511149
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1644511149
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1644511149
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_421
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_433
timestamp 1644511149
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_445
timestamp 1644511149
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_457
timestamp 1644511149
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1644511149
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1644511149
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_480
timestamp 1644511149
transform 1 0 45264 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_487
timestamp 1644511149
transform 1 0 45908 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_512
timestamp 1644511149
transform 1 0 48208 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_7
timestamp 1644511149
transform 1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_32
timestamp 1644511149
transform 1 0 4048 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_44
timestamp 1644511149
transform 1 0 5152 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_205
timestamp 1644511149
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1644511149
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1644511149
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_332
timestamp 1644511149
transform 1 0 31648 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_359
timestamp 1644511149
transform 1 0 34132 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_371
timestamp 1644511149
transform 1 0 35236 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_383
timestamp 1644511149
transform 1 0 36340 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_405
timestamp 1644511149
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_417
timestamp 1644511149
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_429
timestamp 1644511149
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1644511149
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1644511149
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_449
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_461
timestamp 1644511149
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_473
timestamp 1644511149
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_485
timestamp 1644511149
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_500
timestamp 1644511149
transform 1 0 47104 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_505
timestamp 1644511149
transform 1 0 47564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_512
timestamp 1644511149
transform 1 0 48208 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_8
timestamp 1644511149
transform 1 0 1840 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_19
timestamp 1644511149
transform 1 0 2852 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp 1644511149
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_258
timestamp 1644511149
transform 1 0 24840 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_267
timestamp 1644511149
transform 1 0 25668 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_279
timestamp 1644511149
transform 1 0 26772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_291
timestamp 1644511149
transform 1 0 27876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_303
timestamp 1644511149
transform 1 0 28980 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1644511149
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1644511149
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_433
timestamp 1644511149
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_445
timestamp 1644511149
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_457
timestamp 1644511149
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1644511149
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1644511149
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_477
timestamp 1644511149
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_489
timestamp 1644511149
transform 1 0 46092 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_512
timestamp 1644511149
transform 1 0 48208 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_14
timestamp 1644511149
transform 1 0 2392 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_26
timestamp 1644511149
transform 1 0 3496 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_38
timestamp 1644511149
transform 1 0 4600 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_50
timestamp 1644511149
transform 1 0 5704 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1644511149
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1644511149
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_461
timestamp 1644511149
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_473
timestamp 1644511149
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_485
timestamp 1644511149
transform 1 0 45724 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_489
timestamp 1644511149
transform 1 0 46092 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_501
timestamp 1644511149
transform 1 0 47196 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_508
timestamp 1644511149
transform 1 0 47840 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1644511149
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_242
timestamp 1644511149
transform 1 0 23368 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1644511149
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_401
timestamp 1644511149
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1644511149
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1644511149
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_433
timestamp 1644511149
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_445
timestamp 1644511149
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_457
timestamp 1644511149
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1644511149
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1644511149
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_477
timestamp 1644511149
transform 1 0 44988 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_485
timestamp 1644511149
transform 1 0 45724 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_507
timestamp 1644511149
transform 1 0 47748 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_515
timestamp 1644511149
transform 1 0 48484 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7
timestamp 1644511149
transform 1 0 1748 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_11
timestamp 1644511149
transform 1 0 2116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_23
timestamp 1644511149
transform 1 0 3220 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_35
timestamp 1644511149
transform 1 0 4324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_47
timestamp 1644511149
transform 1 0 5428 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_189
timestamp 1644511149
transform 1 0 18492 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_195
timestamp 1644511149
transform 1 0 19044 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_207
timestamp 1644511149
transform 1 0 20148 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_219
timestamp 1644511149
transform 1 0 21252 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_233
timestamp 1644511149
transform 1 0 22540 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_251
timestamp 1644511149
transform 1 0 24196 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_263
timestamp 1644511149
transform 1 0 25300 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_275
timestamp 1644511149
transform 1 0 26404 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_388
timestamp 1644511149
transform 1 0 36800 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_414
timestamp 1644511149
transform 1 0 39192 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_426
timestamp 1644511149
transform 1 0 40296 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_438
timestamp 1644511149
transform 1 0 41400 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_446
timestamp 1644511149
transform 1 0 42136 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_461
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_473
timestamp 1644511149
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_485
timestamp 1644511149
transform 1 0 45724 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_493
timestamp 1644511149
transform 1 0 46460 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_498
timestamp 1644511149
transform 1 0 46920 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_508
timestamp 1644511149
transform 1 0 47840 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_7
timestamp 1644511149
transform 1 0 1748 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_19
timestamp 1644511149
transform 1 0 2852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_185
timestamp 1644511149
transform 1 0 18124 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_191
timestamp 1644511149
transform 1 0 18676 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_218
timestamp 1644511149
transform 1 0 21160 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_238
timestamp 1644511149
transform 1 0 23000 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_247
timestamp 1644511149
transform 1 0 23828 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_261
timestamp 1644511149
transform 1 0 25116 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_270
timestamp 1644511149
transform 1 0 25944 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_276
timestamp 1644511149
transform 1 0 26496 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_285
timestamp 1644511149
transform 1 0 27324 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_297
timestamp 1644511149
transform 1 0 28428 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_305
timestamp 1644511149
transform 1 0 29164 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1644511149
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1644511149
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1644511149
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_457
timestamp 1644511149
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1644511149
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1644511149
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_477
timestamp 1644511149
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_489
timestamp 1644511149
transform 1 0 46092 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_512
timestamp 1644511149
transform 1 0 48208 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_13
timestamp 1644511149
transform 1 0 2300 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_25
timestamp 1644511149
transform 1 0 3404 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_37
timestamp 1644511149
transform 1 0 4508 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_49
timestamp 1644511149
transform 1 0 5612 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_204
timestamp 1644511149
transform 1 0 19872 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_208
timestamp 1644511149
transform 1 0 20240 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_230
timestamp 1644511149
transform 1 0 22264 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_252
timestamp 1644511149
transform 1 0 24288 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_274
timestamp 1644511149
transform 1 0 26312 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_297
timestamp 1644511149
transform 1 0 28428 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_309
timestamp 1644511149
transform 1 0 29532 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_332
timestamp 1644511149
transform 1 0 31648 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_417
timestamp 1644511149
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1644511149
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1644511149
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_449
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_461
timestamp 1644511149
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_473
timestamp 1644511149
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_485
timestamp 1644511149
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1644511149
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1644511149
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_505
timestamp 1644511149
transform 1 0 47564 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_512
timestamp 1644511149
transform 1 0 48208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_213
timestamp 1644511149
transform 1 0 20700 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_222
timestamp 1644511149
transform 1 0 21528 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_226
timestamp 1644511149
transform 1 0 21896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_232
timestamp 1644511149
transform 1 0 22448 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_246
timestamp 1644511149
transform 1 0 23736 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_262
timestamp 1644511149
transform 1 0 25208 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_274
timestamp 1644511149
transform 1 0 26312 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_280
timestamp 1644511149
transform 1 0 26864 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_292
timestamp 1644511149
transform 1 0 27968 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_304
timestamp 1644511149
transform 1 0 29072 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_445
timestamp 1644511149
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_457
timestamp 1644511149
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1644511149
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1644511149
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_477
timestamp 1644511149
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_489
timestamp 1644511149
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_501
timestamp 1644511149
transform 1 0 47196 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_507
timestamp 1644511149
transform 1 0 47748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_512
timestamp 1644511149
transform 1 0 48208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_30
timestamp 1644511149
transform 1 0 3864 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_42
timestamp 1644511149
transform 1 0 4968 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1644511149
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_175
timestamp 1644511149
transform 1 0 17204 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_192
timestamp 1644511149
transform 1 0 18768 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_204
timestamp 1644511149
transform 1 0 19872 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_216
timestamp 1644511149
transform 1 0 20976 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_248
timestamp 1644511149
transform 1 0 23920 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_256
timestamp 1644511149
transform 1 0 24656 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_268
timestamp 1644511149
transform 1 0 25760 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_287
timestamp 1644511149
transform 1 0 27508 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_307
timestamp 1644511149
transform 1 0 29348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_316
timestamp 1644511149
transform 1 0 30176 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_323
timestamp 1644511149
transform 1 0 30820 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1644511149
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_417
timestamp 1644511149
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_429
timestamp 1644511149
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1644511149
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1644511149
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_461
timestamp 1644511149
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_473
timestamp 1644511149
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_485
timestamp 1644511149
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1644511149
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1644511149
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_505
timestamp 1644511149
transform 1 0 47564 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_513
timestamp 1644511149
transform 1 0 48300 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_6
timestamp 1644511149
transform 1 0 1656 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_13
timestamp 1644511149
transform 1 0 2300 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_20
timestamp 1644511149
transform 1 0 2944 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_202
timestamp 1644511149
transform 1 0 19688 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_214
timestamp 1644511149
transform 1 0 20792 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_226
timestamp 1644511149
transform 1 0 21896 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_238
timestamp 1644511149
transform 1 0 23000 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1644511149
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_284
timestamp 1644511149
transform 1 0 27232 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_296
timestamp 1644511149
transform 1 0 28336 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1644511149
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1644511149
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_433
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_445
timestamp 1644511149
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_457
timestamp 1644511149
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1644511149
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1644511149
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_477
timestamp 1644511149
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_489
timestamp 1644511149
transform 1 0 46092 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_512
timestamp 1644511149
transform 1 0 48208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_28
timestamp 1644511149
transform 1 0 3680 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_40
timestamp 1644511149
transform 1 0 4784 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1644511149
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_188
timestamp 1644511149
transform 1 0 18400 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_200
timestamp 1644511149
transform 1 0 19504 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_220
timestamp 1644511149
transform 1 0 21344 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_245
timestamp 1644511149
transform 1 0 23644 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_257
timestamp 1644511149
transform 1 0 24748 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_265
timestamp 1644511149
transform 1 0 25484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_277
timestamp 1644511149
transform 1 0 26588 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_327
timestamp 1644511149
transform 1 0 31188 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_417
timestamp 1644511149
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_429
timestamp 1644511149
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1644511149
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1644511149
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_461
timestamp 1644511149
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_473
timestamp 1644511149
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_485
timestamp 1644511149
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1644511149
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1644511149
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_505
timestamp 1644511149
transform 1 0 47564 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_512
timestamp 1644511149
transform 1 0 48208 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_11
timestamp 1644511149
transform 1 0 2116 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_18
timestamp 1644511149
transform 1 0 2760 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1644511149
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_134
timestamp 1644511149
transform 1 0 13432 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_173
timestamp 1644511149
transform 1 0 17020 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1644511149
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_207
timestamp 1644511149
transform 1 0 20148 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_215
timestamp 1644511149
transform 1 0 20884 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_234
timestamp 1644511149
transform 1 0 22632 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_246
timestamp 1644511149
transform 1 0 23736 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_269
timestamp 1644511149
transform 1 0 25852 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_282
timestamp 1644511149
transform 1 0 27048 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_290
timestamp 1644511149
transform 1 0 27784 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_296
timestamp 1644511149
transform 1 0 28336 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_303
timestamp 1644511149
transform 1 0 28980 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_315
timestamp 1644511149
transform 1 0 30084 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_335
timestamp 1644511149
transform 1 0 31924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_347
timestamp 1644511149
transform 1 0 33028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_359
timestamp 1644511149
transform 1 0 34132 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_396
timestamp 1644511149
transform 1 0 37536 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_408
timestamp 1644511149
transform 1 0 38640 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_433
timestamp 1644511149
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_445
timestamp 1644511149
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_457
timestamp 1644511149
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1644511149
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1644511149
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_477
timestamp 1644511149
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_489
timestamp 1644511149
transform 1 0 46092 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_497
timestamp 1644511149
transform 1 0 46828 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_503
timestamp 1644511149
transform 1 0 47380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_510
timestamp 1644511149
transform 1 0 48024 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1644511149
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_187
timestamp 1644511149
transform 1 0 18308 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_190
timestamp 1644511149
transform 1 0 18584 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_202
timestamp 1644511149
transform 1 0 19688 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_206
timestamp 1644511149
transform 1 0 20056 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_212
timestamp 1644511149
transform 1 0 20608 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_234
timestamp 1644511149
transform 1 0 22632 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_244
timestamp 1644511149
transform 1 0 23552 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_248
timestamp 1644511149
transform 1 0 23920 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_258
timestamp 1644511149
transform 1 0 24840 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_264
timestamp 1644511149
transform 1 0 25392 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_274
timestamp 1644511149
transform 1 0 26312 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_285
timestamp 1644511149
transform 1 0 27324 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_305
timestamp 1644511149
transform 1 0 29164 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_313
timestamp 1644511149
transform 1 0 29900 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_322
timestamp 1644511149
transform 1 0 30728 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_331
timestamp 1644511149
transform 1 0 31556 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1644511149
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_414
timestamp 1644511149
transform 1 0 39192 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_426
timestamp 1644511149
transform 1 0 40296 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_438
timestamp 1644511149
transform 1 0 41400 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_446
timestamp 1644511149
transform 1 0 42136 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_449
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_461
timestamp 1644511149
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_473
timestamp 1644511149
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_485
timestamp 1644511149
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1644511149
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1644511149
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_505
timestamp 1644511149
transform 1 0 47564 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_513
timestamp 1644511149
transform 1 0 48300 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_113
timestamp 1644511149
transform 1 0 11500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_117
timestamp 1644511149
transform 1 0 11868 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_129
timestamp 1644511149
transform 1 0 12972 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_137
timestamp 1644511149
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_177
timestamp 1644511149
transform 1 0 17388 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_185
timestamp 1644511149
transform 1 0 18124 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_191
timestamp 1644511149
transform 1 0 18676 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_205
timestamp 1644511149
transform 1 0 19964 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_217
timestamp 1644511149
transform 1 0 21068 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_221
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_231
timestamp 1644511149
transform 1 0 22356 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_243
timestamp 1644511149
transform 1 0 23460 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_248
timestamp 1644511149
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_263
timestamp 1644511149
transform 1 0 25300 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_274
timestamp 1644511149
transform 1 0 26312 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_282
timestamp 1644511149
transform 1 0 27048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_292
timestamp 1644511149
transform 1 0 27968 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_300
timestamp 1644511149
transform 1 0 28704 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_325
timestamp 1644511149
transform 1 0 31004 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_337
timestamp 1644511149
transform 1 0 32108 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_349
timestamp 1644511149
transform 1 0 33212 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_361
timestamp 1644511149
transform 1 0 34316 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1644511149
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1644511149
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_421
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_433
timestamp 1644511149
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_445
timestamp 1644511149
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_457
timestamp 1644511149
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1644511149
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1644511149
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_477
timestamp 1644511149
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_489
timestamp 1644511149
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_501
timestamp 1644511149
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_513
timestamp 1644511149
transform 1 0 48300 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_13
timestamp 1644511149
transform 1 0 2300 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_25
timestamp 1644511149
transform 1 0 3404 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_37
timestamp 1644511149
transform 1 0 4508 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_49
timestamp 1644511149
transform 1 0 5612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_89
timestamp 1644511149
transform 1 0 9292 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_108
timestamp 1644511149
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_142
timestamp 1644511149
transform 1 0 14168 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_154
timestamp 1644511149
transform 1 0 15272 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1644511149
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_186
timestamp 1644511149
transform 1 0 18216 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_198
timestamp 1644511149
transform 1 0 19320 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_210
timestamp 1644511149
transform 1 0 20424 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_220
timestamp 1644511149
transform 1 0 21344 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_234
timestamp 1644511149
transform 1 0 22632 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_246
timestamp 1644511149
transform 1 0 23736 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_250
timestamp 1644511149
transform 1 0 24104 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_255
timestamp 1644511149
transform 1 0 24564 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_266
timestamp 1644511149
transform 1 0 25576 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_276
timestamp 1644511149
transform 1 0 26496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_294
timestamp 1644511149
transform 1 0 28152 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_303
timestamp 1644511149
transform 1 0 28980 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_315
timestamp 1644511149
transform 1 0 30084 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_327
timestamp 1644511149
transform 1 0 31188 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_342
timestamp 1644511149
transform 1 0 32568 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_354
timestamp 1644511149
transform 1 0 33672 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_366
timestamp 1644511149
transform 1 0 34776 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_378
timestamp 1644511149
transform 1 0 35880 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_390
timestamp 1644511149
transform 1 0 36984 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_417
timestamp 1644511149
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_429
timestamp 1644511149
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1644511149
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1644511149
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_461
timestamp 1644511149
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_473
timestamp 1644511149
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_485
timestamp 1644511149
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1644511149
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1644511149
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_505
timestamp 1644511149
transform 1 0 47564 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_513
timestamp 1644511149
transform 1 0 48300 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_24
timestamp 1644511149
transform 1 0 3312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_162
timestamp 1644511149
transform 1 0 16008 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_170
timestamp 1644511149
transform 1 0 16744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_187
timestamp 1644511149
transform 1 0 18308 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_213
timestamp 1644511149
transform 1 0 20700 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_223
timestamp 1644511149
transform 1 0 21620 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_235
timestamp 1644511149
transform 1 0 22724 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_244
timestamp 1644511149
transform 1 0 23552 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_265
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_273
timestamp 1644511149
transform 1 0 26220 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_281
timestamp 1644511149
transform 1 0 26956 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_287
timestamp 1644511149
transform 1 0 27508 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_297
timestamp 1644511149
transform 1 0 28428 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_305
timestamp 1644511149
transform 1 0 29164 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_317
timestamp 1644511149
transform 1 0 30268 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_322
timestamp 1644511149
transform 1 0 30728 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_342
timestamp 1644511149
transform 1 0 32568 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_354
timestamp 1644511149
transform 1 0 33672 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_362
timestamp 1644511149
transform 1 0 34408 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_401
timestamp 1644511149
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1644511149
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1644511149
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_433
timestamp 1644511149
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_445
timestamp 1644511149
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_457
timestamp 1644511149
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1644511149
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1644511149
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_477
timestamp 1644511149
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_489
timestamp 1644511149
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_501
timestamp 1644511149
transform 1 0 47196 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_507
timestamp 1644511149
transform 1 0 47748 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_515
timestamp 1644511149
transform 1 0 48484 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_9
timestamp 1644511149
transform 1 0 1932 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_13
timestamp 1644511149
transform 1 0 2300 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_20
timestamp 1644511149
transform 1 0 2944 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_32
timestamp 1644511149
transform 1 0 4048 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_44
timestamp 1644511149
transform 1 0 5152 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1644511149
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1644511149
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_182
timestamp 1644511149
transform 1 0 17848 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_202
timestamp 1644511149
transform 1 0 19688 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_208
timestamp 1644511149
transform 1 0 20240 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1644511149
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1644511149
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_234
timestamp 1644511149
transform 1 0 22632 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_256
timestamp 1644511149
transform 1 0 24656 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_268
timestamp 1644511149
transform 1 0 25760 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_288
timestamp 1644511149
transform 1 0 27600 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_308
timestamp 1644511149
transform 1 0 29440 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_320
timestamp 1644511149
transform 1 0 30544 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_330
timestamp 1644511149
transform 1 0 31464 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_359
timestamp 1644511149
transform 1 0 34132 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_371
timestamp 1644511149
transform 1 0 35236 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_383
timestamp 1644511149
transform 1 0 36340 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_417
timestamp 1644511149
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_429
timestamp 1644511149
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1644511149
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1644511149
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_461
timestamp 1644511149
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_473
timestamp 1644511149
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_485
timestamp 1644511149
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1644511149
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1644511149
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_505
timestamp 1644511149
transform 1 0 47564 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_512
timestamp 1644511149
transform 1 0 48208 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1644511149
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_153
timestamp 1644511149
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_165
timestamp 1644511149
transform 1 0 16284 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_173
timestamp 1644511149
transform 1 0 17020 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_178
timestamp 1644511149
transform 1 0 17480 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_186
timestamp 1644511149
transform 1 0 18216 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1644511149
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_200
timestamp 1644511149
transform 1 0 19504 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_212
timestamp 1644511149
transform 1 0 20608 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_225
timestamp 1644511149
transform 1 0 21804 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_238
timestamp 1644511149
transform 1 0 23000 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_246
timestamp 1644511149
transform 1 0 23736 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_257
timestamp 1644511149
transform 1 0 24748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_265
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_275
timestamp 1644511149
transform 1 0 26404 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_290
timestamp 1644511149
transform 1 0 27784 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_297
timestamp 1644511149
transform 1 0 28428 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_305
timestamp 1644511149
transform 1 0 29164 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_321
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_329
timestamp 1644511149
transform 1 0 31372 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_345
timestamp 1644511149
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1644511149
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_401
timestamp 1644511149
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1644511149
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1644511149
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_433
timestamp 1644511149
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_445
timestamp 1644511149
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_457
timestamp 1644511149
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1644511149
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1644511149
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_477
timestamp 1644511149
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_489
timestamp 1644511149
transform 1 0 46092 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_512
timestamp 1644511149
transform 1 0 48208 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1644511149
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1644511149
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1644511149
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1644511149
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_177
timestamp 1644511149
transform 1 0 17388 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_183
timestamp 1644511149
transform 1 0 17940 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_199
timestamp 1644511149
transform 1 0 19412 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_212
timestamp 1644511149
transform 1 0 20608 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_216
timestamp 1644511149
transform 1 0 20976 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1644511149
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_230
timestamp 1644511149
transform 1 0 22264 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_237
timestamp 1644511149
transform 1 0 22908 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_241
timestamp 1644511149
transform 1 0 23276 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_250
timestamp 1644511149
transform 1 0 24104 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_258
timestamp 1644511149
transform 1 0 24840 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_265
timestamp 1644511149
transform 1 0 25484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_277
timestamp 1644511149
transform 1 0 26588 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_289
timestamp 1644511149
transform 1 0 27692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_301
timestamp 1644511149
transform 1 0 28796 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_313
timestamp 1644511149
transform 1 0 29900 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_321
timestamp 1644511149
transform 1 0 30636 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_332
timestamp 1644511149
transform 1 0 31648 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_342
timestamp 1644511149
transform 1 0 32568 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_354
timestamp 1644511149
transform 1 0 33672 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_366
timestamp 1644511149
transform 1 0 34776 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_378
timestamp 1644511149
transform 1 0 35880 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_390
timestamp 1644511149
transform 1 0 36984 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_417
timestamp 1644511149
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_429
timestamp 1644511149
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1644511149
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1644511149
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_461
timestamp 1644511149
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_473
timestamp 1644511149
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_485
timestamp 1644511149
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_500
timestamp 1644511149
transform 1 0 47104 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_508
timestamp 1644511149
transform 1 0 47840 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1644511149
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1644511149
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_153
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_165
timestamp 1644511149
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_177
timestamp 1644511149
transform 1 0 17388 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1644511149
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_207
timestamp 1644511149
transform 1 0 20148 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_218
timestamp 1644511149
transform 1 0 21160 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_230
timestamp 1644511149
transform 1 0 22264 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_236
timestamp 1644511149
transform 1 0 22816 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_248
timestamp 1644511149
transform 1 0 23920 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_265
timestamp 1644511149
transform 1 0 25484 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_273
timestamp 1644511149
transform 1 0 26220 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_281
timestamp 1644511149
transform 1 0 26956 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_290
timestamp 1644511149
transform 1 0 27784 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_294
timestamp 1644511149
transform 1 0 28152 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_304
timestamp 1644511149
transform 1 0 29072 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_325
timestamp 1644511149
transform 1 0 31004 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_329
timestamp 1644511149
transform 1 0 31372 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_346
timestamp 1644511149
transform 1 0 32936 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_358
timestamp 1644511149
transform 1 0 34040 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1644511149
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1644511149
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_433
timestamp 1644511149
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_445
timestamp 1644511149
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_457
timestamp 1644511149
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1644511149
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1644511149
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_477
timestamp 1644511149
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_489
timestamp 1644511149
transform 1 0 46092 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_512
timestamp 1644511149
transform 1 0 48208 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1644511149
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1644511149
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1644511149
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1644511149
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_134
timestamp 1644511149
transform 1 0 13432 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_142
timestamp 1644511149
transform 1 0 14168 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_150
timestamp 1644511149
transform 1 0 14904 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_158
timestamp 1644511149
transform 1 0 15640 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_164
timestamp 1644511149
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_190
timestamp 1644511149
transform 1 0 18584 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_210
timestamp 1644511149
transform 1 0 20424 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_214
timestamp 1644511149
transform 1 0 20792 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_219
timestamp 1644511149
transform 1 0 21252 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_237
timestamp 1644511149
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_249
timestamp 1644511149
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_265
timestamp 1644511149
transform 1 0 25484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_277
timestamp 1644511149
transform 1 0 26588 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_287
timestamp 1644511149
transform 1 0 27508 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_304
timestamp 1644511149
transform 1 0 29072 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_312
timestamp 1644511149
transform 1 0 29808 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_320
timestamp 1644511149
transform 1 0 30544 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_332
timestamp 1644511149
transform 1 0 31648 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_353
timestamp 1644511149
transform 1 0 33580 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_365
timestamp 1644511149
transform 1 0 34684 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_377
timestamp 1644511149
transform 1 0 35788 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_389
timestamp 1644511149
transform 1 0 36892 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_417
timestamp 1644511149
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_429
timestamp 1644511149
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1644511149
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1644511149
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_461
timestamp 1644511149
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_473
timestamp 1644511149
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_485
timestamp 1644511149
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1644511149
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1644511149
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_508
timestamp 1644511149
transform 1 0 47840 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_11
timestamp 1644511149
transform 1 0 2116 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_23
timestamp 1644511149
transform 1 0 3220 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_108
timestamp 1644511149
transform 1 0 11040 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_128
timestamp 1644511149
transform 1 0 12880 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_160
timestamp 1644511149
transform 1 0 15824 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_172
timestamp 1644511149
transform 1 0 16928 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_178
timestamp 1644511149
transform 1 0 17480 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_190
timestamp 1644511149
transform 1 0 18584 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_207
timestamp 1644511149
transform 1 0 20148 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_217
timestamp 1644511149
transform 1 0 21068 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_225
timestamp 1644511149
transform 1 0 21804 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_237
timestamp 1644511149
transform 1 0 22908 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_249
timestamp 1644511149
transform 1 0 24012 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_269
timestamp 1644511149
transform 1 0 25852 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_281
timestamp 1644511149
transform 1 0 26956 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_289
timestamp 1644511149
transform 1 0 27692 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_302
timestamp 1644511149
transform 1 0 28888 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_318
timestamp 1644511149
transform 1 0 30360 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_330
timestamp 1644511149
transform 1 0 31464 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_336
timestamp 1644511149
transform 1 0 32016 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_348
timestamp 1644511149
transform 1 0 33120 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_360
timestamp 1644511149
transform 1 0 34224 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_401
timestamp 1644511149
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1644511149
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1644511149
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_421
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_433
timestamp 1644511149
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_445
timestamp 1644511149
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_457
timestamp 1644511149
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1644511149
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1644511149
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_477
timestamp 1644511149
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_489
timestamp 1644511149
transform 1 0 46092 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_512
timestamp 1644511149
transform 1 0 48208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_28
timestamp 1644511149
transform 1 0 3680 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_40
timestamp 1644511149
transform 1 0 4784 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 1644511149
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_86
timestamp 1644511149
transform 1 0 9016 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_94
timestamp 1644511149
transform 1 0 9752 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_99
timestamp 1644511149
transform 1 0 10212 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_108
timestamp 1644511149
transform 1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_122
timestamp 1644511149
transform 1 0 12328 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_136
timestamp 1644511149
transform 1 0 13616 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_150
timestamp 1644511149
transform 1 0 14904 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_162
timestamp 1644511149
transform 1 0 16008 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_187
timestamp 1644511149
transform 1 0 18308 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_195
timestamp 1644511149
transform 1 0 19044 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_199
timestamp 1644511149
transform 1 0 19412 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_216
timestamp 1644511149
transform 1 0 20976 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_232
timestamp 1644511149
transform 1 0 22448 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_236
timestamp 1644511149
transform 1 0 22816 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_243
timestamp 1644511149
transform 1 0 23460 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_248
timestamp 1644511149
transform 1 0 23920 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_252
timestamp 1644511149
transform 1 0 24288 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_260
timestamp 1644511149
transform 1 0 25024 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_268
timestamp 1644511149
transform 1 0 25760 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_287
timestamp 1644511149
transform 1 0 27508 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_296
timestamp 1644511149
transform 1 0 28336 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_300
timestamp 1644511149
transform 1 0 28704 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_317
timestamp 1644511149
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1644511149
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1644511149
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_371
timestamp 1644511149
transform 1 0 35236 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_383
timestamp 1644511149
transform 1 0 36340 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1644511149
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_417
timestamp 1644511149
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_429
timestamp 1644511149
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1644511149
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1644511149
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_449
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_461
timestamp 1644511149
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_473
timestamp 1644511149
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_485
timestamp 1644511149
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1644511149
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1644511149
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_508
timestamp 1644511149
transform 1 0 47840 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_6
timestamp 1644511149
transform 1 0 1656 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_13
timestamp 1644511149
transform 1 0 2300 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_20
timestamp 1644511149
transform 1 0 2944 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_80
timestamp 1644511149
transform 1 0 8464 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_93
timestamp 1644511149
transform 1 0 9660 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_116
timestamp 1644511149
transform 1 0 11776 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_124
timestamp 1644511149
transform 1 0 12512 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp 1644511149
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_163
timestamp 1644511149
transform 1 0 16100 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_171
timestamp 1644511149
transform 1 0 16836 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1644511149
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_201
timestamp 1644511149
transform 1 0 19596 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_213
timestamp 1644511149
transform 1 0 20700 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_217
timestamp 1644511149
transform 1 0 21068 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_224
timestamp 1644511149
transform 1 0 21712 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_232
timestamp 1644511149
transform 1 0 22448 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_246
timestamp 1644511149
transform 1 0 23736 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_258
timestamp 1644511149
transform 1 0 24840 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_265
timestamp 1644511149
transform 1 0 25484 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_275
timestamp 1644511149
transform 1 0 26404 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_284
timestamp 1644511149
transform 1 0 27232 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_293
timestamp 1644511149
transform 1 0 28060 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1644511149
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1644511149
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_321
timestamp 1644511149
transform 1 0 30636 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_325
timestamp 1644511149
transform 1 0 31004 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_350
timestamp 1644511149
transform 1 0 33304 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1644511149
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1644511149
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_368
timestamp 1644511149
transform 1 0 34960 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_380
timestamp 1644511149
transform 1 0 36064 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_392
timestamp 1644511149
transform 1 0 37168 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_404
timestamp 1644511149
transform 1 0 38272 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_416
timestamp 1644511149
transform 1 0 39376 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_421
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_433
timestamp 1644511149
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_445
timestamp 1644511149
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_457
timestamp 1644511149
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1644511149
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1644511149
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_477
timestamp 1644511149
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_489
timestamp 1644511149
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_501
timestamp 1644511149
transform 1 0 47196 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_507
timestamp 1644511149
transform 1 0 47748 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_515
timestamp 1644511149
transform 1 0 48484 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_28
timestamp 1644511149
transform 1 0 3680 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_35
timestamp 1644511149
transform 1 0 4324 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_47
timestamp 1644511149
transform 1 0 5428 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_125
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_143
timestamp 1644511149
transform 1 0 14260 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_155
timestamp 1644511149
transform 1 0 15364 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 1644511149
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_175
timestamp 1644511149
transform 1 0 17204 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_183
timestamp 1644511149
transform 1 0 17940 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_189
timestamp 1644511149
transform 1 0 18492 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_193
timestamp 1644511149
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_205
timestamp 1644511149
transform 1 0 19964 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1644511149
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_232
timestamp 1644511149
transform 1 0 22448 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_238
timestamp 1644511149
transform 1 0 23000 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_244
timestamp 1644511149
transform 1 0 23552 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_252
timestamp 1644511149
transform 1 0 24288 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_262
timestamp 1644511149
transform 1 0 25208 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_270
timestamp 1644511149
transform 1 0 25944 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1644511149
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_291
timestamp 1644511149
transform 1 0 27876 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_305
timestamp 1644511149
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_317
timestamp 1644511149
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1644511149
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1644511149
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_366
timestamp 1644511149
transform 1 0 34776 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_378
timestamp 1644511149
transform 1 0 35880 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_390
timestamp 1644511149
transform 1 0 36984 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_405
timestamp 1644511149
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_417
timestamp 1644511149
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_429
timestamp 1644511149
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1644511149
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1644511149
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_449
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_461
timestamp 1644511149
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_473
timestamp 1644511149
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_485
timestamp 1644511149
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1644511149
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1644511149
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_505
timestamp 1644511149
transform 1 0 47564 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_513
timestamp 1644511149
transform 1 0 48300 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_24
timestamp 1644511149
transform 1 0 3312 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_91
timestamp 1644511149
transform 1 0 9476 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_100
timestamp 1644511149
transform 1 0 10304 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_108
timestamp 1644511149
transform 1 0 11040 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_126
timestamp 1644511149
transform 1 0 12696 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_135
timestamp 1644511149
transform 1 0 13524 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_149
timestamp 1644511149
transform 1 0 14812 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_157
timestamp 1644511149
transform 1 0 15548 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_174
timestamp 1644511149
transform 1 0 17112 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_181
timestamp 1644511149
transform 1 0 17756 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_193
timestamp 1644511149
transform 1 0 18860 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_205
timestamp 1644511149
transform 1 0 19964 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_214
timestamp 1644511149
transform 1 0 20792 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_224
timestamp 1644511149
transform 1 0 21712 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_231
timestamp 1644511149
transform 1 0 22356 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_239
timestamp 1644511149
transform 1 0 23092 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_246
timestamp 1644511149
transform 1 0 23736 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_258
timestamp 1644511149
transform 1 0 24840 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_266
timestamp 1644511149
transform 1 0 25576 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_277
timestamp 1644511149
transform 1 0 26588 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_288
timestamp 1644511149
transform 1 0 27600 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_292
timestamp 1644511149
transform 1 0 27968 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_302
timestamp 1644511149
transform 1 0 28888 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_321
timestamp 1644511149
transform 1 0 30636 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_339
timestamp 1644511149
transform 1 0 32292 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_351
timestamp 1644511149
transform 1 0 33396 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1644511149
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_389
timestamp 1644511149
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_401
timestamp 1644511149
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1644511149
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1644511149
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_421
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_433
timestamp 1644511149
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_445
timestamp 1644511149
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_457
timestamp 1644511149
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1644511149
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1644511149
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_477
timestamp 1644511149
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_489
timestamp 1644511149
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_501
timestamp 1644511149
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_513
timestamp 1644511149
transform 1 0 48300 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_7
timestamp 1644511149
transform 1 0 1748 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_14
timestamp 1644511149
transform 1 0 2392 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_26
timestamp 1644511149
transform 1 0 3496 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_38
timestamp 1644511149
transform 1 0 4600 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_50
timestamp 1644511149
transform 1 0 5704 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_103
timestamp 1644511149
transform 1 0 10580 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_121
timestamp 1644511149
transform 1 0 12236 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_143
timestamp 1644511149
transform 1 0 14260 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_155
timestamp 1644511149
transform 1 0 15364 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_163
timestamp 1644511149
transform 1 0 16100 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1644511149
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_172
timestamp 1644511149
transform 1 0 16928 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_182
timestamp 1644511149
transform 1 0 17848 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_194
timestamp 1644511149
transform 1 0 18952 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_206
timestamp 1644511149
transform 1 0 20056 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_216
timestamp 1644511149
transform 1 0 20976 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_232
timestamp 1644511149
transform 1 0 22448 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_238
timestamp 1644511149
transform 1 0 23000 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_243
timestamp 1644511149
transform 1 0 23460 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_251
timestamp 1644511149
transform 1 0 24196 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_265
timestamp 1644511149
transform 1 0 25484 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_276
timestamp 1644511149
transform 1 0 26496 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_285
timestamp 1644511149
transform 1 0 27324 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_295
timestamp 1644511149
transform 1 0 28244 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_315
timestamp 1644511149
transform 1 0 30084 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_332
timestamp 1644511149
transform 1 0 31648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_353
timestamp 1644511149
transform 1 0 33580 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_365
timestamp 1644511149
transform 1 0 34684 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_377
timestamp 1644511149
transform 1 0 35788 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_389
timestamp 1644511149
transform 1 0 36892 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_417
timestamp 1644511149
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_429
timestamp 1644511149
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1644511149
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1644511149
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_449
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_461
timestamp 1644511149
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_473
timestamp 1644511149
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_485
timestamp 1644511149
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_500
timestamp 1644511149
transform 1 0 47104 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_505
timestamp 1644511149
transform 1 0 47564 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_512
timestamp 1644511149
transform 1 0 48208 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1644511149
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_57
timestamp 1644511149
transform 1 0 6348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_79
timestamp 1644511149
transform 1 0 8372 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_93
timestamp 1644511149
transform 1 0 9660 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_108
timestamp 1644511149
transform 1 0 11040 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_120
timestamp 1644511149
transform 1 0 12144 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_132
timestamp 1644511149
transform 1 0 13248 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_146
timestamp 1644511149
transform 1 0 14536 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_158
timestamp 1644511149
transform 1 0 15640 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_170
timestamp 1644511149
transform 1 0 16744 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1644511149
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_213
timestamp 1644511149
transform 1 0 20700 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_226
timestamp 1644511149
transform 1 0 21896 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_237
timestamp 1644511149
transform 1 0 22908 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1644511149
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1644511149
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_267
timestamp 1644511149
transform 1 0 25668 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_279
timestamp 1644511149
transform 1 0 26772 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_290
timestamp 1644511149
transform 1 0 27784 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_302
timestamp 1644511149
transform 1 0 28888 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_327
timestamp 1644511149
transform 1 0 31188 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_339
timestamp 1644511149
transform 1 0 32292 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_351
timestamp 1644511149
transform 1 0 33396 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1644511149
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_389
timestamp 1644511149
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_401
timestamp 1644511149
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1644511149
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1644511149
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_421
timestamp 1644511149
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_433
timestamp 1644511149
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_445
timestamp 1644511149
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_457
timestamp 1644511149
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1644511149
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1644511149
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_477
timestamp 1644511149
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_489
timestamp 1644511149
transform 1 0 46092 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_512
timestamp 1644511149
transform 1 0 48208 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_47
timestamp 1644511149
transform 1 0 5428 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_52
timestamp 1644511149
transform 1 0 5888 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_78
timestamp 1644511149
transform 1 0 8280 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_98
timestamp 1644511149
transform 1 0 10120 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_107
timestamp 1644511149
transform 1 0 10948 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_125
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_131
timestamp 1644511149
transform 1 0 13156 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_135
timestamp 1644511149
transform 1 0 13524 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_147
timestamp 1644511149
transform 1 0 14628 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_159
timestamp 1644511149
transform 1 0 15732 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_164
timestamp 1644511149
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_179
timestamp 1644511149
transform 1 0 17572 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_191
timestamp 1644511149
transform 1 0 18676 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_200
timestamp 1644511149
transform 1 0 19504 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_206
timestamp 1644511149
transform 1 0 20056 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_211
timestamp 1644511149
transform 1 0 20516 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_220
timestamp 1644511149
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_234
timestamp 1644511149
transform 1 0 22632 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_240
timestamp 1644511149
transform 1 0 23184 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_245
timestamp 1644511149
transform 1 0 23644 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_251
timestamp 1644511149
transform 1 0 24196 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_256
timestamp 1644511149
transform 1 0 24656 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_266
timestamp 1644511149
transform 1 0 25576 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_274
timestamp 1644511149
transform 1 0 26312 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_285
timestamp 1644511149
transform 1 0 27324 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_295
timestamp 1644511149
transform 1 0 28244 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_305
timestamp 1644511149
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_317
timestamp 1644511149
transform 1 0 30268 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_324
timestamp 1644511149
transform 1 0 30912 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_342
timestamp 1644511149
transform 1 0 32568 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_354
timestamp 1644511149
transform 1 0 33672 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_360
timestamp 1644511149
transform 1 0 34224 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_364
timestamp 1644511149
transform 1 0 34592 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_376
timestamp 1644511149
transform 1 0 35696 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_388
timestamp 1644511149
transform 1 0 36800 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_417
timestamp 1644511149
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_429
timestamp 1644511149
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1644511149
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1644511149
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_449
timestamp 1644511149
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_461
timestamp 1644511149
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_473
timestamp 1644511149
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_485
timestamp 1644511149
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1644511149
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1644511149
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_508
timestamp 1644511149
transform 1 0 47840 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_59
timestamp 1644511149
transform 1 0 6532 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_63
timestamp 1644511149
transform 1 0 6900 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1644511149
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_101
timestamp 1644511149
transform 1 0 10396 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_110
timestamp 1644511149
transform 1 0 11224 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_122
timestamp 1644511149
transform 1 0 12328 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_134
timestamp 1644511149
transform 1 0 13432 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_159
timestamp 1644511149
transform 1 0 15732 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_171
timestamp 1644511149
transform 1 0 16836 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1644511149
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1644511149
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_209
timestamp 1644511149
transform 1 0 20332 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_215
timestamp 1644511149
transform 1 0 20884 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_220
timestamp 1644511149
transform 1 0 21344 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_231
timestamp 1644511149
transform 1 0 22356 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_241
timestamp 1644511149
transform 1 0 23276 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_248
timestamp 1644511149
transform 1 0 23920 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_265
timestamp 1644511149
transform 1 0 25484 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_273
timestamp 1644511149
transform 1 0 26220 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_280
timestamp 1644511149
transform 1 0 26864 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_304
timestamp 1644511149
transform 1 0 29072 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_317
timestamp 1644511149
transform 1 0 30268 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_329
timestamp 1644511149
transform 1 0 31372 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_333
timestamp 1644511149
transform 1 0 31740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_339
timestamp 1644511149
transform 1 0 32292 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_359
timestamp 1644511149
transform 1 0 34132 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1644511149
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_368
timestamp 1644511149
transform 1 0 34960 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_380
timestamp 1644511149
transform 1 0 36064 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_392
timestamp 1644511149
transform 1 0 37168 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_404
timestamp 1644511149
transform 1 0 38272 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_416
timestamp 1644511149
transform 1 0 39376 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_421
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_433
timestamp 1644511149
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_445
timestamp 1644511149
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_457
timestamp 1644511149
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1644511149
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1644511149
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_477
timestamp 1644511149
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_489
timestamp 1644511149
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_501
timestamp 1644511149
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_513
timestamp 1644511149
transform 1 0 48300 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_63
timestamp 1644511149
transform 1 0 6900 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_75
timestamp 1644511149
transform 1 0 8004 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_87
timestamp 1644511149
transform 1 0 9108 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_96
timestamp 1644511149
transform 1 0 9936 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_108
timestamp 1644511149
transform 1 0 11040 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_122
timestamp 1644511149
transform 1 0 12328 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_131
timestamp 1644511149
transform 1 0 13156 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_137
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_159
timestamp 1644511149
transform 1 0 15732 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1644511149
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_186
timestamp 1644511149
transform 1 0 18216 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_195
timestamp 1644511149
transform 1 0 19044 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_207
timestamp 1644511149
transform 1 0 20148 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_219
timestamp 1644511149
transform 1 0 21252 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1644511149
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_229
timestamp 1644511149
transform 1 0 22172 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_239
timestamp 1644511149
transform 1 0 23092 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_254
timestamp 1644511149
transform 1 0 24472 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_258
timestamp 1644511149
transform 1 0 24840 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_275
timestamp 1644511149
transform 1 0 26404 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1644511149
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_293
timestamp 1644511149
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_305
timestamp 1644511149
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_317
timestamp 1644511149
transform 1 0 30268 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_323
timestamp 1644511149
transform 1 0 30820 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_332
timestamp 1644511149
transform 1 0 31648 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_337
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_357
timestamp 1644511149
transform 1 0 33948 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_384
timestamp 1644511149
transform 1 0 36432 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_417
timestamp 1644511149
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_429
timestamp 1644511149
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1644511149
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1644511149
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_449
timestamp 1644511149
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_461
timestamp 1644511149
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_473
timestamp 1644511149
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_485
timestamp 1644511149
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1644511149
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1644511149
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_505
timestamp 1644511149
transform 1 0 47564 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_513
timestamp 1644511149
transform 1 0 48300 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_57
timestamp 1644511149
transform 1 0 6348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_79
timestamp 1644511149
transform 1 0 8372 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_93
timestamp 1644511149
transform 1 0 9660 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_99
timestamp 1644511149
transform 1 0 10212 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_104
timestamp 1644511149
transform 1 0 10672 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_112
timestamp 1644511149
transform 1 0 11408 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_130
timestamp 1644511149
transform 1 0 13064 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1644511149
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_153
timestamp 1644511149
transform 1 0 15180 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_162
timestamp 1644511149
transform 1 0 16008 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_170
timestamp 1644511149
transform 1 0 16744 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_182
timestamp 1644511149
transform 1 0 17848 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_188
timestamp 1644511149
transform 1 0 18400 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_36_205
timestamp 1644511149
transform 1 0 19964 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_213
timestamp 1644511149
transform 1 0 20700 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_217
timestamp 1644511149
transform 1 0 21068 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_230
timestamp 1644511149
transform 1 0 22264 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_242
timestamp 1644511149
transform 1 0 23368 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1644511149
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_257
timestamp 1644511149
transform 1 0 24748 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_269
timestamp 1644511149
transform 1 0 25852 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_281
timestamp 1644511149
transform 1 0 26956 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_293
timestamp 1644511149
transform 1 0 28060 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_305
timestamp 1644511149
transform 1 0 29164 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_317
timestamp 1644511149
transform 1 0 30268 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_326
timestamp 1644511149
transform 1 0 31096 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_338
timestamp 1644511149
transform 1 0 32200 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_347
timestamp 1644511149
transform 1 0 33028 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_356
timestamp 1644511149
transform 1 0 33856 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_386
timestamp 1644511149
transform 1 0 36616 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_398
timestamp 1644511149
transform 1 0 37720 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_410
timestamp 1644511149
transform 1 0 38824 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_418
timestamp 1644511149
transform 1 0 39560 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_421
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_433
timestamp 1644511149
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_445
timestamp 1644511149
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_457
timestamp 1644511149
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1644511149
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1644511149
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_477
timestamp 1644511149
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_489
timestamp 1644511149
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_501
timestamp 1644511149
transform 1 0 47196 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_507
timestamp 1644511149
transform 1 0 47748 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_512
timestamp 1644511149
transform 1 0 48208 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_7
timestamp 1644511149
transform 1 0 1748 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_11
timestamp 1644511149
transform 1 0 2116 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_65
timestamp 1644511149
transform 1 0 7084 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_82
timestamp 1644511149
transform 1 0 8648 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_91
timestamp 1644511149
transform 1 0 9476 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_107
timestamp 1644511149
transform 1 0 10948 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_129
timestamp 1644511149
transform 1 0 12972 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_138
timestamp 1644511149
transform 1 0 13800 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_150
timestamp 1644511149
transform 1 0 14904 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_154
timestamp 1644511149
transform 1 0 15272 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_164
timestamp 1644511149
transform 1 0 16192 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_174
timestamp 1644511149
transform 1 0 17112 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_194
timestamp 1644511149
transform 1 0 18952 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_214
timestamp 1644511149
transform 1 0 20792 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1644511149
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_241
timestamp 1644511149
transform 1 0 23276 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_249
timestamp 1644511149
transform 1 0 24012 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_256
timestamp 1644511149
transform 1 0 24656 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_266
timestamp 1644511149
transform 1 0 25576 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1644511149
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1644511149
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_286
timestamp 1644511149
transform 1 0 27416 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_294
timestamp 1644511149
transform 1 0 28152 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_302
timestamp 1644511149
transform 1 0 28888 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_322
timestamp 1644511149
transform 1 0 30728 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_334
timestamp 1644511149
transform 1 0 31832 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_353
timestamp 1644511149
transform 1 0 33580 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_365
timestamp 1644511149
transform 1 0 34684 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_377
timestamp 1644511149
transform 1 0 35788 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_389
timestamp 1644511149
transform 1 0 36892 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_417
timestamp 1644511149
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_429
timestamp 1644511149
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1644511149
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1644511149
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_449
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_461
timestamp 1644511149
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_473
timestamp 1644511149
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_485
timestamp 1644511149
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1644511149
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1644511149
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_505
timestamp 1644511149
transform 1 0 47564 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_512
timestamp 1644511149
transform 1 0 48208 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_24
timestamp 1644511149
transform 1 0 3312 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_73
timestamp 1644511149
transform 1 0 7820 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_80
timestamp 1644511149
transform 1 0 8464 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_93
timestamp 1644511149
transform 1 0 9660 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_105
timestamp 1644511149
transform 1 0 10764 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_113
timestamp 1644511149
transform 1 0 11500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_122
timestamp 1644511149
transform 1 0 12328 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_131
timestamp 1644511149
transform 1 0 13156 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_157
timestamp 1644511149
transform 1 0 15548 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_177
timestamp 1644511149
transform 1 0 17388 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1644511149
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1644511149
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_200
timestamp 1644511149
transform 1 0 19504 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_212
timestamp 1644511149
transform 1 0 20608 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_230
timestamp 1644511149
transform 1 0 22264 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_238
timestamp 1644511149
transform 1 0 23000 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_248
timestamp 1644511149
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_262
timestamp 1644511149
transform 1 0 25208 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_276
timestamp 1644511149
transform 1 0 26496 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_282
timestamp 1644511149
transform 1 0 27048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_288
timestamp 1644511149
transform 1 0 27600 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_304
timestamp 1644511149
transform 1 0 29072 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_317
timestamp 1644511149
transform 1 0 30268 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_329
timestamp 1644511149
transform 1 0 31372 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_341
timestamp 1644511149
transform 1 0 32476 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_347
timestamp 1644511149
transform 1 0 33028 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_351
timestamp 1644511149
transform 1 0 33396 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1644511149
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_377
timestamp 1644511149
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_389
timestamp 1644511149
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_401
timestamp 1644511149
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1644511149
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1644511149
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_421
timestamp 1644511149
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_433
timestamp 1644511149
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_445
timestamp 1644511149
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_457
timestamp 1644511149
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1644511149
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1644511149
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_477
timestamp 1644511149
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_489
timestamp 1644511149
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_501
timestamp 1644511149
transform 1 0 47196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_512
timestamp 1644511149
transform 1 0 48208 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_7
timestamp 1644511149
transform 1 0 1748 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_11
timestamp 1644511149
transform 1 0 2116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_23
timestamp 1644511149
transform 1 0 3220 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_35
timestamp 1644511149
transform 1 0 4324 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_47
timestamp 1644511149
transform 1 0 5428 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_89
timestamp 1644511149
transform 1 0 9292 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_101
timestamp 1644511149
transform 1 0 10396 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_109
timestamp 1644511149
transform 1 0 11132 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_129
timestamp 1644511149
transform 1 0 12972 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_134
timestamp 1644511149
transform 1 0 13432 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_142
timestamp 1644511149
transform 1 0 14168 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_146
timestamp 1644511149
transform 1 0 14536 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_150
timestamp 1644511149
transform 1 0 14904 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_162
timestamp 1644511149
transform 1 0 16008 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_173
timestamp 1644511149
transform 1 0 17020 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_178
timestamp 1644511149
transform 1 0 17480 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_194
timestamp 1644511149
transform 1 0 18952 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_201
timestamp 1644511149
transform 1 0 19596 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_213
timestamp 1644511149
transform 1 0 20700 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_221
timestamp 1644511149
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_237
timestamp 1644511149
transform 1 0 22908 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_241
timestamp 1644511149
transform 1 0 23276 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_248
timestamp 1644511149
transform 1 0 23920 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_252
timestamp 1644511149
transform 1 0 24288 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_259
timestamp 1644511149
transform 1 0 24932 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1644511149
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1644511149
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_297
timestamp 1644511149
transform 1 0 28428 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_301
timestamp 1644511149
transform 1 0 28796 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_307
timestamp 1644511149
transform 1 0 29348 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_327
timestamp 1644511149
transform 1 0 31188 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1644511149
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_370
timestamp 1644511149
transform 1 0 35144 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_382
timestamp 1644511149
transform 1 0 36248 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_390
timestamp 1644511149
transform 1 0 36984 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_397
timestamp 1644511149
transform 1 0 37628 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_409
timestamp 1644511149
transform 1 0 38732 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_421
timestamp 1644511149
transform 1 0 39836 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_433
timestamp 1644511149
transform 1 0 40940 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_445
timestamp 1644511149
transform 1 0 42044 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_449
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_461
timestamp 1644511149
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_473
timestamp 1644511149
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_485
timestamp 1644511149
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1644511149
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1644511149
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_505
timestamp 1644511149
transform 1 0 47564 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_513
timestamp 1644511149
transform 1 0 48300 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_7
timestamp 1644511149
transform 1 0 1748 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_19
timestamp 1644511149
transform 1 0 2852 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_24
timestamp 1644511149
transform 1 0 3312 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_50
timestamp 1644511149
transform 1 0 5704 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_62
timestamp 1644511149
transform 1 0 6808 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_74
timestamp 1644511149
transform 1 0 7912 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1644511149
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_93
timestamp 1644511149
transform 1 0 9660 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_102
timestamp 1644511149
transform 1 0 10488 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_114
timestamp 1644511149
transform 1 0 11592 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_125
timestamp 1644511149
transform 1 0 12604 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_136
timestamp 1644511149
transform 1 0 13616 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_146
timestamp 1644511149
transform 1 0 14536 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_158
timestamp 1644511149
transform 1 0 15640 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_170
timestamp 1644511149
transform 1 0 16744 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1644511149
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_203
timestamp 1644511149
transform 1 0 19780 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_209
timestamp 1644511149
transform 1 0 20332 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_217
timestamp 1644511149
transform 1 0 21068 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_240
timestamp 1644511149
transform 1 0 23184 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_263
timestamp 1644511149
transform 1 0 25300 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_275
timestamp 1644511149
transform 1 0 26404 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_295
timestamp 1644511149
transform 1 0 28244 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_304
timestamp 1644511149
transform 1 0 29072 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_325
timestamp 1644511149
transform 1 0 31004 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_337
timestamp 1644511149
transform 1 0 32108 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_360
timestamp 1644511149
transform 1 0 34224 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_368
timestamp 1644511149
transform 1 0 34960 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_380
timestamp 1644511149
transform 1 0 36064 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_392
timestamp 1644511149
transform 1 0 37168 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_414
timestamp 1644511149
transform 1 0 39192 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_421
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_433
timestamp 1644511149
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_445
timestamp 1644511149
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_457
timestamp 1644511149
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1644511149
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1644511149
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_477
timestamp 1644511149
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_489
timestamp 1644511149
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_501
timestamp 1644511149
transform 1 0 47196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_512
timestamp 1644511149
transform 1 0 48208 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_74
timestamp 1644511149
transform 1 0 7912 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_99
timestamp 1644511149
transform 1 0 10212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_134
timestamp 1644511149
transform 1 0 13432 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_142
timestamp 1644511149
transform 1 0 14168 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_154
timestamp 1644511149
transform 1 0 15272 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1644511149
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_180
timestamp 1644511149
transform 1 0 17664 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_189
timestamp 1644511149
transform 1 0 18492 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_201
timestamp 1644511149
transform 1 0 19596 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_205
timestamp 1644511149
transform 1 0 19964 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_214
timestamp 1644511149
transform 1 0 20792 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1644511149
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_233
timestamp 1644511149
transform 1 0 22540 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_245
timestamp 1644511149
transform 1 0 23644 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_249
timestamp 1644511149
transform 1 0 24012 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_261
timestamp 1644511149
transform 1 0 25116 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_268
timestamp 1644511149
transform 1 0 25760 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_289
timestamp 1644511149
transform 1 0 27692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_301
timestamp 1644511149
transform 1 0 28796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_313
timestamp 1644511149
transform 1 0 29900 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_321
timestamp 1644511149
transform 1 0 30636 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_325
timestamp 1644511149
transform 1 0 31004 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_331
timestamp 1644511149
transform 1 0 31556 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1644511149
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_341
timestamp 1644511149
transform 1 0 32476 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_345
timestamp 1644511149
transform 1 0 32844 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_41_374
timestamp 1644511149
transform 1 0 35512 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_382
timestamp 1644511149
transform 1 0 36248 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_388
timestamp 1644511149
transform 1 0 36800 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_414
timestamp 1644511149
transform 1 0 39192 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_426
timestamp 1644511149
transform 1 0 40296 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_438
timestamp 1644511149
transform 1 0 41400 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_446
timestamp 1644511149
transform 1 0 42136 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_449
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_461
timestamp 1644511149
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_473
timestamp 1644511149
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_485
timestamp 1644511149
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1644511149
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1644511149
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_505
timestamp 1644511149
transform 1 0 47564 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_512
timestamp 1644511149
transform 1 0 48208 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1644511149
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_61
timestamp 1644511149
transform 1 0 6716 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_66
timestamp 1644511149
transform 1 0 7176 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_78
timestamp 1644511149
transform 1 0 8280 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_90
timestamp 1644511149
transform 1 0 9384 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_99
timestamp 1644511149
transform 1 0 10212 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_110
timestamp 1644511149
transform 1 0 11224 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_118
timestamp 1644511149
transform 1 0 11960 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_125
timestamp 1644511149
transform 1 0 12604 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_132
timestamp 1644511149
transform 1 0 13248 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_146
timestamp 1644511149
transform 1 0 14536 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_158
timestamp 1644511149
transform 1 0 15640 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_170
timestamp 1644511149
transform 1 0 16744 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_174
timestamp 1644511149
transform 1 0 17112 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_191
timestamp 1644511149
transform 1 0 18676 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1644511149
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_202
timestamp 1644511149
transform 1 0 19688 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_223
timestamp 1644511149
transform 1 0 21620 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_231
timestamp 1644511149
transform 1 0 22356 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_239
timestamp 1644511149
transform 1 0 23092 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_248
timestamp 1644511149
transform 1 0 23920 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_257
timestamp 1644511149
transform 1 0 24748 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_264
timestamp 1644511149
transform 1 0 25392 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_276
timestamp 1644511149
transform 1 0 26496 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_288
timestamp 1644511149
transform 1 0 27600 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_300
timestamp 1644511149
transform 1 0 28704 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_321
timestamp 1644511149
transform 1 0 30636 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_325
timestamp 1644511149
transform 1 0 31004 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_338
timestamp 1644511149
transform 1 0 32200 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_348
timestamp 1644511149
transform 1 0 33120 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_360
timestamp 1644511149
transform 1 0 34224 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_377
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_389
timestamp 1644511149
transform 1 0 36892 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_399
timestamp 1644511149
transform 1 0 37812 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_408
timestamp 1644511149
transform 1 0 38640 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_421
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_433
timestamp 1644511149
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_445
timestamp 1644511149
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_457
timestamp 1644511149
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1644511149
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1644511149
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_477
timestamp 1644511149
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_489
timestamp 1644511149
transform 1 0 46092 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_512
timestamp 1644511149
transform 1 0 48208 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_6
timestamp 1644511149
transform 1 0 1656 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_10
timestamp 1644511149
transform 1 0 2024 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_14
timestamp 1644511149
transform 1 0 2392 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_26
timestamp 1644511149
transform 1 0 3496 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_38
timestamp 1644511149
transform 1 0 4600 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_50
timestamp 1644511149
transform 1 0 5704 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_61
timestamp 1644511149
transform 1 0 6716 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_83
timestamp 1644511149
transform 1 0 8740 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_95
timestamp 1644511149
transform 1 0 9844 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_106
timestamp 1644511149
transform 1 0 10856 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_119
timestamp 1644511149
transform 1 0 12052 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_126
timestamp 1644511149
transform 1 0 12696 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_134
timestamp 1644511149
transform 1 0 13432 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_142
timestamp 1644511149
transform 1 0 14168 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_152
timestamp 1644511149
transform 1 0 15088 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1644511149
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_186
timestamp 1644511149
transform 1 0 18216 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_190
timestamp 1644511149
transform 1 0 18584 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_200
timestamp 1644511149
transform 1 0 19504 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_214
timestamp 1644511149
transform 1 0 20792 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1644511149
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_235
timestamp 1644511149
transform 1 0 22724 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_243
timestamp 1644511149
transform 1 0 23460 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_253
timestamp 1644511149
transform 1 0 24380 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_263
timestamp 1644511149
transform 1 0 25300 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_271
timestamp 1644511149
transform 1 0 26036 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_275
timestamp 1644511149
transform 1 0 26404 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1644511149
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_293
timestamp 1644511149
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_305
timestamp 1644511149
transform 1 0 29164 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_319
timestamp 1644511149
transform 1 0 30452 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_332
timestamp 1644511149
transform 1 0 31648 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_355
timestamp 1644511149
transform 1 0 33764 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_359
timestamp 1644511149
transform 1 0 34132 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_376
timestamp 1644511149
transform 1 0 35696 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_388
timestamp 1644511149
transform 1 0 36800 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_401
timestamp 1644511149
transform 1 0 37996 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_423
timestamp 1644511149
transform 1 0 40020 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_435
timestamp 1644511149
transform 1 0 41124 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1644511149
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_449
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_461
timestamp 1644511149
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_473
timestamp 1644511149
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_485
timestamp 1644511149
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_500
timestamp 1644511149
transform 1 0 47104 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_508
timestamp 1644511149
transform 1 0 47840 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_24
timestamp 1644511149
transform 1 0 3312 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_49
timestamp 1644511149
transform 1 0 5612 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_62
timestamp 1644511149
transform 1 0 6808 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_74
timestamp 1644511149
transform 1 0 7912 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_82
timestamp 1644511149
transform 1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_95
timestamp 1644511149
transform 1 0 9844 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_104
timestamp 1644511149
transform 1 0 10672 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_116
timestamp 1644511149
transform 1 0 11776 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_123
timestamp 1644511149
transform 1 0 12420 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_135
timestamp 1644511149
transform 1 0 13524 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_145
timestamp 1644511149
transform 1 0 14444 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_155
timestamp 1644511149
transform 1 0 15364 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_167
timestamp 1644511149
transform 1 0 16468 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_187
timestamp 1644511149
transform 1 0 18308 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1644511149
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_203
timestamp 1644511149
transform 1 0 19780 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_223
timestamp 1644511149
transform 1 0 21620 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_235
timestamp 1644511149
transform 1 0 22724 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_247
timestamp 1644511149
transform 1 0 23828 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1644511149
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_265
timestamp 1644511149
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_277
timestamp 1644511149
transform 1 0 26588 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_281
timestamp 1644511149
transform 1 0 26956 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_285
timestamp 1644511149
transform 1 0 27324 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_297
timestamp 1644511149
transform 1 0 28428 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_305
timestamp 1644511149
transform 1 0 29164 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_44_315
timestamp 1644511149
transform 1 0 30084 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_330
timestamp 1644511149
transform 1 0 31464 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_344
timestamp 1644511149
transform 1 0 32752 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_352
timestamp 1644511149
transform 1 0 33488 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_360
timestamp 1644511149
transform 1 0 34224 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_365
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_371
timestamp 1644511149
transform 1 0 35236 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_388
timestamp 1644511149
transform 1 0 36800 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_400
timestamp 1644511149
transform 1 0 37904 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_405
timestamp 1644511149
transform 1 0 38364 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1644511149
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1644511149
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_421
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_433
timestamp 1644511149
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_445
timestamp 1644511149
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_457
timestamp 1644511149
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1644511149
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1644511149
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_477
timestamp 1644511149
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_489
timestamp 1644511149
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_501
timestamp 1644511149
transform 1 0 47196 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_507
timestamp 1644511149
transform 1 0 47748 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_512
timestamp 1644511149
transform 1 0 48208 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_6
timestamp 1644511149
transform 1 0 1656 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_13
timestamp 1644511149
transform 1 0 2300 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_20
timestamp 1644511149
transform 1 0 2944 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_32
timestamp 1644511149
transform 1 0 4048 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_44
timestamp 1644511149
transform 1 0 5152 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_88
timestamp 1644511149
transform 1 0 9200 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_100
timestamp 1644511149
transform 1 0 10304 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_107
timestamp 1644511149
transform 1 0 10948 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_137
timestamp 1644511149
transform 1 0 13708 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_145
timestamp 1644511149
transform 1 0 14444 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_153
timestamp 1644511149
transform 1 0 15180 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_165
timestamp 1644511149
transform 1 0 16284 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_181
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_193
timestamp 1644511149
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_205
timestamp 1644511149
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1644511149
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1644511149
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_245
timestamp 1644511149
transform 1 0 23644 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_257
timestamp 1644511149
transform 1 0 24748 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_269
timestamp 1644511149
transform 1 0 25852 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_277
timestamp 1644511149
transform 1 0 26588 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_303
timestamp 1644511149
transform 1 0 28980 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_332
timestamp 1644511149
transform 1 0 31648 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_348
timestamp 1644511149
transform 1 0 33120 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_362
timestamp 1644511149
transform 1 0 34408 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_374
timestamp 1644511149
transform 1 0 35512 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_383
timestamp 1644511149
transform 1 0 36340 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1644511149
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_417
timestamp 1644511149
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_429
timestamp 1644511149
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1644511149
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1644511149
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_461
timestamp 1644511149
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_473
timestamp 1644511149
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_485
timestamp 1644511149
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1644511149
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1644511149
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_505
timestamp 1644511149
transform 1 0 47564 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_513
timestamp 1644511149
transform 1 0 48300 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_24
timestamp 1644511149
transform 1 0 3312 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_99
timestamp 1644511149
transform 1 0 10212 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_110
timestamp 1644511149
transform 1 0 11224 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_118
timestamp 1644511149
transform 1 0 11960 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_136
timestamp 1644511149
transform 1 0 13616 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_165
timestamp 1644511149
transform 1 0 16284 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_173
timestamp 1644511149
transform 1 0 17020 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_180
timestamp 1644511149
transform 1 0 17664 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1644511149
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_205
timestamp 1644511149
transform 1 0 19964 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_214
timestamp 1644511149
transform 1 0 20792 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_226
timestamp 1644511149
transform 1 0 21896 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_248
timestamp 1644511149
transform 1 0 23920 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_257
timestamp 1644511149
transform 1 0 24748 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_269
timestamp 1644511149
transform 1 0 25852 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_286
timestamp 1644511149
transform 1 0 27416 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_295
timestamp 1644511149
transform 1 0 28244 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_304
timestamp 1644511149
transform 1 0 29072 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_325
timestamp 1644511149
transform 1 0 31004 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_333
timestamp 1644511149
transform 1 0 31740 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_344
timestamp 1644511149
transform 1 0 32752 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_353
timestamp 1644511149
transform 1 0 33580 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_361
timestamp 1644511149
transform 1 0 34316 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_374
timestamp 1644511149
transform 1 0 35512 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_394
timestamp 1644511149
transform 1 0 37352 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_406
timestamp 1644511149
transform 1 0 38456 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_418
timestamp 1644511149
transform 1 0 39560 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_421
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_433
timestamp 1644511149
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_445
timestamp 1644511149
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_457
timestamp 1644511149
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1644511149
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1644511149
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_477
timestamp 1644511149
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_489
timestamp 1644511149
transform 1 0 46092 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_512
timestamp 1644511149
transform 1 0 48208 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_9
timestamp 1644511149
transform 1 0 1932 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_13
timestamp 1644511149
transform 1 0 2300 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_25
timestamp 1644511149
transform 1 0 3404 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_37
timestamp 1644511149
transform 1 0 4508 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_49
timestamp 1644511149
transform 1 0 5612 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_89
timestamp 1644511149
transform 1 0 9292 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_97
timestamp 1644511149
transform 1 0 10028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_109
timestamp 1644511149
transform 1 0 11132 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_120
timestamp 1644511149
transform 1 0 12144 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_131
timestamp 1644511149
transform 1 0 13156 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_143
timestamp 1644511149
transform 1 0 14260 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_151
timestamp 1644511149
transform 1 0 14996 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_164
timestamp 1644511149
transform 1 0 16192 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_172
timestamp 1644511149
transform 1 0 16928 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_183
timestamp 1644511149
transform 1 0 17940 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_191
timestamp 1644511149
transform 1 0 18676 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_203
timestamp 1644511149
transform 1 0 19780 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_220
timestamp 1644511149
transform 1 0 21344 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_237
timestamp 1644511149
transform 1 0 22908 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_259
timestamp 1644511149
transform 1 0 24932 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_267
timestamp 1644511149
transform 1 0 25668 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_276
timestamp 1644511149
transform 1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_297
timestamp 1644511149
transform 1 0 28428 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_303
timestamp 1644511149
transform 1 0 28980 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_312
timestamp 1644511149
transform 1 0 29808 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_324
timestamp 1644511149
transform 1 0 30912 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_341
timestamp 1644511149
transform 1 0 32476 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_358
timestamp 1644511149
transform 1 0 34040 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_366
timestamp 1644511149
transform 1 0 34776 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_376
timestamp 1644511149
transform 1 0 35696 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_388
timestamp 1644511149
transform 1 0 36800 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_405
timestamp 1644511149
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_417
timestamp 1644511149
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_429
timestamp 1644511149
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1644511149
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1644511149
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_449
timestamp 1644511149
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_461
timestamp 1644511149
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_473
timestamp 1644511149
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_485
timestamp 1644511149
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_500
timestamp 1644511149
transform 1 0 47104 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_47_505
timestamp 1644511149
transform 1 0 47564 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_512
timestamp 1644511149
transform 1 0 48208 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_24
timestamp 1644511149
transform 1 0 3312 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_61
timestamp 1644511149
transform 1 0 6716 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_80
timestamp 1644511149
transform 1 0 8464 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_93
timestamp 1644511149
transform 1 0 9660 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_101
timestamp 1644511149
transform 1 0 10396 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_113
timestamp 1644511149
transform 1 0 11500 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_125
timestamp 1644511149
transform 1 0 12604 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_137
timestamp 1644511149
transform 1 0 13708 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_148
timestamp 1644511149
transform 1 0 14720 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_156
timestamp 1644511149
transform 1 0 15456 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_163
timestamp 1644511149
transform 1 0 16100 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_183
timestamp 1644511149
transform 1 0 17940 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_192
timestamp 1644511149
transform 1 0 18768 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_205
timestamp 1644511149
transform 1 0 19964 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_211
timestamp 1644511149
transform 1 0 20516 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_223
timestamp 1644511149
transform 1 0 21620 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_235
timestamp 1644511149
transform 1 0 22724 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_241
timestamp 1644511149
transform 1 0 23276 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_249
timestamp 1644511149
transform 1 0 24012 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_265
timestamp 1644511149
transform 1 0 25484 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_272
timestamp 1644511149
transform 1 0 26128 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_285
timestamp 1644511149
transform 1 0 27324 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_297
timestamp 1644511149
transform 1 0 28428 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_305
timestamp 1644511149
transform 1 0 29164 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_321
timestamp 1644511149
transform 1 0 30636 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_330
timestamp 1644511149
transform 1 0 31464 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_350
timestamp 1644511149
transform 1 0 33304 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_359
timestamp 1644511149
transform 1 0 34132 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1644511149
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_375
timestamp 1644511149
transform 1 0 35604 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_382
timestamp 1644511149
transform 1 0 36248 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_407
timestamp 1644511149
transform 1 0 38548 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1644511149
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_421
timestamp 1644511149
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_433
timestamp 1644511149
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_445
timestamp 1644511149
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_457
timestamp 1644511149
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1644511149
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1644511149
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_477
timestamp 1644511149
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_489
timestamp 1644511149
transform 1 0 46092 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_512
timestamp 1644511149
transform 1 0 48208 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_7
timestamp 1644511149
transform 1 0 1748 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_11
timestamp 1644511149
transform 1 0 2116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_23
timestamp 1644511149
transform 1 0 3220 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_35
timestamp 1644511149
transform 1 0 4324 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_47
timestamp 1644511149
transform 1 0 5428 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_65
timestamp 1644511149
transform 1 0 7084 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_82
timestamp 1644511149
transform 1 0 8648 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_94
timestamp 1644511149
transform 1 0 9752 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_106
timestamp 1644511149
transform 1 0 10856 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_121
timestamp 1644511149
transform 1 0 12236 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_132
timestamp 1644511149
transform 1 0 13248 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_154
timestamp 1644511149
transform 1 0 15272 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_162
timestamp 1644511149
transform 1 0 16008 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_173
timestamp 1644511149
transform 1 0 17020 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_181
timestamp 1644511149
transform 1 0 17756 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_187
timestamp 1644511149
transform 1 0 18308 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_205
timestamp 1644511149
transform 1 0 19964 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_212
timestamp 1644511149
transform 1 0 20608 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_230
timestamp 1644511149
transform 1 0 22264 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_238
timestamp 1644511149
transform 1 0 23000 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_243
timestamp 1644511149
transform 1 0 23460 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_251
timestamp 1644511149
transform 1 0 24196 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_263
timestamp 1644511149
transform 1 0 25300 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_270
timestamp 1644511149
transform 1 0 25944 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_278
timestamp 1644511149
transform 1 0 26680 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_285
timestamp 1644511149
transform 1 0 27324 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_290
timestamp 1644511149
transform 1 0 27784 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_310
timestamp 1644511149
transform 1 0 29624 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_322
timestamp 1644511149
transform 1 0 30728 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_332
timestamp 1644511149
transform 1 0 31648 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_49_352
timestamp 1644511149
transform 1 0 33488 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_360
timestamp 1644511149
transform 1 0 34224 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_366
timestamp 1644511149
transform 1 0 34776 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_386
timestamp 1644511149
transform 1 0 36616 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_417
timestamp 1644511149
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_429
timestamp 1644511149
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1644511149
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1644511149
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_449
timestamp 1644511149
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_461
timestamp 1644511149
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_473
timestamp 1644511149
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_485
timestamp 1644511149
transform 1 0 45724 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_49_494
timestamp 1644511149
transform 1 0 46552 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_502
timestamp 1644511149
transform 1 0 47288 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_508
timestamp 1644511149
transform 1 0 47840 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_9
timestamp 1644511149
transform 1 0 1932 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_13
timestamp 1644511149
transform 1 0 2300 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_17
timestamp 1644511149
transform 1 0 2668 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_21
timestamp 1644511149
transform 1 0 3036 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_73
timestamp 1644511149
transform 1 0 7820 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_80
timestamp 1644511149
transform 1 0 8464 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_90
timestamp 1644511149
transform 1 0 9384 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_102
timestamp 1644511149
transform 1 0 10488 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_122
timestamp 1644511149
transform 1 0 12328 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_136
timestamp 1644511149
transform 1 0 13616 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_156
timestamp 1644511149
transform 1 0 15456 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_164
timestamp 1644511149
transform 1 0 16192 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_172
timestamp 1644511149
transform 1 0 16928 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_178
timestamp 1644511149
transform 1 0 17480 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_190
timestamp 1644511149
transform 1 0 18584 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_50_200
timestamp 1644511149
transform 1 0 19504 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_206
timestamp 1644511149
transform 1 0 20056 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_226
timestamp 1644511149
transform 1 0 21896 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_236
timestamp 1644511149
transform 1 0 22816 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_248
timestamp 1644511149
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_269
timestamp 1644511149
transform 1 0 25852 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_277
timestamp 1644511149
transform 1 0 26588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_282
timestamp 1644511149
transform 1 0 27048 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_291
timestamp 1644511149
transform 1 0 27876 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_299
timestamp 1644511149
transform 1 0 28612 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_304
timestamp 1644511149
transform 1 0 29072 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_318
timestamp 1644511149
transform 1 0 30360 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_330
timestamp 1644511149
transform 1 0 31464 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_339
timestamp 1644511149
transform 1 0 32292 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_351
timestamp 1644511149
transform 1 0 33396 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1644511149
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_374
timestamp 1644511149
transform 1 0 35512 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_386
timestamp 1644511149
transform 1 0 36616 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_398
timestamp 1644511149
transform 1 0 37720 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_410
timestamp 1644511149
transform 1 0 38824 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_418
timestamp 1644511149
transform 1 0 39560 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_421
timestamp 1644511149
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_433
timestamp 1644511149
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_445
timestamp 1644511149
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_457
timestamp 1644511149
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1644511149
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1644511149
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_477
timestamp 1644511149
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_489
timestamp 1644511149
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_501
timestamp 1644511149
transform 1 0 47196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_512
timestamp 1644511149
transform 1 0 48208 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_30
timestamp 1644511149
transform 1 0 3864 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_42
timestamp 1644511149
transform 1 0 4968 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_54
timestamp 1644511149
transform 1 0 6072 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_101
timestamp 1644511149
transform 1 0 10396 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_121
timestamp 1644511149
transform 1 0 12236 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_129
timestamp 1644511149
transform 1 0 12972 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_135
timestamp 1644511149
transform 1 0 13524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_141
timestamp 1644511149
transform 1 0 14076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_149
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_156
timestamp 1644511149
transform 1 0 15456 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_173
timestamp 1644511149
transform 1 0 17020 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_184
timestamp 1644511149
transform 1 0 18032 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_196
timestamp 1644511149
transform 1 0 19136 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_211
timestamp 1644511149
transform 1 0 20516 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_215
timestamp 1644511149
transform 1 0 20884 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_220
timestamp 1644511149
transform 1 0 21344 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_229
timestamp 1644511149
transform 1 0 22172 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_241
timestamp 1644511149
transform 1 0 23276 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_253
timestamp 1644511149
transform 1 0 24380 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_257
timestamp 1644511149
transform 1 0 24748 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_266
timestamp 1644511149
transform 1 0 25576 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_274
timestamp 1644511149
transform 1 0 26312 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_285
timestamp 1644511149
transform 1 0 27324 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_294
timestamp 1644511149
transform 1 0 28152 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_314
timestamp 1644511149
transform 1 0 29992 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_322
timestamp 1644511149
transform 1 0 30728 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_334
timestamp 1644511149
transform 1 0 31832 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_346
timestamp 1644511149
transform 1 0 32936 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_352
timestamp 1644511149
transform 1 0 33488 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_361
timestamp 1644511149
transform 1 0 34316 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_372
timestamp 1644511149
transform 1 0 35328 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_384
timestamp 1644511149
transform 1 0 36432 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_417
timestamp 1644511149
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_429
timestamp 1644511149
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1644511149
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1644511149
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_449
timestamp 1644511149
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_461
timestamp 1644511149
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_473
timestamp 1644511149
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_485
timestamp 1644511149
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1644511149
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1644511149
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_505
timestamp 1644511149
transform 1 0 47564 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_513
timestamp 1644511149
transform 1 0 48300 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_9
timestamp 1644511149
transform 1 0 1932 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_13
timestamp 1644511149
transform 1 0 2300 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_17
timestamp 1644511149
transform 1 0 2668 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_21
timestamp 1644511149
transform 1 0 3036 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_104
timestamp 1644511149
transform 1 0 10672 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_118
timestamp 1644511149
transform 1 0 11960 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_131
timestamp 1644511149
transform 1 0 13156 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_145
timestamp 1644511149
transform 1 0 14444 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_155
timestamp 1644511149
transform 1 0 15364 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_170
timestamp 1644511149
transform 1 0 16744 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_179
timestamp 1644511149
transform 1 0 17572 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_187
timestamp 1644511149
transform 1 0 18308 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1644511149
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_205
timestamp 1644511149
transform 1 0 19964 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_213
timestamp 1644511149
transform 1 0 20700 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_225
timestamp 1644511149
transform 1 0 21804 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_233
timestamp 1644511149
transform 1 0 22540 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_244
timestamp 1644511149
transform 1 0 23552 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_52_258
timestamp 1644511149
transform 1 0 24840 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_52_280
timestamp 1644511149
transform 1 0 26864 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_290
timestamp 1644511149
transform 1 0 27784 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_298
timestamp 1644511149
transform 1 0 28520 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_306
timestamp 1644511149
transform 1 0 29256 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_317
timestamp 1644511149
transform 1 0 30268 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_321
timestamp 1644511149
transform 1 0 30636 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_331
timestamp 1644511149
transform 1 0 31556 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_351
timestamp 1644511149
transform 1 0 33396 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1644511149
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_381
timestamp 1644511149
transform 1 0 36156 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_393
timestamp 1644511149
transform 1 0 37260 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_405
timestamp 1644511149
transform 1 0 38364 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_417
timestamp 1644511149
transform 1 0 39468 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_421
timestamp 1644511149
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_433
timestamp 1644511149
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_445
timestamp 1644511149
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_457
timestamp 1644511149
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1644511149
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1644511149
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_477
timestamp 1644511149
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_489
timestamp 1644511149
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_501
timestamp 1644511149
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_513
timestamp 1644511149
transform 1 0 48300 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_30
timestamp 1644511149
transform 1 0 3864 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_42
timestamp 1644511149
transform 1 0 4968 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_54
timestamp 1644511149
transform 1 0 6072 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_101
timestamp 1644511149
transform 1 0 10396 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_108
timestamp 1644511149
transform 1 0 11040 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_117
timestamp 1644511149
transform 1 0 11868 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_123
timestamp 1644511149
transform 1 0 12420 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_131
timestamp 1644511149
transform 1 0 13156 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_136
timestamp 1644511149
transform 1 0 13616 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_146
timestamp 1644511149
transform 1 0 14536 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_154
timestamp 1644511149
transform 1 0 15272 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_166
timestamp 1644511149
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_177
timestamp 1644511149
transform 1 0 17388 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_186
timestamp 1644511149
transform 1 0 18216 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_190
timestamp 1644511149
transform 1 0 18584 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_212
timestamp 1644511149
transform 1 0 20608 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_220
timestamp 1644511149
transform 1 0 21344 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_235
timestamp 1644511149
transform 1 0 22724 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_244
timestamp 1644511149
transform 1 0 23552 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_259
timestamp 1644511149
transform 1 0 24932 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_271
timestamp 1644511149
transform 1 0 26036 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1644511149
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_289
timestamp 1644511149
transform 1 0 27692 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_295
timestamp 1644511149
transform 1 0 28244 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_303
timestamp 1644511149
transform 1 0 28980 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_311
timestamp 1644511149
transform 1 0 29716 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_324
timestamp 1644511149
transform 1 0 30912 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_342
timestamp 1644511149
transform 1 0 32568 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_354
timestamp 1644511149
transform 1 0 33672 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_366
timestamp 1644511149
transform 1 0 34776 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_378
timestamp 1644511149
transform 1 0 35880 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_382
timestamp 1644511149
transform 1 0 36248 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_390
timestamp 1644511149
transform 1 0 36984 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_405
timestamp 1644511149
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_417
timestamp 1644511149
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_429
timestamp 1644511149
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1644511149
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1644511149
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_449
timestamp 1644511149
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_461
timestamp 1644511149
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_473
timestamp 1644511149
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_485
timestamp 1644511149
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1644511149
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1644511149
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_505
timestamp 1644511149
transform 1 0 47564 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_513
timestamp 1644511149
transform 1 0 48300 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_11
timestamp 1644511149
transform 1 0 2116 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_54_22
timestamp 1644511149
transform 1 0 3128 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_96
timestamp 1644511149
transform 1 0 9936 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_108
timestamp 1644511149
transform 1 0 11040 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_112
timestamp 1644511149
transform 1 0 11408 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_117
timestamp 1644511149
transform 1 0 11868 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_129
timestamp 1644511149
transform 1 0 12972 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_136
timestamp 1644511149
transform 1 0 13616 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_153
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_159
timestamp 1644511149
transform 1 0 15732 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_168
timestamp 1644511149
transform 1 0 16560 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_188
timestamp 1644511149
transform 1 0 18400 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_218
timestamp 1644511149
transform 1 0 21160 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_226
timestamp 1644511149
transform 1 0 21896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_235
timestamp 1644511149
transform 1 0 22724 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_247
timestamp 1644511149
transform 1 0 23828 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1644511149
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_259
timestamp 1644511149
transform 1 0 24932 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_263
timestamp 1644511149
transform 1 0 25300 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_280
timestamp 1644511149
transform 1 0 26864 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_300
timestamp 1644511149
transform 1 0 28704 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_313
timestamp 1644511149
transform 1 0 29900 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_320
timestamp 1644511149
transform 1 0 30544 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_329
timestamp 1644511149
transform 1 0 31372 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_341
timestamp 1644511149
transform 1 0 32476 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_345
timestamp 1644511149
transform 1 0 32844 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_355
timestamp 1644511149
transform 1 0 33764 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1644511149
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_377
timestamp 1644511149
transform 1 0 35788 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_400
timestamp 1644511149
transform 1 0 37904 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_412
timestamp 1644511149
transform 1 0 39008 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_421
timestamp 1644511149
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_433
timestamp 1644511149
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_445
timestamp 1644511149
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_457
timestamp 1644511149
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1644511149
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1644511149
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_477
timestamp 1644511149
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_489
timestamp 1644511149
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_501
timestamp 1644511149
transform 1 0 47196 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_507
timestamp 1644511149
transform 1 0 47748 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_512
timestamp 1644511149
transform 1 0 48208 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_9
timestamp 1644511149
transform 1 0 1932 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_31
timestamp 1644511149
transform 1 0 3956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_43
timestamp 1644511149
transform 1 0 5060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_97
timestamp 1644511149
transform 1 0 10028 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_106
timestamp 1644511149
transform 1 0 10856 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_122
timestamp 1644511149
transform 1 0 12328 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_133
timestamp 1644511149
transform 1 0 13340 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_146
timestamp 1644511149
transform 1 0 14536 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_155
timestamp 1644511149
transform 1 0 15364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_188
timestamp 1644511149
transform 1 0 18400 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_196
timestamp 1644511149
transform 1 0 19136 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_208
timestamp 1644511149
transform 1 0 20240 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_220
timestamp 1644511149
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_243
timestamp 1644511149
transform 1 0 23460 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_256
timestamp 1644511149
transform 1 0 24656 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_269
timestamp 1644511149
transform 1 0 25852 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_277
timestamp 1644511149
transform 1 0 26588 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_288
timestamp 1644511149
transform 1 0 27600 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_301
timestamp 1644511149
transform 1 0 28796 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_309
timestamp 1644511149
transform 1 0 29532 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_320
timestamp 1644511149
transform 1 0 30544 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1644511149
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1644511149
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_359
timestamp 1644511149
transform 1 0 34132 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_371
timestamp 1644511149
transform 1 0 35236 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_383
timestamp 1644511149
transform 1 0 36340 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1644511149
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_405
timestamp 1644511149
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_417
timestamp 1644511149
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_429
timestamp 1644511149
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1644511149
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1644511149
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_449
timestamp 1644511149
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_461
timestamp 1644511149
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_473
timestamp 1644511149
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_485
timestamp 1644511149
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1644511149
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1644511149
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_505
timestamp 1644511149
transform 1 0 47564 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_512
timestamp 1644511149
transform 1 0 48208 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_9
timestamp 1644511149
transform 1 0 1932 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_13
timestamp 1644511149
transform 1 0 2300 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_20
timestamp 1644511149
transform 1 0 2944 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_102
timestamp 1644511149
transform 1 0 10488 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_111
timestamp 1644511149
transform 1 0 11316 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_117
timestamp 1644511149
transform 1 0 11868 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_128
timestamp 1644511149
transform 1 0 12880 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_136
timestamp 1644511149
transform 1 0 13616 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_155
timestamp 1644511149
transform 1 0 15364 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_167
timestamp 1644511149
transform 1 0 16468 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_179
timestamp 1644511149
transform 1 0 17572 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_187
timestamp 1644511149
transform 1 0 18308 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_192
timestamp 1644511149
transform 1 0 18768 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_200
timestamp 1644511149
transform 1 0 19504 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_208
timestamp 1644511149
transform 1 0 20240 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_218
timestamp 1644511149
transform 1 0 21160 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_226
timestamp 1644511149
transform 1 0 21896 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1644511149
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1644511149
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_265
timestamp 1644511149
transform 1 0 25484 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_276
timestamp 1644511149
transform 1 0 26496 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_284
timestamp 1644511149
transform 1 0 27232 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_56_298
timestamp 1644511149
transform 1 0 28520 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_306
timestamp 1644511149
transform 1 0 29256 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_320
timestamp 1644511149
transform 1 0 30544 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_326
timestamp 1644511149
transform 1 0 31096 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_343
timestamp 1644511149
transform 1 0 32660 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_355
timestamp 1644511149
transform 1 0 33764 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1644511149
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_377
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_389
timestamp 1644511149
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_401
timestamp 1644511149
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1644511149
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1644511149
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_421
timestamp 1644511149
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_433
timestamp 1644511149
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_445
timestamp 1644511149
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_457
timestamp 1644511149
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1644511149
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1644511149
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_477
timestamp 1644511149
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_489
timestamp 1644511149
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_501
timestamp 1644511149
transform 1 0 47196 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_507
timestamp 1644511149
transform 1 0 47748 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_515
timestamp 1644511149
transform 1 0 48484 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_7
timestamp 1644511149
transform 1 0 1748 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_29
timestamp 1644511149
transform 1 0 3772 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_41
timestamp 1644511149
transform 1 0 4876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_53
timestamp 1644511149
transform 1 0 5980 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_77
timestamp 1644511149
transform 1 0 8188 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_95
timestamp 1644511149
transform 1 0 9844 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_99
timestamp 1644511149
transform 1 0 10212 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_108
timestamp 1644511149
transform 1 0 11040 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_122
timestamp 1644511149
transform 1 0 12328 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_130
timestamp 1644511149
transform 1 0 13064 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_139
timestamp 1644511149
transform 1 0 13892 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_159
timestamp 1644511149
transform 1 0 15732 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_173
timestamp 1644511149
transform 1 0 17020 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_179
timestamp 1644511149
transform 1 0 17572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_191
timestamp 1644511149
transform 1 0 18676 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_197
timestamp 1644511149
transform 1 0 19228 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_203
timestamp 1644511149
transform 1 0 19780 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_220
timestamp 1644511149
transform 1 0 21344 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_231
timestamp 1644511149
transform 1 0 22356 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_243
timestamp 1644511149
transform 1 0 23460 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_248
timestamp 1644511149
transform 1 0 23920 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_260
timestamp 1644511149
transform 1 0 25024 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_276
timestamp 1644511149
transform 1 0 26496 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_292
timestamp 1644511149
transform 1 0 27968 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_312
timestamp 1644511149
transform 1 0 29808 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_57_326
timestamp 1644511149
transform 1 0 31096 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_334
timestamp 1644511149
transform 1 0 31832 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_357
timestamp 1644511149
transform 1 0 33948 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_369
timestamp 1644511149
transform 1 0 35052 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_380
timestamp 1644511149
transform 1 0 36064 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_417
timestamp 1644511149
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_429
timestamp 1644511149
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1644511149
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1644511149
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_449
timestamp 1644511149
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_461
timestamp 1644511149
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_473
timestamp 1644511149
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_485
timestamp 1644511149
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_500
timestamp 1644511149
transform 1 0 47104 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_57_505
timestamp 1644511149
transform 1 0 47564 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_512
timestamp 1644511149
transform 1 0 48208 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_24
timestamp 1644511149
transform 1 0 3312 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_96
timestamp 1644511149
transform 1 0 9936 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_116
timestamp 1644511149
transform 1 0 11776 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_124
timestamp 1644511149
transform 1 0 12512 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_136
timestamp 1644511149
transform 1 0 13616 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_147
timestamp 1644511149
transform 1 0 14628 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_58_163
timestamp 1644511149
transform 1 0 16100 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_171
timestamp 1644511149
transform 1 0 16836 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_192
timestamp 1644511149
transform 1 0 18768 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_209
timestamp 1644511149
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_221
timestamp 1644511149
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_233
timestamp 1644511149
transform 1 0 22540 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_240
timestamp 1644511149
transform 1 0 23184 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_261
timestamp 1644511149
transform 1 0 25116 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_273
timestamp 1644511149
transform 1 0 26220 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_283
timestamp 1644511149
transform 1 0 27140 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_58_300
timestamp 1644511149
transform 1 0 28704 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_317
timestamp 1644511149
transform 1 0 30268 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_325
timestamp 1644511149
transform 1 0 31004 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_337
timestamp 1644511149
transform 1 0 32108 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_349
timestamp 1644511149
transform 1 0 33212 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_361
timestamp 1644511149
transform 1 0 34316 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_398
timestamp 1644511149
transform 1 0 37720 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_410
timestamp 1644511149
transform 1 0 38824 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_418
timestamp 1644511149
transform 1 0 39560 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_421
timestamp 1644511149
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_433
timestamp 1644511149
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_445
timestamp 1644511149
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_457
timestamp 1644511149
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1644511149
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1644511149
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_477
timestamp 1644511149
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_489
timestamp 1644511149
transform 1 0 46092 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_512
timestamp 1644511149
transform 1 0 48208 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_6
timestamp 1644511149
transform 1 0 1656 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_13
timestamp 1644511149
transform 1 0 2300 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_20
timestamp 1644511149
transform 1 0 2944 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_32
timestamp 1644511149
transform 1 0 4048 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_44
timestamp 1644511149
transform 1 0 5152 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_119
timestamp 1644511149
transform 1 0 12052 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_128
timestamp 1644511149
transform 1 0 12880 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_59_139
timestamp 1644511149
transform 1 0 13892 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_59_150
timestamp 1644511149
transform 1 0 14904 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_158
timestamp 1644511149
transform 1 0 15640 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_163
timestamp 1644511149
transform 1 0 16100 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_177
timestamp 1644511149
transform 1 0 17388 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_181
timestamp 1644511149
transform 1 0 17756 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_186
timestamp 1644511149
transform 1 0 18216 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_194
timestamp 1644511149
transform 1 0 18952 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_209
timestamp 1644511149
transform 1 0 20332 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_219
timestamp 1644511149
transform 1 0 21252 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_231
timestamp 1644511149
transform 1 0 22356 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_237
timestamp 1644511149
transform 1 0 22908 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_247
timestamp 1644511149
transform 1 0 23828 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_256
timestamp 1644511149
transform 1 0 24656 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_265
timestamp 1644511149
transform 1 0 25484 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_269
timestamp 1644511149
transform 1 0 25852 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_276
timestamp 1644511149
transform 1 0 26496 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_285
timestamp 1644511149
transform 1 0 27324 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_295
timestamp 1644511149
transform 1 0 28244 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_307
timestamp 1644511149
transform 1 0 29348 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_314
timestamp 1644511149
transform 1 0 29992 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_323
timestamp 1644511149
transform 1 0 30820 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1644511149
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_349
timestamp 1644511149
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_361
timestamp 1644511149
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_373
timestamp 1644511149
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1644511149
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1644511149
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_417
timestamp 1644511149
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_429
timestamp 1644511149
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1644511149
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1644511149
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_449
timestamp 1644511149
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_461
timestamp 1644511149
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_473
timestamp 1644511149
transform 1 0 44620 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_500
timestamp 1644511149
transform 1 0 47104 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_508
timestamp 1644511149
transform 1 0 47840 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_11
timestamp 1644511149
transform 1 0 2116 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_23
timestamp 1644511149
transform 1 0 3220 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_117
timestamp 1644511149
transform 1 0 11868 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_136
timestamp 1644511149
transform 1 0 13616 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_159
timestamp 1644511149
transform 1 0 15732 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_168
timestamp 1644511149
transform 1 0 16560 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_179
timestamp 1644511149
transform 1 0 17572 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_192
timestamp 1644511149
transform 1 0 18768 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_201
timestamp 1644511149
transform 1 0 19596 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_205
timestamp 1644511149
transform 1 0 19964 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_222
timestamp 1644511149
transform 1 0 21528 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_235
timestamp 1644511149
transform 1 0 22724 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_239
timestamp 1644511149
transform 1 0 23092 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_243
timestamp 1644511149
transform 1 0 23460 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1644511149
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_261
timestamp 1644511149
transform 1 0 25116 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_269
timestamp 1644511149
transform 1 0 25852 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_275
timestamp 1644511149
transform 1 0 26404 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_280
timestamp 1644511149
transform 1 0 26864 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_289
timestamp 1644511149
transform 1 0 27692 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_296
timestamp 1644511149
transform 1 0 28336 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_304
timestamp 1644511149
transform 1 0 29072 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_60_321
timestamp 1644511149
transform 1 0 30636 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_60_329
timestamp 1644511149
transform 1 0 31372 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_339
timestamp 1644511149
transform 1 0 32292 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_343
timestamp 1644511149
transform 1 0 32660 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_360
timestamp 1644511149
transform 1 0 34224 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_401
timestamp 1644511149
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1644511149
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1644511149
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_421
timestamp 1644511149
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_433
timestamp 1644511149
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_445
timestamp 1644511149
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_457
timestamp 1644511149
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1644511149
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1644511149
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_477
timestamp 1644511149
transform 1 0 44988 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_483
timestamp 1644511149
transform 1 0 45540 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_487
timestamp 1644511149
transform 1 0 45908 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_512
timestamp 1644511149
transform 1 0 48208 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_9
timestamp 1644511149
transform 1 0 1932 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_31
timestamp 1644511149
transform 1 0 3956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_43
timestamp 1644511149
transform 1 0 5060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1644511149
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_85
timestamp 1644511149
transform 1 0 8924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_89
timestamp 1644511149
transform 1 0 9292 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_101
timestamp 1644511149
transform 1 0 10396 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_109
timestamp 1644511149
transform 1 0 11132 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_155
timestamp 1644511149
transform 1 0 15364 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_164
timestamp 1644511149
transform 1 0 16192 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_187
timestamp 1644511149
transform 1 0 18308 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_195
timestamp 1644511149
transform 1 0 19044 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_208
timestamp 1644511149
transform 1 0 20240 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_220
timestamp 1644511149
transform 1 0 21344 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_228
timestamp 1644511149
transform 1 0 22080 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_236
timestamp 1644511149
transform 1 0 22816 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_245
timestamp 1644511149
transform 1 0 23644 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_255
timestamp 1644511149
transform 1 0 24564 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_259
timestamp 1644511149
transform 1 0 24932 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_269
timestamp 1644511149
transform 1 0 25852 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_276
timestamp 1644511149
transform 1 0 26496 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_293
timestamp 1644511149
transform 1 0 28060 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_298
timestamp 1644511149
transform 1 0 28520 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_306
timestamp 1644511149
transform 1 0 29256 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_315
timestamp 1644511149
transform 1 0 30084 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_328
timestamp 1644511149
transform 1 0 31280 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_353
timestamp 1644511149
transform 1 0 33580 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_365
timestamp 1644511149
transform 1 0 34684 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_377
timestamp 1644511149
transform 1 0 35788 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_389
timestamp 1644511149
transform 1 0 36892 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_417
timestamp 1644511149
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_429
timestamp 1644511149
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1644511149
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1644511149
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_449
timestamp 1644511149
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_461
timestamp 1644511149
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_473
timestamp 1644511149
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_485
timestamp 1644511149
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_500
timestamp 1644511149
transform 1 0 47104 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_61_505
timestamp 1644511149
transform 1 0 47564 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_512
timestamp 1644511149
transform 1 0 48208 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_15
timestamp 1644511149
transform 1 0 2484 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_19
timestamp 1644511149
transform 1 0 2852 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_23
timestamp 1644511149
transform 1 0 3220 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1644511149
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_115
timestamp 1644511149
transform 1 0 11684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_127
timestamp 1644511149
transform 1 0 12788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_149
timestamp 1644511149
transform 1 0 14812 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_168
timestamp 1644511149
transform 1 0 16560 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_180
timestamp 1644511149
transform 1 0 17664 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_192
timestamp 1644511149
transform 1 0 18768 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_201
timestamp 1644511149
transform 1 0 19596 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_205
timestamp 1644511149
transform 1 0 19964 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_227
timestamp 1644511149
transform 1 0 21988 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_241
timestamp 1644511149
transform 1 0 23276 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_249
timestamp 1644511149
transform 1 0 24012 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_257
timestamp 1644511149
transform 1 0 24748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_270
timestamp 1644511149
transform 1 0 25944 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_282
timestamp 1644511149
transform 1 0 27048 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_290
timestamp 1644511149
transform 1 0 27784 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_302
timestamp 1644511149
transform 1 0 28888 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_62_309
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_321
timestamp 1644511149
transform 1 0 30636 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_331
timestamp 1644511149
transform 1 0 31556 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_343
timestamp 1644511149
transform 1 0 32660 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_355
timestamp 1644511149
transform 1 0 33764 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1644511149
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_401
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1644511149
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1644511149
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_421
timestamp 1644511149
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_433
timestamp 1644511149
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_445
timestamp 1644511149
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_457
timestamp 1644511149
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1644511149
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1644511149
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_477
timestamp 1644511149
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_489
timestamp 1644511149
transform 1 0 46092 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_512
timestamp 1644511149
transform 1 0 48208 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_14
timestamp 1644511149
transform 1 0 2392 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_26
timestamp 1644511149
transform 1 0 3496 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_38
timestamp 1644511149
transform 1 0 4600 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_50
timestamp 1644511149
transform 1 0 5704 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_134
timestamp 1644511149
transform 1 0 13432 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_63_158
timestamp 1644511149
transform 1 0 15640 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_166
timestamp 1644511149
transform 1 0 16376 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_185
timestamp 1644511149
transform 1 0 18124 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_201
timestamp 1644511149
transform 1 0 19596 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_209
timestamp 1644511149
transform 1 0 20332 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_220
timestamp 1644511149
transform 1 0 21344 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_231
timestamp 1644511149
transform 1 0 22356 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_251
timestamp 1644511149
transform 1 0 24196 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_255
timestamp 1644511149
transform 1 0 24564 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_265
timestamp 1644511149
transform 1 0 25484 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_274
timestamp 1644511149
transform 1 0 26312 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_297
timestamp 1644511149
transform 1 0 28428 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_318
timestamp 1644511149
transform 1 0 30360 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_327
timestamp 1644511149
transform 1 0 31188 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1644511149
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_361
timestamp 1644511149
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1644511149
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_417
timestamp 1644511149
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_429
timestamp 1644511149
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1644511149
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1644511149
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_449
timestamp 1644511149
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_461
timestamp 1644511149
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_473
timestamp 1644511149
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_485
timestamp 1644511149
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1644511149
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1644511149
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_508
timestamp 1644511149
transform 1 0 47840 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_13
timestamp 1644511149
transform 1 0 2300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_25
timestamp 1644511149
transform 1 0 3404 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_106
timestamp 1644511149
transform 1 0 10856 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_118
timestamp 1644511149
transform 1 0 11960 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_130
timestamp 1644511149
transform 1 0 13064 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_138
timestamp 1644511149
transform 1 0 13800 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_149
timestamp 1644511149
transform 1 0 14812 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_173
timestamp 1644511149
transform 1 0 17020 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1644511149
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1644511149
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_213
timestamp 1644511149
transform 1 0 20700 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_233
timestamp 1644511149
transform 1 0 22540 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_248
timestamp 1644511149
transform 1 0 23920 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_261
timestamp 1644511149
transform 1 0 25116 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_275
timestamp 1644511149
transform 1 0 26404 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_295
timestamp 1644511149
transform 1 0 28244 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_304
timestamp 1644511149
transform 1 0 29072 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_315
timestamp 1644511149
transform 1 0 30084 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_325
timestamp 1644511149
transform 1 0 31004 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_329
timestamp 1644511149
transform 1 0 31372 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_346
timestamp 1644511149
transform 1 0 32936 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_358
timestamp 1644511149
transform 1 0 34040 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_377
timestamp 1644511149
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_389
timestamp 1644511149
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_401
timestamp 1644511149
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1644511149
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1644511149
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_421
timestamp 1644511149
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_433
timestamp 1644511149
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_445
timestamp 1644511149
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_457
timestamp 1644511149
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1644511149
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1644511149
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_477
timestamp 1644511149
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_489
timestamp 1644511149
transform 1 0 46092 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_497
timestamp 1644511149
transform 1 0 46828 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_503
timestamp 1644511149
transform 1 0 47380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_510
timestamp 1644511149
transform 1 0 48024 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_11
timestamp 1644511149
transform 1 0 2116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_23
timestamp 1644511149
transform 1 0 3220 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_35
timestamp 1644511149
transform 1 0 4324 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_47
timestamp 1644511149
transform 1 0 5428 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_88
timestamp 1644511149
transform 1 0 9200 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_100
timestamp 1644511149
transform 1 0 10304 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_149
timestamp 1644511149
transform 1 0 14812 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_157
timestamp 1644511149
transform 1 0 15548 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_164
timestamp 1644511149
transform 1 0 16192 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_185
timestamp 1644511149
transform 1 0 18124 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_205
timestamp 1644511149
transform 1 0 19964 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_218
timestamp 1644511149
transform 1 0 21160 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_233
timestamp 1644511149
transform 1 0 22540 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_237
timestamp 1644511149
transform 1 0 22908 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_243
timestamp 1644511149
transform 1 0 23460 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_255
timestamp 1644511149
transform 1 0 24564 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_263
timestamp 1644511149
transform 1 0 25300 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_269
timestamp 1644511149
transform 1 0 25852 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_277
timestamp 1644511149
transform 1 0 26588 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_65_281
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_289
timestamp 1644511149
transform 1 0 27692 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_299
timestamp 1644511149
transform 1 0 28612 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_312
timestamp 1644511149
transform 1 0 29808 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_320
timestamp 1644511149
transform 1 0 30544 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1644511149
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1644511149
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_353
timestamp 1644511149
transform 1 0 33580 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_365
timestamp 1644511149
transform 1 0 34684 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_377
timestamp 1644511149
transform 1 0 35788 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_389
timestamp 1644511149
transform 1 0 36892 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_393
timestamp 1644511149
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_405
timestamp 1644511149
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_417
timestamp 1644511149
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_429
timestamp 1644511149
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1644511149
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1644511149
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_449
timestamp 1644511149
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_461
timestamp 1644511149
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_473
timestamp 1644511149
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_485
timestamp 1644511149
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1644511149
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1644511149
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_65_505
timestamp 1644511149
transform 1 0 47564 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_512
timestamp 1644511149
transform 1 0 48208 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_15
timestamp 1644511149
transform 1 0 2484 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_22
timestamp 1644511149
transform 1 0 3128 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1644511149
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_157
timestamp 1644511149
transform 1 0 15548 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_161
timestamp 1644511149
transform 1 0 15916 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_186
timestamp 1644511149
transform 1 0 18216 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_194
timestamp 1644511149
transform 1 0 18952 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_218
timestamp 1644511149
transform 1 0 21160 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_222
timestamp 1644511149
transform 1 0 21528 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_227
timestamp 1644511149
transform 1 0 21988 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_237
timestamp 1644511149
transform 1 0 22908 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_247
timestamp 1644511149
transform 1 0 23828 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1644511149
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_253
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_265
timestamp 1644511149
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_277
timestamp 1644511149
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_289
timestamp 1644511149
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1644511149
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1644511149
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_325
timestamp 1644511149
transform 1 0 31004 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_337
timestamp 1644511149
transform 1 0 32108 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_349
timestamp 1644511149
transform 1 0 33212 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_361
timestamp 1644511149
transform 1 0 34316 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_365
timestamp 1644511149
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_377
timestamp 1644511149
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_389
timestamp 1644511149
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_401
timestamp 1644511149
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1644511149
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1644511149
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_421
timestamp 1644511149
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_433
timestamp 1644511149
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_445
timestamp 1644511149
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_457
timestamp 1644511149
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1644511149
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1644511149
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_477
timestamp 1644511149
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_489
timestamp 1644511149
transform 1 0 46092 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_512
timestamp 1644511149
transform 1 0 48208 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_9
timestamp 1644511149
transform 1 0 1932 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_31
timestamp 1644511149
transform 1 0 3956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_43
timestamp 1644511149
transform 1 0 5060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1644511149
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1644511149
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_149
timestamp 1644511149
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1644511149
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1644511149
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_173
timestamp 1644511149
transform 1 0 17020 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_180
timestamp 1644511149
transform 1 0 17664 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_188
timestamp 1644511149
transform 1 0 18400 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_198
timestamp 1644511149
transform 1 0 19320 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_202
timestamp 1644511149
transform 1 0 19688 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_206
timestamp 1644511149
transform 1 0 20056 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_218
timestamp 1644511149
transform 1 0 21160 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_225
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_229
timestamp 1644511149
transform 1 0 22172 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_236
timestamp 1644511149
transform 1 0 22816 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_248
timestamp 1644511149
transform 1 0 23920 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_276
timestamp 1644511149
transform 1 0 26496 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_289
timestamp 1644511149
transform 1 0 27692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_301
timestamp 1644511149
transform 1 0 28796 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_313
timestamp 1644511149
transform 1 0 29900 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_317
timestamp 1644511149
transform 1 0 30268 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_323
timestamp 1644511149
transform 1 0 30820 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1644511149
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_337
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_349
timestamp 1644511149
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_361
timestamp 1644511149
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_373
timestamp 1644511149
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1644511149
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1644511149
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_393
timestamp 1644511149
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_405
timestamp 1644511149
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_417
timestamp 1644511149
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_429
timestamp 1644511149
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1644511149
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1644511149
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_449
timestamp 1644511149
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_461
timestamp 1644511149
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_473
timestamp 1644511149
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_485
timestamp 1644511149
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1644511149
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1644511149
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_67_505
timestamp 1644511149
transform 1 0 47564 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_512
timestamp 1644511149
transform 1 0 48208 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_3
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_9
timestamp 1644511149
transform 1 0 1932 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_13
timestamp 1644511149
transform 1 0 2300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_25
timestamp 1644511149
transform 1 0 3404 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_41
timestamp 1644511149
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_53
timestamp 1644511149
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_65
timestamp 1644511149
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1644511149
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1644511149
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_109
timestamp 1644511149
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_121
timestamp 1644511149
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1644511149
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1644511149
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1644511149
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_165
timestamp 1644511149
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_181
timestamp 1644511149
transform 1 0 17756 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_68_190
timestamp 1644511149
transform 1 0 18584 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_68_197
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_209
timestamp 1644511149
transform 1 0 20332 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_226
timestamp 1644511149
transform 1 0 21896 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_238
timestamp 1644511149
transform 1 0 23000 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_247
timestamp 1644511149
transform 1 0 23828 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1644511149
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_269
timestamp 1644511149
transform 1 0 25852 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_277
timestamp 1644511149
transform 1 0 26588 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_296
timestamp 1644511149
transform 1 0 28336 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_321
timestamp 1644511149
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_333
timestamp 1644511149
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_345
timestamp 1644511149
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1644511149
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1644511149
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_365
timestamp 1644511149
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_377
timestamp 1644511149
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_389
timestamp 1644511149
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_401
timestamp 1644511149
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1644511149
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1644511149
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_421
timestamp 1644511149
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_433
timestamp 1644511149
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_445
timestamp 1644511149
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_457
timestamp 1644511149
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1644511149
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1644511149
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_477
timestamp 1644511149
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_489
timestamp 1644511149
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_501
timestamp 1644511149
transform 1 0 47196 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_68_507
timestamp 1644511149
transform 1 0 47748 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_515
timestamp 1644511149
transform 1 0 48484 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1644511149
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1644511149
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_39
timestamp 1644511149
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1644511149
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1644511149
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1644511149
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1644511149
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_93
timestamp 1644511149
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1644511149
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1644511149
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_113
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_125
timestamp 1644511149
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_137
timestamp 1644511149
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_149
timestamp 1644511149
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1644511149
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1644511149
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_169
timestamp 1644511149
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_181
timestamp 1644511149
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_193
timestamp 1644511149
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_205
timestamp 1644511149
transform 1 0 19964 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_213
timestamp 1644511149
transform 1 0 20700 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_220
timestamp 1644511149
transform 1 0 21344 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_241
timestamp 1644511149
transform 1 0 23276 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_261
timestamp 1644511149
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1644511149
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1644511149
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_281
timestamp 1644511149
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_293
timestamp 1644511149
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_305
timestamp 1644511149
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_317
timestamp 1644511149
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1644511149
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1644511149
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_337
timestamp 1644511149
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_349
timestamp 1644511149
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_361
timestamp 1644511149
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_373
timestamp 1644511149
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1644511149
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1644511149
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_393
timestamp 1644511149
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_405
timestamp 1644511149
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_417
timestamp 1644511149
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_429
timestamp 1644511149
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1644511149
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1644511149
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_449
timestamp 1644511149
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_461
timestamp 1644511149
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_473
timestamp 1644511149
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_485
timestamp 1644511149
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1644511149
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1644511149
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_508
timestamp 1644511149
transform 1 0 47840 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_7
timestamp 1644511149
transform 1 0 1748 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_19
timestamp 1644511149
transform 1 0 2852 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1644511149
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1644511149
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1644511149
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1644511149
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1644511149
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1644511149
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_97
timestamp 1644511149
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_109
timestamp 1644511149
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_121
timestamp 1644511149
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1644511149
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1644511149
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_153
timestamp 1644511149
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_165
timestamp 1644511149
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_177
timestamp 1644511149
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1644511149
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1644511149
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_197
timestamp 1644511149
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_209
timestamp 1644511149
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_221
timestamp 1644511149
transform 1 0 21436 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_229
timestamp 1644511149
transform 1 0 22172 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_239
timestamp 1644511149
transform 1 0 23092 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1644511149
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_253
timestamp 1644511149
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_265
timestamp 1644511149
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_277
timestamp 1644511149
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_289
timestamp 1644511149
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1644511149
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1644511149
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_309
timestamp 1644511149
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_321
timestamp 1644511149
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_333
timestamp 1644511149
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_345
timestamp 1644511149
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1644511149
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1644511149
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_365
timestamp 1644511149
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_377
timestamp 1644511149
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_389
timestamp 1644511149
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_401
timestamp 1644511149
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1644511149
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1644511149
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_421
timestamp 1644511149
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_433
timestamp 1644511149
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_445
timestamp 1644511149
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_457
timestamp 1644511149
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1644511149
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1644511149
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_477
timestamp 1644511149
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_489
timestamp 1644511149
transform 1 0 46092 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_512
timestamp 1644511149
transform 1 0 48208 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_3
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_11
timestamp 1644511149
transform 1 0 2116 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_18
timestamp 1644511149
transform 1 0 2760 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_30
timestamp 1644511149
transform 1 0 3864 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_42
timestamp 1644511149
transform 1 0 4968 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_54
timestamp 1644511149
transform 1 0 6072 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1644511149
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_93
timestamp 1644511149
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1644511149
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1644511149
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_125
timestamp 1644511149
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_137
timestamp 1644511149
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_149
timestamp 1644511149
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1644511149
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1644511149
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_169
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_181
timestamp 1644511149
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_193
timestamp 1644511149
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_205
timestamp 1644511149
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1644511149
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1644511149
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_225
timestamp 1644511149
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_237
timestamp 1644511149
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_249
timestamp 1644511149
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_261
timestamp 1644511149
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1644511149
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1644511149
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_281
timestamp 1644511149
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_293
timestamp 1644511149
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_305
timestamp 1644511149
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_317
timestamp 1644511149
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1644511149
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1644511149
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_337
timestamp 1644511149
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_349
timestamp 1644511149
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_361
timestamp 1644511149
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_373
timestamp 1644511149
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1644511149
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1644511149
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_393
timestamp 1644511149
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_405
timestamp 1644511149
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_417
timestamp 1644511149
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_429
timestamp 1644511149
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1644511149
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1644511149
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_449
timestamp 1644511149
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_461
timestamp 1644511149
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_473
timestamp 1644511149
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_485
timestamp 1644511149
transform 1 0 45724 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_489
timestamp 1644511149
transform 1 0 46092 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_500
timestamp 1644511149
transform 1 0 47104 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_508
timestamp 1644511149
transform 1 0 47840 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_72_24
timestamp 1644511149
transform 1 0 3312 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1644511149
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1644511149
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1644511149
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1644511149
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1644511149
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1644511149
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_97
timestamp 1644511149
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_109
timestamp 1644511149
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_121
timestamp 1644511149
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1644511149
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1644511149
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1644511149
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_153
timestamp 1644511149
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_165
timestamp 1644511149
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_177
timestamp 1644511149
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1644511149
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1644511149
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_197
timestamp 1644511149
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_209
timestamp 1644511149
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_221
timestamp 1644511149
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_233
timestamp 1644511149
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1644511149
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1644511149
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_253
timestamp 1644511149
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_265
timestamp 1644511149
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_277
timestamp 1644511149
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_289
timestamp 1644511149
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1644511149
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1644511149
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_309
timestamp 1644511149
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_321
timestamp 1644511149
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_333
timestamp 1644511149
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_345
timestamp 1644511149
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1644511149
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1644511149
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_365
timestamp 1644511149
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_377
timestamp 1644511149
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_389
timestamp 1644511149
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_401
timestamp 1644511149
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1644511149
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1644511149
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_421
timestamp 1644511149
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_433
timestamp 1644511149
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_445
timestamp 1644511149
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_457
timestamp 1644511149
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1644511149
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1644511149
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_477
timestamp 1644511149
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_489
timestamp 1644511149
transform 1 0 46092 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_512
timestamp 1644511149
transform 1 0 48208 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_3
timestamp 1644511149
transform 1 0 1380 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_7
timestamp 1644511149
transform 1 0 1748 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_11
timestamp 1644511149
transform 1 0 2116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_23
timestamp 1644511149
transform 1 0 3220 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_35
timestamp 1644511149
transform 1 0 4324 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_47
timestamp 1644511149
transform 1 0 5428 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1644511149
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1644511149
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_93
timestamp 1644511149
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1644511149
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1644511149
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1644511149
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1644511149
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_137
timestamp 1644511149
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_149
timestamp 1644511149
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1644511149
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1644511149
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_169
timestamp 1644511149
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_181
timestamp 1644511149
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_193
timestamp 1644511149
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_205
timestamp 1644511149
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1644511149
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1644511149
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_225
timestamp 1644511149
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_237
timestamp 1644511149
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_249
timestamp 1644511149
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_261
timestamp 1644511149
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1644511149
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1644511149
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_281
timestamp 1644511149
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_293
timestamp 1644511149
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_305
timestamp 1644511149
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_317
timestamp 1644511149
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1644511149
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1644511149
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_337
timestamp 1644511149
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_349
timestamp 1644511149
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_361
timestamp 1644511149
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_373
timestamp 1644511149
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1644511149
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1644511149
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_393
timestamp 1644511149
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_405
timestamp 1644511149
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_417
timestamp 1644511149
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_429
timestamp 1644511149
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1644511149
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1644511149
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_449
timestamp 1644511149
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_461
timestamp 1644511149
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_473
timestamp 1644511149
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_485
timestamp 1644511149
transform 1 0 45724 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_493
timestamp 1644511149
transform 1 0 46460 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_499
timestamp 1644511149
transform 1 0 47012 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1644511149
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_508
timestamp 1644511149
transform 1 0 47840 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1644511149
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1644511149
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1644511149
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1644511149
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1644511149
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_53
timestamp 1644511149
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_65
timestamp 1644511149
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1644511149
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1644511149
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_85
timestamp 1644511149
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_97
timestamp 1644511149
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_109
timestamp 1644511149
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_121
timestamp 1644511149
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1644511149
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1644511149
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1644511149
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_153
timestamp 1644511149
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_165
timestamp 1644511149
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_177
timestamp 1644511149
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1644511149
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1644511149
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_197
timestamp 1644511149
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_209
timestamp 1644511149
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_221
timestamp 1644511149
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_233
timestamp 1644511149
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1644511149
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1644511149
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_253
timestamp 1644511149
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_265
timestamp 1644511149
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_277
timestamp 1644511149
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_289
timestamp 1644511149
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1644511149
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1644511149
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_309
timestamp 1644511149
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_321
timestamp 1644511149
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_333
timestamp 1644511149
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_345
timestamp 1644511149
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1644511149
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1644511149
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_365
timestamp 1644511149
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_377
timestamp 1644511149
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_389
timestamp 1644511149
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_401
timestamp 1644511149
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1644511149
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1644511149
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_421
timestamp 1644511149
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_433
timestamp 1644511149
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_445
timestamp 1644511149
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_457
timestamp 1644511149
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1644511149
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1644511149
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_477
timestamp 1644511149
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_489
timestamp 1644511149
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_504
timestamp 1644511149
transform 1 0 47472 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_512
timestamp 1644511149
transform 1 0 48208 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_3
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_13
timestamp 1644511149
transform 1 0 2300 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_25
timestamp 1644511149
transform 1 0 3404 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_37
timestamp 1644511149
transform 1 0 4508 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_49
timestamp 1644511149
transform 1 0 5612 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1644511149
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1644511149
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1644511149
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_93
timestamp 1644511149
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1644511149
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1644511149
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_113
timestamp 1644511149
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_125
timestamp 1644511149
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_137
timestamp 1644511149
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_149
timestamp 1644511149
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1644511149
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1644511149
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_169
timestamp 1644511149
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_181
timestamp 1644511149
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_193
timestamp 1644511149
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_205
timestamp 1644511149
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1644511149
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1644511149
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_225
timestamp 1644511149
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_237
timestamp 1644511149
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_249
timestamp 1644511149
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_261
timestamp 1644511149
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1644511149
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1644511149
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_281
timestamp 1644511149
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_293
timestamp 1644511149
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_305
timestamp 1644511149
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_317
timestamp 1644511149
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1644511149
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1644511149
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_337
timestamp 1644511149
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_349
timestamp 1644511149
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_361
timestamp 1644511149
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_373
timestamp 1644511149
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1644511149
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1644511149
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_393
timestamp 1644511149
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_405
timestamp 1644511149
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_417
timestamp 1644511149
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_429
timestamp 1644511149
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1644511149
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1644511149
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_449
timestamp 1644511149
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_461
timestamp 1644511149
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_473
timestamp 1644511149
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_485
timestamp 1644511149
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_500
timestamp 1644511149
transform 1 0 47104 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_75_505
timestamp 1644511149
transform 1 0 47564 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_512
timestamp 1644511149
transform 1 0 48208 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_3
timestamp 1644511149
transform 1 0 1380 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_13
timestamp 1644511149
transform 1 0 2300 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_20
timestamp 1644511149
transform 1 0 2944 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1644511149
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1644511149
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1644511149
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_65
timestamp 1644511149
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1644511149
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1644511149
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_85
timestamp 1644511149
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_97
timestamp 1644511149
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_109
timestamp 1644511149
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_121
timestamp 1644511149
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1644511149
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1644511149
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_141
timestamp 1644511149
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_153
timestamp 1644511149
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_165
timestamp 1644511149
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_177
timestamp 1644511149
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1644511149
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1644511149
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_197
timestamp 1644511149
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_209
timestamp 1644511149
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_221
timestamp 1644511149
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_233
timestamp 1644511149
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1644511149
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1644511149
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_253
timestamp 1644511149
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_265
timestamp 1644511149
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_277
timestamp 1644511149
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_289
timestamp 1644511149
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1644511149
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1644511149
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_309
timestamp 1644511149
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_321
timestamp 1644511149
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_333
timestamp 1644511149
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_345
timestamp 1644511149
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1644511149
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1644511149
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_365
timestamp 1644511149
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_377
timestamp 1644511149
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_389
timestamp 1644511149
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_401
timestamp 1644511149
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1644511149
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1644511149
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_421
timestamp 1644511149
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_433
timestamp 1644511149
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_445
timestamp 1644511149
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_457
timestamp 1644511149
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1644511149
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1644511149
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_477
timestamp 1644511149
transform 1 0 44988 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_483
timestamp 1644511149
transform 1 0 45540 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_487
timestamp 1644511149
transform 1 0 45908 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_512
timestamp 1644511149
transform 1 0 48208 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_3
timestamp 1644511149
transform 1 0 1380 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_7
timestamp 1644511149
transform 1 0 1748 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_29
timestamp 1644511149
transform 1 0 3772 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_41
timestamp 1644511149
transform 1 0 4876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_53
timestamp 1644511149
transform 1 0 5980 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1644511149
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1644511149
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1644511149
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_93
timestamp 1644511149
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1644511149
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1644511149
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_113
timestamp 1644511149
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_125
timestamp 1644511149
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_137
timestamp 1644511149
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_149
timestamp 1644511149
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1644511149
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1644511149
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_169
timestamp 1644511149
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_181
timestamp 1644511149
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_193
timestamp 1644511149
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_205
timestamp 1644511149
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1644511149
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1644511149
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_225
timestamp 1644511149
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_237
timestamp 1644511149
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_249
timestamp 1644511149
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_261
timestamp 1644511149
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1644511149
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1644511149
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_281
timestamp 1644511149
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_293
timestamp 1644511149
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_305
timestamp 1644511149
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_317
timestamp 1644511149
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1644511149
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1644511149
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_337
timestamp 1644511149
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_349
timestamp 1644511149
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_361
timestamp 1644511149
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_373
timestamp 1644511149
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1644511149
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1644511149
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_393
timestamp 1644511149
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_405
timestamp 1644511149
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_417
timestamp 1644511149
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_429
timestamp 1644511149
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1644511149
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1644511149
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_449
timestamp 1644511149
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_461
timestamp 1644511149
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_473
timestamp 1644511149
transform 1 0 44620 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_77_500
timestamp 1644511149
transform 1 0 47104 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_508
timestamp 1644511149
transform 1 0 47840 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_78_24
timestamp 1644511149
transform 1 0 3312 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_32
timestamp 1644511149
transform 1 0 4048 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_44
timestamp 1644511149
transform 1 0 5152 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_56
timestamp 1644511149
transform 1 0 6256 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_68
timestamp 1644511149
transform 1 0 7360 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_80
timestamp 1644511149
transform 1 0 8464 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_85
timestamp 1644511149
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_97
timestamp 1644511149
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_109
timestamp 1644511149
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_121
timestamp 1644511149
transform 1 0 12236 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_78_132
timestamp 1644511149
transform 1 0 13248 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1644511149
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_153
timestamp 1644511149
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_165
timestamp 1644511149
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_177
timestamp 1644511149
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1644511149
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1644511149
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_197
timestamp 1644511149
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_209
timestamp 1644511149
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_221
timestamp 1644511149
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_233
timestamp 1644511149
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1644511149
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1644511149
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_253
timestamp 1644511149
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_265
timestamp 1644511149
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_277
timestamp 1644511149
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_289
timestamp 1644511149
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1644511149
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1644511149
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_309
timestamp 1644511149
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_321
timestamp 1644511149
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_333
timestamp 1644511149
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_345
timestamp 1644511149
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1644511149
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1644511149
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_365
timestamp 1644511149
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_377
timestamp 1644511149
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_389
timestamp 1644511149
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_401
timestamp 1644511149
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1644511149
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1644511149
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_421
timestamp 1644511149
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_433
timestamp 1644511149
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_445
timestamp 1644511149
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_457
timestamp 1644511149
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1644511149
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1644511149
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_480
timestamp 1644511149
transform 1 0 45264 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_487
timestamp 1644511149
transform 1 0 45908 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_512
timestamp 1644511149
transform 1 0 48208 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_6
timestamp 1644511149
transform 1 0 1656 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_13
timestamp 1644511149
transform 1 0 2300 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_38
timestamp 1644511149
transform 1 0 4600 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_50
timestamp 1644511149
transform 1 0 5704 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1644511149
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1644511149
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_81
timestamp 1644511149
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_93
timestamp 1644511149
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1644511149
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1644511149
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_113
timestamp 1644511149
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_125
timestamp 1644511149
transform 1 0 12604 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_149
timestamp 1644511149
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1644511149
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1644511149
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_169
timestamp 1644511149
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_181
timestamp 1644511149
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_202
timestamp 1644511149
transform 1 0 19688 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_214
timestamp 1644511149
transform 1 0 20792 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_222
timestamp 1644511149
transform 1 0 21528 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_225
timestamp 1644511149
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_237
timestamp 1644511149
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_249
timestamp 1644511149
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_261
timestamp 1644511149
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1644511149
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1644511149
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_281
timestamp 1644511149
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_293
timestamp 1644511149
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_305
timestamp 1644511149
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_317
timestamp 1644511149
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1644511149
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1644511149
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_337
timestamp 1644511149
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_349
timestamp 1644511149
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_361
timestamp 1644511149
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_373
timestamp 1644511149
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1644511149
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1644511149
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_393
timestamp 1644511149
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_405
timestamp 1644511149
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_417
timestamp 1644511149
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_429
timestamp 1644511149
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1644511149
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1644511149
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_449
timestamp 1644511149
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_461
timestamp 1644511149
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_476
timestamp 1644511149
transform 1 0 44896 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_483
timestamp 1644511149
transform 1 0 45540 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_489
timestamp 1644511149
transform 1 0 46092 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_493
timestamp 1644511149
transform 1 0 46460 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_500
timestamp 1644511149
transform 1 0 47104 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_508
timestamp 1644511149
transform 1 0 47840 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_80_7
timestamp 1644511149
transform 1 0 1748 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_13
timestamp 1644511149
transform 1 0 2300 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_17
timestamp 1644511149
transform 1 0 2668 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_24
timestamp 1644511149
transform 1 0 3312 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_32
timestamp 1644511149
transform 1 0 4048 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_44
timestamp 1644511149
transform 1 0 5152 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_56
timestamp 1644511149
transform 1 0 6256 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_68
timestamp 1644511149
transform 1 0 7360 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_80
timestamp 1644511149
transform 1 0 8464 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_85
timestamp 1644511149
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_97
timestamp 1644511149
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_109
timestamp 1644511149
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_121
timestamp 1644511149
transform 1 0 12236 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_129
timestamp 1644511149
transform 1 0 12972 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_135
timestamp 1644511149
transform 1 0 13524 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1644511149
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_141
timestamp 1644511149
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_153
timestamp 1644511149
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_165
timestamp 1644511149
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_177
timestamp 1644511149
transform 1 0 17388 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_185
timestamp 1644511149
transform 1 0 18124 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_192
timestamp 1644511149
transform 1 0 18768 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_209
timestamp 1644511149
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_221
timestamp 1644511149
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_233
timestamp 1644511149
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1644511149
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1644511149
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_253
timestamp 1644511149
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_265
timestamp 1644511149
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_277
timestamp 1644511149
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_289
timestamp 1644511149
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1644511149
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1644511149
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_309
timestamp 1644511149
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_321
timestamp 1644511149
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_333
timestamp 1644511149
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_345
timestamp 1644511149
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1644511149
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1644511149
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_365
timestamp 1644511149
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_377
timestamp 1644511149
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_389
timestamp 1644511149
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_401
timestamp 1644511149
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_413
timestamp 1644511149
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1644511149
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_421
timestamp 1644511149
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_433
timestamp 1644511149
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_445
timestamp 1644511149
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_457
timestamp 1644511149
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_472
timestamp 1644511149
transform 1 0 44528 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_477
timestamp 1644511149
transform 1 0 44988 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_481
timestamp 1644511149
transform 1 0 45356 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_489
timestamp 1644511149
transform 1 0 46092 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_512
timestamp 1644511149
transform 1 0 48208 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_3
timestamp 1644511149
transform 1 0 1380 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_81_30
timestamp 1644511149
transform 1 0 3864 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_42
timestamp 1644511149
transform 1 0 4968 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_54
timestamp 1644511149
transform 1 0 6072 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1644511149
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_69
timestamp 1644511149
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_81
timestamp 1644511149
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_93
timestamp 1644511149
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1644511149
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1644511149
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_113
timestamp 1644511149
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_125
timestamp 1644511149
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_137
timestamp 1644511149
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_149
timestamp 1644511149
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1644511149
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1644511149
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_169
timestamp 1644511149
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_181
timestamp 1644511149
transform 1 0 17756 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_189
timestamp 1644511149
transform 1 0 18492 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_209
timestamp 1644511149
transform 1 0 20332 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_221
timestamp 1644511149
transform 1 0 21436 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_225
timestamp 1644511149
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_237
timestamp 1644511149
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_249
timestamp 1644511149
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_261
timestamp 1644511149
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1644511149
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1644511149
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_281
timestamp 1644511149
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_293
timestamp 1644511149
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_305
timestamp 1644511149
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_317
timestamp 1644511149
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1644511149
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1644511149
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_337
timestamp 1644511149
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_349
timestamp 1644511149
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_361
timestamp 1644511149
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_373
timestamp 1644511149
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1644511149
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1644511149
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_393
timestamp 1644511149
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_405
timestamp 1644511149
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_417
timestamp 1644511149
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_429
timestamp 1644511149
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1644511149
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1644511149
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_449
timestamp 1644511149
transform 1 0 42412 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_454
timestamp 1644511149
transform 1 0 42872 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_461
timestamp 1644511149
transform 1 0 43516 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_468
timestamp 1644511149
transform 1 0 44160 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_475
timestamp 1644511149
transform 1 0 44804 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_500
timestamp 1644511149
transform 1 0 47104 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_508
timestamp 1644511149
transform 1 0 47840 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_82_7
timestamp 1644511149
transform 1 0 1748 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_13
timestamp 1644511149
transform 1 0 2300 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_17
timestamp 1644511149
transform 1 0 2668 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_24
timestamp 1644511149
transform 1 0 3312 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_32
timestamp 1644511149
transform 1 0 4048 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_44
timestamp 1644511149
transform 1 0 5152 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_56
timestamp 1644511149
transform 1 0 6256 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_68
timestamp 1644511149
transform 1 0 7360 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_73
timestamp 1644511149
transform 1 0 7820 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_81
timestamp 1644511149
transform 1 0 8556 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_85
timestamp 1644511149
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_97
timestamp 1644511149
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_109
timestamp 1644511149
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_121
timestamp 1644511149
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1644511149
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1644511149
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_141
timestamp 1644511149
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_153
timestamp 1644511149
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_165
timestamp 1644511149
transform 1 0 16284 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_82_174
timestamp 1644511149
transform 1 0 17112 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_186
timestamp 1644511149
transform 1 0 18216 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_194
timestamp 1644511149
transform 1 0 18952 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_209
timestamp 1644511149
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_221
timestamp 1644511149
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_233
timestamp 1644511149
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1644511149
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1644511149
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_253
timestamp 1644511149
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_265
timestamp 1644511149
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_277
timestamp 1644511149
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_289
timestamp 1644511149
transform 1 0 27692 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_296
timestamp 1644511149
transform 1 0 28336 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_309
timestamp 1644511149
transform 1 0 29532 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_317
timestamp 1644511149
transform 1 0 30268 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_322
timestamp 1644511149
transform 1 0 30728 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_334
timestamp 1644511149
transform 1 0 31832 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_346
timestamp 1644511149
transform 1 0 32936 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_358
timestamp 1644511149
transform 1 0 34040 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_82_365
timestamp 1644511149
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_377
timestamp 1644511149
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_389
timestamp 1644511149
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_401
timestamp 1644511149
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1644511149
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1644511149
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_421
timestamp 1644511149
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_433
timestamp 1644511149
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_445
timestamp 1644511149
transform 1 0 42044 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_449
timestamp 1644511149
transform 1 0 42412 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_457
timestamp 1644511149
transform 1 0 43148 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_461
timestamp 1644511149
transform 1 0 43516 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1644511149
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1644511149
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_498
timestamp 1644511149
transform 1 0 46920 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_506
timestamp 1644511149
transform 1 0 47656 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_512
timestamp 1644511149
transform 1 0 48208 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_83_3
timestamp 1644511149
transform 1 0 1380 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_83_30
timestamp 1644511149
transform 1 0 3864 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_36
timestamp 1644511149
transform 1 0 4416 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_40
timestamp 1644511149
transform 1 0 4784 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_44
timestamp 1644511149
transform 1 0 5152 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_48
timestamp 1644511149
transform 1 0 5520 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_57
timestamp 1644511149
transform 1 0 6348 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_61
timestamp 1644511149
transform 1 0 6716 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_83_86
timestamp 1644511149
transform 1 0 9016 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_98
timestamp 1644511149
transform 1 0 10120 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_83_110
timestamp 1644511149
transform 1 0 11224 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_83_116
timestamp 1644511149
transform 1 0 11776 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_83_123
timestamp 1644511149
transform 1 0 12420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_135
timestamp 1644511149
transform 1 0 13524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_141
timestamp 1644511149
transform 1 0 14076 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_145
timestamp 1644511149
transform 1 0 14444 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_157
timestamp 1644511149
transform 1 0 15548 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_164
timestamp 1644511149
transform 1 0 16192 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_169
timestamp 1644511149
transform 1 0 16652 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_191
timestamp 1644511149
transform 1 0 18676 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_83_198
timestamp 1644511149
transform 1 0 19320 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_83_209
timestamp 1644511149
transform 1 0 20332 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_83_221
timestamp 1644511149
transform 1 0 21436 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_83_228
timestamp 1644511149
transform 1 0 22080 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_83_235
timestamp 1644511149
transform 1 0 22724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_83_247
timestamp 1644511149
transform 1 0 23828 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_251
timestamp 1644511149
transform 1 0 24196 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_263
timestamp 1644511149
transform 1 0 25300 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_275
timestamp 1644511149
transform 1 0 26404 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_279
timestamp 1644511149
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_284
timestamp 1644511149
transform 1 0 27232 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_288
timestamp 1644511149
transform 1 0 27600 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_310
timestamp 1644511149
transform 1 0 29624 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_83_317
timestamp 1644511149
transform 1 0 30268 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_325
timestamp 1644511149
transform 1 0 31004 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 1644511149
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1644511149
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_340
timestamp 1644511149
transform 1 0 32384 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_348
timestamp 1644511149
transform 1 0 33120 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_83_371
timestamp 1644511149
transform 1 0 35236 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_83_380
timestamp 1644511149
transform 1 0 36064 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_393
timestamp 1644511149
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_405
timestamp 1644511149
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_417
timestamp 1644511149
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_429
timestamp 1644511149
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_444
timestamp 1644511149
transform 1 0 41952 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_83_449
timestamp 1644511149
transform 1 0 42412 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_83_454
timestamp 1644511149
transform 1 0 42872 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_479
timestamp 1644511149
transform 1 0 45172 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_486
timestamp 1644511149
transform 1 0 45816 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_493
timestamp 1644511149
transform 1 0 46460 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_500
timestamp 1644511149
transform 1 0 47104 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_505
timestamp 1644511149
transform 1 0 47564 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_512
timestamp 1644511149
transform 1 0 48208 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_24
timestamp 1644511149
transform 1 0 3312 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_32
timestamp 1644511149
transform 1 0 4048 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_57
timestamp 1644511149
transform 1 0 6348 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_64
timestamp 1644511149
transform 1 0 6992 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_84_71
timestamp 1644511149
transform 1 0 7636 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1644511149
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_85
timestamp 1644511149
transform 1 0 8924 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_84_92
timestamp 1644511149
transform 1 0 9568 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_100
timestamp 1644511149
transform 1 0 10304 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_84_123
timestamp 1644511149
transform 1 0 12420 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_84_131
timestamp 1644511149
transform 1 0 13156 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1644511149
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_141
timestamp 1644511149
transform 1 0 14076 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_84_148
timestamp 1644511149
transform 1 0 14720 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_160
timestamp 1644511149
transform 1 0 15824 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_164
timestamp 1644511149
transform 1 0 16192 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1644511149
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1644511149
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_200
timestamp 1644511149
transform 1 0 19504 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_84_229
timestamp 1644511149
transform 1 0 22172 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_236
timestamp 1644511149
transform 1 0 22816 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_84_243
timestamp 1644511149
transform 1 0 23460 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1644511149
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_256
timestamp 1644511149
transform 1 0 24656 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_263
timestamp 1644511149
transform 1 0 25300 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_270
timestamp 1644511149
transform 1 0 25944 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_295
timestamp 1644511149
transform 1 0 28244 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_84_302
timestamp 1644511149
transform 1 0 28888 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_84_309
timestamp 1644511149
transform 1 0 29532 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_84_314
timestamp 1644511149
transform 1 0 29992 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_321
timestamp 1644511149
transform 1 0 30636 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_346
timestamp 1644511149
transform 1 0 32936 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_84_353
timestamp 1644511149
transform 1 0 33580 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_84_361
timestamp 1644511149
transform 1 0 34316 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_84_365
timestamp 1644511149
transform 1 0 34684 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_84_370
timestamp 1644511149
transform 1 0 35144 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_84_395
timestamp 1644511149
transform 1 0 37444 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_407
timestamp 1644511149
transform 1 0 38548 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1644511149
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_424
timestamp 1644511149
transform 1 0 40112 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_432
timestamp 1644511149
transform 1 0 40848 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_84_437
timestamp 1644511149
transform 1 0 41308 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_447
timestamp 1644511149
transform 1 0 42228 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_472
timestamp 1644511149
transform 1 0 44528 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_84_481
timestamp 1644511149
transform 1 0 45356 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_489
timestamp 1644511149
transform 1 0 46092 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_84_512
timestamp 1644511149
transform 1 0 48208 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_6
timestamp 1644511149
transform 1 0 1656 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_31
timestamp 1644511149
transform 1 0 3956 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_39
timestamp 1644511149
transform 1 0 4692 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_85_46
timestamp 1644511149
transform 1 0 5336 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_85_54
timestamp 1644511149
transform 1 0 6072 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_85_78
timestamp 1644511149
transform 1 0 8280 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_84
timestamp 1644511149
transform 1 0 8832 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_85_106
timestamp 1644511149
transform 1 0 10856 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_85_134
timestamp 1644511149
transform 1 0 13432 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_85_163
timestamp 1644511149
transform 1 0 16100 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1644511149
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_85_169
timestamp 1644511149
transform 1 0 16652 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_85_193
timestamp 1644511149
transform 1 0 18860 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_85_218
timestamp 1644511149
transform 1 0 21160 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_225
timestamp 1644511149
transform 1 0 21804 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_230
timestamp 1644511149
transform 1 0 22264 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_85_255
timestamp 1644511149
transform 1 0 24564 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_261
timestamp 1644511149
transform 1 0 25116 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_265
timestamp 1644511149
transform 1 0 25484 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_85_273
timestamp 1644511149
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1644511149
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_281
timestamp 1644511149
transform 1 0 26956 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_306
timestamp 1644511149
transform 1 0 29256 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_331
timestamp 1644511149
transform 1 0 31556 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1644511149
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_85_358
timestamp 1644511149
transform 1 0 34040 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_85_366
timestamp 1644511149
transform 1 0 34776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_388
timestamp 1644511149
transform 1 0 36800 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_393
timestamp 1644511149
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_405
timestamp 1644511149
transform 1 0 38364 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_85_414
timestamp 1644511149
transform 1 0 39192 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_85_439
timestamp 1644511149
transform 1 0 41492 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1644511149
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_85_470
timestamp 1644511149
transform 1 0 44344 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_85_478
timestamp 1644511149
transform 1 0 45080 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_500
timestamp 1644511149
transform 1 0 47104 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_505
timestamp 1644511149
transform 1 0 47564 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_512
timestamp 1644511149
transform 1 0 48208 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_3
timestamp 1644511149
transform 1 0 1380 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_13
timestamp 1644511149
transform 1 0 2300 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_21
timestamp 1644511149
transform 1 0 3036 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1644511149
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_29
timestamp 1644511149
transform 1 0 3772 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_39
timestamp 1644511149
transform 1 0 4692 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_86_47
timestamp 1644511149
transform 1 0 5428 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_55
timestamp 1644511149
transform 1 0 6164 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_57
timestamp 1644511149
transform 1 0 6348 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_65
timestamp 1644511149
transform 1 0 7084 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_86_72
timestamp 1644511149
transform 1 0 7728 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_88
timestamp 1644511149
transform 1 0 9200 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_96
timestamp 1644511149
transform 1 0 9936 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_86_101
timestamp 1644511149
transform 1 0 10396 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_108
timestamp 1644511149
transform 1 0 11040 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_113
timestamp 1644511149
transform 1 0 11500 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_86_121
timestamp 1644511149
transform 1 0 12236 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_86_129
timestamp 1644511149
transform 1 0 12972 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_86_136
timestamp 1644511149
transform 1 0 13616 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_141
timestamp 1644511149
transform 1 0 14076 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_86_153
timestamp 1644511149
transform 1 0 15180 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_86_164
timestamp 1644511149
transform 1 0 16192 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_169
timestamp 1644511149
transform 1 0 16652 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_177
timestamp 1644511149
transform 1 0 17388 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_181
timestamp 1644511149
transform 1 0 17756 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_192
timestamp 1644511149
transform 1 0 18768 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_197
timestamp 1644511149
transform 1 0 19228 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_202
timestamp 1644511149
transform 1 0 19688 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_210
timestamp 1644511149
transform 1 0 20424 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_217
timestamp 1644511149
transform 1 0 21068 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_223
timestamp 1644511149
transform 1 0 21620 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_86_225
timestamp 1644511149
transform 1 0 21804 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_86_248
timestamp 1644511149
transform 1 0 23920 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_274
timestamp 1644511149
transform 1 0 26312 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_86_281
timestamp 1644511149
transform 1 0 26956 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_289
timestamp 1644511149
transform 1 0 27692 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_296
timestamp 1644511149
transform 1 0 28336 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_304
timestamp 1644511149
transform 1 0 29072 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_309
timestamp 1644511149
transform 1 0 29532 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_86_332
timestamp 1644511149
transform 1 0 31648 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_86_340
timestamp 1644511149
transform 1 0 32384 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_86_348
timestamp 1644511149
transform 1 0 33120 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_86_354
timestamp 1644511149
transform 1 0 33672 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_362
timestamp 1644511149
transform 1 0 34408 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_86_365
timestamp 1644511149
transform 1 0 34684 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_373
timestamp 1644511149
transform 1 0 35420 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_86_378
timestamp 1644511149
transform 1 0 35880 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_385
timestamp 1644511149
transform 1 0 36524 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_391
timestamp 1644511149
transform 1 0 37076 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_393
timestamp 1644511149
transform 1 0 37260 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_401
timestamp 1644511149
transform 1 0 37996 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_406
timestamp 1644511149
transform 1 0 38456 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_86_418
timestamp 1644511149
transform 1 0 39560 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_86_421
timestamp 1644511149
transform 1 0 39836 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_429
timestamp 1644511149
transform 1 0 40572 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_440
timestamp 1644511149
transform 1 0 41584 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_449
timestamp 1644511149
transform 1 0 42412 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_86_472
timestamp 1644511149
transform 1 0 44528 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_477
timestamp 1644511149
transform 1 0 44988 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_86_500
timestamp 1644511149
transform 1 0 47104 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_505
timestamp 1644511149
transform 1 0 47564 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_512
timestamp 1644511149
transform 1 0 48208 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 48852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 48852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 48852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 48852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 48852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 48852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 48852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 48852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 48852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 48852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 48852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 48852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 48852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 48852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 48852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 48852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 48852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 48852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 48852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 48852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 48852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 48852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 48852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 48852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 48852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 48852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 48852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 48852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 48852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 48852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 48852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 48852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 48852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 48852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 48852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 48852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 48852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 48852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 48852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 48852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 48852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 48852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 48852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 48852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 48852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 48852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 48852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 48852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 48852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 48852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 48852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 48852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 48852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 48852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 48852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 48852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 48852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 48852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 48852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 48852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 48852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 48852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 48852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 48852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 48852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 48852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 48852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 48852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 48852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 48852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 48852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 48852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 48852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 48852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 48852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 48852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1644511149
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1644511149
transform -1 0 48852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1644511149
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1644511149
transform -1 0 48852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1644511149
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1644511149
transform -1 0 48852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1644511149
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1644511149
transform -1 0 48852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1644511149
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1644511149
transform -1 0 48852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1644511149
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1644511149
transform -1 0 48852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1644511149
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1644511149
transform -1 0 48852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1644511149
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1644511149
transform -1 0 48852 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1644511149
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1644511149
transform -1 0 48852 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1644511149
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1644511149
transform -1 0 48852 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1644511149
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1644511149
transform -1 0 48852 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1644511149
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1644511149
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1644511149
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1644511149
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1644511149
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1644511149
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1644511149
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1644511149
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1644511149
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1644511149
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1644511149
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1644511149
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1644511149
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1644511149
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1644511149
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1644511149
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1644511149
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1644511149
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1644511149
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1644511149
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1644511149
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1644511149
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1644511149
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1644511149
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1644511149
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1644511149
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1644511149
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1644511149
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1644511149
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1644511149
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1644511149
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1644511149
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1644511149
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1644511149
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1644511149
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1644511149
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1644511149
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1644511149
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1644511149
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1644511149
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1644511149
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1644511149
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1644511149
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1644511149
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1644511149
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1644511149
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1644511149
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1644511149
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1644511149
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1644511149
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1644511149
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1644511149
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1644511149
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1644511149
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1644511149
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1644511149
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1644511149
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1644511149
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1644511149
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1644511149
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1644511149
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1644511149
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1644511149
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1644511149
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1644511149
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1644511149
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1644511149
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1644511149
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1644511149
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1644511149
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1644511149
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1644511149
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1644511149
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1644511149
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1644511149
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1644511149
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1644511149
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1644511149
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1644511149
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1644511149
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1644511149
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1644511149
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1644511149
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1644511149
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1644511149
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1644511149
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1644511149
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1644511149
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1644511149
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1644511149
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1644511149
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1644511149
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1644511149
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1644511149
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1644511149
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1644511149
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1644511149
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1644511149
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1644511149
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1644511149
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1644511149
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1644511149
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1644511149
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1644511149
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1644511149
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1644511149
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1644511149
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1644511149
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1644511149
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1644511149
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1644511149
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1644511149
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1644511149
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1644511149
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1644511149
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1644511149
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1644511149
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1644511149
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1644511149
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1644511149
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1644511149
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1644511149
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1644511149
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1644511149
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1644511149
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1644511149
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1644511149
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1644511149
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1644511149
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1644511149
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1644511149
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1644511149
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1644511149
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1644511149
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1644511149
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1644511149
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1644511149
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1644511149
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1644511149
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1644511149
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1644511149
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1644511149
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1644511149
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1644511149
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1644511149
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1644511149
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1644511149
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1644511149
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1644511149
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1644511149
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1644511149
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1644511149
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1644511149
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1644511149
transform 1 0 6256 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1644511149
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1644511149
transform 1 0 11408 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1644511149
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1644511149
transform 1 0 16560 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1644511149
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1644511149
transform 1 0 21712 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1644511149
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1644511149
transform 1 0 26864 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1644511149
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1644511149
transform 1 0 32016 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1644511149
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1644511149
transform 1 0 37168 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1644511149
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1644511149
transform 1 0 42320 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1644511149
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1644511149
transform 1 0 47472 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0851_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 46828 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0852_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0853_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17756 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  _0854_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9568 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0855_
timestamp 1644511149
transform 1 0 44988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0856_
timestamp 1644511149
transform 1 0 6716 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0857_
timestamp 1644511149
transform 1 0 46828 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0858_
timestamp 1644511149
transform 1 0 7544 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0859_
timestamp 1644511149
transform 1 0 46828 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0860_
timestamp 1644511149
transform 1 0 18216 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  _0861_
timestamp 1644511149
transform 1 0 18492 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0862_
timestamp 1644511149
transform 1 0 46828 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0863_
timestamp 1644511149
transform 1 0 2116 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0864_
timestamp 1644511149
transform 1 0 2484 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0865_
timestamp 1644511149
transform 1 0 36156 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0866_
timestamp 1644511149
transform 1 0 47196 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0867_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18492 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0868_
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0869_
timestamp 1644511149
transform 1 0 45540 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0870_
timestamp 1644511149
transform 1 0 2116 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0871_
timestamp 1644511149
transform 1 0 46184 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0872_
timestamp 1644511149
transform 1 0 24380 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _0873_
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0874_
timestamp 1644511149
transform 1 0 2208 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0875_
timestamp 1644511149
transform 1 0 47564 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0876_
timestamp 1644511149
transform 1 0 3772 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0877_
timestamp 1644511149
transform 1 0 11868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0878_
timestamp 1644511149
transform 1 0 46828 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0879_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18492 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0880_
timestamp 1644511149
transform 1 0 2024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0881_
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0882_
timestamp 1644511149
transform 1 0 21804 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0883_
timestamp 1644511149
transform 1 0 2024 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0884_
timestamp 1644511149
transform 1 0 2024 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0885_
timestamp 1644511149
transform 1 0 20332 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0886_
timestamp 1644511149
transform 1 0 37996 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0887_
timestamp 1644511149
transform 1 0 2852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0888_
timestamp 1644511149
transform 1 0 8924 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0889_
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0890_
timestamp 1644511149
transform 1 0 37260 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0891_
timestamp 1644511149
transform 1 0 18676 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0892_
timestamp 1644511149
transform 1 0 19596 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0893_
timestamp 1644511149
transform 1 0 18400 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0894_
timestamp 1644511149
transform 1 0 18768 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0895_
timestamp 1644511149
transform 1 0 29900 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0896_
timestamp 1644511149
transform 1 0 31464 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0897_
timestamp 1644511149
transform 1 0 30544 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0898_
timestamp 1644511149
transform 1 0 19596 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0899_
timestamp 1644511149
transform 1 0 33672 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0900_
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0901_
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0902_
timestamp 1644511149
transform 1 0 30728 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0903_
timestamp 1644511149
transform 1 0 34316 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _0904_
timestamp 1644511149
transform 1 0 18952 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0905_
timestamp 1644511149
transform 1 0 40848 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0906_
timestamp 1644511149
transform 1 0 47564 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0907_
timestamp 1644511149
transform 1 0 2392 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0908_
timestamp 1644511149
transform 1 0 41032 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0909_
timestamp 1644511149
transform 1 0 2668 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0910_
timestamp 1644511149
transform 1 0 18308 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0911_
timestamp 1644511149
transform 1 0 2760 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0912_
timestamp 1644511149
transform 1 0 17664 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0913_
timestamp 1644511149
transform 1 0 20056 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0914_
timestamp 1644511149
transform 1 0 14996 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0915_
timestamp 1644511149
transform 1 0 28704 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0916_
timestamp 1644511149
transform 1 0 17664 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0917_
timestamp 1644511149
transform 1 0 2760 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0918_
timestamp 1644511149
transform 1 0 46828 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0919_
timestamp 1644511149
transform 1 0 46276 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0920_
timestamp 1644511149
transform 1 0 7636 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0921_
timestamp 1644511149
transform 1 0 12604 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0922_
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _0923_
timestamp 1644511149
transform 1 0 17940 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0924_
timestamp 1644511149
transform 1 0 46828 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0925_
timestamp 1644511149
transform 1 0 45080 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0926_
timestamp 1644511149
transform 1 0 39836 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0927_
timestamp 1644511149
transform 1 0 11500 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0928_
timestamp 1644511149
transform 1 0 46828 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0929_
timestamp 1644511149
transform 1 0 20700 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0930_
timestamp 1644511149
transform 1 0 27048 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0931_
timestamp 1644511149
transform 1 0 23000 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0932_
timestamp 1644511149
transform 1 0 35972 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0933_
timestamp 1644511149
transform 1 0 35972 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0934_
timestamp 1644511149
transform 1 0 35788 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0935_
timestamp 1644511149
transform 1 0 19228 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0936_
timestamp 1644511149
transform 1 0 20240 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0937_
timestamp 1644511149
transform 1 0 2944 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0938_
timestamp 1644511149
transform 1 0 29716 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0939_
timestamp 1644511149
transform 1 0 34868 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0940_
timestamp 1644511149
transform 1 0 12144 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0941_
timestamp 1644511149
transform 1 0 19136 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0942_
timestamp 1644511149
transform 1 0 25300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0943_
timestamp 1644511149
transform 1 0 23552 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0944_
timestamp 1644511149
transform 1 0 19228 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0945_
timestamp 1644511149
transform 1 0 47564 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0946_
timestamp 1644511149
transform 1 0 28612 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0947_
timestamp 1644511149
transform 1 0 21896 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0948_
timestamp 1644511149
transform 1 0 4876 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0949_
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0950_
timestamp 1644511149
transform 1 0 9936 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0951_
timestamp 1644511149
transform 1 0 30360 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0952_
timestamp 1644511149
transform 1 0 29716 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0953_
timestamp 1644511149
transform 1 0 17388 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  _0954_
timestamp 1644511149
transform 1 0 17020 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0955_
timestamp 1644511149
transform 1 0 2668 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0956_
timestamp 1644511149
transform 1 0 22540 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0957_
timestamp 1644511149
transform 1 0 2024 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0958_
timestamp 1644511149
transform 1 0 47564 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0959_
timestamp 1644511149
transform 1 0 1380 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0960_
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0961_
timestamp 1644511149
transform 1 0 46736 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0962_
timestamp 1644511149
transform 1 0 45816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0963_
timestamp 1644511149
transform 1 0 3772 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0964_
timestamp 1644511149
transform 1 0 11408 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0965_
timestamp 1644511149
transform 1 0 45816 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0966_
timestamp 1644511149
transform 1 0 17112 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0967_
timestamp 1644511149
transform 1 0 18308 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0968_
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0969_
timestamp 1644511149
transform 1 0 18492 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0970_
timestamp 1644511149
transform 1 0 15640 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1644511149
transform 1 0 2852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0972_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15640 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0973_
timestamp 1644511149
transform 1 0 6624 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0974_
timestamp 1644511149
transform 1 0 6624 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0975_
timestamp 1644511149
transform 1 0 6900 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0976_
timestamp 1644511149
transform 1 0 15916 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0977_
timestamp 1644511149
transform 1 0 5612 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0978_
timestamp 1644511149
transform 1 0 17020 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0979_
timestamp 1644511149
transform 1 0 30728 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0980_
timestamp 1644511149
transform 1 0 2668 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0981_
timestamp 1644511149
transform 1 0 3036 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0982_
timestamp 1644511149
transform 1 0 6440 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0983_
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0984_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31188 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  _0985_
timestamp 1644511149
transform 1 0 31096 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0986_
timestamp 1644511149
transform 1 0 2668 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0987_
timestamp 1644511149
transform 1 0 10764 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0988_
timestamp 1644511149
transform 1 0 9292 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0989_
timestamp 1644511149
transform 1 0 15916 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0990_
timestamp 1644511149
transform 1 0 32108 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0991_
timestamp 1644511149
transform 1 0 32568 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0992_
timestamp 1644511149
transform 1 0 14628 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0993_
timestamp 1644511149
transform 1 0 36524 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0994_
timestamp 1644511149
transform 1 0 38088 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0995_
timestamp 1644511149
transform 1 0 37352 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0996_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 38732 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _0997_
timestamp 1644511149
transform 1 0 29900 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0998_
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0999_
timestamp 1644511149
transform 1 0 33120 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1000_
timestamp 1644511149
transform 1 0 13248 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1001_
timestamp 1644511149
transform 1 0 32568 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1002_
timestamp 1644511149
transform 1 0 15088 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1003_
timestamp 1644511149
transform 1 0 30820 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1004_
timestamp 1644511149
transform 1 0 29808 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1005_
timestamp 1644511149
transform 1 0 12972 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1006_
timestamp 1644511149
transform 1 0 16836 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1007_
timestamp 1644511149
transform 1 0 33304 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1008_
timestamp 1644511149
transform 1 0 14444 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1009_
timestamp 1644511149
transform 1 0 30636 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1010_
timestamp 1644511149
transform 1 0 2668 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1011_
timestamp 1644511149
transform 1 0 2024 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1012_
timestamp 1644511149
transform 1 0 2024 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1013_
timestamp 1644511149
transform 1 0 46644 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1014_
timestamp 1644511149
transform 1 0 43792 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1015_
timestamp 1644511149
transform 1 0 18400 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  _1016_
timestamp 1644511149
transform 1 0 18860 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1017_
timestamp 1644511149
transform 1 0 2944 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1018_
timestamp 1644511149
transform 1 0 28060 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1019_
timestamp 1644511149
transform 1 0 47564 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1020_
timestamp 1644511149
transform 1 0 41676 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1021_
timestamp 1644511149
transform 1 0 47104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1022_
timestamp 1644511149
transform 1 0 17940 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1023_
timestamp 1644511149
transform 1 0 5244 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1024_
timestamp 1644511149
transform 1 0 13248 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1025_
timestamp 1644511149
transform 1 0 26956 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1026_
timestamp 1644511149
transform 1 0 42596 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1027_
timestamp 1644511149
transform 1 0 41676 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1028_
timestamp 1644511149
transform 1 0 18860 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1029_
timestamp 1644511149
transform 1 0 2392 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1030_
timestamp 1644511149
transform 1 0 46828 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1031_
timestamp 1644511149
transform 1 0 2024 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1032_
timestamp 1644511149
transform 1 0 47104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1033_
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1034_
timestamp 1644511149
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1035_
timestamp 1644511149
transform 1 0 47564 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1036_
timestamp 1644511149
transform 1 0 44528 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1037_
timestamp 1644511149
transform 1 0 7452 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1038_
timestamp 1644511149
transform 1 0 35788 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1039_
timestamp 1644511149
transform 1 0 47564 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1040_
timestamp 1644511149
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1041_
timestamp 1644511149
transform 1 0 2116 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1042_
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1043_
timestamp 1644511149
transform 1 0 2208 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1044_
timestamp 1644511149
transform 1 0 19044 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1045_
timestamp 1644511149
transform 1 0 29992 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1046_
timestamp 1644511149
transform 1 0 13892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1047_
timestamp 1644511149
transform 1 0 8740 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1048_
timestamp 1644511149
transform 1 0 11592 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1049_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26128 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1050_
timestamp 1644511149
transform 1 0 25208 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1051_
timestamp 1644511149
transform 1 0 24840 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1052_
timestamp 1644511149
transform 1 0 20884 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1053_
timestamp 1644511149
transform 1 0 17112 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1054_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24748 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1055_
timestamp 1644511149
transform 1 0 23276 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1056_
timestamp 1644511149
transform 1 0 21988 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1057_
timestamp 1644511149
transform 1 0 25392 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1058_
timestamp 1644511149
transform 1 0 23276 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1059_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23092 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1060_
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1061_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25944 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1062_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21988 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1063_
timestamp 1644511149
transform 1 0 23092 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1064_
timestamp 1644511149
transform 1 0 28612 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1065_
timestamp 1644511149
transform 1 0 21896 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1066_
timestamp 1644511149
transform 1 0 23184 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1067_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1068_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23644 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1069_
timestamp 1644511149
transform 1 0 15272 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__or3b_2  _1070_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17296 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1071_
timestamp 1644511149
transform 1 0 12696 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1072_
timestamp 1644511149
transform 1 0 13156 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__and2_2  _1073_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22264 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1074_
timestamp 1644511149
transform 1 0 23184 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1075_
timestamp 1644511149
transform 1 0 22908 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1076_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15824 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1077_
timestamp 1644511149
transform 1 0 15640 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1078_
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1079_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1080_
timestamp 1644511149
transform 1 0 15180 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1081_
timestamp 1644511149
transform 1 0 14168 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1082_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17112 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1083_
timestamp 1644511149
transform 1 0 17296 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1084_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20240 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1085_
timestamp 1644511149
transform 1 0 20148 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1086_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17480 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1087_
timestamp 1644511149
transform 1 0 23920 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1088_
timestamp 1644511149
transform 1 0 22908 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1089_
timestamp 1644511149
transform 1 0 17572 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1090_
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1091_
timestamp 1644511149
transform 1 0 11040 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1092_
timestamp 1644511149
transform 1 0 14076 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1093_
timestamp 1644511149
transform 1 0 13984 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1094_
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1095_
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1096_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14444 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1097_
timestamp 1644511149
transform 1 0 18584 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1098_
timestamp 1644511149
transform 1 0 24104 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_2  _1099_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 47288 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__or4_2  _1100_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25024 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1101_
timestamp 1644511149
transform 1 0 24472 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1102_
timestamp 1644511149
transform 1 0 25024 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1103_
timestamp 1644511149
transform 1 0 37996 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _1104_
timestamp 1644511149
transform 1 0 6164 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1105_
timestamp 1644511149
transform 1 0 23828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1106_
timestamp 1644511149
transform 1 0 22908 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1107_
timestamp 1644511149
transform 1 0 24748 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1108_
timestamp 1644511149
transform 1 0 25116 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1109_
timestamp 1644511149
transform 1 0 24380 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1110_
timestamp 1644511149
transform 1 0 24656 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1111_
timestamp 1644511149
transform 1 0 19596 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1112_
timestamp 1644511149
transform 1 0 25484 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1113_
timestamp 1644511149
transform 1 0 23736 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_4  _1114_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1115_
timestamp 1644511149
transform 1 0 18768 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1116_
timestamp 1644511149
transform 1 0 17940 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1117_
timestamp 1644511149
transform 1 0 23644 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1118_
timestamp 1644511149
transform 1 0 25024 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1119_
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1120_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18768 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1121_
timestamp 1644511149
transform 1 0 21068 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1122_
timestamp 1644511149
transform 1 0 20332 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1123_
timestamp 1644511149
transform 1 0 20148 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1124_
timestamp 1644511149
transform 1 0 20056 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1125_
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1126_
timestamp 1644511149
transform 1 0 19136 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1127_
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1128_
timestamp 1644511149
transform 1 0 19412 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1129_
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1130_
timestamp 1644511149
transform 1 0 30452 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1131_
timestamp 1644511149
transform 1 0 29624 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1132_
timestamp 1644511149
transform 1 0 30084 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1133_
timestamp 1644511149
transform 1 0 29992 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1134_
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1135_
timestamp 1644511149
transform 1 0 30728 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1136_
timestamp 1644511149
transform 1 0 31096 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1137_
timestamp 1644511149
transform 1 0 31372 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1138_
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1139_
timestamp 1644511149
transform 1 0 30912 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1140_
timestamp 1644511149
transform 1 0 31556 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1141_
timestamp 1644511149
transform 1 0 30912 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1142_
timestamp 1644511149
transform 1 0 30452 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1143_
timestamp 1644511149
transform 1 0 30636 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1144_
timestamp 1644511149
transform 1 0 32568 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1145_
timestamp 1644511149
transform 1 0 30268 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1146_
timestamp 1644511149
transform 1 0 31464 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1147_
timestamp 1644511149
transform 1 0 31188 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1148_
timestamp 1644511149
transform 1 0 31556 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1149_
timestamp 1644511149
transform 1 0 31832 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1150_
timestamp 1644511149
transform 1 0 30912 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1151_
timestamp 1644511149
transform 1 0 33396 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1152_
timestamp 1644511149
transform 1 0 30360 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1153_
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1154_
timestamp 1644511149
transform 1 0 32660 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1155_
timestamp 1644511149
transform 1 0 12696 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1156_
timestamp 1644511149
transform 1 0 12696 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1157_
timestamp 1644511149
transform 1 0 15732 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1158_
timestamp 1644511149
transform 1 0 13984 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1159_
timestamp 1644511149
transform 1 0 14628 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1160_
timestamp 1644511149
transform 1 0 13064 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1161_
timestamp 1644511149
transform 1 0 13064 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1162_
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1163_
timestamp 1644511149
transform 1 0 13800 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1164_
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1165_
timestamp 1644511149
transform 1 0 14628 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1166_
timestamp 1644511149
transform 1 0 14444 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1167_
timestamp 1644511149
transform 1 0 15272 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1168_
timestamp 1644511149
transform 1 0 10580 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1169_
timestamp 1644511149
transform 1 0 11592 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1170_
timestamp 1644511149
transform 1 0 10304 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1171_
timestamp 1644511149
transform 1 0 10028 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1172_
timestamp 1644511149
transform 1 0 8004 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1173_
timestamp 1644511149
transform 1 0 10120 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1174_
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1175_
timestamp 1644511149
transform 1 0 10764 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1176_
timestamp 1644511149
transform 1 0 9200 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1177_
timestamp 1644511149
transform 1 0 8004 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1178_
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1179_
timestamp 1644511149
transform 1 0 9016 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1180_
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1181_
timestamp 1644511149
transform 1 0 10488 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1182_
timestamp 1644511149
transform 1 0 9568 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1183_
timestamp 1644511149
transform 1 0 23368 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1184_
timestamp 1644511149
transform 1 0 23368 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1185_
timestamp 1644511149
transform 1 0 16744 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1186_
timestamp 1644511149
transform 1 0 22632 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1187_
timestamp 1644511149
transform 1 0 15916 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1188_
timestamp 1644511149
transform 1 0 24288 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1189_
timestamp 1644511149
transform 1 0 16376 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1190_
timestamp 1644511149
transform 1 0 13892 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and4_2  _1191_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1192_
timestamp 1644511149
transform 1 0 17848 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1193_
timestamp 1644511149
transform 1 0 12696 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1194_
timestamp 1644511149
transform 1 0 11592 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1195_
timestamp 1644511149
transform 1 0 13340 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1196_
timestamp 1644511149
transform 1 0 14168 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1197_
timestamp 1644511149
transform 1 0 15548 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1198_
timestamp 1644511149
transform 1 0 15456 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1199_
timestamp 1644511149
transform 1 0 12696 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1200_
timestamp 1644511149
transform 1 0 11592 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1201_
timestamp 1644511149
transform 1 0 17848 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1202_
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1203_
timestamp 1644511149
transform 1 0 19320 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1204_
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1205_
timestamp 1644511149
transform 1 0 18032 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1206_
timestamp 1644511149
transform 1 0 20056 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1207_
timestamp 1644511149
transform 1 0 18032 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1208_
timestamp 1644511149
transform 1 0 18768 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1209_
timestamp 1644511149
transform 1 0 17204 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1210_
timestamp 1644511149
transform 1 0 17572 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1211_
timestamp 1644511149
transform 1 0 19320 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1212_
timestamp 1644511149
transform 1 0 20056 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1213_
timestamp 1644511149
transform 1 0 19872 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1214_
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1215_
timestamp 1644511149
transform 1 0 24288 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1216_
timestamp 1644511149
transform 1 0 23000 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1217_
timestamp 1644511149
transform 1 0 23368 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1218_
timestamp 1644511149
transform 1 0 22816 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1219_
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1220_
timestamp 1644511149
transform 1 0 26404 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1221_
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1222_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1223_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17204 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1224_
timestamp 1644511149
transform 1 0 21988 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1225_
timestamp 1644511149
transform 1 0 22632 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1226_
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1227_
timestamp 1644511149
transform 1 0 24472 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1228_
timestamp 1644511149
transform 1 0 27048 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1229_
timestamp 1644511149
transform 1 0 27232 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1230_
timestamp 1644511149
transform 1 0 25300 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1231_
timestamp 1644511149
transform 1 0 25944 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1232_
timestamp 1644511149
transform 1 0 28612 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1233_
timestamp 1644511149
transform 1 0 25576 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1234_
timestamp 1644511149
transform 1 0 29164 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1235_
timestamp 1644511149
transform 1 0 28888 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1236_
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1237_
timestamp 1644511149
transform 1 0 28428 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1238_
timestamp 1644511149
transform 1 0 28336 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1239_
timestamp 1644511149
transform 1 0 27140 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1240_
timestamp 1644511149
transform 1 0 25668 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1241_
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1242_
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1243_
timestamp 1644511149
transform 1 0 17940 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1244_
timestamp 1644511149
transform 1 0 17112 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1245_
timestamp 1644511149
transform 1 0 17756 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1246_
timestamp 1644511149
transform 1 0 17756 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1247_
timestamp 1644511149
transform 1 0 16836 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1248_
timestamp 1644511149
transform 1 0 19044 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1249_
timestamp 1644511149
transform 1 0 17940 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1250_
timestamp 1644511149
transform 1 0 18584 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1251_
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _1252_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23368 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1253_
timestamp 1644511149
transform 1 0 9016 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1254_
timestamp 1644511149
transform 1 0 23828 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1255_
timestamp 1644511149
transform 1 0 24932 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1256_
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1257_
timestamp 1644511149
transform 1 0 25208 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1258_
timestamp 1644511149
transform 1 0 21436 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _1259_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23276 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1260_
timestamp 1644511149
transform 1 0 25116 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1261_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_1  _1262_
timestamp 1644511149
transform 1 0 23000 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1263_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21528 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1264_
timestamp 1644511149
transform 1 0 22172 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1265_
timestamp 1644511149
transform 1 0 22632 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1266_
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1267_
timestamp 1644511149
transform 1 0 22356 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1268_
timestamp 1644511149
transform 1 0 25944 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1269_
timestamp 1644511149
transform 1 0 25576 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1270_
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1271_
timestamp 1644511149
transform 1 0 22172 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1272_
timestamp 1644511149
transform 1 0 22080 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1273_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23368 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1274_
timestamp 1644511149
transform 1 0 20976 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1275_
timestamp 1644511149
transform 1 0 21068 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1276_
timestamp 1644511149
transform 1 0 20056 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1277_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20516 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1278_
timestamp 1644511149
transform 1 0 19780 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1279_
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1280_
timestamp 1644511149
transform 1 0 25116 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1281_
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__or4_2  _1282_
timestamp 1644511149
transform 1 0 21988 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1283_
timestamp 1644511149
transform 1 0 25116 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1284_
timestamp 1644511149
transform 1 0 21252 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1285_
timestamp 1644511149
transform 1 0 26036 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1286_
timestamp 1644511149
transform 1 0 23368 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1287_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20332 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1288_
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1289_
timestamp 1644511149
transform 1 0 24196 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1290_
timestamp 1644511149
transform 1 0 23552 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1291_
timestamp 1644511149
transform 1 0 23920 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1292_
timestamp 1644511149
transform 1 0 25484 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1293_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24748 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1294_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25116 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1295_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25668 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1296_
timestamp 1644511149
transform 1 0 26220 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1297_
timestamp 1644511149
transform 1 0 27324 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1298_
timestamp 1644511149
transform 1 0 28520 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1299_
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1300_
timestamp 1644511149
transform 1 0 28704 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1301_
timestamp 1644511149
transform 1 0 27140 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1302_
timestamp 1644511149
transform 1 0 27600 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or4_2  _1303_
timestamp 1644511149
transform 1 0 26312 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1304_
timestamp 1644511149
transform 1 0 28152 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1305_
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1306_
timestamp 1644511149
transform 1 0 27140 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1307_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27140 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1308_
timestamp 1644511149
transform 1 0 28244 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1309_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1310_
timestamp 1644511149
transform 1 0 26404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1311_
timestamp 1644511149
transform 1 0 27324 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1312_
timestamp 1644511149
transform 1 0 28244 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1313_
timestamp 1644511149
transform 1 0 28060 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1314_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27048 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1315_
timestamp 1644511149
transform 1 0 27876 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1316_
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1317_
timestamp 1644511149
transform 1 0 27048 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1318_
timestamp 1644511149
transform 1 0 26772 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1319_
timestamp 1644511149
transform 1 0 27416 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1320_
timestamp 1644511149
transform 1 0 27600 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1321_
timestamp 1644511149
transform 1 0 26956 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1322_
timestamp 1644511149
transform 1 0 27232 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1323_
timestamp 1644511149
transform 1 0 28060 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1324_
timestamp 1644511149
transform 1 0 27416 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1325_
timestamp 1644511149
transform 1 0 26036 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _1326_
timestamp 1644511149
transform 1 0 25944 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1327_
timestamp 1644511149
transform 1 0 24564 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1328_
timestamp 1644511149
transform 1 0 26588 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1329_
timestamp 1644511149
transform 1 0 26220 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1330_
timestamp 1644511149
transform 1 0 28612 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1331_
timestamp 1644511149
transform 1 0 27140 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1332_
timestamp 1644511149
transform 1 0 23644 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1333_
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1334_
timestamp 1644511149
transform 1 0 23092 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1335_
timestamp 1644511149
transform 1 0 24656 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1336_
timestamp 1644511149
transform 1 0 22264 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1337_
timestamp 1644511149
transform 1 0 22724 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1338_
timestamp 1644511149
transform 1 0 22172 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1339_
timestamp 1644511149
transform 1 0 20976 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1340_
timestamp 1644511149
transform 1 0 21712 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1341_
timestamp 1644511149
transform 1 0 21436 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1342_
timestamp 1644511149
transform 1 0 20792 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1343_
timestamp 1644511149
transform 1 0 21068 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1344_
timestamp 1644511149
transform 1 0 20884 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1345_
timestamp 1644511149
transform 1 0 20148 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1346_
timestamp 1644511149
transform 1 0 25852 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1347_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22264 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1348_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20240 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1349_
timestamp 1644511149
transform 1 0 20516 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1350_
timestamp 1644511149
transform 1 0 22080 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1351_
timestamp 1644511149
transform 1 0 21160 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _1352_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20240 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1353_
timestamp 1644511149
transform 1 0 21160 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1354_
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1355_
timestamp 1644511149
transform 1 0 20516 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1356_
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1357_
timestamp 1644511149
transform 1 0 15548 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1358_
timestamp 1644511149
transform 1 0 24196 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1359_
timestamp 1644511149
transform 1 0 24012 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1360_
timestamp 1644511149
transform 1 0 24564 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1361_
timestamp 1644511149
transform 1 0 25024 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1362_
timestamp 1644511149
transform 1 0 29440 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1363_
timestamp 1644511149
transform 1 0 24748 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1364_
timestamp 1644511149
transform 1 0 26220 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1365_
timestamp 1644511149
transform 1 0 29992 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1366_
timestamp 1644511149
transform 1 0 25944 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1367_
timestamp 1644511149
transform 1 0 26588 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_2  _1368_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25484 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1369_
timestamp 1644511149
transform 1 0 26128 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1370_
timestamp 1644511149
transform 1 0 23828 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1371_
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1372_
timestamp 1644511149
transform 1 0 22908 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _1373_
timestamp 1644511149
transform 1 0 12972 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1374_
timestamp 1644511149
transform 1 0 9752 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1375_
timestamp 1644511149
transform 1 0 9936 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1376_
timestamp 1644511149
transform 1 0 9016 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _1377_
timestamp 1644511149
transform 1 0 9476 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _1378_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9292 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1379_
timestamp 1644511149
transform 1 0 10212 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1380_
timestamp 1644511149
transform 1 0 10672 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1381_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8648 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1382_
timestamp 1644511149
transform 1 0 9568 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1383_
timestamp 1644511149
transform 1 0 9384 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1384_
timestamp 1644511149
transform 1 0 10580 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1385_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1386_
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1387_
timestamp 1644511149
transform 1 0 12328 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1388_
timestamp 1644511149
transform 1 0 12144 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1389_
timestamp 1644511149
transform 1 0 12052 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1390_
timestamp 1644511149
transform 1 0 9844 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1391_
timestamp 1644511149
transform 1 0 10580 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1392_
timestamp 1644511149
transform 1 0 13800 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1393_
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1394_
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _1395_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14168 0 1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1396_
timestamp 1644511149
transform 1 0 13524 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _1397_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14812 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1398_
timestamp 1644511149
transform 1 0 14812 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1399_
timestamp 1644511149
transform 1 0 14536 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1400_
timestamp 1644511149
transform 1 0 12144 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1401_
timestamp 1644511149
transform 1 0 12972 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1402_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12512 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_2  _1403_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17112 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _1404_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14168 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1405_
timestamp 1644511149
transform 1 0 13248 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1406_
timestamp 1644511149
transform 1 0 13616 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1407_
timestamp 1644511149
transform 1 0 13432 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1408_
timestamp 1644511149
transform 1 0 20884 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1409_
timestamp 1644511149
transform 1 0 19872 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1410_
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1411_
timestamp 1644511149
transform 1 0 11960 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1412_
timestamp 1644511149
transform 1 0 13248 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1413_
timestamp 1644511149
transform 1 0 13064 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1414_
timestamp 1644511149
transform 1 0 12696 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1415_
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1416_
timestamp 1644511149
transform 1 0 12696 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1417_
timestamp 1644511149
transform 1 0 12144 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1418_
timestamp 1644511149
transform 1 0 14904 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _1419_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14628 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1420_
timestamp 1644511149
transform 1 0 12328 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1421_
timestamp 1644511149
transform 1 0 14168 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1422_
timestamp 1644511149
transform 1 0 14904 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1423_
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1424_
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1425_
timestamp 1644511149
transform 1 0 12052 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1426_
timestamp 1644511149
transform 1 0 11960 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _1427_
timestamp 1644511149
transform 1 0 12328 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1428_
timestamp 1644511149
transform 1 0 10212 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1429_
timestamp 1644511149
transform 1 0 11500 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1430_
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1431_
timestamp 1644511149
transform 1 0 10304 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _1432_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11592 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1433_
timestamp 1644511149
transform 1 0 10488 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1434_
timestamp 1644511149
transform 1 0 9660 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1435_
timestamp 1644511149
transform 1 0 10120 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1436_
timestamp 1644511149
transform 1 0 10212 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1437_
timestamp 1644511149
transform 1 0 10856 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _1438_
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1439_
timestamp 1644511149
transform 1 0 9292 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1440_
timestamp 1644511149
transform 1 0 10304 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _1441_
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1442_
timestamp 1644511149
transform 1 0 20976 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1443_
timestamp 1644511149
transform 1 0 27416 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1444_
timestamp 1644511149
transform 1 0 20976 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1445_
timestamp 1644511149
transform 1 0 30360 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1446_
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1447_
timestamp 1644511149
transform 1 0 27416 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1448_
timestamp 1644511149
transform 1 0 28152 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1449_
timestamp 1644511149
transform 1 0 27416 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1450_
timestamp 1644511149
transform 1 0 25944 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1451_
timestamp 1644511149
transform 1 0 25576 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1452_
timestamp 1644511149
transform 1 0 26496 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1453_
timestamp 1644511149
transform 1 0 25668 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1454_
timestamp 1644511149
transform 1 0 25760 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1455_
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1456_
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1457_
timestamp 1644511149
transform 1 0 30820 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1458_
timestamp 1644511149
transform 1 0 30820 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1459_
timestamp 1644511149
transform 1 0 31004 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1460_
timestamp 1644511149
transform 1 0 31556 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1461_
timestamp 1644511149
transform 1 0 32660 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1462_
timestamp 1644511149
transform 1 0 33672 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1463_
timestamp 1644511149
transform 1 0 32016 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1464_
timestamp 1644511149
transform 1 0 28152 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1465_
timestamp 1644511149
transform 1 0 32936 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1466_
timestamp 1644511149
transform 1 0 30912 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1467_
timestamp 1644511149
transform 1 0 28888 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1468_
timestamp 1644511149
transform 1 0 31556 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1469_
timestamp 1644511149
transform 1 0 28060 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1470_
timestamp 1644511149
transform 1 0 28704 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1471_
timestamp 1644511149
transform 1 0 30176 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1472_
timestamp 1644511149
transform 1 0 30360 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1473_
timestamp 1644511149
transform 1 0 30636 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1474_
timestamp 1644511149
transform 1 0 30452 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1475_
timestamp 1644511149
transform 1 0 29624 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1476_
timestamp 1644511149
transform 1 0 30820 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1477_
timestamp 1644511149
transform 1 0 28980 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1478_
timestamp 1644511149
transform 1 0 28612 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1479_
timestamp 1644511149
transform 1 0 27876 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1480_
timestamp 1644511149
transform 1 0 29532 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1481_
timestamp 1644511149
transform 1 0 30728 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1482_
timestamp 1644511149
transform 1 0 31372 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1483_
timestamp 1644511149
transform 1 0 26864 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1484_
timestamp 1644511149
transform 1 0 29808 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1485_
timestamp 1644511149
transform 1 0 30360 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1486_
timestamp 1644511149
transform 1 0 27876 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1487_
timestamp 1644511149
transform 1 0 30360 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1488_
timestamp 1644511149
transform 1 0 26220 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1489_
timestamp 1644511149
transform 1 0 29900 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1490_
timestamp 1644511149
transform 1 0 27968 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1491_
timestamp 1644511149
transform 1 0 27140 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1492_
timestamp 1644511149
transform 1 0 27968 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1493_
timestamp 1644511149
transform 1 0 29716 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1494_
timestamp 1644511149
transform 1 0 30912 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1495_
timestamp 1644511149
transform 1 0 33028 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1496_
timestamp 1644511149
transform 1 0 29716 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1497_
timestamp 1644511149
transform 1 0 30452 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1498_
timestamp 1644511149
transform 1 0 31740 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1499_
timestamp 1644511149
transform 1 0 27876 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1500_
timestamp 1644511149
transform 1 0 27508 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1501_
timestamp 1644511149
transform 1 0 27784 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1502_
timestamp 1644511149
transform 1 0 27416 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1503_
timestamp 1644511149
transform 1 0 27416 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1504_
timestamp 1644511149
transform 1 0 27232 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1505_
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1506_
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1507_
timestamp 1644511149
transform 1 0 23184 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1508_
timestamp 1644511149
transform 1 0 25484 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1509_
timestamp 1644511149
transform 1 0 24656 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1510_
timestamp 1644511149
transform 1 0 24656 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1511_
timestamp 1644511149
transform 1 0 24748 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1512_
timestamp 1644511149
transform 1 0 25116 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1513_
timestamp 1644511149
transform 1 0 25852 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1514_
timestamp 1644511149
transform 1 0 25668 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1515_
timestamp 1644511149
transform 1 0 25024 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1516_
timestamp 1644511149
transform 1 0 25392 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1517_
timestamp 1644511149
transform 1 0 26312 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1518_
timestamp 1644511149
transform 1 0 23092 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1519_
timestamp 1644511149
transform 1 0 23000 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1520_
timestamp 1644511149
transform 1 0 22908 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1521_
timestamp 1644511149
transform 1 0 22632 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1522_
timestamp 1644511149
transform 1 0 23000 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1523_
timestamp 1644511149
transform 1 0 22724 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1524_
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1525_
timestamp 1644511149
transform 1 0 21988 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1526_
timestamp 1644511149
transform 1 0 23828 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1527_
timestamp 1644511149
transform 1 0 23092 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1528_
timestamp 1644511149
transform 1 0 23092 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1529_
timestamp 1644511149
transform 1 0 24104 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1530_
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1531_
timestamp 1644511149
transform 1 0 24840 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1532_
timestamp 1644511149
transform 1 0 25024 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1533_
timestamp 1644511149
transform 1 0 24472 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1534_
timestamp 1644511149
transform 1 0 25300 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1535_
timestamp 1644511149
transform 1 0 23368 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1536_
timestamp 1644511149
transform 1 0 23644 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1537_
timestamp 1644511149
transform 1 0 21620 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1538_
timestamp 1644511149
transform 1 0 22356 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1539_
timestamp 1644511149
transform 1 0 23276 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1540_
timestamp 1644511149
transform 1 0 20424 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1541_
timestamp 1644511149
transform 1 0 23184 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1542_
timestamp 1644511149
transform 1 0 22264 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1543_
timestamp 1644511149
transform 1 0 23092 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1544_
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1545_
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1546_
timestamp 1644511149
transform 1 0 20792 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1547_
timestamp 1644511149
transform 1 0 20424 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1548_
timestamp 1644511149
transform 1 0 22356 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1549_
timestamp 1644511149
transform 1 0 22356 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1550_
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1551_
timestamp 1644511149
transform 1 0 19412 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1552_
timestamp 1644511149
transform 1 0 20424 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1553_
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1554_
timestamp 1644511149
transform 1 0 20608 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1555_
timestamp 1644511149
transform 1 0 26680 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1556_
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1557_
timestamp 1644511149
transform 1 0 28612 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1558_
timestamp 1644511149
transform 1 0 29072 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1559_
timestamp 1644511149
transform 1 0 27784 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1560_
timestamp 1644511149
transform 1 0 27692 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1561_
timestamp 1644511149
transform 1 0 34868 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1562_
timestamp 1644511149
transform 1 0 33580 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1563_
timestamp 1644511149
transform 1 0 31832 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1564_
timestamp 1644511149
transform 1 0 33764 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1565_
timestamp 1644511149
transform 1 0 33672 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1566_
timestamp 1644511149
transform 1 0 35052 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1567_
timestamp 1644511149
transform 1 0 34960 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1568_
timestamp 1644511149
transform 1 0 35880 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1569_
timestamp 1644511149
transform 1 0 34776 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1570_
timestamp 1644511149
transform 1 0 34316 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1571_
timestamp 1644511149
transform 1 0 34776 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1572_
timestamp 1644511149
transform 1 0 33120 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1573_
timestamp 1644511149
transform 1 0 32384 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1574_
timestamp 1644511149
transform 1 0 17112 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1575_
timestamp 1644511149
transform 1 0 16468 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1576_
timestamp 1644511149
transform 1 0 15732 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1577_
timestamp 1644511149
transform 1 0 15824 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1578_
timestamp 1644511149
transform 1 0 17112 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1579_
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1580_
timestamp 1644511149
transform 1 0 17112 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1581_
timestamp 1644511149
transform 1 0 16928 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1582_
timestamp 1644511149
transform 1 0 17756 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1583_
timestamp 1644511149
transform 1 0 19596 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1584_
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1585_
timestamp 1644511149
transform 1 0 17112 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1586_
timestamp 1644511149
transform 1 0 15824 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1587_
timestamp 1644511149
transform 1 0 18308 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1588_
timestamp 1644511149
transform 1 0 17848 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1589_
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1590_
timestamp 1644511149
transform 1 0 9016 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1591_
timestamp 1644511149
transform 1 0 8004 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1592_
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1593_
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1594_
timestamp 1644511149
transform 1 0 20332 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1595_
timestamp 1644511149
transform 1 0 19688 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1596_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14168 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1597_
timestamp 1644511149
transform 1 0 15640 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1598_
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1599_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17204 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1600_
timestamp 1644511149
transform 1 0 17296 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1601_
timestamp 1644511149
transform 1 0 21528 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1602_
timestamp 1644511149
transform 1 0 19872 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1603_
timestamp 1644511149
transform 1 0 17296 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1604_
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1605_
timestamp 1644511149
transform 1 0 29716 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1606_
timestamp 1644511149
transform 1 0 31096 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1607_
timestamp 1644511149
transform 1 0 30452 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1608_
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1609_
timestamp 1644511149
transform 1 0 31464 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1610_
timestamp 1644511149
transform 1 0 32476 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1611_
timestamp 1644511149
transform 1 0 30820 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1612_
timestamp 1644511149
transform 1 0 32660 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1613_
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1614_
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1615_
timestamp 1644511149
transform 1 0 14628 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1616_
timestamp 1644511149
transform 1 0 11224 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1617_
timestamp 1644511149
transform 1 0 12788 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1618_
timestamp 1644511149
transform 1 0 14352 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1619_
timestamp 1644511149
transform 1 0 11408 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1620_
timestamp 1644511149
transform 1 0 7820 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1621_
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1622_
timestamp 1644511149
transform 1 0 8648 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1623_
timestamp 1644511149
transform 1 0 7176 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1624_
timestamp 1644511149
transform 1 0 9108 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1625_
timestamp 1644511149
transform 1 0 14168 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1626_
timestamp 1644511149
transform 1 0 11592 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1627_
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1628_
timestamp 1644511149
transform 1 0 15916 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1629_
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1630_
timestamp 1644511149
transform 1 0 20056 0 1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1631_
timestamp 1644511149
transform 1 0 17204 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1632_
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1633_
timestamp 1644511149
transform 1 0 20148 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1634_
timestamp 1644511149
transform 1 0 20792 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1635_
timestamp 1644511149
transform 1 0 22724 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1636_
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1637_
timestamp 1644511149
transform 1 0 16836 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1638_
timestamp 1644511149
transform 1 0 22816 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1639_
timestamp 1644511149
transform 1 0 24840 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1640_
timestamp 1644511149
transform 1 0 27876 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1641_
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1642_
timestamp 1644511149
transform 1 0 29716 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1643_
timestamp 1644511149
transform 1 0 29256 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1644_
timestamp 1644511149
transform 1 0 26772 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1645_
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1646_
timestamp 1644511149
transform 1 0 17480 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1647_
timestamp 1644511149
transform 1 0 17020 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1648_
timestamp 1644511149
transform 1 0 17296 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1649_
timestamp 1644511149
transform 1 0 19320 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1650_
timestamp 1644511149
transform 1 0 8188 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1651_
timestamp 1644511149
transform 1 0 21160 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1652_
timestamp 1644511149
transform 1 0 23184 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1653_
timestamp 1644511149
transform 1 0 18216 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1654_
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1655_
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1656_
timestamp 1644511149
transform 1 0 25760 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1657_
timestamp 1644511149
transform 1 0 27692 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1658_
timestamp 1644511149
transform 1 0 27968 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1659_
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1660_
timestamp 1644511149
transform 1 0 28796 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1661_
timestamp 1644511149
transform 1 0 28612 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1662_
timestamp 1644511149
transform 1 0 27600 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1663_
timestamp 1644511149
transform 1 0 24932 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1664_
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1665_
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1666_
timestamp 1644511149
transform 1 0 19504 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1667_
timestamp 1644511149
transform 1 0 16468 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1668_
timestamp 1644511149
transform 1 0 22448 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1669_
timestamp 1644511149
transform 1 0 14260 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1670_
timestamp 1644511149
transform 1 0 12144 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1671_
timestamp 1644511149
transform 1 0 12144 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1672_
timestamp 1644511149
transform 1 0 10856 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1673_
timestamp 1644511149
transform 1 0 8924 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1674_
timestamp 1644511149
transform 1 0 7084 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1675_
timestamp 1644511149
transform 1 0 8372 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1676_
timestamp 1644511149
transform 1 0 10304 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1677_
timestamp 1644511149
transform 1 0 28152 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1678_
timestamp 1644511149
transform 1 0 25944 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1679_
timestamp 1644511149
transform 1 0 31924 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1680_
timestamp 1644511149
transform 1 0 31832 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1681_
timestamp 1644511149
transform 1 0 32568 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1682_
timestamp 1644511149
transform 1 0 32752 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1683_
timestamp 1644511149
transform 1 0 32108 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1684_
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1685_
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1686_
timestamp 1644511149
transform 1 0 31464 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1687_
timestamp 1644511149
transform 1 0 31188 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1688_
timestamp 1644511149
transform 1 0 28520 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1689_
timestamp 1644511149
transform 1 0 32476 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1690_
timestamp 1644511149
transform 1 0 32660 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1691_
timestamp 1644511149
transform 1 0 28336 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1692_
timestamp 1644511149
transform 1 0 26864 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1693_
timestamp 1644511149
transform 1 0 25024 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1694_
timestamp 1644511149
transform 1 0 26772 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1695_
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1696_
timestamp 1644511149
transform 1 0 22724 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1697_
timestamp 1644511149
transform 1 0 22172 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1698_
timestamp 1644511149
transform 1 0 21988 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1699_
timestamp 1644511149
transform 1 0 25392 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1700_
timestamp 1644511149
transform 1 0 25392 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1701_
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1702_
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1703_
timestamp 1644511149
transform 1 0 23644 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1704_
timestamp 1644511149
transform 1 0 21068 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1705_
timestamp 1644511149
transform 1 0 20424 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1706_
timestamp 1644511149
transform 1 0 21804 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1707_
timestamp 1644511149
transform 1 0 19872 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1708_
timestamp 1644511149
transform 1 0 20056 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1709_
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1710_
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1711_
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1712_
timestamp 1644511149
transform 1 0 34224 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1713_
timestamp 1644511149
transform 1 0 35880 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1714_
timestamp 1644511149
transform 1 0 35328 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1715_
timestamp 1644511149
transform 1 0 35144 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1716_
timestamp 1644511149
transform 1 0 32292 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1717_
timestamp 1644511149
transform 1 0 15088 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1718_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17020 0 1 33728
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1719_
timestamp 1644511149
transform 1 0 16836 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1720_
timestamp 1644511149
transform 1 0 16928 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1721_
timestamp 1644511149
transform 1 0 16928 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1722_
timestamp 1644511149
transform 1 0 18400 0 -1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1723_
timestamp 1644511149
transform 1 0 7176 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1724_
timestamp 1644511149
transform 1 0 6992 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1725_
timestamp 1644511149
transform 1 0 20148 0 1 29376
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1726_
timestamp 1644511149
transform 1 0 13800 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1727_
timestamp 1644511149
transform 1 0 19872 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1728_
timestamp 1644511149
transform 1 0 14812 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1729__200 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 39928 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1730__201
timestamp 1644511149
transform 1 0 32108 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1731__202
timestamp 1644511149
transform 1 0 8924 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1732__203
timestamp 1644511149
transform 1 0 2668 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1733__96
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1734__97
timestamp 1644511149
transform 1 0 28060 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1735__98
timestamp 1644511149
transform 1 0 15916 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1736__99
timestamp 1644511149
transform 1 0 26036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1737__100
timestamp 1644511149
transform 1 0 35604 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1738__101
timestamp 1644511149
transform 1 0 2116 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1739__102
timestamp 1644511149
transform 1 0 47472 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1740__103
timestamp 1644511149
transform 1 0 1472 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1741__104
timestamp 1644511149
transform 1 0 1472 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1742__105
timestamp 1644511149
transform 1 0 2024 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1743__106
timestamp 1644511149
transform 1 0 30452 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1744__107
timestamp 1644511149
transform 1 0 15916 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1745__108
timestamp 1644511149
transform 1 0 2024 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1746__109
timestamp 1644511149
transform 1 0 31096 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1747__110
timestamp 1644511149
transform 1 0 4232 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1748__111
timestamp 1644511149
transform 1 0 47472 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1749__112
timestamp 1644511149
transform 1 0 22908 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1750__113
timestamp 1644511149
transform 1 0 10764 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1751__114
timestamp 1644511149
transform 1 0 29992 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1752__115
timestamp 1644511149
transform 1 0 19964 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1753__116
timestamp 1644511149
transform 1 0 41032 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1754__117
timestamp 1644511149
transform 1 0 45632 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1755__118
timestamp 1644511149
transform 1 0 5060 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1756__119
timestamp 1644511149
transform 1 0 42136 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1757__120
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1758__121
timestamp 1644511149
transform 1 0 2024 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1759__122
timestamp 1644511149
transform 1 0 17020 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1760__123
timestamp 1644511149
transform 1 0 20792 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1761__124
timestamp 1644511149
transform 1 0 14352 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1762__125
timestamp 1644511149
transform 1 0 29348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1763__126
timestamp 1644511149
transform 1 0 2024 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1764__127
timestamp 1644511149
transform 1 0 47564 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1765__128
timestamp 1644511149
transform 1 0 30452 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1766__129
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1767__130
timestamp 1644511149
transform 1 0 23184 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1768__131
timestamp 1644511149
transform 1 0 1840 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1769__132
timestamp 1644511149
transform 1 0 46184 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1770__133
timestamp 1644511149
transform 1 0 6716 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1771__134
timestamp 1644511149
transform 1 0 47564 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1772__135
timestamp 1644511149
transform 1 0 45172 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1773__136
timestamp 1644511149
transform 1 0 47564 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1774__137
timestamp 1644511149
transform 1 0 3036 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1775__138
timestamp 1644511149
transform 1 0 36248 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1776__139
timestamp 1644511149
transform 1 0 12236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1777__140
timestamp 1644511149
transform 1 0 47564 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1778__141
timestamp 1644511149
transform 1 0 45264 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1779__142
timestamp 1644511149
transform 1 0 38916 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1780__143
timestamp 1644511149
transform 1 0 10120 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1781__144
timestamp 1644511149
transform 1 0 7360 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1782__145
timestamp 1644511149
transform 1 0 47472 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1783__146
timestamp 1644511149
transform 1 0 33396 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1784__147
timestamp 1644511149
transform 1 0 14168 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1785__148
timestamp 1644511149
transform 1 0 1380 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1786__149
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1787__150
timestamp 1644511149
transform 1 0 2668 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1788__151
timestamp 1644511149
transform 1 0 47564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1789__152
timestamp 1644511149
transform 1 0 44068 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1790__153
timestamp 1644511149
transform 1 0 1564 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1791__154
timestamp 1644511149
transform 1 0 25208 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1792__155
timestamp 1644511149
transform 1 0 47564 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1793__156
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1794__157
timestamp 1644511149
transform 1 0 47748 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1795__158
timestamp 1644511149
transform 1 0 4508 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1796__159
timestamp 1644511149
transform 1 0 12972 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1797__160
timestamp 1644511149
transform 1 0 25668 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1798__161
timestamp 1644511149
transform 1 0 43240 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1799__162
timestamp 1644511149
transform 1 0 7912 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1800__163
timestamp 1644511149
transform 1 0 42596 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1801__164
timestamp 1644511149
transform 1 0 3036 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1802__165
timestamp 1644511149
transform 1 0 45632 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1803__166
timestamp 1644511149
transform 1 0 3772 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1804__167
timestamp 1644511149
transform 1 0 47748 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1805__168
timestamp 1644511149
transform 1 0 19780 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1806__169
timestamp 1644511149
transform 1 0 47472 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1807__170
timestamp 1644511149
transform 1 0 43884 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1808__171
timestamp 1644511149
transform 1 0 47564 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1809__172
timestamp 1644511149
transform 1 0 47564 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1810__173
timestamp 1644511149
transform 1 0 44988 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1811__174
timestamp 1644511149
transform 1 0 5612 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1812__175
timestamp 1644511149
transform 1 0 45632 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1813__176
timestamp 1644511149
transform 1 0 7452 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1814__177
timestamp 1644511149
transform 1 0 45632 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1815__178
timestamp 1644511149
transform 1 0 47564 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1816__179
timestamp 1644511149
transform 1 0 1840 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1817__180
timestamp 1644511149
transform 1 0 1840 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1818__181
timestamp 1644511149
transform 1 0 36340 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1819__182
timestamp 1644511149
transform 1 0 44988 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1820__183
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1821__184
timestamp 1644511149
transform 1 0 44252 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1822__185
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1823__186
timestamp 1644511149
transform 1 0 44620 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1824__187
timestamp 1644511149
transform 1 0 25024 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1825__188
timestamp 1644511149
transform 1 0 1840 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1826__189
timestamp 1644511149
transform 1 0 46828 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1827__190
timestamp 1644511149
transform 1 0 3772 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1828__191
timestamp 1644511149
transform 1 0 11592 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1829__192
timestamp 1644511149
transform 1 0 43240 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1830__193
timestamp 1644511149
transform 1 0 3312 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1831__194
timestamp 1644511149
transform 1 0 32752 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1832__195
timestamp 1644511149
transform 1 0 22448 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1833__196
timestamp 1644511149
transform 1 0 4048 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1834__197
timestamp 1644511149
transform 1 0 2668 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1835__198
timestamp 1644511149
transform 1 0 38732 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1836__199
timestamp 1644511149
transform 1 0 2024 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1837_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1838_
timestamp 1644511149
transform 1 0 11500 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1839_
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1840_
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1841_
timestamp 1644511149
transform 1 0 17940 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1842_
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1843_
timestamp 1644511149
transform 1 0 29808 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1844_
timestamp 1644511149
transform 1 0 32200 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1845_
timestamp 1644511149
transform 1 0 29716 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1846_
timestamp 1644511149
transform 1 0 33304 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1847_
timestamp 1644511149
transform 1 0 32844 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1848_
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1849_
timestamp 1644511149
transform 1 0 31372 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1850_
timestamp 1644511149
transform 1 0 34500 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1851_
timestamp 1644511149
transform 1 0 33212 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1852_
timestamp 1644511149
transform 1 0 32200 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1853_
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1854_
timestamp 1644511149
transform 1 0 12328 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1855_
timestamp 1644511149
transform 1 0 13800 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1856_
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1857_
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1858_
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1859_
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1860_
timestamp 1644511149
transform 1 0 6440 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1861_
timestamp 1644511149
transform 1 0 6440 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1862_
timestamp 1644511149
transform 1 0 9844 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1863_
timestamp 1644511149
transform 1 0 3312 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1864_
timestamp 1644511149
transform 1 0 27324 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1865_
timestamp 1644511149
transform 1 0 16928 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1866_
timestamp 1644511149
transform 1 0 25944 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1867_
timestamp 1644511149
transform 1 0 35512 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1868_
timestamp 1644511149
transform 1 0 2024 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1869_
timestamp 1644511149
transform 1 0 46276 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_2  _1870_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7636 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_8  _1871_
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1872_
timestamp 1644511149
transform 1 0 29624 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1873_
timestamp 1644511149
transform 1 0 19228 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1874_
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1875_
timestamp 1644511149
transform 1 0 39928 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1876_
timestamp 1644511149
transform 1 0 32108 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1877_
timestamp 1644511149
transform 1 0 8924 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1878_
timestamp 1644511149
transform 1 0 1840 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1879_
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1880_
timestamp 1644511149
transform 1 0 1932 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1881_
timestamp 1644511149
transform 1 0 31096 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1882_
timestamp 1644511149
transform 1 0 16560 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1883_
timestamp 1644511149
transform 1 0 2024 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1884_
timestamp 1644511149
transform 1 0 31004 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1885_
timestamp 1644511149
transform 1 0 4416 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1886_
timestamp 1644511149
transform 1 0 46276 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1887_
timestamp 1644511149
transform 1 0 23184 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1888_
timestamp 1644511149
transform 1 0 11500 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1889_
timestamp 1644511149
transform 1 0 29716 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1890_
timestamp 1644511149
transform 1 0 19964 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1891_
timestamp 1644511149
transform 1 0 41492 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1892_
timestamp 1644511149
transform 1 0 46276 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1893_
timestamp 1644511149
transform 1 0 2024 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1894_
timestamp 1644511149
transform 1 0 42412 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1895_
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1896_
timestamp 1644511149
transform 1 0 1932 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1897_
timestamp 1644511149
transform 1 0 17296 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1898_
timestamp 1644511149
transform 1 0 20240 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1899_
timestamp 1644511149
transform 1 0 14260 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1900_
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1901_
timestamp 1644511149
transform 1 0 1932 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1902_
timestamp 1644511149
transform 1 0 46276 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1903_
timestamp 1644511149
transform 1 0 29716 0 1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1904_
timestamp 1644511149
transform 1 0 1748 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1905_
timestamp 1644511149
transform 1 0 22632 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1906_
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1907_
timestamp 1644511149
transform 1 0 46276 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1908_
timestamp 1644511149
transform 1 0 1932 0 -1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1909_
timestamp 1644511149
transform 1 0 46276 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1910_
timestamp 1644511149
transform 1 0 46000 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1911_
timestamp 1644511149
transform 1 0 46276 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1912_
timestamp 1644511149
transform 1 0 2668 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1913_
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1914_
timestamp 1644511149
transform 1 0 45816 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1915_
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1916_
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1917_
timestamp 1644511149
transform 1 0 18676 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1918_
timestamp 1644511149
transform 1 0 46276 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1919_
timestamp 1644511149
transform 1 0 8280 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1920_
timestamp 1644511149
transform 1 0 6808 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1921_
timestamp 1644511149
transform 1 0 34868 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1922_
timestamp 1644511149
transform 1 0 11960 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1923_
timestamp 1644511149
transform 1 0 46276 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1924_
timestamp 1644511149
transform 1 0 45172 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1925_
timestamp 1644511149
transform 1 0 39560 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1926_
timestamp 1644511149
transform 1 0 10488 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1927_
timestamp 1644511149
transform 1 0 6348 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1928_
timestamp 1644511149
transform 1 0 45172 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1929_
timestamp 1644511149
transform 1 0 27048 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1930_
timestamp 1644511149
transform 1 0 23000 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1931_
timestamp 1644511149
transform 1 0 35972 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1932_
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1933_
timestamp 1644511149
transform 1 0 38088 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1934_
timestamp 1644511149
transform 1 0 37260 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1935_
timestamp 1644511149
transform 1 0 36616 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1936_
timestamp 1644511149
transform 1 0 33580 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1937_
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1938_
timestamp 1644511149
transform 1 0 32292 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1939_
timestamp 1644511149
transform 1 0 15088 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1940_
timestamp 1644511149
transform 1 0 29716 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1941_
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1942_
timestamp 1644511149
transform 1 0 16744 0 -1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1943_
timestamp 1644511149
transform 1 0 33304 0 -1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1944_
timestamp 1644511149
transform 1 0 14168 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1945_
timestamp 1644511149
transform 1 0 1380 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1946_
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1947_
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1948_
timestamp 1644511149
transform 1 0 46276 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1949_
timestamp 1644511149
transform 1 0 43976 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1950_
timestamp 1644511149
transform 1 0 2116 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1951_
timestamp 1644511149
transform 1 0 27692 0 -1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1952_
timestamp 1644511149
transform 1 0 46276 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1953_
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1954_
timestamp 1644511149
transform 1 0 46276 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1955_
timestamp 1644511149
transform 1 0 4416 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1956_
timestamp 1644511149
transform 1 0 12880 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1957_
timestamp 1644511149
transform 1 0 26312 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1958_
timestamp 1644511149
transform 1 0 43240 0 -1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1959_
timestamp 1644511149
transform 1 0 6624 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1960_
timestamp 1644511149
transform 1 0 42596 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1961_
timestamp 1644511149
transform 1 0 1932 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1962_
timestamp 1644511149
transform 1 0 46276 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1963_
timestamp 1644511149
transform 1 0 1840 0 -1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1964_
timestamp 1644511149
transform 1 0 46276 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1965_
timestamp 1644511149
transform 1 0 20056 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1966_
timestamp 1644511149
transform 1 0 46276 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1967_
timestamp 1644511149
transform 1 0 45172 0 1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1968_
timestamp 1644511149
transform 1 0 46276 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1969_
timestamp 1644511149
transform 1 0 46276 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1970_
timestamp 1644511149
transform 1 0 44988 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1971_
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1972_
timestamp 1644511149
transform 1 0 46276 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1973_
timestamp 1644511149
transform 1 0 7084 0 -1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1974_
timestamp 1644511149
transform 1 0 46276 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1975_
timestamp 1644511149
transform 1 0 46276 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1976_
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1977_
timestamp 1644511149
transform 1 0 1380 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1978_
timestamp 1644511149
transform 1 0 36340 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1979_
timestamp 1644511149
transform 1 0 45172 0 -1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1980_
timestamp 1644511149
transform 1 0 1748 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1981_
timestamp 1644511149
transform 1 0 44988 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1982_
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1983_
timestamp 1644511149
transform 1 0 42596 0 1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1984_
timestamp 1644511149
transform 1 0 24380 0 1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1985_
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1986_
timestamp 1644511149
transform 1 0 46276 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1987_
timestamp 1644511149
transform 1 0 1380 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1988_
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1989_
timestamp 1644511149
transform 1 0 45172 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1990_
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1991_
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1992_
timestamp 1644511149
transform 1 0 21988 0 1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1993_
timestamp 1644511149
transform 1 0 1748 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1994_
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1995_
timestamp 1644511149
transform 1 0 38732 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1996_
timestamp 1644511149
transform 1 0 2024 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21344 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 20976 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 23552 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 18216 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 26036 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 18768 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 28612 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 17572 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 16468 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 28336 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 29440 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_4_0_wb_clk_i
timestamp 1644511149
transform 1 0 17940 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_5_0_wb_clk_i
timestamp 1644511149
transform 1 0 17848 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_6_0_wb_clk_i
timestamp 1644511149
transform 1 0 28704 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_7_0_wb_clk_i
timestamp 1644511149
transform 1 0 29348 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 17112 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 18308 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 15732 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 17480 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_4_0_wb_clk_i
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_5_0_wb_clk_i
timestamp 1644511149
transform 1 0 27968 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_6_0_wb_clk_i
timestamp 1644511149
transform 1 0 28428 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_7_0_wb_clk_i
timestamp 1644511149
transform 1 0 30176 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_8_0_wb_clk_i
timestamp 1644511149
transform 1 0 14996 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_9_0_wb_clk_i
timestamp 1644511149
transform 1 0 18308 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_10_0_wb_clk_i
timestamp 1644511149
transform 1 0 15732 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_11_0_wb_clk_i
timestamp 1644511149
transform 1 0 18860 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_12_0_wb_clk_i
timestamp 1644511149
transform 1 0 27416 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_13_0_wb_clk_i
timestamp 1644511149
transform 1 0 30268 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_14_0_wb_clk_i
timestamp 1644511149
transform 1 0 26496 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_15_0_wb_clk_i
timestamp 1644511149
transform 1 0 30636 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  hold1
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input1
timestamp 1644511149
transform 1 0 47656 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input2
timestamp 1644511149
transform 1 0 1748 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 1644511149
transform 1 0 13248 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 1644511149
transform 1 0 22632 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input6
timestamp 1644511149
transform 1 0 47656 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input7
timestamp 1644511149
transform 1 0 47840 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1644511149
transform 1 0 21896 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1644511149
transform 1 0 12788 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1644511149
transform 1 0 17848 0 1 48960
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input11
timestamp 1644511149
transform 1 0 27048 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input12
timestamp 1644511149
transform 1 0 32936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1644511149
transform 1 0 1748 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input14
timestamp 1644511149
transform 1 0 8924 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input15
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1644511149
transform 1 0 17020 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input17
timestamp 1644511149
transform 1 0 47656 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1644511149
transform 1 0 47840 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1644511149
transform 1 0 47840 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1644511149
transform 1 0 47840 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1644511149
transform 1 0 23920 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1644511149
transform 1 0 2668 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1644511149
transform 1 0 47840 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input25
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input26
timestamp 1644511149
transform 1 0 47656 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1644511149
transform 1 0 14260 0 1 48960
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 1644511149
transform 1 0 47288 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input29
timestamp 1644511149
transform 1 0 47288 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input30
timestamp 1644511149
transform 1 0 1380 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input31
timestamp 1644511149
transform 1 0 5060 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input32
timestamp 1644511149
transform 1 0 20056 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1644511149
transform 1 0 1748 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input34
timestamp 1644511149
transform 1 0 40664 0 1 48960
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1644511149
transform 1 0 27324 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1644511149
transform 1 0 1748 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1644511149
transform 1 0 38088 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input38
timestamp 1644511149
transform 1 0 20056 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1644511149
transform 1 0 6716 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input41
timestamp 1644511149
transform 1 0 47840 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1644511149
transform 1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input43
timestamp 1644511149
transform 1 0 27784 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input44
timestamp 1644511149
transform 1 0 1748 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1644511149
transform 1 0 1748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1644511149
transform 1 0 43240 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input47
timestamp 1644511149
transform 1 0 44988 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input48
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1644511149
transform 1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1644511149
transform 1 0 36156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1644511149
transform 1 0 47840 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1644511149
transform 1 0 19320 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input53
timestamp 1644511149
transform 1 0 24564 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input54
timestamp 1644511149
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1644511149
transform 1 0 28704 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1644511149
transform 1 0 47932 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1644511149
transform 1 0 46184 0 -1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input58
timestamp 1644511149
transform 1 0 17480 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1644511149
transform 1 0 47840 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1644511149
transform 1 0 46828 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input61
timestamp 1644511149
transform 1 0 34868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input62
timestamp 1644511149
transform 1 0 47656 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1644511149
transform 1 0 33856 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 1644511149
transform 1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input65
timestamp 1644511149
transform 1 0 1380 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input66
timestamp 1644511149
transform 1 0 46276 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1644511149
transform 1 0 47840 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1644511149
transform 1 0 25852 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input69
timestamp 1644511149
transform 1 0 47840 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input70
timestamp 1644511149
transform 1 0 1748 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input71
timestamp 1644511149
transform 1 0 4140 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input72
timestamp 1644511149
transform 1 0 4324 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input73
timestamp 1644511149
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1644511149
transform 1 0 10212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input75
timestamp 1644511149
transform 1 0 47840 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input76
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input77
timestamp 1644511149
transform 1 0 41676 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input78
timestamp 1644511149
transform 1 0 47656 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input79
timestamp 1644511149
transform 1 0 11868 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input80
timestamp 1644511149
transform 1 0 7176 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input81
timestamp 1644511149
transform 1 0 47840 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input82
timestamp 1644511149
transform 1 0 47656 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input83
timestamp 1644511149
transform 1 0 1748 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input84
timestamp 1644511149
transform 1 0 47840 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input85
timestamp 1644511149
transform 1 0 1748 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input86
timestamp 1644511149
transform 1 0 38456 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input87
timestamp 1644511149
transform 1 0 47840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input88
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1644511149
transform 1 0 23368 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input90
timestamp 1644511149
transform 1 0 47840 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input91
timestamp 1644511149
transform 1 0 43884 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input92
timestamp 1644511149
transform 1 0 47840 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input93
timestamp 1644511149
transform 1 0 47840 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input94
timestamp 1644511149
transform 1 0 1748 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input95
timestamp 1644511149
transform 1 0 47840 0 -1 25024
box -38 -48 406 592
<< labels >>
rlabel metal3 s 49200 31968 50000 32088 6 active
port 0 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 25134 51200 25190 52000 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 49200 15648 50000 15768 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 21270 51200 21326 52000 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 49200 2048 50000 2168 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 io_in[18]
port 10 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 49200 18368 50000 18488 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 0 30608 800 30728 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 49200 21088 50000 21208 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 49200 32648 50000 32768 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 49200 23128 50000 23248 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 2594 51200 2650 52000 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 46386 51200 46442 52000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 9034 51200 9090 52000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 31574 51200 31630 52000 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 49200 47608 50000 47728 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 49200 20408 50000 20528 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 35438 51200 35494 52000 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 49200 2728 50000 2848 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 3882 51200 3938 52000 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 io_oeb[0]
port 39 nsew signal tristate
rlabel metal3 s 49200 24488 50000 24608 6 io_oeb[10]
port 40 nsew signal tristate
rlabel metal2 s 45098 0 45154 800 6 io_oeb[11]
port 41 nsew signal tristate
rlabel metal2 s 5814 0 5870 800 6 io_oeb[12]
port 42 nsew signal tristate
rlabel metal2 s 48318 0 48374 800 6 io_oeb[13]
port 43 nsew signal tristate
rlabel metal2 s 7746 51200 7802 52000 6 io_oeb[14]
port 44 nsew signal tristate
rlabel metal3 s 49200 43528 50000 43648 6 io_oeb[15]
port 45 nsew signal tristate
rlabel metal3 s 49200 4768 50000 4888 6 io_oeb[16]
port 46 nsew signal tristate
rlabel metal3 s 0 6808 800 6928 6 io_oeb[17]
port 47 nsew signal tristate
rlabel metal3 s 0 41488 800 41608 6 io_oeb[18]
port 48 nsew signal tristate
rlabel metal2 s 36726 0 36782 800 6 io_oeb[19]
port 49 nsew signal tristate
rlabel metal2 s 43166 51200 43222 52000 6 io_oeb[1]
port 50 nsew signal tristate
rlabel metal3 s 49200 46928 50000 47048 6 io_oeb[20]
port 51 nsew signal tristate
rlabel metal3 s 0 9528 800 9648 6 io_oeb[21]
port 52 nsew signal tristate
rlabel metal2 s 45098 51200 45154 52000 6 io_oeb[22]
port 53 nsew signal tristate
rlabel metal3 s 0 26528 800 26648 6 io_oeb[23]
port 54 nsew signal tristate
rlabel metal3 s 49200 51688 50000 51808 6 io_oeb[24]
port 55 nsew signal tristate
rlabel metal2 s 24490 51200 24546 52000 6 io_oeb[25]
port 56 nsew signal tristate
rlabel metal3 s 0 23128 800 23248 6 io_oeb[26]
port 57 nsew signal tristate
rlabel metal3 s 49200 28568 50000 28688 6 io_oeb[27]
port 58 nsew signal tristate
rlabel metal2 s 1306 51200 1362 52000 6 io_oeb[28]
port 59 nsew signal tristate
rlabel metal2 s 12254 0 12310 800 6 io_oeb[29]
port 60 nsew signal tristate
rlabel metal3 s 0 51688 800 51808 6 io_oeb[2]
port 61 nsew signal tristate
rlabel metal2 s 49606 51200 49662 52000 6 io_oeb[30]
port 62 nsew signal tristate
rlabel metal3 s 0 3408 800 3528 6 io_oeb[31]
port 63 nsew signal tristate
rlabel metal2 s 33506 0 33562 800 6 io_oeb[32]
port 64 nsew signal tristate
rlabel metal2 s 22558 51200 22614 52000 6 io_oeb[33]
port 65 nsew signal tristate
rlabel metal3 s 0 17688 800 17808 6 io_oeb[34]
port 66 nsew signal tristate
rlabel metal3 s 0 13608 800 13728 6 io_oeb[35]
port 67 nsew signal tristate
rlabel metal2 s 39946 0 40002 800 6 io_oeb[36]
port 68 nsew signal tristate
rlabel metal3 s 0 39448 800 39568 6 io_oeb[37]
port 69 nsew signal tristate
rlabel metal3 s 49200 45568 50000 45688 6 io_oeb[3]
port 70 nsew signal tristate
rlabel metal3 s 0 44888 800 45008 6 io_oeb[4]
port 71 nsew signal tristate
rlabel metal3 s 49200 36728 50000 36848 6 io_oeb[5]
port 72 nsew signal tristate
rlabel metal2 s 21270 0 21326 800 6 io_oeb[6]
port 73 nsew signal tristate
rlabel metal3 s 49200 17008 50000 17128 6 io_oeb[7]
port 74 nsew signal tristate
rlabel metal3 s 49200 49648 50000 49768 6 io_oeb[8]
port 75 nsew signal tristate
rlabel metal3 s 49200 16328 50000 16448 6 io_oeb[9]
port 76 nsew signal tristate
rlabel metal2 s 36082 51200 36138 52000 6 io_out[0]
port 77 nsew signal tristate
rlabel metal3 s 49200 44208 50000 44328 6 io_out[10]
port 78 nsew signal tristate
rlabel metal3 s 49200 9528 50000 9648 6 io_out[11]
port 79 nsew signal tristate
rlabel metal2 s 48962 0 49018 800 6 io_out[12]
port 80 nsew signal tristate
rlabel metal2 s 47030 0 47086 800 6 io_out[13]
port 81 nsew signal tristate
rlabel metal3 s 49200 12248 50000 12368 6 io_out[14]
port 82 nsew signal tristate
rlabel metal2 s 37370 0 37426 800 6 io_out[15]
port 83 nsew signal tristate
rlabel metal2 s 37370 51200 37426 52000 6 io_out[16]
port 84 nsew signal tristate
rlabel metal2 s 38658 51200 38714 52000 6 io_out[17]
port 85 nsew signal tristate
rlabel metal2 s 15474 51200 15530 52000 6 io_out[18]
port 86 nsew signal tristate
rlabel metal3 s 49200 3408 50000 3528 6 io_out[19]
port 87 nsew signal tristate
rlabel metal2 s 12898 0 12954 800 6 io_out[1]
port 88 nsew signal tristate
rlabel metal2 s 11610 0 11666 800 6 io_out[20]
port 89 nsew signal tristate
rlabel metal3 s 0 48288 800 48408 6 io_out[21]
port 90 nsew signal tristate
rlabel metal2 s 34794 51200 34850 52000 6 io_out[22]
port 91 nsew signal tristate
rlabel metal2 s 14830 51200 14886 52000 6 io_out[23]
port 92 nsew signal tristate
rlabel metal3 s 0 46248 800 46368 6 io_out[24]
port 93 nsew signal tristate
rlabel metal3 s 0 34008 800 34128 6 io_out[25]
port 94 nsew signal tristate
rlabel metal3 s 0 27208 800 27328 6 io_out[26]
port 95 nsew signal tristate
rlabel metal3 s 49200 7488 50000 7608 6 io_out[27]
port 96 nsew signal tristate
rlabel metal2 s 44454 0 44510 800 6 io_out[28]
port 97 nsew signal tristate
rlabel metal3 s 0 5448 800 5568 6 io_out[29]
port 98 nsew signal tristate
rlabel metal3 s 49200 35368 50000 35488 6 io_out[2]
port 99 nsew signal tristate
rlabel metal2 s 28354 51200 28410 52000 6 io_out[30]
port 100 nsew signal tristate
rlabel metal3 s 49200 46248 50000 46368 6 io_out[31]
port 101 nsew signal tristate
rlabel metal2 s 42522 0 42578 800 6 io_out[32]
port 102 nsew signal tristate
rlabel metal3 s 49200 10888 50000 11008 6 io_out[33]
port 103 nsew signal tristate
rlabel metal3 s 0 51008 800 51128 6 io_out[34]
port 104 nsew signal tristate
rlabel metal2 s 13542 0 13598 800 6 io_out[35]
port 105 nsew signal tristate
rlabel metal2 s 27066 51200 27122 52000 6 io_out[36]
port 106 nsew signal tristate
rlabel metal2 s 48318 51200 48374 52000 6 io_out[37]
port 107 nsew signal tristate
rlabel metal2 s 45742 51200 45798 52000 6 io_out[3]
port 108 nsew signal tristate
rlabel metal2 s 39946 51200 40002 52000 6 io_out[4]
port 109 nsew signal tristate
rlabel metal2 s 10322 51200 10378 52000 6 io_out[5]
port 110 nsew signal tristate
rlabel metal2 s 7102 51200 7158 52000 6 io_out[6]
port 111 nsew signal tristate
rlabel metal3 s 49200 34008 50000 34128 6 io_out[7]
port 112 nsew signal tristate
rlabel metal2 s 2594 0 2650 800 6 io_out[8]
port 113 nsew signal tristate
rlabel metal2 s 8390 51200 8446 52000 6 io_out[9]
port 114 nsew signal tristate
rlabel metal3 s 0 8168 800 8288 6 rambus_wb_ack_i
port 115 nsew signal input
rlabel metal3 s 49200 40128 50000 40248 6 rambus_wb_adr_o[0]
port 116 nsew signal tristate
rlabel metal3 s 0 46928 800 47048 6 rambus_wb_adr_o[1]
port 117 nsew signal tristate
rlabel metal2 s 10966 51200 11022 52000 6 rambus_wb_adr_o[2]
port 118 nsew signal tristate
rlabel metal3 s 49200 6128 50000 6248 6 rambus_wb_adr_o[3]
port 119 nsew signal tristate
rlabel metal3 s 49200 51008 50000 51128 6 rambus_wb_adr_o[4]
port 120 nsew signal tristate
rlabel metal3 s 49200 17688 50000 17808 6 rambus_wb_adr_o[5]
port 121 nsew signal tristate
rlabel metal3 s 49200 6808 50000 6928 6 rambus_wb_adr_o[6]
port 122 nsew signal tristate
rlabel metal3 s 49200 29248 50000 29368 6 rambus_wb_adr_o[7]
port 123 nsew signal tristate
rlabel metal2 s 9034 0 9090 800 6 rambus_wb_adr_o[8]
port 124 nsew signal tristate
rlabel metal3 s 0 2048 800 2168 6 rambus_wb_adr_o[9]
port 125 nsew signal tristate
rlabel metal3 s 0 18368 800 18488 6 rambus_wb_clk_o
port 126 nsew signal tristate
rlabel metal2 s 5170 51200 5226 52000 6 rambus_wb_cyc_o
port 127 nsew signal tristate
rlabel metal2 s 13542 51200 13598 52000 6 rambus_wb_dat_i[0]
port 128 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 rambus_wb_dat_i[10]
port 129 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 rambus_wb_dat_i[11]
port 130 nsew signal input
rlabel metal3 s 49200 688 50000 808 6 rambus_wb_dat_i[12]
port 131 nsew signal input
rlabel metal3 s 49200 13608 50000 13728 6 rambus_wb_dat_i[13]
port 132 nsew signal input
rlabel metal2 s 21914 51200 21970 52000 6 rambus_wb_dat_i[14]
port 133 nsew signal input
rlabel metal2 s 12898 51200 12954 52000 6 rambus_wb_dat_i[15]
port 134 nsew signal input
rlabel metal2 s 18050 51200 18106 52000 6 rambus_wb_dat_i[16]
port 135 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 rambus_wb_dat_i[17]
port 136 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 rambus_wb_dat_i[18]
port 137 nsew signal input
rlabel metal3 s 0 34688 800 34808 6 rambus_wb_dat_i[19]
port 138 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 rambus_wb_dat_i[1]
port 139 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 rambus_wb_dat_i[20]
port 140 nsew signal input
rlabel metal2 s 16118 51200 16174 52000 6 rambus_wb_dat_i[21]
port 141 nsew signal input
rlabel metal3 s 49200 8168 50000 8288 6 rambus_wb_dat_i[22]
port 142 nsew signal input
rlabel metal3 s 49200 31288 50000 31408 6 rambus_wb_dat_i[23]
port 143 nsew signal input
rlabel metal3 s 49200 33328 50000 33448 6 rambus_wb_dat_i[24]
port 144 nsew signal input
rlabel metal3 s 49200 38768 50000 38888 6 rambus_wb_dat_i[25]
port 145 nsew signal input
rlabel metal2 s 23846 51200 23902 52000 6 rambus_wb_dat_i[26]
port 146 nsew signal input
rlabel metal3 s 0 36728 800 36848 6 rambus_wb_dat_i[27]
port 147 nsew signal input
rlabel metal2 s 18 51200 74 52000 6 rambus_wb_dat_i[28]
port 148 nsew signal input
rlabel metal3 s 49200 42168 50000 42288 6 rambus_wb_dat_i[29]
port 149 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 rambus_wb_dat_i[2]
port 150 nsew signal input
rlabel metal3 s 49200 10208 50000 10328 6 rambus_wb_dat_i[30]
port 151 nsew signal input
rlabel metal2 s 14186 51200 14242 52000 6 rambus_wb_dat_i[31]
port 152 nsew signal input
rlabel metal3 s 49200 29928 50000 30048 6 rambus_wb_dat_i[3]
port 153 nsew signal input
rlabel metal3 s 49200 23808 50000 23928 6 rambus_wb_dat_i[4]
port 154 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 rambus_wb_dat_i[5]
port 155 nsew signal input
rlabel metal2 s 4526 51200 4582 52000 6 rambus_wb_dat_i[6]
port 156 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 rambus_wb_dat_i[7]
port 157 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 rambus_wb_dat_i[8]
port 158 nsew signal input
rlabel metal2 s 40590 51200 40646 52000 6 rambus_wb_dat_i[9]
port 159 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 rambus_wb_dat_o[0]
port 160 nsew signal tristate
rlabel metal2 s 30286 0 30342 800 6 rambus_wb_dat_o[10]
port 161 nsew signal tristate
rlabel metal2 s 20626 0 20682 800 6 rambus_wb_dat_o[11]
port 162 nsew signal tristate
rlabel metal2 s 41878 0 41934 800 6 rambus_wb_dat_o[12]
port 163 nsew signal tristate
rlabel metal3 s 49200 34688 50000 34808 6 rambus_wb_dat_o[13]
port 164 nsew signal tristate
rlabel metal3 s 0 50328 800 50448 6 rambus_wb_dat_o[14]
port 165 nsew signal tristate
rlabel metal2 s 42522 51200 42578 52000 6 rambus_wb_dat_o[15]
port 166 nsew signal tristate
rlabel metal2 s 1306 0 1362 800 6 rambus_wb_dat_o[16]
port 167 nsew signal tristate
rlabel metal3 s 0 29928 800 30048 6 rambus_wb_dat_o[17]
port 168 nsew signal tristate
rlabel metal2 s 18050 0 18106 800 6 rambus_wb_dat_o[18]
port 169 nsew signal tristate
rlabel metal2 s 20626 51200 20682 52000 6 rambus_wb_dat_o[19]
port 170 nsew signal tristate
rlabel metal3 s 0 10208 800 10328 6 rambus_wb_dat_o[1]
port 171 nsew signal tristate
rlabel metal2 s 15474 0 15530 800 6 rambus_wb_dat_o[20]
port 172 nsew signal tristate
rlabel metal2 s 30930 0 30986 800 6 rambus_wb_dat_o[21]
port 173 nsew signal tristate
rlabel metal3 s 0 31968 800 32088 6 rambus_wb_dat_o[22]
port 174 nsew signal tristate
rlabel metal3 s 49200 19728 50000 19848 6 rambus_wb_dat_o[23]
port 175 nsew signal tristate
rlabel metal2 s 30930 51200 30986 52000 6 rambus_wb_dat_o[24]
port 176 nsew signal tristate
rlabel metal3 s 0 16328 800 16448 6 rambus_wb_dat_o[25]
port 177 nsew signal tristate
rlabel metal2 s 23202 51200 23258 52000 6 rambus_wb_dat_o[26]
port 178 nsew signal tristate
rlabel metal3 s 0 28568 800 28688 6 rambus_wb_dat_o[27]
port 179 nsew signal tristate
rlabel metal3 s 49200 50328 50000 50448 6 rambus_wb_dat_o[28]
port 180 nsew signal tristate
rlabel metal3 s 0 48968 800 49088 6 rambus_wb_dat_o[29]
port 181 nsew signal tristate
rlabel metal2 s 31574 0 31630 800 6 rambus_wb_dat_o[2]
port 182 nsew signal tristate
rlabel metal3 s 49200 41488 50000 41608 6 rambus_wb_dat_o[30]
port 183 nsew signal tristate
rlabel metal2 s 46386 0 46442 800 6 rambus_wb_dat_o[31]
port 184 nsew signal tristate
rlabel metal2 s 17406 51200 17462 52000 6 rambus_wb_dat_o[3]
port 185 nsew signal tristate
rlabel metal3 s 0 32648 800 32768 6 rambus_wb_dat_o[4]
port 186 nsew signal tristate
rlabel metal2 s 32218 51200 32274 52000 6 rambus_wb_dat_o[5]
port 187 nsew signal tristate
rlabel metal2 s 5170 0 5226 800 6 rambus_wb_dat_o[6]
port 188 nsew signal tristate
rlabel metal3 s 49200 14288 50000 14408 6 rambus_wb_dat_o[7]
port 189 nsew signal tristate
rlabel metal2 s 23846 0 23902 800 6 rambus_wb_dat_o[8]
port 190 nsew signal tristate
rlabel metal2 s 12254 51200 12310 52000 6 rambus_wb_dat_o[9]
port 191 nsew signal tristate
rlabel metal3 s 0 8848 800 8968 6 rambus_wb_rst_o
port 192 nsew signal tristate
rlabel metal2 s 41234 0 41290 800 6 rambus_wb_sel_o[0]
port 193 nsew signal tristate
rlabel metal2 s 32862 51200 32918 52000 6 rambus_wb_sel_o[1]
port 194 nsew signal tristate
rlabel metal2 s 9678 51200 9734 52000 6 rambus_wb_sel_o[2]
port 195 nsew signal tristate
rlabel metal3 s 0 33328 800 33448 6 rambus_wb_sel_o[3]
port 196 nsew signal tristate
rlabel metal2 s 29642 51200 29698 52000 6 rambus_wb_stb_o
port 197 nsew signal tristate
rlabel metal3 s 0 4768 800 4888 6 rambus_wb_we_o
port 198 nsew signal tristate
rlabel metal4 s 4208 2128 4528 49552 6 vccd1
port 199 nsew power input
rlabel metal4 s 34928 2128 35248 49552 6 vccd1
port 199 nsew power input
rlabel metal4 s 19568 2128 19888 49552 6 vssd1
port 200 nsew ground input
rlabel metal3 s 49200 1368 50000 1488 6 wb_clk_i
port 201 nsew signal input
rlabel metal2 s 26422 51200 26478 52000 6 wb_rst_i
port 202 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 wbs_ack_o
port 203 nsew signal tristate
rlabel metal3 s 0 31288 800 31408 6 wbs_adr_i[0]
port 204 nsew signal input
rlabel metal2 s 38014 51200 38070 52000 6 wbs_adr_i[10]
port 205 nsew signal input
rlabel metal2 s 19982 51200 20038 52000 6 wbs_adr_i[11]
port 206 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 wbs_adr_i[12]
port 207 nsew signal input
rlabel metal2 s 6458 51200 6514 52000 6 wbs_adr_i[13]
port 208 nsew signal input
rlabel metal3 s 49200 27888 50000 28008 6 wbs_adr_i[14]
port 209 nsew signal input
rlabel metal3 s 0 688 800 808 6 wbs_adr_i[15]
port 210 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 wbs_adr_i[16]
port 211 nsew signal input
rlabel metal3 s 0 44208 800 44328 6 wbs_adr_i[17]
port 212 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 wbs_adr_i[18]
port 213 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 wbs_adr_i[19]
port 214 nsew signal input
rlabel metal2 s 44454 51200 44510 52000 6 wbs_adr_i[1]
port 215 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 wbs_adr_i[20]
port 216 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 wbs_adr_i[21]
port 217 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wbs_adr_i[22]
port 218 nsew signal input
rlabel metal3 s 49200 5448 50000 5568 6 wbs_adr_i[23]
port 219 nsew signal input
rlabel metal2 s 19338 51200 19394 52000 6 wbs_adr_i[24]
port 220 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_adr_i[25]
port 221 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_adr_i[26]
port 222 nsew signal input
rlabel metal2 s 28998 51200 29054 52000 6 wbs_adr_i[27]
port 223 nsew signal input
rlabel metal3 s 49200 22448 50000 22568 6 wbs_adr_i[28]
port 224 nsew signal input
rlabel metal3 s 49200 40808 50000 40928 6 wbs_adr_i[29]
port 225 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_adr_i[2]
port 226 nsew signal input
rlabel metal2 s 48962 51200 49018 52000 6 wbs_adr_i[30]
port 227 nsew signal input
rlabel metal3 s 49200 14968 50000 15088 6 wbs_adr_i[31]
port 228 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 wbs_adr_i[3]
port 229 nsew signal input
rlabel metal2 s 47674 51200 47730 52000 6 wbs_adr_i[4]
port 230 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 wbs_adr_i[5]
port 231 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 wbs_adr_i[6]
port 232 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 wbs_adr_i[7]
port 233 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 wbs_adr_i[8]
port 234 nsew signal input
rlabel metal3 s 49200 8848 50000 8968 6 wbs_adr_i[9]
port 235 nsew signal input
rlabel metal2 s 25778 51200 25834 52000 6 wbs_cyc_i
port 236 nsew signal input
rlabel metal3 s 49200 38088 50000 38208 6 wbs_dat_i[0]
port 237 nsew signal input
rlabel metal2 s 662 51200 718 52000 6 wbs_dat_i[10]
port 238 nsew signal input
rlabel metal2 s 3238 51200 3294 52000 6 wbs_dat_i[11]
port 239 nsew signal input
rlabel metal2 s 1950 51200 2006 52000 6 wbs_dat_i[12]
port 240 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wbs_dat_i[13]
port 241 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 wbs_dat_i[14]
port 242 nsew signal input
rlabel metal3 s 49200 21768 50000 21888 6 wbs_dat_i[15]
port 243 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 wbs_dat_i[16]
port 244 nsew signal input
rlabel metal2 s 41878 51200 41934 52000 6 wbs_dat_i[17]
port 245 nsew signal input
rlabel metal3 s 49200 48968 50000 49088 6 wbs_dat_i[18]
port 246 nsew signal input
rlabel metal2 s 11610 51200 11666 52000 6 wbs_dat_i[19]
port 247 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_dat_i[1]
port 248 nsew signal input
rlabel metal3 s 49200 25848 50000 25968 6 wbs_dat_i[20]
port 249 nsew signal input
rlabel metal3 s 49200 48288 50000 48408 6 wbs_dat_i[21]
port 250 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 wbs_dat_i[22]
port 251 nsew signal input
rlabel metal3 s 49200 36048 50000 36168 6 wbs_dat_i[23]
port 252 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 wbs_dat_i[24]
port 253 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 wbs_dat_i[25]
port 254 nsew signal input
rlabel metal2 s 47030 51200 47086 52000 6 wbs_dat_i[26]
port 255 nsew signal input
rlabel metal2 s 18694 51200 18750 52000 6 wbs_dat_i[27]
port 256 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_i[28]
port 257 nsew signal input
rlabel metal3 s 49200 27208 50000 27328 6 wbs_dat_i[29]
port 258 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 wbs_dat_i[2]
port 259 nsew signal input
rlabel metal3 s 49200 11568 50000 11688 6 wbs_dat_i[30]
port 260 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 wbs_dat_i[31]
port 261 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 wbs_dat_i[3]
port 262 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_dat_i[4]
port 263 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 wbs_dat_i[5]
port 264 nsew signal input
rlabel metal3 s 49200 19048 50000 19168 6 wbs_dat_i[6]
port 265 nsew signal input
rlabel metal2 s 43810 51200 43866 52000 6 wbs_dat_i[7]
port 266 nsew signal input
rlabel metal3 s 49200 42848 50000 42968 6 wbs_dat_i[8]
port 267 nsew signal input
rlabel metal3 s 49200 8 50000 128 6 wbs_dat_i[9]
port 268 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_o[0]
port 269 nsew signal tristate
rlabel metal3 s 49200 26528 50000 26648 6 wbs_dat_o[10]
port 270 nsew signal tristate
rlabel metal2 s 662 0 718 800 6 wbs_dat_o[11]
port 271 nsew signal tristate
rlabel metal3 s 49200 44888 50000 45008 6 wbs_dat_o[12]
port 272 nsew signal tristate
rlabel metal2 s 41234 51200 41290 52000 6 wbs_dat_o[13]
port 273 nsew signal tristate
rlabel metal3 s 49200 4088 50000 4208 6 wbs_dat_o[14]
port 274 nsew signal tristate
rlabel metal2 s 39302 51200 39358 52000 6 wbs_dat_o[15]
port 275 nsew signal tristate
rlabel metal3 s 0 19728 800 19848 6 wbs_dat_o[16]
port 276 nsew signal tristate
rlabel metal3 s 0 21768 800 21888 6 wbs_dat_o[17]
port 277 nsew signal tristate
rlabel metal2 s 32218 0 32274 800 6 wbs_dat_o[18]
port 278 nsew signal tristate
rlabel metal2 s 18 0 74 800 6 wbs_dat_o[19]
port 279 nsew signal tristate
rlabel metal2 s 38014 0 38070 800 6 wbs_dat_o[1]
port 280 nsew signal tristate
rlabel metal3 s 0 29248 800 29368 6 wbs_dat_o[20]
port 281 nsew signal tristate
rlabel metal3 s 0 4088 800 4208 6 wbs_dat_o[21]
port 282 nsew signal tristate
rlabel metal3 s 0 12928 800 13048 6 wbs_dat_o[22]
port 283 nsew signal tristate
rlabel metal3 s 0 21088 800 21208 6 wbs_dat_o[23]
port 284 nsew signal tristate
rlabel metal2 s 10322 0 10378 800 6 wbs_dat_o[24]
port 285 nsew signal tristate
rlabel metal2 s 3238 0 3294 800 6 wbs_dat_o[25]
port 286 nsew signal tristate
rlabel metal2 s 27710 51200 27766 52000 6 wbs_dat_o[26]
port 287 nsew signal tristate
rlabel metal2 s 16762 51200 16818 52000 6 wbs_dat_o[27]
port 288 nsew signal tristate
rlabel metal2 s 26422 0 26478 800 6 wbs_dat_o[28]
port 289 nsew signal tristate
rlabel metal2 s 36726 51200 36782 52000 6 wbs_dat_o[29]
port 290 nsew signal tristate
rlabel metal3 s 49200 12928 50000 13048 6 wbs_dat_o[2]
port 291 nsew signal tristate
rlabel metal3 s 0 36048 800 36168 6 wbs_dat_o[30]
port 292 nsew signal tristate
rlabel metal3 s 49200 39448 50000 39568 6 wbs_dat_o[31]
port 293 nsew signal tristate
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_o[3]
port 294 nsew signal tristate
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_o[4]
port 295 nsew signal tristate
rlabel metal3 s 0 6128 800 6248 6 wbs_dat_o[5]
port 296 nsew signal tristate
rlabel metal3 s 49200 37408 50000 37528 6 wbs_dat_o[6]
port 297 nsew signal tristate
rlabel metal2 s 29642 0 29698 800 6 wbs_dat_o[7]
port 298 nsew signal tristate
rlabel metal2 s 34150 51200 34206 52000 6 wbs_dat_o[8]
port 299 nsew signal tristate
rlabel metal2 s 33506 51200 33562 52000 6 wbs_dat_o[9]
port 300 nsew signal tristate
rlabel metal3 s 0 49648 800 49768 6 wbs_sel_i[0]
port 301 nsew signal input
rlabel metal2 s 5814 51200 5870 52000 6 wbs_sel_i[1]
port 302 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 wbs_sel_i[2]
port 303 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 wbs_sel_i[3]
port 304 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 wbs_stb_i
port 305 nsew signal input
rlabel metal3 s 49200 25168 50000 25288 6 wbs_we_i
port 306 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 50000 52000
<< end >>
