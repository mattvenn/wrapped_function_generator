magic
tech sky130A
magscale 1 2
timestamp 1651661546
<< obsli1 >>
rect 1104 2159 48852 49521
<< obsm1 >>
rect 14 1844 49666 50244
<< metal2 >>
rect 18 51200 74 52000
rect 662 51200 718 52000
rect 1306 51200 1362 52000
rect 1950 51200 2006 52000
rect 2594 51200 2650 52000
rect 3238 51200 3294 52000
rect 3882 51200 3938 52000
rect 4526 51200 4582 52000
rect 5170 51200 5226 52000
rect 5814 51200 5870 52000
rect 6458 51200 6514 52000
rect 7102 51200 7158 52000
rect 7746 51200 7802 52000
rect 8390 51200 8446 52000
rect 9034 51200 9090 52000
rect 9678 51200 9734 52000
rect 10322 51200 10378 52000
rect 10966 51200 11022 52000
rect 11610 51200 11666 52000
rect 12254 51200 12310 52000
rect 12898 51200 12954 52000
rect 13542 51200 13598 52000
rect 14186 51200 14242 52000
rect 14830 51200 14886 52000
rect 15474 51200 15530 52000
rect 16118 51200 16174 52000
rect 16762 51200 16818 52000
rect 17406 51200 17462 52000
rect 18050 51200 18106 52000
rect 18694 51200 18750 52000
rect 19338 51200 19394 52000
rect 19982 51200 20038 52000
rect 20626 51200 20682 52000
rect 21270 51200 21326 52000
rect 21914 51200 21970 52000
rect 22558 51200 22614 52000
rect 23202 51200 23258 52000
rect 23846 51200 23902 52000
rect 24490 51200 24546 52000
rect 25134 51200 25190 52000
rect 25778 51200 25834 52000
rect 26422 51200 26478 52000
rect 27066 51200 27122 52000
rect 27710 51200 27766 52000
rect 28354 51200 28410 52000
rect 28998 51200 29054 52000
rect 29642 51200 29698 52000
rect 30930 51200 30986 52000
rect 31574 51200 31630 52000
rect 32218 51200 32274 52000
rect 32862 51200 32918 52000
rect 33506 51200 33562 52000
rect 34150 51200 34206 52000
rect 34794 51200 34850 52000
rect 35438 51200 35494 52000
rect 36082 51200 36138 52000
rect 36726 51200 36782 52000
rect 37370 51200 37426 52000
rect 38014 51200 38070 52000
rect 38658 51200 38714 52000
rect 39302 51200 39358 52000
rect 39946 51200 40002 52000
rect 40590 51200 40646 52000
rect 41234 51200 41290 52000
rect 41878 51200 41934 52000
rect 42522 51200 42578 52000
rect 43166 51200 43222 52000
rect 43810 51200 43866 52000
rect 44454 51200 44510 52000
rect 45098 51200 45154 52000
rect 45742 51200 45798 52000
rect 46386 51200 46442 52000
rect 47030 51200 47086 52000
rect 47674 51200 47730 52000
rect 48318 51200 48374 52000
rect 48962 51200 49018 52000
rect 49606 51200 49662 52000
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 1950 0 2006 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 23846 0 23902 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 25778 0 25834 800
rect 26422 0 26478 800
rect 27066 0 27122 800
rect 27710 0 27766 800
rect 28354 0 28410 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30286 0 30342 800
rect 30930 0 30986 800
rect 31574 0 31630 800
rect 32218 0 32274 800
rect 32862 0 32918 800
rect 33506 0 33562 800
rect 34150 0 34206 800
rect 34794 0 34850 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 36726 0 36782 800
rect 37370 0 37426 800
rect 38014 0 38070 800
rect 38658 0 38714 800
rect 39946 0 40002 800
rect 40590 0 40646 800
rect 41234 0 41290 800
rect 41878 0 41934 800
rect 42522 0 42578 800
rect 43166 0 43222 800
rect 43810 0 43866 800
rect 44454 0 44510 800
rect 45098 0 45154 800
rect 45742 0 45798 800
rect 46386 0 46442 800
rect 47030 0 47086 800
rect 47674 0 47730 800
rect 48318 0 48374 800
rect 48962 0 49018 800
rect 49606 0 49662 800
<< obsm2 >>
rect 130 51144 606 51785
rect 774 51144 1250 51785
rect 1418 51144 1894 51785
rect 2062 51144 2538 51785
rect 2706 51144 3182 51785
rect 3350 51144 3826 51785
rect 3994 51144 4470 51785
rect 4638 51144 5114 51785
rect 5282 51144 5758 51785
rect 5926 51144 6402 51785
rect 6570 51144 7046 51785
rect 7214 51144 7690 51785
rect 7858 51144 8334 51785
rect 8502 51144 8978 51785
rect 9146 51144 9622 51785
rect 9790 51144 10266 51785
rect 10434 51144 10910 51785
rect 11078 51144 11554 51785
rect 11722 51144 12198 51785
rect 12366 51144 12842 51785
rect 13010 51144 13486 51785
rect 13654 51144 14130 51785
rect 14298 51144 14774 51785
rect 14942 51144 15418 51785
rect 15586 51144 16062 51785
rect 16230 51144 16706 51785
rect 16874 51144 17350 51785
rect 17518 51144 17994 51785
rect 18162 51144 18638 51785
rect 18806 51144 19282 51785
rect 19450 51144 19926 51785
rect 20094 51144 20570 51785
rect 20738 51144 21214 51785
rect 21382 51144 21858 51785
rect 22026 51144 22502 51785
rect 22670 51144 23146 51785
rect 23314 51144 23790 51785
rect 23958 51144 24434 51785
rect 24602 51144 25078 51785
rect 25246 51144 25722 51785
rect 25890 51144 26366 51785
rect 26534 51144 27010 51785
rect 27178 51144 27654 51785
rect 27822 51144 28298 51785
rect 28466 51144 28942 51785
rect 29110 51144 29586 51785
rect 29754 51144 30874 51785
rect 31042 51144 31518 51785
rect 31686 51144 32162 51785
rect 32330 51144 32806 51785
rect 32974 51144 33450 51785
rect 33618 51144 34094 51785
rect 34262 51144 34738 51785
rect 34906 51144 35382 51785
rect 35550 51144 36026 51785
rect 36194 51144 36670 51785
rect 36838 51144 37314 51785
rect 37482 51144 37958 51785
rect 38126 51144 38602 51785
rect 38770 51144 39246 51785
rect 39414 51144 39890 51785
rect 40058 51144 40534 51785
rect 40702 51144 41178 51785
rect 41346 51144 41822 51785
rect 41990 51144 42466 51785
rect 42634 51144 43110 51785
rect 43278 51144 43754 51785
rect 43922 51144 44398 51785
rect 44566 51144 45042 51785
rect 45210 51144 45686 51785
rect 45854 51144 46330 51785
rect 46498 51144 46974 51785
rect 47142 51144 47618 51785
rect 47786 51144 48262 51785
rect 48430 51144 48906 51785
rect 49074 51144 49550 51785
rect 20 856 49660 51144
rect 130 31 606 856
rect 774 31 1250 856
rect 1418 31 1894 856
rect 2062 31 2538 856
rect 2706 31 3182 856
rect 3350 31 3826 856
rect 3994 31 4470 856
rect 4638 31 5114 856
rect 5282 31 5758 856
rect 5926 31 6402 856
rect 6570 31 7046 856
rect 7214 31 7690 856
rect 7858 31 8334 856
rect 8502 31 8978 856
rect 9146 31 9622 856
rect 9790 31 10266 856
rect 10434 31 10910 856
rect 11078 31 11554 856
rect 11722 31 12198 856
rect 12366 31 12842 856
rect 13010 31 13486 856
rect 13654 31 14130 856
rect 14298 31 14774 856
rect 14942 31 15418 856
rect 15586 31 16062 856
rect 16230 31 16706 856
rect 16874 31 17350 856
rect 17518 31 17994 856
rect 18162 31 18638 856
rect 18806 31 19282 856
rect 19450 31 19926 856
rect 20094 31 20570 856
rect 20738 31 21214 856
rect 21382 31 21858 856
rect 22026 31 22502 856
rect 22670 31 23146 856
rect 23314 31 23790 856
rect 23958 31 24434 856
rect 24602 31 25078 856
rect 25246 31 25722 856
rect 25890 31 26366 856
rect 26534 31 27010 856
rect 27178 31 27654 856
rect 27822 31 28298 856
rect 28466 31 28942 856
rect 29110 31 29586 856
rect 29754 31 30230 856
rect 30398 31 30874 856
rect 31042 31 31518 856
rect 31686 31 32162 856
rect 32330 31 32806 856
rect 32974 31 33450 856
rect 33618 31 34094 856
rect 34262 31 34738 856
rect 34906 31 35382 856
rect 35550 31 36026 856
rect 36194 31 36670 856
rect 36838 31 37314 856
rect 37482 31 37958 856
rect 38126 31 38602 856
rect 38770 31 39890 856
rect 40058 31 40534 856
rect 40702 31 41178 856
rect 41346 31 41822 856
rect 41990 31 42466 856
rect 42634 31 43110 856
rect 43278 31 43754 856
rect 43922 31 44398 856
rect 44566 31 45042 856
rect 45210 31 45686 856
rect 45854 31 46330 856
rect 46498 31 46974 856
rect 47142 31 47618 856
rect 47786 31 48262 856
rect 48430 31 48906 856
rect 49074 31 49550 856
<< metal3 >>
rect 0 51688 800 51808
rect 49200 51688 50000 51808
rect 0 51008 800 51128
rect 49200 51008 50000 51128
rect 0 50328 800 50448
rect 49200 50328 50000 50448
rect 0 49648 800 49768
rect 49200 49648 50000 49768
rect 0 48968 800 49088
rect 49200 48968 50000 49088
rect 0 48288 800 48408
rect 49200 48288 50000 48408
rect 0 47608 800 47728
rect 49200 47608 50000 47728
rect 0 46928 800 47048
rect 49200 46928 50000 47048
rect 0 46248 800 46368
rect 49200 46248 50000 46368
rect 0 45568 800 45688
rect 49200 45568 50000 45688
rect 0 44888 800 45008
rect 49200 44888 50000 45008
rect 0 44208 800 44328
rect 49200 44208 50000 44328
rect 0 43528 800 43648
rect 49200 43528 50000 43648
rect 0 42848 800 42968
rect 49200 42848 50000 42968
rect 49200 42168 50000 42288
rect 0 41488 800 41608
rect 49200 41488 50000 41608
rect 0 40808 800 40928
rect 49200 40808 50000 40928
rect 0 40128 800 40248
rect 49200 40128 50000 40248
rect 0 39448 800 39568
rect 49200 39448 50000 39568
rect 0 38768 800 38888
rect 49200 38768 50000 38888
rect 0 38088 800 38208
rect 49200 38088 50000 38208
rect 0 37408 800 37528
rect 49200 37408 50000 37528
rect 0 36728 800 36848
rect 49200 36728 50000 36848
rect 0 36048 800 36168
rect 49200 36048 50000 36168
rect 0 35368 800 35488
rect 49200 35368 50000 35488
rect 0 34688 800 34808
rect 49200 34688 50000 34808
rect 0 34008 800 34128
rect 49200 34008 50000 34128
rect 0 33328 800 33448
rect 49200 33328 50000 33448
rect 0 32648 800 32768
rect 49200 32648 50000 32768
rect 0 31968 800 32088
rect 49200 31968 50000 32088
rect 0 31288 800 31408
rect 49200 31288 50000 31408
rect 0 30608 800 30728
rect 0 29928 800 30048
rect 49200 29928 50000 30048
rect 0 29248 800 29368
rect 49200 29248 50000 29368
rect 0 28568 800 28688
rect 49200 28568 50000 28688
rect 0 27888 800 28008
rect 49200 27888 50000 28008
rect 0 27208 800 27328
rect 49200 27208 50000 27328
rect 0 26528 800 26648
rect 49200 26528 50000 26648
rect 0 25848 800 25968
rect 49200 25848 50000 25968
rect 0 25168 800 25288
rect 49200 25168 50000 25288
rect 0 24488 800 24608
rect 49200 24488 50000 24608
rect 0 23808 800 23928
rect 49200 23808 50000 23928
rect 0 23128 800 23248
rect 49200 23128 50000 23248
rect 0 22448 800 22568
rect 49200 22448 50000 22568
rect 0 21768 800 21888
rect 49200 21768 50000 21888
rect 0 21088 800 21208
rect 49200 21088 50000 21208
rect 0 20408 800 20528
rect 49200 20408 50000 20528
rect 0 19728 800 19848
rect 49200 19728 50000 19848
rect 0 19048 800 19168
rect 49200 19048 50000 19168
rect 0 18368 800 18488
rect 49200 18368 50000 18488
rect 0 17688 800 17808
rect 49200 17688 50000 17808
rect 0 17008 800 17128
rect 49200 17008 50000 17128
rect 0 16328 800 16448
rect 49200 16328 50000 16448
rect 0 15648 800 15768
rect 49200 15648 50000 15768
rect 0 14968 800 15088
rect 49200 14968 50000 15088
rect 0 14288 800 14408
rect 49200 14288 50000 14408
rect 0 13608 800 13728
rect 49200 13608 50000 13728
rect 0 12928 800 13048
rect 49200 12928 50000 13048
rect 0 12248 800 12368
rect 49200 12248 50000 12368
rect 0 11568 800 11688
rect 49200 11568 50000 11688
rect 0 10888 800 11008
rect 49200 10888 50000 11008
rect 0 10208 800 10328
rect 49200 10208 50000 10328
rect 0 9528 800 9648
rect 49200 9528 50000 9648
rect 0 8848 800 8968
rect 49200 8848 50000 8968
rect 0 8168 800 8288
rect 49200 8168 50000 8288
rect 0 7488 800 7608
rect 49200 7488 50000 7608
rect 0 6808 800 6928
rect 49200 6808 50000 6928
rect 0 6128 800 6248
rect 49200 6128 50000 6248
rect 0 5448 800 5568
rect 49200 5448 50000 5568
rect 0 4768 800 4888
rect 49200 4768 50000 4888
rect 0 4088 800 4208
rect 49200 4088 50000 4208
rect 0 3408 800 3528
rect 49200 3408 50000 3528
rect 0 2728 800 2848
rect 49200 2728 50000 2848
rect 0 2048 800 2168
rect 49200 2048 50000 2168
rect 0 1368 800 1488
rect 49200 1368 50000 1488
rect 0 688 800 808
rect 49200 688 50000 808
rect 49200 8 50000 128
<< obsm3 >>
rect 880 51608 49120 51781
rect 800 51208 49200 51608
rect 880 50928 49120 51208
rect 800 50528 49200 50928
rect 880 50248 49120 50528
rect 800 49848 49200 50248
rect 880 49568 49120 49848
rect 800 49168 49200 49568
rect 880 48888 49120 49168
rect 800 48488 49200 48888
rect 880 48208 49120 48488
rect 800 47808 49200 48208
rect 880 47528 49120 47808
rect 800 47128 49200 47528
rect 880 46848 49120 47128
rect 800 46448 49200 46848
rect 880 46168 49120 46448
rect 800 45768 49200 46168
rect 880 45488 49120 45768
rect 800 45088 49200 45488
rect 880 44808 49120 45088
rect 800 44408 49200 44808
rect 880 44128 49120 44408
rect 800 43728 49200 44128
rect 880 43448 49120 43728
rect 800 43048 49200 43448
rect 880 42768 49120 43048
rect 800 42368 49200 42768
rect 800 42088 49120 42368
rect 800 41688 49200 42088
rect 880 41408 49120 41688
rect 800 41008 49200 41408
rect 880 40728 49120 41008
rect 800 40328 49200 40728
rect 880 40048 49120 40328
rect 800 39648 49200 40048
rect 880 39368 49120 39648
rect 800 38968 49200 39368
rect 880 38688 49120 38968
rect 800 38288 49200 38688
rect 880 38008 49120 38288
rect 800 37608 49200 38008
rect 880 37328 49120 37608
rect 800 36928 49200 37328
rect 880 36648 49120 36928
rect 800 36248 49200 36648
rect 880 35968 49120 36248
rect 800 35568 49200 35968
rect 880 35288 49120 35568
rect 800 34888 49200 35288
rect 880 34608 49120 34888
rect 800 34208 49200 34608
rect 880 33928 49120 34208
rect 800 33528 49200 33928
rect 880 33248 49120 33528
rect 800 32848 49200 33248
rect 880 32568 49120 32848
rect 800 32168 49200 32568
rect 880 31888 49120 32168
rect 800 31488 49200 31888
rect 880 31208 49120 31488
rect 800 30808 49200 31208
rect 880 30528 49200 30808
rect 800 30128 49200 30528
rect 880 29848 49120 30128
rect 800 29448 49200 29848
rect 880 29168 49120 29448
rect 800 28768 49200 29168
rect 880 28488 49120 28768
rect 800 28088 49200 28488
rect 880 27808 49120 28088
rect 800 27408 49200 27808
rect 880 27128 49120 27408
rect 800 26728 49200 27128
rect 880 26448 49120 26728
rect 800 26048 49200 26448
rect 880 25768 49120 26048
rect 800 25368 49200 25768
rect 880 25088 49120 25368
rect 800 24688 49200 25088
rect 880 24408 49120 24688
rect 800 24008 49200 24408
rect 880 23728 49120 24008
rect 800 23328 49200 23728
rect 880 23048 49120 23328
rect 800 22648 49200 23048
rect 880 22368 49120 22648
rect 800 21968 49200 22368
rect 880 21688 49120 21968
rect 800 21288 49200 21688
rect 880 21008 49120 21288
rect 800 20608 49200 21008
rect 880 20328 49120 20608
rect 800 19928 49200 20328
rect 880 19648 49120 19928
rect 800 19248 49200 19648
rect 880 18968 49120 19248
rect 800 18568 49200 18968
rect 880 18288 49120 18568
rect 800 17888 49200 18288
rect 880 17608 49120 17888
rect 800 17208 49200 17608
rect 880 16928 49120 17208
rect 800 16528 49200 16928
rect 880 16248 49120 16528
rect 800 15848 49200 16248
rect 880 15568 49120 15848
rect 800 15168 49200 15568
rect 880 14888 49120 15168
rect 800 14488 49200 14888
rect 880 14208 49120 14488
rect 800 13808 49200 14208
rect 880 13528 49120 13808
rect 800 13128 49200 13528
rect 880 12848 49120 13128
rect 800 12448 49200 12848
rect 880 12168 49120 12448
rect 800 11768 49200 12168
rect 880 11488 49120 11768
rect 800 11088 49200 11488
rect 880 10808 49120 11088
rect 800 10408 49200 10808
rect 880 10128 49120 10408
rect 800 9728 49200 10128
rect 880 9448 49120 9728
rect 800 9048 49200 9448
rect 880 8768 49120 9048
rect 800 8368 49200 8768
rect 880 8088 49120 8368
rect 800 7688 49200 8088
rect 880 7408 49120 7688
rect 800 7008 49200 7408
rect 880 6728 49120 7008
rect 800 6328 49200 6728
rect 880 6048 49120 6328
rect 800 5648 49200 6048
rect 880 5368 49120 5648
rect 800 4968 49200 5368
rect 880 4688 49120 4968
rect 800 4288 49200 4688
rect 880 4008 49120 4288
rect 800 3608 49200 4008
rect 880 3328 49120 3608
rect 800 2928 49200 3328
rect 880 2648 49120 2928
rect 800 2248 49200 2648
rect 880 1968 49120 2248
rect 800 1568 49200 1968
rect 880 1288 49120 1568
rect 800 888 49200 1288
rect 880 608 49120 888
rect 800 208 49200 608
rect 800 35 49120 208
<< metal4 >>
rect 4208 2128 4528 49552
rect 19568 2128 19888 49552
rect 34928 2128 35248 49552
<< obsm4 >>
rect 20115 2347 32693 21997
<< labels >>
rlabel metal3 s 49200 31968 50000 32088 6 active
port 1 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 io_in[0]
port 2 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 io_in[10]
port 3 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 io_in[11]
port 4 nsew signal input
rlabel metal2 s 25134 51200 25190 52000 6 io_in[12]
port 5 nsew signal input
rlabel metal3 s 49200 15648 50000 15768 6 io_in[13]
port 6 nsew signal input
rlabel metal2 s 21270 51200 21326 52000 6 io_in[14]
port 7 nsew signal input
rlabel metal3 s 49200 2048 50000 2168 6 io_in[15]
port 8 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 io_in[16]
port 9 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 io_in[17]
port 10 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 io_in[18]
port 11 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 io_in[19]
port 12 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 io_in[1]
port 13 nsew signal input
rlabel metal3 s 49200 18368 50000 18488 6 io_in[20]
port 14 nsew signal input
rlabel metal3 s 0 30608 800 30728 6 io_in[21]
port 15 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 io_in[22]
port 16 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 io_in[23]
port 17 nsew signal input
rlabel metal3 s 49200 21088 50000 21208 6 io_in[24]
port 18 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 io_in[25]
port 19 nsew signal input
rlabel metal3 s 49200 32648 50000 32768 6 io_in[26]
port 20 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 io_in[27]
port 21 nsew signal input
rlabel metal3 s 49200 23128 50000 23248 6 io_in[28]
port 22 nsew signal input
rlabel metal2 s 2594 51200 2650 52000 6 io_in[29]
port 23 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 io_in[2]
port 24 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 io_in[30]
port 25 nsew signal input
rlabel metal2 s 46386 51200 46442 52000 6 io_in[31]
port 26 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 io_in[32]
port 27 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 io_in[33]
port 28 nsew signal input
rlabel metal2 s 9034 51200 9090 52000 6 io_in[34]
port 29 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 io_in[35]
port 30 nsew signal input
rlabel metal2 s 31574 51200 31630 52000 6 io_in[36]
port 31 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 io_in[37]
port 32 nsew signal input
rlabel metal3 s 49200 47608 50000 47728 6 io_in[3]
port 33 nsew signal input
rlabel metal3 s 49200 20408 50000 20528 6 io_in[4]
port 34 nsew signal input
rlabel metal2 s 35438 51200 35494 52000 6 io_in[5]
port 35 nsew signal input
rlabel metal3 s 49200 2728 50000 2848 6 io_in[6]
port 36 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 io_in[7]
port 37 nsew signal input
rlabel metal2 s 3882 51200 3938 52000 6 io_in[8]
port 38 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 io_in[9]
port 39 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 io_oeb[0]
port 40 nsew signal bidirectional
rlabel metal3 s 49200 24488 50000 24608 6 io_oeb[10]
port 41 nsew signal bidirectional
rlabel metal2 s 45098 0 45154 800 6 io_oeb[11]
port 42 nsew signal bidirectional
rlabel metal2 s 5814 0 5870 800 6 io_oeb[12]
port 43 nsew signal bidirectional
rlabel metal2 s 48318 0 48374 800 6 io_oeb[13]
port 44 nsew signal bidirectional
rlabel metal2 s 7746 51200 7802 52000 6 io_oeb[14]
port 45 nsew signal bidirectional
rlabel metal3 s 49200 43528 50000 43648 6 io_oeb[15]
port 46 nsew signal bidirectional
rlabel metal3 s 49200 4768 50000 4888 6 io_oeb[16]
port 47 nsew signal bidirectional
rlabel metal3 s 0 6808 800 6928 6 io_oeb[17]
port 48 nsew signal bidirectional
rlabel metal3 s 0 41488 800 41608 6 io_oeb[18]
port 49 nsew signal bidirectional
rlabel metal2 s 36726 0 36782 800 6 io_oeb[19]
port 50 nsew signal bidirectional
rlabel metal2 s 43166 51200 43222 52000 6 io_oeb[1]
port 51 nsew signal bidirectional
rlabel metal3 s 49200 46928 50000 47048 6 io_oeb[20]
port 52 nsew signal bidirectional
rlabel metal3 s 0 9528 800 9648 6 io_oeb[21]
port 53 nsew signal bidirectional
rlabel metal2 s 45098 51200 45154 52000 6 io_oeb[22]
port 54 nsew signal bidirectional
rlabel metal3 s 0 26528 800 26648 6 io_oeb[23]
port 55 nsew signal bidirectional
rlabel metal3 s 49200 51688 50000 51808 6 io_oeb[24]
port 56 nsew signal bidirectional
rlabel metal2 s 24490 51200 24546 52000 6 io_oeb[25]
port 57 nsew signal bidirectional
rlabel metal3 s 0 23128 800 23248 6 io_oeb[26]
port 58 nsew signal bidirectional
rlabel metal3 s 49200 28568 50000 28688 6 io_oeb[27]
port 59 nsew signal bidirectional
rlabel metal2 s 1306 51200 1362 52000 6 io_oeb[28]
port 60 nsew signal bidirectional
rlabel metal2 s 12254 0 12310 800 6 io_oeb[29]
port 61 nsew signal bidirectional
rlabel metal3 s 0 51688 800 51808 6 io_oeb[2]
port 62 nsew signal bidirectional
rlabel metal2 s 49606 51200 49662 52000 6 io_oeb[30]
port 63 nsew signal bidirectional
rlabel metal3 s 0 3408 800 3528 6 io_oeb[31]
port 64 nsew signal bidirectional
rlabel metal2 s 33506 0 33562 800 6 io_oeb[32]
port 65 nsew signal bidirectional
rlabel metal2 s 22558 51200 22614 52000 6 io_oeb[33]
port 66 nsew signal bidirectional
rlabel metal3 s 0 17688 800 17808 6 io_oeb[34]
port 67 nsew signal bidirectional
rlabel metal3 s 0 13608 800 13728 6 io_oeb[35]
port 68 nsew signal bidirectional
rlabel metal2 s 39946 0 40002 800 6 io_oeb[36]
port 69 nsew signal bidirectional
rlabel metal3 s 0 39448 800 39568 6 io_oeb[37]
port 70 nsew signal bidirectional
rlabel metal3 s 49200 45568 50000 45688 6 io_oeb[3]
port 71 nsew signal bidirectional
rlabel metal3 s 0 44888 800 45008 6 io_oeb[4]
port 72 nsew signal bidirectional
rlabel metal3 s 49200 36728 50000 36848 6 io_oeb[5]
port 73 nsew signal bidirectional
rlabel metal2 s 21270 0 21326 800 6 io_oeb[6]
port 74 nsew signal bidirectional
rlabel metal3 s 49200 17008 50000 17128 6 io_oeb[7]
port 75 nsew signal bidirectional
rlabel metal3 s 49200 49648 50000 49768 6 io_oeb[8]
port 76 nsew signal bidirectional
rlabel metal3 s 49200 16328 50000 16448 6 io_oeb[9]
port 77 nsew signal bidirectional
rlabel metal2 s 36082 51200 36138 52000 6 io_out[0]
port 78 nsew signal bidirectional
rlabel metal3 s 49200 44208 50000 44328 6 io_out[10]
port 79 nsew signal bidirectional
rlabel metal3 s 49200 9528 50000 9648 6 io_out[11]
port 80 nsew signal bidirectional
rlabel metal2 s 48962 0 49018 800 6 io_out[12]
port 81 nsew signal bidirectional
rlabel metal2 s 47030 0 47086 800 6 io_out[13]
port 82 nsew signal bidirectional
rlabel metal3 s 49200 12248 50000 12368 6 io_out[14]
port 83 nsew signal bidirectional
rlabel metal2 s 37370 0 37426 800 6 io_out[15]
port 84 nsew signal bidirectional
rlabel metal2 s 37370 51200 37426 52000 6 io_out[16]
port 85 nsew signal bidirectional
rlabel metal2 s 38658 51200 38714 52000 6 io_out[17]
port 86 nsew signal bidirectional
rlabel metal2 s 15474 51200 15530 52000 6 io_out[18]
port 87 nsew signal bidirectional
rlabel metal3 s 49200 3408 50000 3528 6 io_out[19]
port 88 nsew signal bidirectional
rlabel metal2 s 12898 0 12954 800 6 io_out[1]
port 89 nsew signal bidirectional
rlabel metal2 s 11610 0 11666 800 6 io_out[20]
port 90 nsew signal bidirectional
rlabel metal3 s 0 48288 800 48408 6 io_out[21]
port 91 nsew signal bidirectional
rlabel metal2 s 34794 51200 34850 52000 6 io_out[22]
port 92 nsew signal bidirectional
rlabel metal2 s 14830 51200 14886 52000 6 io_out[23]
port 93 nsew signal bidirectional
rlabel metal3 s 0 46248 800 46368 6 io_out[24]
port 94 nsew signal bidirectional
rlabel metal3 s 0 34008 800 34128 6 io_out[25]
port 95 nsew signal bidirectional
rlabel metal3 s 0 27208 800 27328 6 io_out[26]
port 96 nsew signal bidirectional
rlabel metal3 s 49200 7488 50000 7608 6 io_out[27]
port 97 nsew signal bidirectional
rlabel metal2 s 44454 0 44510 800 6 io_out[28]
port 98 nsew signal bidirectional
rlabel metal3 s 0 5448 800 5568 6 io_out[29]
port 99 nsew signal bidirectional
rlabel metal3 s 49200 35368 50000 35488 6 io_out[2]
port 100 nsew signal bidirectional
rlabel metal2 s 28354 51200 28410 52000 6 io_out[30]
port 101 nsew signal bidirectional
rlabel metal3 s 49200 46248 50000 46368 6 io_out[31]
port 102 nsew signal bidirectional
rlabel metal2 s 42522 0 42578 800 6 io_out[32]
port 103 nsew signal bidirectional
rlabel metal3 s 49200 10888 50000 11008 6 io_out[33]
port 104 nsew signal bidirectional
rlabel metal3 s 0 51008 800 51128 6 io_out[34]
port 105 nsew signal bidirectional
rlabel metal2 s 13542 0 13598 800 6 io_out[35]
port 106 nsew signal bidirectional
rlabel metal2 s 27066 51200 27122 52000 6 io_out[36]
port 107 nsew signal bidirectional
rlabel metal2 s 48318 51200 48374 52000 6 io_out[37]
port 108 nsew signal bidirectional
rlabel metal2 s 45742 51200 45798 52000 6 io_out[3]
port 109 nsew signal bidirectional
rlabel metal2 s 39946 51200 40002 52000 6 io_out[4]
port 110 nsew signal bidirectional
rlabel metal2 s 10322 51200 10378 52000 6 io_out[5]
port 111 nsew signal bidirectional
rlabel metal2 s 7102 51200 7158 52000 6 io_out[6]
port 112 nsew signal bidirectional
rlabel metal3 s 49200 34008 50000 34128 6 io_out[7]
port 113 nsew signal bidirectional
rlabel metal2 s 2594 0 2650 800 6 io_out[8]
port 114 nsew signal bidirectional
rlabel metal2 s 8390 51200 8446 52000 6 io_out[9]
port 115 nsew signal bidirectional
rlabel metal3 s 0 8168 800 8288 6 rambus_wb_ack_i
port 116 nsew signal input
rlabel metal3 s 49200 40128 50000 40248 6 rambus_wb_adr_o[0]
port 117 nsew signal bidirectional
rlabel metal3 s 0 46928 800 47048 6 rambus_wb_adr_o[1]
port 118 nsew signal bidirectional
rlabel metal2 s 10966 51200 11022 52000 6 rambus_wb_adr_o[2]
port 119 nsew signal bidirectional
rlabel metal3 s 49200 6128 50000 6248 6 rambus_wb_adr_o[3]
port 120 nsew signal bidirectional
rlabel metal3 s 49200 51008 50000 51128 6 rambus_wb_adr_o[4]
port 121 nsew signal bidirectional
rlabel metal3 s 49200 17688 50000 17808 6 rambus_wb_adr_o[5]
port 122 nsew signal bidirectional
rlabel metal3 s 49200 6808 50000 6928 6 rambus_wb_adr_o[6]
port 123 nsew signal bidirectional
rlabel metal3 s 49200 29248 50000 29368 6 rambus_wb_adr_o[7]
port 124 nsew signal bidirectional
rlabel metal2 s 9034 0 9090 800 6 rambus_wb_adr_o[8]
port 125 nsew signal bidirectional
rlabel metal3 s 0 2048 800 2168 6 rambus_wb_adr_o[9]
port 126 nsew signal bidirectional
rlabel metal3 s 0 18368 800 18488 6 rambus_wb_clk_o
port 127 nsew signal bidirectional
rlabel metal2 s 5170 51200 5226 52000 6 rambus_wb_cyc_o
port 128 nsew signal bidirectional
rlabel metal2 s 13542 51200 13598 52000 6 rambus_wb_dat_i[0]
port 129 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 rambus_wb_dat_i[10]
port 130 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 rambus_wb_dat_i[11]
port 131 nsew signal input
rlabel metal3 s 49200 688 50000 808 6 rambus_wb_dat_i[12]
port 132 nsew signal input
rlabel metal3 s 49200 13608 50000 13728 6 rambus_wb_dat_i[13]
port 133 nsew signal input
rlabel metal2 s 21914 51200 21970 52000 6 rambus_wb_dat_i[14]
port 134 nsew signal input
rlabel metal2 s 12898 51200 12954 52000 6 rambus_wb_dat_i[15]
port 135 nsew signal input
rlabel metal2 s 18050 51200 18106 52000 6 rambus_wb_dat_i[16]
port 136 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 rambus_wb_dat_i[17]
port 137 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 rambus_wb_dat_i[18]
port 138 nsew signal input
rlabel metal3 s 0 34688 800 34808 6 rambus_wb_dat_i[19]
port 139 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 rambus_wb_dat_i[1]
port 140 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 rambus_wb_dat_i[20]
port 141 nsew signal input
rlabel metal2 s 16118 51200 16174 52000 6 rambus_wb_dat_i[21]
port 142 nsew signal input
rlabel metal3 s 49200 8168 50000 8288 6 rambus_wb_dat_i[22]
port 143 nsew signal input
rlabel metal3 s 49200 31288 50000 31408 6 rambus_wb_dat_i[23]
port 144 nsew signal input
rlabel metal3 s 49200 33328 50000 33448 6 rambus_wb_dat_i[24]
port 145 nsew signal input
rlabel metal3 s 49200 38768 50000 38888 6 rambus_wb_dat_i[25]
port 146 nsew signal input
rlabel metal2 s 23846 51200 23902 52000 6 rambus_wb_dat_i[26]
port 147 nsew signal input
rlabel metal3 s 0 36728 800 36848 6 rambus_wb_dat_i[27]
port 148 nsew signal input
rlabel metal2 s 18 51200 74 52000 6 rambus_wb_dat_i[28]
port 149 nsew signal input
rlabel metal3 s 49200 42168 50000 42288 6 rambus_wb_dat_i[29]
port 150 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 rambus_wb_dat_i[2]
port 151 nsew signal input
rlabel metal3 s 49200 10208 50000 10328 6 rambus_wb_dat_i[30]
port 152 nsew signal input
rlabel metal2 s 14186 51200 14242 52000 6 rambus_wb_dat_i[31]
port 153 nsew signal input
rlabel metal3 s 49200 29928 50000 30048 6 rambus_wb_dat_i[3]
port 154 nsew signal input
rlabel metal3 s 49200 23808 50000 23928 6 rambus_wb_dat_i[4]
port 155 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 rambus_wb_dat_i[5]
port 156 nsew signal input
rlabel metal2 s 4526 51200 4582 52000 6 rambus_wb_dat_i[6]
port 157 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 rambus_wb_dat_i[7]
port 158 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 rambus_wb_dat_i[8]
port 159 nsew signal input
rlabel metal2 s 40590 51200 40646 52000 6 rambus_wb_dat_i[9]
port 160 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 rambus_wb_dat_o[0]
port 161 nsew signal bidirectional
rlabel metal2 s 30286 0 30342 800 6 rambus_wb_dat_o[10]
port 162 nsew signal bidirectional
rlabel metal2 s 20626 0 20682 800 6 rambus_wb_dat_o[11]
port 163 nsew signal bidirectional
rlabel metal2 s 41878 0 41934 800 6 rambus_wb_dat_o[12]
port 164 nsew signal bidirectional
rlabel metal3 s 49200 34688 50000 34808 6 rambus_wb_dat_o[13]
port 165 nsew signal bidirectional
rlabel metal3 s 0 50328 800 50448 6 rambus_wb_dat_o[14]
port 166 nsew signal bidirectional
rlabel metal2 s 42522 51200 42578 52000 6 rambus_wb_dat_o[15]
port 167 nsew signal bidirectional
rlabel metal2 s 1306 0 1362 800 6 rambus_wb_dat_o[16]
port 168 nsew signal bidirectional
rlabel metal3 s 0 29928 800 30048 6 rambus_wb_dat_o[17]
port 169 nsew signal bidirectional
rlabel metal2 s 18050 0 18106 800 6 rambus_wb_dat_o[18]
port 170 nsew signal bidirectional
rlabel metal2 s 20626 51200 20682 52000 6 rambus_wb_dat_o[19]
port 171 nsew signal bidirectional
rlabel metal3 s 0 10208 800 10328 6 rambus_wb_dat_o[1]
port 172 nsew signal bidirectional
rlabel metal2 s 15474 0 15530 800 6 rambus_wb_dat_o[20]
port 173 nsew signal bidirectional
rlabel metal2 s 30930 0 30986 800 6 rambus_wb_dat_o[21]
port 174 nsew signal bidirectional
rlabel metal3 s 0 31968 800 32088 6 rambus_wb_dat_o[22]
port 175 nsew signal bidirectional
rlabel metal3 s 49200 19728 50000 19848 6 rambus_wb_dat_o[23]
port 176 nsew signal bidirectional
rlabel metal2 s 30930 51200 30986 52000 6 rambus_wb_dat_o[24]
port 177 nsew signal bidirectional
rlabel metal3 s 0 16328 800 16448 6 rambus_wb_dat_o[25]
port 178 nsew signal bidirectional
rlabel metal2 s 23202 51200 23258 52000 6 rambus_wb_dat_o[26]
port 179 nsew signal bidirectional
rlabel metal3 s 0 28568 800 28688 6 rambus_wb_dat_o[27]
port 180 nsew signal bidirectional
rlabel metal3 s 49200 50328 50000 50448 6 rambus_wb_dat_o[28]
port 181 nsew signal bidirectional
rlabel metal3 s 0 48968 800 49088 6 rambus_wb_dat_o[29]
port 182 nsew signal bidirectional
rlabel metal2 s 31574 0 31630 800 6 rambus_wb_dat_o[2]
port 183 nsew signal bidirectional
rlabel metal3 s 49200 41488 50000 41608 6 rambus_wb_dat_o[30]
port 184 nsew signal bidirectional
rlabel metal2 s 46386 0 46442 800 6 rambus_wb_dat_o[31]
port 185 nsew signal bidirectional
rlabel metal2 s 17406 51200 17462 52000 6 rambus_wb_dat_o[3]
port 186 nsew signal bidirectional
rlabel metal3 s 0 32648 800 32768 6 rambus_wb_dat_o[4]
port 187 nsew signal bidirectional
rlabel metal2 s 32218 51200 32274 52000 6 rambus_wb_dat_o[5]
port 188 nsew signal bidirectional
rlabel metal2 s 5170 0 5226 800 6 rambus_wb_dat_o[6]
port 189 nsew signal bidirectional
rlabel metal3 s 49200 14288 50000 14408 6 rambus_wb_dat_o[7]
port 190 nsew signal bidirectional
rlabel metal2 s 23846 0 23902 800 6 rambus_wb_dat_o[8]
port 191 nsew signal bidirectional
rlabel metal2 s 12254 51200 12310 52000 6 rambus_wb_dat_o[9]
port 192 nsew signal bidirectional
rlabel metal3 s 0 8848 800 8968 6 rambus_wb_rst_o
port 193 nsew signal bidirectional
rlabel metal2 s 41234 0 41290 800 6 rambus_wb_sel_o[0]
port 194 nsew signal bidirectional
rlabel metal2 s 32862 51200 32918 52000 6 rambus_wb_sel_o[1]
port 195 nsew signal bidirectional
rlabel metal2 s 9678 51200 9734 52000 6 rambus_wb_sel_o[2]
port 196 nsew signal bidirectional
rlabel metal3 s 0 33328 800 33448 6 rambus_wb_sel_o[3]
port 197 nsew signal bidirectional
rlabel metal2 s 29642 51200 29698 52000 6 rambus_wb_stb_o
port 198 nsew signal bidirectional
rlabel metal3 s 0 4768 800 4888 6 rambus_wb_we_o
port 199 nsew signal bidirectional
rlabel metal4 s 4208 2128 4528 49552 6 vccd1
port 200 nsew power input
rlabel metal4 s 34928 2128 35248 49552 6 vccd1
port 200 nsew power input
rlabel metal4 s 19568 2128 19888 49552 6 vssd1
port 201 nsew ground input
rlabel metal3 s 49200 1368 50000 1488 6 wb_clk_i
port 202 nsew signal input
rlabel metal2 s 26422 51200 26478 52000 6 wb_rst_i
port 203 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 wbs_ack_o
port 204 nsew signal bidirectional
rlabel metal3 s 0 31288 800 31408 6 wbs_adr_i[0]
port 205 nsew signal input
rlabel metal2 s 38014 51200 38070 52000 6 wbs_adr_i[10]
port 206 nsew signal input
rlabel metal2 s 19982 51200 20038 52000 6 wbs_adr_i[11]
port 207 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 wbs_adr_i[12]
port 208 nsew signal input
rlabel metal2 s 6458 51200 6514 52000 6 wbs_adr_i[13]
port 209 nsew signal input
rlabel metal3 s 49200 27888 50000 28008 6 wbs_adr_i[14]
port 210 nsew signal input
rlabel metal3 s 0 688 800 808 6 wbs_adr_i[15]
port 211 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 wbs_adr_i[16]
port 212 nsew signal input
rlabel metal3 s 0 44208 800 44328 6 wbs_adr_i[17]
port 213 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 wbs_adr_i[18]
port 214 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 wbs_adr_i[19]
port 215 nsew signal input
rlabel metal2 s 44454 51200 44510 52000 6 wbs_adr_i[1]
port 216 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 wbs_adr_i[20]
port 217 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 wbs_adr_i[21]
port 218 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wbs_adr_i[22]
port 219 nsew signal input
rlabel metal3 s 49200 5448 50000 5568 6 wbs_adr_i[23]
port 220 nsew signal input
rlabel metal2 s 19338 51200 19394 52000 6 wbs_adr_i[24]
port 221 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_adr_i[25]
port 222 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_adr_i[26]
port 223 nsew signal input
rlabel metal2 s 28998 51200 29054 52000 6 wbs_adr_i[27]
port 224 nsew signal input
rlabel metal3 s 49200 22448 50000 22568 6 wbs_adr_i[28]
port 225 nsew signal input
rlabel metal3 s 49200 40808 50000 40928 6 wbs_adr_i[29]
port 226 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_adr_i[2]
port 227 nsew signal input
rlabel metal2 s 48962 51200 49018 52000 6 wbs_adr_i[30]
port 228 nsew signal input
rlabel metal3 s 49200 14968 50000 15088 6 wbs_adr_i[31]
port 229 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 wbs_adr_i[3]
port 230 nsew signal input
rlabel metal2 s 47674 51200 47730 52000 6 wbs_adr_i[4]
port 231 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 wbs_adr_i[5]
port 232 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 wbs_adr_i[6]
port 233 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 wbs_adr_i[7]
port 234 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 wbs_adr_i[8]
port 235 nsew signal input
rlabel metal3 s 49200 8848 50000 8968 6 wbs_adr_i[9]
port 236 nsew signal input
rlabel metal2 s 25778 51200 25834 52000 6 wbs_cyc_i
port 237 nsew signal input
rlabel metal3 s 49200 38088 50000 38208 6 wbs_dat_i[0]
port 238 nsew signal input
rlabel metal2 s 662 51200 718 52000 6 wbs_dat_i[10]
port 239 nsew signal input
rlabel metal2 s 3238 51200 3294 52000 6 wbs_dat_i[11]
port 240 nsew signal input
rlabel metal2 s 1950 51200 2006 52000 6 wbs_dat_i[12]
port 241 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wbs_dat_i[13]
port 242 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 wbs_dat_i[14]
port 243 nsew signal input
rlabel metal3 s 49200 21768 50000 21888 6 wbs_dat_i[15]
port 244 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 wbs_dat_i[16]
port 245 nsew signal input
rlabel metal2 s 41878 51200 41934 52000 6 wbs_dat_i[17]
port 246 nsew signal input
rlabel metal3 s 49200 48968 50000 49088 6 wbs_dat_i[18]
port 247 nsew signal input
rlabel metal2 s 11610 51200 11666 52000 6 wbs_dat_i[19]
port 248 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_dat_i[1]
port 249 nsew signal input
rlabel metal3 s 49200 25848 50000 25968 6 wbs_dat_i[20]
port 250 nsew signal input
rlabel metal3 s 49200 48288 50000 48408 6 wbs_dat_i[21]
port 251 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 wbs_dat_i[22]
port 252 nsew signal input
rlabel metal3 s 49200 36048 50000 36168 6 wbs_dat_i[23]
port 253 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 wbs_dat_i[24]
port 254 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 wbs_dat_i[25]
port 255 nsew signal input
rlabel metal2 s 47030 51200 47086 52000 6 wbs_dat_i[26]
port 256 nsew signal input
rlabel metal2 s 18694 51200 18750 52000 6 wbs_dat_i[27]
port 257 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_i[28]
port 258 nsew signal input
rlabel metal3 s 49200 27208 50000 27328 6 wbs_dat_i[29]
port 259 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 wbs_dat_i[2]
port 260 nsew signal input
rlabel metal3 s 49200 11568 50000 11688 6 wbs_dat_i[30]
port 261 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 wbs_dat_i[31]
port 262 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 wbs_dat_i[3]
port 263 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_dat_i[4]
port 264 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 wbs_dat_i[5]
port 265 nsew signal input
rlabel metal3 s 49200 19048 50000 19168 6 wbs_dat_i[6]
port 266 nsew signal input
rlabel metal2 s 43810 51200 43866 52000 6 wbs_dat_i[7]
port 267 nsew signal input
rlabel metal3 s 49200 42848 50000 42968 6 wbs_dat_i[8]
port 268 nsew signal input
rlabel metal3 s 49200 8 50000 128 6 wbs_dat_i[9]
port 269 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_o[0]
port 270 nsew signal bidirectional
rlabel metal3 s 49200 26528 50000 26648 6 wbs_dat_o[10]
port 271 nsew signal bidirectional
rlabel metal2 s 662 0 718 800 6 wbs_dat_o[11]
port 272 nsew signal bidirectional
rlabel metal3 s 49200 44888 50000 45008 6 wbs_dat_o[12]
port 273 nsew signal bidirectional
rlabel metal2 s 41234 51200 41290 52000 6 wbs_dat_o[13]
port 274 nsew signal bidirectional
rlabel metal3 s 49200 4088 50000 4208 6 wbs_dat_o[14]
port 275 nsew signal bidirectional
rlabel metal2 s 39302 51200 39358 52000 6 wbs_dat_o[15]
port 276 nsew signal bidirectional
rlabel metal3 s 0 19728 800 19848 6 wbs_dat_o[16]
port 277 nsew signal bidirectional
rlabel metal3 s 0 21768 800 21888 6 wbs_dat_o[17]
port 278 nsew signal bidirectional
rlabel metal2 s 32218 0 32274 800 6 wbs_dat_o[18]
port 279 nsew signal bidirectional
rlabel metal2 s 18 0 74 800 6 wbs_dat_o[19]
port 280 nsew signal bidirectional
rlabel metal2 s 38014 0 38070 800 6 wbs_dat_o[1]
port 281 nsew signal bidirectional
rlabel metal3 s 0 29248 800 29368 6 wbs_dat_o[20]
port 282 nsew signal bidirectional
rlabel metal3 s 0 4088 800 4208 6 wbs_dat_o[21]
port 283 nsew signal bidirectional
rlabel metal3 s 0 12928 800 13048 6 wbs_dat_o[22]
port 284 nsew signal bidirectional
rlabel metal3 s 0 21088 800 21208 6 wbs_dat_o[23]
port 285 nsew signal bidirectional
rlabel metal2 s 10322 0 10378 800 6 wbs_dat_o[24]
port 286 nsew signal bidirectional
rlabel metal2 s 3238 0 3294 800 6 wbs_dat_o[25]
port 287 nsew signal bidirectional
rlabel metal2 s 27710 51200 27766 52000 6 wbs_dat_o[26]
port 288 nsew signal bidirectional
rlabel metal2 s 16762 51200 16818 52000 6 wbs_dat_o[27]
port 289 nsew signal bidirectional
rlabel metal2 s 26422 0 26478 800 6 wbs_dat_o[28]
port 290 nsew signal bidirectional
rlabel metal2 s 36726 51200 36782 52000 6 wbs_dat_o[29]
port 291 nsew signal bidirectional
rlabel metal3 s 49200 12928 50000 13048 6 wbs_dat_o[2]
port 292 nsew signal bidirectional
rlabel metal3 s 0 36048 800 36168 6 wbs_dat_o[30]
port 293 nsew signal bidirectional
rlabel metal3 s 49200 39448 50000 39568 6 wbs_dat_o[31]
port 294 nsew signal bidirectional
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_o[3]
port 295 nsew signal bidirectional
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_o[4]
port 296 nsew signal bidirectional
rlabel metal3 s 0 6128 800 6248 6 wbs_dat_o[5]
port 297 nsew signal bidirectional
rlabel metal3 s 49200 37408 50000 37528 6 wbs_dat_o[6]
port 298 nsew signal bidirectional
rlabel metal2 s 29642 0 29698 800 6 wbs_dat_o[7]
port 299 nsew signal bidirectional
rlabel metal2 s 34150 51200 34206 52000 6 wbs_dat_o[8]
port 300 nsew signal bidirectional
rlabel metal2 s 33506 51200 33562 52000 6 wbs_dat_o[9]
port 301 nsew signal bidirectional
rlabel metal3 s 0 49648 800 49768 6 wbs_sel_i[0]
port 302 nsew signal input
rlabel metal2 s 5814 51200 5870 52000 6 wbs_sel_i[1]
port 303 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 wbs_sel_i[2]
port 304 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 wbs_sel_i[3]
port 305 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 wbs_stb_i
port 306 nsew signal input
rlabel metal3 s 49200 25168 50000 25288 6 wbs_we_i
port 307 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 50000 52000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3880846
string GDS_FILE /openlane/designs/wrapped_function_generator/runs/RUN_2022.05.04_10.50.24/results/finishing/wrapped_function_generator.magic.gds
string GDS_START 432158
<< end >>

